
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module LoadUnit(
  input          clock,
                 reset,
                 lsuRequest_valid,
  input  [2:0]   lsuRequest_bits_instructionInformation_nf,
  input          lsuRequest_bits_instructionInformation_mew,
  input  [1:0]   lsuRequest_bits_instructionInformation_mop,
  input  [4:0]   lsuRequest_bits_instructionInformation_lumop,
  input  [1:0]   lsuRequest_bits_instructionInformation_eew,
  input  [4:0]   lsuRequest_bits_instructionInformation_vs3,
  input          lsuRequest_bits_instructionInformation_isStore,
                 lsuRequest_bits_instructionInformation_maskedLoadStore,
  input  [31:0]  lsuRequest_bits_rs1Data,
                 lsuRequest_bits_rs2Data,
  input  [2:0]   lsuRequest_bits_instructionIndex,
  input  [10:0]  csrInterface_vl,
                 csrInterface_vStart,
  input  [2:0]   csrInterface_vlmul,
  input  [1:0]   csrInterface_vSew,
                 csrInterface_vxrm,
  input          csrInterface_vta,
                 csrInterface_vma,
  input  [63:0]  maskInput,
  output         maskSelect_valid,
  output [3:0]   maskSelect_bits,
  input          addressConflict,
                 memRequest_ready,
  output         memRequest_valid,
  output [4:0]   memRequest_bits_src,
  output [31:0]  memRequest_bits_address,
  output         memResponse_ready,
  input          memResponse_valid,
  input  [511:0] memResponse_bits_data,
  input  [4:0]   memResponse_bits_index,
  output         status_idle,
                 status_last,
  output [2:0]   status_instructionIndex,
  output         status_changeMaskGroup,
  output [31:0]  status_startAddress,
                 status_endAddress,
  input          vrfWritePort_0_ready,
  output         vrfWritePort_0_valid,
  output [4:0]   vrfWritePort_0_bits_vd,
  output         vrfWritePort_0_bits_offset,
  output [3:0]   vrfWritePort_0_bits_mask,
  output [31:0]  vrfWritePort_0_bits_data,
  output [2:0]   vrfWritePort_0_bits_instructionIndex,
  input          vrfWritePort_1_ready,
  output         vrfWritePort_1_valid,
  output [4:0]   vrfWritePort_1_bits_vd,
  output         vrfWritePort_1_bits_offset,
  output [3:0]   vrfWritePort_1_bits_mask,
  output [31:0]  vrfWritePort_1_bits_data,
  output [2:0]   vrfWritePort_1_bits_instructionIndex,
  input          vrfWritePort_2_ready,
  output         vrfWritePort_2_valid,
  output [4:0]   vrfWritePort_2_bits_vd,
  output         vrfWritePort_2_bits_offset,
  output [3:0]   vrfWritePort_2_bits_mask,
  output [31:0]  vrfWritePort_2_bits_data,
  output [2:0]   vrfWritePort_2_bits_instructionIndex,
  input          vrfWritePort_3_ready,
  output         vrfWritePort_3_valid,
  output [4:0]   vrfWritePort_3_bits_vd,
  output         vrfWritePort_3_bits_offset,
  output [3:0]   vrfWritePort_3_bits_mask,
  output [31:0]  vrfWritePort_3_bits_data,
  output [2:0]   vrfWritePort_3_bits_instructionIndex,
  input          vrfWritePort_4_ready,
  output         vrfWritePort_4_valid,
  output [4:0]   vrfWritePort_4_bits_vd,
  output         vrfWritePort_4_bits_offset,
  output [3:0]   vrfWritePort_4_bits_mask,
  output [31:0]  vrfWritePort_4_bits_data,
  output [2:0]   vrfWritePort_4_bits_instructionIndex,
  input          vrfWritePort_5_ready,
  output         vrfWritePort_5_valid,
  output [4:0]   vrfWritePort_5_bits_vd,
  output         vrfWritePort_5_bits_offset,
  output [3:0]   vrfWritePort_5_bits_mask,
  output [31:0]  vrfWritePort_5_bits_data,
  output [2:0]   vrfWritePort_5_bits_instructionIndex,
  input          vrfWritePort_6_ready,
  output         vrfWritePort_6_valid,
  output [4:0]   vrfWritePort_6_bits_vd,
  output         vrfWritePort_6_bits_offset,
  output [3:0]   vrfWritePort_6_bits_mask,
  output [31:0]  vrfWritePort_6_bits_data,
  output [2:0]   vrfWritePort_6_bits_instructionIndex,
  input          vrfWritePort_7_ready,
  output         vrfWritePort_7_valid,
  output [4:0]   vrfWritePort_7_bits_vd,
  output         vrfWritePort_7_bits_offset,
  output [3:0]   vrfWritePort_7_bits_mask,
  output [31:0]  vrfWritePort_7_bits_data,
  output [2:0]   vrfWritePort_7_bits_instructionIndex,
  input          vrfWritePort_8_ready,
  output         vrfWritePort_8_valid,
  output [4:0]   vrfWritePort_8_bits_vd,
  output         vrfWritePort_8_bits_offset,
  output [3:0]   vrfWritePort_8_bits_mask,
  output [31:0]  vrfWritePort_8_bits_data,
  output [2:0]   vrfWritePort_8_bits_instructionIndex,
  input          vrfWritePort_9_ready,
  output         vrfWritePort_9_valid,
  output [4:0]   vrfWritePort_9_bits_vd,
  output         vrfWritePort_9_bits_offset,
  output [3:0]   vrfWritePort_9_bits_mask,
  output [31:0]  vrfWritePort_9_bits_data,
  output [2:0]   vrfWritePort_9_bits_instructionIndex,
  input          vrfWritePort_10_ready,
  output         vrfWritePort_10_valid,
  output [4:0]   vrfWritePort_10_bits_vd,
  output         vrfWritePort_10_bits_offset,
  output [3:0]   vrfWritePort_10_bits_mask,
  output [31:0]  vrfWritePort_10_bits_data,
  output [2:0]   vrfWritePort_10_bits_instructionIndex,
  input          vrfWritePort_11_ready,
  output         vrfWritePort_11_valid,
  output [4:0]   vrfWritePort_11_bits_vd,
  output         vrfWritePort_11_bits_offset,
  output [3:0]   vrfWritePort_11_bits_mask,
  output [31:0]  vrfWritePort_11_bits_data,
  output [2:0]   vrfWritePort_11_bits_instructionIndex,
  input          vrfWritePort_12_ready,
  output         vrfWritePort_12_valid,
  output [4:0]   vrfWritePort_12_bits_vd,
  output         vrfWritePort_12_bits_offset,
  output [3:0]   vrfWritePort_12_bits_mask,
  output [31:0]  vrfWritePort_12_bits_data,
  output [2:0]   vrfWritePort_12_bits_instructionIndex,
  input          vrfWritePort_13_ready,
  output         vrfWritePort_13_valid,
  output [4:0]   vrfWritePort_13_bits_vd,
  output         vrfWritePort_13_bits_offset,
  output [3:0]   vrfWritePort_13_bits_mask,
  output [31:0]  vrfWritePort_13_bits_data,
  output [2:0]   vrfWritePort_13_bits_instructionIndex,
  input          vrfWritePort_14_ready,
  output         vrfWritePort_14_valid,
  output [4:0]   vrfWritePort_14_bits_vd,
  output         vrfWritePort_14_bits_offset,
  output [3:0]   vrfWritePort_14_bits_mask,
  output [31:0]  vrfWritePort_14_bits_data,
  output [2:0]   vrfWritePort_14_bits_instructionIndex,
  input          vrfWritePort_15_ready,
  output         vrfWritePort_15_valid,
  output [4:0]   vrfWritePort_15_bits_vd,
  output         vrfWritePort_15_bits_offset,
  output [3:0]   vrfWritePort_15_bits_mask,
  output [31:0]  vrfWritePort_15_bits_data,
  output [2:0]   vrfWritePort_15_bits_instructionIndex
);

  wire          memRequest_ready_0 = memRequest_ready;
  wire          memResponse_valid_0 = memResponse_valid;
  wire [511:0]  memResponse_bits_data_0 = memResponse_bits_data;
  wire [4:0]    memResponse_bits_index_0 = memResponse_bits_index;
  wire          vrfWritePort_0_ready_0 = vrfWritePort_0_ready;
  wire          vrfWritePort_1_ready_0 = vrfWritePort_1_ready;
  wire          vrfWritePort_2_ready_0 = vrfWritePort_2_ready;
  wire          vrfWritePort_3_ready_0 = vrfWritePort_3_ready;
  wire          vrfWritePort_4_ready_0 = vrfWritePort_4_ready;
  wire          vrfWritePort_5_ready_0 = vrfWritePort_5_ready;
  wire          vrfWritePort_6_ready_0 = vrfWritePort_6_ready;
  wire          vrfWritePort_7_ready_0 = vrfWritePort_7_ready;
  wire          vrfWritePort_8_ready_0 = vrfWritePort_8_ready;
  wire          vrfWritePort_9_ready_0 = vrfWritePort_9_ready;
  wire          vrfWritePort_10_ready_0 = vrfWritePort_10_ready;
  wire          vrfWritePort_11_ready_0 = vrfWritePort_11_ready;
  wire          vrfWritePort_12_ready_0 = vrfWritePort_12_ready;
  wire          vrfWritePort_13_ready_0 = vrfWritePort_13_ready;
  wire          vrfWritePort_14_ready_0 = vrfWritePort_14_ready;
  wire          vrfWritePort_15_ready_0 = vrfWritePort_15_ready;
  wire [2047:0] hi = 2048'h0;
  wire [2047:0] hi_1 = 2048'h0;
  wire [2047:0] hi_2 = 2048'h0;
  wire [2047:0] hi_3 = 2048'h0;
  wire [2047:0] hi_8 = 2048'h0;
  wire [2047:0] hi_9 = 2048'h0;
  wire [2047:0] hi_10 = 2048'h0;
  wire [2047:0] hi_11 = 2048'h0;
  wire [2047:0] hi_16 = 2048'h0;
  wire [2047:0] hi_17 = 2048'h0;
  wire [2047:0] hi_18 = 2048'h0;
  wire [2047:0] hi_19 = 2048'h0;
  wire [1023:0] lo_hi = 1024'h0;
  wire [1023:0] hi_lo = 1024'h0;
  wire [1023:0] hi_hi = 1024'h0;
  wire [1023:0] lo_hi_1 = 1024'h0;
  wire [1023:0] hi_lo_1 = 1024'h0;
  wire [1023:0] hi_hi_1 = 1024'h0;
  wire [1023:0] hi_lo_2 = 1024'h0;
  wire [1023:0] hi_hi_2 = 1024'h0;
  wire [1023:0] hi_lo_3 = 1024'h0;
  wire [1023:0] hi_hi_3 = 1024'h0;
  wire [1023:0] hi_hi_4 = 1024'h0;
  wire [1023:0] hi_hi_5 = 1024'h0;
  wire [1023:0] lo_hi_8 = 1024'h0;
  wire [1023:0] hi_lo_8 = 1024'h0;
  wire [1023:0] hi_hi_8 = 1024'h0;
  wire [1023:0] lo_hi_9 = 1024'h0;
  wire [1023:0] hi_lo_9 = 1024'h0;
  wire [1023:0] hi_hi_9 = 1024'h0;
  wire [1023:0] hi_lo_10 = 1024'h0;
  wire [1023:0] hi_hi_10 = 1024'h0;
  wire [1023:0] hi_lo_11 = 1024'h0;
  wire [1023:0] hi_hi_11 = 1024'h0;
  wire [1023:0] hi_hi_12 = 1024'h0;
  wire [1023:0] hi_hi_13 = 1024'h0;
  wire [1023:0] lo_hi_16 = 1024'h0;
  wire [1023:0] hi_lo_16 = 1024'h0;
  wire [1023:0] hi_hi_16 = 1024'h0;
  wire [1023:0] lo_hi_17 = 1024'h0;
  wire [1023:0] hi_lo_17 = 1024'h0;
  wire [1023:0] hi_hi_17 = 1024'h0;
  wire [1023:0] hi_lo_18 = 1024'h0;
  wire [1023:0] hi_hi_18 = 1024'h0;
  wire [1023:0] hi_lo_19 = 1024'h0;
  wire [1023:0] hi_hi_19 = 1024'h0;
  wire [1023:0] hi_hi_20 = 1024'h0;
  wire [1023:0] hi_hi_21 = 1024'h0;
  wire [511:0]  res_1 = 512'h0;
  wire [511:0]  res_2 = 512'h0;
  wire [511:0]  res_3 = 512'h0;
  wire [511:0]  res_4 = 512'h0;
  wire [511:0]  res_5 = 512'h0;
  wire [511:0]  res_6 = 512'h0;
  wire [511:0]  res_7 = 512'h0;
  wire [511:0]  res_10 = 512'h0;
  wire [511:0]  res_11 = 512'h0;
  wire [511:0]  res_12 = 512'h0;
  wire [511:0]  res_13 = 512'h0;
  wire [511:0]  res_14 = 512'h0;
  wire [511:0]  res_15 = 512'h0;
  wire [511:0]  res_19 = 512'h0;
  wire [511:0]  res_20 = 512'h0;
  wire [511:0]  res_21 = 512'h0;
  wire [511:0]  res_22 = 512'h0;
  wire [511:0]  res_23 = 512'h0;
  wire [511:0]  res_28 = 512'h0;
  wire [511:0]  res_29 = 512'h0;
  wire [511:0]  res_30 = 512'h0;
  wire [511:0]  res_31 = 512'h0;
  wire [511:0]  res_37 = 512'h0;
  wire [511:0]  res_38 = 512'h0;
  wire [511:0]  res_39 = 512'h0;
  wire [511:0]  res_46 = 512'h0;
  wire [511:0]  res_47 = 512'h0;
  wire [511:0]  res_55 = 512'h0;
  wire [511:0]  res_65 = 512'h0;
  wire [511:0]  res_66 = 512'h0;
  wire [511:0]  res_67 = 512'h0;
  wire [511:0]  res_68 = 512'h0;
  wire [511:0]  res_69 = 512'h0;
  wire [511:0]  res_70 = 512'h0;
  wire [511:0]  res_71 = 512'h0;
  wire [511:0]  res_74 = 512'h0;
  wire [511:0]  res_75 = 512'h0;
  wire [511:0]  res_76 = 512'h0;
  wire [511:0]  res_77 = 512'h0;
  wire [511:0]  res_78 = 512'h0;
  wire [511:0]  res_79 = 512'h0;
  wire [511:0]  res_83 = 512'h0;
  wire [511:0]  res_84 = 512'h0;
  wire [511:0]  res_85 = 512'h0;
  wire [511:0]  res_86 = 512'h0;
  wire [511:0]  res_87 = 512'h0;
  wire [511:0]  res_92 = 512'h0;
  wire [511:0]  res_93 = 512'h0;
  wire [511:0]  res_94 = 512'h0;
  wire [511:0]  res_95 = 512'h0;
  wire [511:0]  res_101 = 512'h0;
  wire [511:0]  res_102 = 512'h0;
  wire [511:0]  res_103 = 512'h0;
  wire [511:0]  res_110 = 512'h0;
  wire [511:0]  res_111 = 512'h0;
  wire [511:0]  res_119 = 512'h0;
  wire [511:0]  res_129 = 512'h0;
  wire [511:0]  res_130 = 512'h0;
  wire [511:0]  res_131 = 512'h0;
  wire [511:0]  res_132 = 512'h0;
  wire [511:0]  res_133 = 512'h0;
  wire [511:0]  res_134 = 512'h0;
  wire [511:0]  res_135 = 512'h0;
  wire [511:0]  res_138 = 512'h0;
  wire [511:0]  res_139 = 512'h0;
  wire [511:0]  res_140 = 512'h0;
  wire [511:0]  res_141 = 512'h0;
  wire [511:0]  res_142 = 512'h0;
  wire [511:0]  res_143 = 512'h0;
  wire [511:0]  res_147 = 512'h0;
  wire [511:0]  res_148 = 512'h0;
  wire [511:0]  res_149 = 512'h0;
  wire [511:0]  res_150 = 512'h0;
  wire [511:0]  res_151 = 512'h0;
  wire [511:0]  res_156 = 512'h0;
  wire [511:0]  res_157 = 512'h0;
  wire [511:0]  res_158 = 512'h0;
  wire [511:0]  res_159 = 512'h0;
  wire [511:0]  res_165 = 512'h0;
  wire [511:0]  res_166 = 512'h0;
  wire [511:0]  res_167 = 512'h0;
  wire [511:0]  res_174 = 512'h0;
  wire [511:0]  res_175 = 512'h0;
  wire [511:0]  res_183 = 512'h0;
  wire          vrfWritePort_0_bits_last = 1'h0;
  wire          vrfWritePort_1_bits_last = 1'h0;
  wire          vrfWritePort_2_bits_last = 1'h0;
  wire          vrfWritePort_3_bits_last = 1'h0;
  wire          vrfWritePort_4_bits_last = 1'h0;
  wire          vrfWritePort_5_bits_last = 1'h0;
  wire          vrfWritePort_6_bits_last = 1'h0;
  wire          vrfWritePort_7_bits_last = 1'h0;
  wire          vrfWritePort_8_bits_last = 1'h0;
  wire          vrfWritePort_9_bits_last = 1'h0;
  wire          vrfWritePort_10_bits_last = 1'h0;
  wire          vrfWritePort_11_bits_last = 1'h0;
  wire          vrfWritePort_12_bits_last = 1'h0;
  wire          vrfWritePort_13_bits_last = 1'h0;
  wire          vrfWritePort_14_bits_last = 1'h0;
  wire          vrfWritePort_15_bits_last = 1'h0;
  wire [31:0]   requestAddress;
  wire          unalignedEnqueueReady;
  reg  [2:0]    lsuRequestReg_instructionInformation_nf;
  reg           lsuRequestReg_instructionInformation_mew;
  reg  [1:0]    lsuRequestReg_instructionInformation_mop;
  reg  [4:0]    lsuRequestReg_instructionInformation_lumop;
  reg  [1:0]    lsuRequestReg_instructionInformation_eew;
  reg  [4:0]    lsuRequestReg_instructionInformation_vs3;
  reg           lsuRequestReg_instructionInformation_isStore;
  reg           lsuRequestReg_instructionInformation_maskedLoadStore;
  reg  [31:0]   lsuRequestReg_rs1Data;
  reg  [31:0]   lsuRequestReg_rs2Data;
  reg  [2:0]    lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_0_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_1_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_2_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_3_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_4_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_5_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_6_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_7_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_8_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_9_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_10_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_11_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_12_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_13_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_14_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_15_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  reg  [10:0]   csrInterfaceReg_vl;
  reg  [10:0]   csrInterfaceReg_vStart;
  reg  [2:0]    csrInterfaceReg_vlmul;
  reg  [1:0]    csrInterfaceReg_vSew;
  reg  [1:0]    csrInterfaceReg_vxrm;
  reg           csrInterfaceReg_vta;
  reg           csrInterfaceReg_vma;
  reg           requestFireNext;
  reg  [1:0]    dataEEW;
  wire [3:0]    _dataEEWOH_T = 4'h1 << dataEEW;
  wire [2:0]    dataEEWOH = _dataEEWOH_T[2:0];
  wire          isMaskType = lsuRequest_valid ? lsuRequest_bits_instructionInformation_maskedLoadStore : lsuRequestReg_instructionInformation_maskedLoadStore;
  wire [63:0]   maskAmend = isMaskType ? maskInput : 64'hFFFFFFFFFFFFFFFF;
  reg  [63:0]   maskReg;
  wire [63:0]   _lastMaskAmend_T_1 = 64'h1 << csrInterface_vl[5:0];
  wire [61:0]   _GEN = _lastMaskAmend_T_1[62:1] | _lastMaskAmend_T_1[63:2];
  wire [60:0]   _GEN_0 = _GEN[60:0] | {_lastMaskAmend_T_1[63], _GEN[61:2]};
  wire [58:0]   _GEN_1 = _GEN_0[58:0] | {_lastMaskAmend_T_1[63], _GEN[61], _GEN_0[60:4]};
  wire [54:0]   _GEN_2 = _GEN_1[54:0] | {_lastMaskAmend_T_1[63], _GEN[61], _GEN_0[60:59], _GEN_1[58:8]};
  wire [46:0]   _GEN_3 = _GEN_2[46:0] | {_lastMaskAmend_T_1[63], _GEN[61], _GEN_0[60:59], _GEN_1[58:55], _GEN_2[54:16]};
  wire [62:0]   lastMaskAmend = {_lastMaskAmend_T_1[63], _GEN[61], _GEN_0[60:59], _GEN_1[58:55], _GEN_2[54:47], _GEN_3[46:31], _GEN_3[30:0] | {_lastMaskAmend_T_1[63], _GEN[61], _GEN_0[60:59], _GEN_1[58:55], _GEN_2[54:47], _GEN_3[46:32]}};
  reg           needAmend;
  reg  [62:0]   lastMaskAmendReg;
  wire [1:0]    countEndForGroup = {1'h0, dataEEWOH[1]} | {2{dataEEWOH[2]}};
  reg  [3:0]    maskGroupCounter;
  wire [3:0]    nextMaskGroup = maskGroupCounter + 4'h1;
  reg  [1:0]    maskCounterInGroup;
  wire [1:0]    nextMaskCount = maskCounterInGroup + 2'h1;
  wire          isLastDataGroup = maskCounterInGroup == countEndForGroup;
  wire [3:0]    _maskSelect_bits_output = lsuRequest_valid ? 4'h0 : nextMaskGroup;
  reg  [63:0]   maskForGroup;
  reg           isLastMaskGroup;
  wire [63:0]   maskWire = maskReg & (needAmend & isLastMaskGroup ? {1'h0, lastMaskAmendReg} : 64'hFFFFFFFFFFFFFFFF);
  wire [3:0]    maskForGroupWire_lo_lo_lo_lo_lo = {{2{maskWire[1]}}, {2{maskWire[0]}}};
  wire [3:0]    maskForGroupWire_lo_lo_lo_lo_hi = {{2{maskWire[3]}}, {2{maskWire[2]}}};
  wire [7:0]    maskForGroupWire_lo_lo_lo_lo = {maskForGroupWire_lo_lo_lo_lo_hi, maskForGroupWire_lo_lo_lo_lo_lo};
  wire [3:0]    maskForGroupWire_lo_lo_lo_hi_lo = {{2{maskWire[5]}}, {2{maskWire[4]}}};
  wire [3:0]    maskForGroupWire_lo_lo_lo_hi_hi = {{2{maskWire[7]}}, {2{maskWire[6]}}};
  wire [7:0]    maskForGroupWire_lo_lo_lo_hi = {maskForGroupWire_lo_lo_lo_hi_hi, maskForGroupWire_lo_lo_lo_hi_lo};
  wire [15:0]   maskForGroupWire_lo_lo_lo = {maskForGroupWire_lo_lo_lo_hi, maskForGroupWire_lo_lo_lo_lo};
  wire [3:0]    maskForGroupWire_lo_lo_hi_lo_lo = {{2{maskWire[9]}}, {2{maskWire[8]}}};
  wire [3:0]    maskForGroupWire_lo_lo_hi_lo_hi = {{2{maskWire[11]}}, {2{maskWire[10]}}};
  wire [7:0]    maskForGroupWire_lo_lo_hi_lo = {maskForGroupWire_lo_lo_hi_lo_hi, maskForGroupWire_lo_lo_hi_lo_lo};
  wire [3:0]    maskForGroupWire_lo_lo_hi_hi_lo = {{2{maskWire[13]}}, {2{maskWire[12]}}};
  wire [3:0]    maskForGroupWire_lo_lo_hi_hi_hi = {{2{maskWire[15]}}, {2{maskWire[14]}}};
  wire [7:0]    maskForGroupWire_lo_lo_hi_hi = {maskForGroupWire_lo_lo_hi_hi_hi, maskForGroupWire_lo_lo_hi_hi_lo};
  wire [15:0]   maskForGroupWire_lo_lo_hi = {maskForGroupWire_lo_lo_hi_hi, maskForGroupWire_lo_lo_hi_lo};
  wire [31:0]   maskForGroupWire_lo_lo = {maskForGroupWire_lo_lo_hi, maskForGroupWire_lo_lo_lo};
  wire [3:0]    maskForGroupWire_lo_hi_lo_lo_lo = {{2{maskWire[17]}}, {2{maskWire[16]}}};
  wire [3:0]    maskForGroupWire_lo_hi_lo_lo_hi = {{2{maskWire[19]}}, {2{maskWire[18]}}};
  wire [7:0]    maskForGroupWire_lo_hi_lo_lo = {maskForGroupWire_lo_hi_lo_lo_hi, maskForGroupWire_lo_hi_lo_lo_lo};
  wire [3:0]    maskForGroupWire_lo_hi_lo_hi_lo = {{2{maskWire[21]}}, {2{maskWire[20]}}};
  wire [3:0]    maskForGroupWire_lo_hi_lo_hi_hi = {{2{maskWire[23]}}, {2{maskWire[22]}}};
  wire [7:0]    maskForGroupWire_lo_hi_lo_hi = {maskForGroupWire_lo_hi_lo_hi_hi, maskForGroupWire_lo_hi_lo_hi_lo};
  wire [15:0]   maskForGroupWire_lo_hi_lo = {maskForGroupWire_lo_hi_lo_hi, maskForGroupWire_lo_hi_lo_lo};
  wire [3:0]    maskForGroupWire_lo_hi_hi_lo_lo = {{2{maskWire[25]}}, {2{maskWire[24]}}};
  wire [3:0]    maskForGroupWire_lo_hi_hi_lo_hi = {{2{maskWire[27]}}, {2{maskWire[26]}}};
  wire [7:0]    maskForGroupWire_lo_hi_hi_lo = {maskForGroupWire_lo_hi_hi_lo_hi, maskForGroupWire_lo_hi_hi_lo_lo};
  wire [3:0]    maskForGroupWire_lo_hi_hi_hi_lo = {{2{maskWire[29]}}, {2{maskWire[28]}}};
  wire [3:0]    maskForGroupWire_lo_hi_hi_hi_hi = {{2{maskWire[31]}}, {2{maskWire[30]}}};
  wire [7:0]    maskForGroupWire_lo_hi_hi_hi = {maskForGroupWire_lo_hi_hi_hi_hi, maskForGroupWire_lo_hi_hi_hi_lo};
  wire [15:0]   maskForGroupWire_lo_hi_hi = {maskForGroupWire_lo_hi_hi_hi, maskForGroupWire_lo_hi_hi_lo};
  wire [31:0]   maskForGroupWire_lo_hi = {maskForGroupWire_lo_hi_hi, maskForGroupWire_lo_hi_lo};
  wire [63:0]   maskForGroupWire_lo = {maskForGroupWire_lo_hi, maskForGroupWire_lo_lo};
  wire [3:0]    maskForGroupWire_hi_lo_lo_lo_lo = {{2{maskWire[33]}}, {2{maskWire[32]}}};
  wire [3:0]    maskForGroupWire_hi_lo_lo_lo_hi = {{2{maskWire[35]}}, {2{maskWire[34]}}};
  wire [7:0]    maskForGroupWire_hi_lo_lo_lo = {maskForGroupWire_hi_lo_lo_lo_hi, maskForGroupWire_hi_lo_lo_lo_lo};
  wire [3:0]    maskForGroupWire_hi_lo_lo_hi_lo = {{2{maskWire[37]}}, {2{maskWire[36]}}};
  wire [3:0]    maskForGroupWire_hi_lo_lo_hi_hi = {{2{maskWire[39]}}, {2{maskWire[38]}}};
  wire [7:0]    maskForGroupWire_hi_lo_lo_hi = {maskForGroupWire_hi_lo_lo_hi_hi, maskForGroupWire_hi_lo_lo_hi_lo};
  wire [15:0]   maskForGroupWire_hi_lo_lo = {maskForGroupWire_hi_lo_lo_hi, maskForGroupWire_hi_lo_lo_lo};
  wire [3:0]    maskForGroupWire_hi_lo_hi_lo_lo = {{2{maskWire[41]}}, {2{maskWire[40]}}};
  wire [3:0]    maskForGroupWire_hi_lo_hi_lo_hi = {{2{maskWire[43]}}, {2{maskWire[42]}}};
  wire [7:0]    maskForGroupWire_hi_lo_hi_lo = {maskForGroupWire_hi_lo_hi_lo_hi, maskForGroupWire_hi_lo_hi_lo_lo};
  wire [3:0]    maskForGroupWire_hi_lo_hi_hi_lo = {{2{maskWire[45]}}, {2{maskWire[44]}}};
  wire [3:0]    maskForGroupWire_hi_lo_hi_hi_hi = {{2{maskWire[47]}}, {2{maskWire[46]}}};
  wire [7:0]    maskForGroupWire_hi_lo_hi_hi = {maskForGroupWire_hi_lo_hi_hi_hi, maskForGroupWire_hi_lo_hi_hi_lo};
  wire [15:0]   maskForGroupWire_hi_lo_hi = {maskForGroupWire_hi_lo_hi_hi, maskForGroupWire_hi_lo_hi_lo};
  wire [31:0]   maskForGroupWire_hi_lo = {maskForGroupWire_hi_lo_hi, maskForGroupWire_hi_lo_lo};
  wire [3:0]    maskForGroupWire_hi_hi_lo_lo_lo = {{2{maskWire[49]}}, {2{maskWire[48]}}};
  wire [3:0]    maskForGroupWire_hi_hi_lo_lo_hi = {{2{maskWire[51]}}, {2{maskWire[50]}}};
  wire [7:0]    maskForGroupWire_hi_hi_lo_lo = {maskForGroupWire_hi_hi_lo_lo_hi, maskForGroupWire_hi_hi_lo_lo_lo};
  wire [3:0]    maskForGroupWire_hi_hi_lo_hi_lo = {{2{maskWire[53]}}, {2{maskWire[52]}}};
  wire [3:0]    maskForGroupWire_hi_hi_lo_hi_hi = {{2{maskWire[55]}}, {2{maskWire[54]}}};
  wire [7:0]    maskForGroupWire_hi_hi_lo_hi = {maskForGroupWire_hi_hi_lo_hi_hi, maskForGroupWire_hi_hi_lo_hi_lo};
  wire [15:0]   maskForGroupWire_hi_hi_lo = {maskForGroupWire_hi_hi_lo_hi, maskForGroupWire_hi_hi_lo_lo};
  wire [3:0]    maskForGroupWire_hi_hi_hi_lo_lo = {{2{maskWire[57]}}, {2{maskWire[56]}}};
  wire [3:0]    maskForGroupWire_hi_hi_hi_lo_hi = {{2{maskWire[59]}}, {2{maskWire[58]}}};
  wire [7:0]    maskForGroupWire_hi_hi_hi_lo = {maskForGroupWire_hi_hi_hi_lo_hi, maskForGroupWire_hi_hi_hi_lo_lo};
  wire [3:0]    maskForGroupWire_hi_hi_hi_hi_lo = {{2{maskWire[61]}}, {2{maskWire[60]}}};
  wire [3:0]    maskForGroupWire_hi_hi_hi_hi_hi = {{2{maskWire[63]}}, {2{maskWire[62]}}};
  wire [7:0]    maskForGroupWire_hi_hi_hi_hi = {maskForGroupWire_hi_hi_hi_hi_hi, maskForGroupWire_hi_hi_hi_hi_lo};
  wire [15:0]   maskForGroupWire_hi_hi_hi = {maskForGroupWire_hi_hi_hi_hi, maskForGroupWire_hi_hi_hi_lo};
  wire [31:0]   maskForGroupWire_hi_hi = {maskForGroupWire_hi_hi_hi, maskForGroupWire_hi_hi_lo};
  wire [63:0]   maskForGroupWire_hi = {maskForGroupWire_hi_hi, maskForGroupWire_hi_lo};
  wire [3:0]    maskForGroupWire_lo_lo_lo_lo_lo_1 = {{2{maskWire[1]}}, {2{maskWire[0]}}};
  wire [3:0]    maskForGroupWire_lo_lo_lo_lo_hi_1 = {{2{maskWire[3]}}, {2{maskWire[2]}}};
  wire [7:0]    maskForGroupWire_lo_lo_lo_lo_1 = {maskForGroupWire_lo_lo_lo_lo_hi_1, maskForGroupWire_lo_lo_lo_lo_lo_1};
  wire [3:0]    maskForGroupWire_lo_lo_lo_hi_lo_1 = {{2{maskWire[5]}}, {2{maskWire[4]}}};
  wire [3:0]    maskForGroupWire_lo_lo_lo_hi_hi_1 = {{2{maskWire[7]}}, {2{maskWire[6]}}};
  wire [7:0]    maskForGroupWire_lo_lo_lo_hi_1 = {maskForGroupWire_lo_lo_lo_hi_hi_1, maskForGroupWire_lo_lo_lo_hi_lo_1};
  wire [15:0]   maskForGroupWire_lo_lo_lo_1 = {maskForGroupWire_lo_lo_lo_hi_1, maskForGroupWire_lo_lo_lo_lo_1};
  wire [3:0]    maskForGroupWire_lo_lo_hi_lo_lo_1 = {{2{maskWire[9]}}, {2{maskWire[8]}}};
  wire [3:0]    maskForGroupWire_lo_lo_hi_lo_hi_1 = {{2{maskWire[11]}}, {2{maskWire[10]}}};
  wire [7:0]    maskForGroupWire_lo_lo_hi_lo_1 = {maskForGroupWire_lo_lo_hi_lo_hi_1, maskForGroupWire_lo_lo_hi_lo_lo_1};
  wire [3:0]    maskForGroupWire_lo_lo_hi_hi_lo_1 = {{2{maskWire[13]}}, {2{maskWire[12]}}};
  wire [3:0]    maskForGroupWire_lo_lo_hi_hi_hi_1 = {{2{maskWire[15]}}, {2{maskWire[14]}}};
  wire [7:0]    maskForGroupWire_lo_lo_hi_hi_1 = {maskForGroupWire_lo_lo_hi_hi_hi_1, maskForGroupWire_lo_lo_hi_hi_lo_1};
  wire [15:0]   maskForGroupWire_lo_lo_hi_1 = {maskForGroupWire_lo_lo_hi_hi_1, maskForGroupWire_lo_lo_hi_lo_1};
  wire [31:0]   maskForGroupWire_lo_lo_1 = {maskForGroupWire_lo_lo_hi_1, maskForGroupWire_lo_lo_lo_1};
  wire [3:0]    maskForGroupWire_lo_hi_lo_lo_lo_1 = {{2{maskWire[17]}}, {2{maskWire[16]}}};
  wire [3:0]    maskForGroupWire_lo_hi_lo_lo_hi_1 = {{2{maskWire[19]}}, {2{maskWire[18]}}};
  wire [7:0]    maskForGroupWire_lo_hi_lo_lo_1 = {maskForGroupWire_lo_hi_lo_lo_hi_1, maskForGroupWire_lo_hi_lo_lo_lo_1};
  wire [3:0]    maskForGroupWire_lo_hi_lo_hi_lo_1 = {{2{maskWire[21]}}, {2{maskWire[20]}}};
  wire [3:0]    maskForGroupWire_lo_hi_lo_hi_hi_1 = {{2{maskWire[23]}}, {2{maskWire[22]}}};
  wire [7:0]    maskForGroupWire_lo_hi_lo_hi_1 = {maskForGroupWire_lo_hi_lo_hi_hi_1, maskForGroupWire_lo_hi_lo_hi_lo_1};
  wire [15:0]   maskForGroupWire_lo_hi_lo_1 = {maskForGroupWire_lo_hi_lo_hi_1, maskForGroupWire_lo_hi_lo_lo_1};
  wire [3:0]    maskForGroupWire_lo_hi_hi_lo_lo_1 = {{2{maskWire[25]}}, {2{maskWire[24]}}};
  wire [3:0]    maskForGroupWire_lo_hi_hi_lo_hi_1 = {{2{maskWire[27]}}, {2{maskWire[26]}}};
  wire [7:0]    maskForGroupWire_lo_hi_hi_lo_1 = {maskForGroupWire_lo_hi_hi_lo_hi_1, maskForGroupWire_lo_hi_hi_lo_lo_1};
  wire [3:0]    maskForGroupWire_lo_hi_hi_hi_lo_1 = {{2{maskWire[29]}}, {2{maskWire[28]}}};
  wire [3:0]    maskForGroupWire_lo_hi_hi_hi_hi_1 = {{2{maskWire[31]}}, {2{maskWire[30]}}};
  wire [7:0]    maskForGroupWire_lo_hi_hi_hi_1 = {maskForGroupWire_lo_hi_hi_hi_hi_1, maskForGroupWire_lo_hi_hi_hi_lo_1};
  wire [15:0]   maskForGroupWire_lo_hi_hi_1 = {maskForGroupWire_lo_hi_hi_hi_1, maskForGroupWire_lo_hi_hi_lo_1};
  wire [31:0]   maskForGroupWire_lo_hi_1 = {maskForGroupWire_lo_hi_hi_1, maskForGroupWire_lo_hi_lo_1};
  wire [63:0]   maskForGroupWire_lo_1 = {maskForGroupWire_lo_hi_1, maskForGroupWire_lo_lo_1};
  wire [3:0]    maskForGroupWire_hi_lo_lo_lo_lo_1 = {{2{maskWire[33]}}, {2{maskWire[32]}}};
  wire [3:0]    maskForGroupWire_hi_lo_lo_lo_hi_1 = {{2{maskWire[35]}}, {2{maskWire[34]}}};
  wire [7:0]    maskForGroupWire_hi_lo_lo_lo_1 = {maskForGroupWire_hi_lo_lo_lo_hi_1, maskForGroupWire_hi_lo_lo_lo_lo_1};
  wire [3:0]    maskForGroupWire_hi_lo_lo_hi_lo_1 = {{2{maskWire[37]}}, {2{maskWire[36]}}};
  wire [3:0]    maskForGroupWire_hi_lo_lo_hi_hi_1 = {{2{maskWire[39]}}, {2{maskWire[38]}}};
  wire [7:0]    maskForGroupWire_hi_lo_lo_hi_1 = {maskForGroupWire_hi_lo_lo_hi_hi_1, maskForGroupWire_hi_lo_lo_hi_lo_1};
  wire [15:0]   maskForGroupWire_hi_lo_lo_1 = {maskForGroupWire_hi_lo_lo_hi_1, maskForGroupWire_hi_lo_lo_lo_1};
  wire [3:0]    maskForGroupWire_hi_lo_hi_lo_lo_1 = {{2{maskWire[41]}}, {2{maskWire[40]}}};
  wire [3:0]    maskForGroupWire_hi_lo_hi_lo_hi_1 = {{2{maskWire[43]}}, {2{maskWire[42]}}};
  wire [7:0]    maskForGroupWire_hi_lo_hi_lo_1 = {maskForGroupWire_hi_lo_hi_lo_hi_1, maskForGroupWire_hi_lo_hi_lo_lo_1};
  wire [3:0]    maskForGroupWire_hi_lo_hi_hi_lo_1 = {{2{maskWire[45]}}, {2{maskWire[44]}}};
  wire [3:0]    maskForGroupWire_hi_lo_hi_hi_hi_1 = {{2{maskWire[47]}}, {2{maskWire[46]}}};
  wire [7:0]    maskForGroupWire_hi_lo_hi_hi_1 = {maskForGroupWire_hi_lo_hi_hi_hi_1, maskForGroupWire_hi_lo_hi_hi_lo_1};
  wire [15:0]   maskForGroupWire_hi_lo_hi_1 = {maskForGroupWire_hi_lo_hi_hi_1, maskForGroupWire_hi_lo_hi_lo_1};
  wire [31:0]   maskForGroupWire_hi_lo_1 = {maskForGroupWire_hi_lo_hi_1, maskForGroupWire_hi_lo_lo_1};
  wire [3:0]    maskForGroupWire_hi_hi_lo_lo_lo_1 = {{2{maskWire[49]}}, {2{maskWire[48]}}};
  wire [3:0]    maskForGroupWire_hi_hi_lo_lo_hi_1 = {{2{maskWire[51]}}, {2{maskWire[50]}}};
  wire [7:0]    maskForGroupWire_hi_hi_lo_lo_1 = {maskForGroupWire_hi_hi_lo_lo_hi_1, maskForGroupWire_hi_hi_lo_lo_lo_1};
  wire [3:0]    maskForGroupWire_hi_hi_lo_hi_lo_1 = {{2{maskWire[53]}}, {2{maskWire[52]}}};
  wire [3:0]    maskForGroupWire_hi_hi_lo_hi_hi_1 = {{2{maskWire[55]}}, {2{maskWire[54]}}};
  wire [7:0]    maskForGroupWire_hi_hi_lo_hi_1 = {maskForGroupWire_hi_hi_lo_hi_hi_1, maskForGroupWire_hi_hi_lo_hi_lo_1};
  wire [15:0]   maskForGroupWire_hi_hi_lo_1 = {maskForGroupWire_hi_hi_lo_hi_1, maskForGroupWire_hi_hi_lo_lo_1};
  wire [3:0]    maskForGroupWire_hi_hi_hi_lo_lo_1 = {{2{maskWire[57]}}, {2{maskWire[56]}}};
  wire [3:0]    maskForGroupWire_hi_hi_hi_lo_hi_1 = {{2{maskWire[59]}}, {2{maskWire[58]}}};
  wire [7:0]    maskForGroupWire_hi_hi_hi_lo_1 = {maskForGroupWire_hi_hi_hi_lo_hi_1, maskForGroupWire_hi_hi_hi_lo_lo_1};
  wire [3:0]    maskForGroupWire_hi_hi_hi_hi_lo_1 = {{2{maskWire[61]}}, {2{maskWire[60]}}};
  wire [3:0]    maskForGroupWire_hi_hi_hi_hi_hi_1 = {{2{maskWire[63]}}, {2{maskWire[62]}}};
  wire [7:0]    maskForGroupWire_hi_hi_hi_hi_1 = {maskForGroupWire_hi_hi_hi_hi_hi_1, maskForGroupWire_hi_hi_hi_hi_lo_1};
  wire [15:0]   maskForGroupWire_hi_hi_hi_1 = {maskForGroupWire_hi_hi_hi_hi_1, maskForGroupWire_hi_hi_hi_lo_1};
  wire [31:0]   maskForGroupWire_hi_hi_1 = {maskForGroupWire_hi_hi_hi_1, maskForGroupWire_hi_hi_lo_1};
  wire [63:0]   maskForGroupWire_hi_1 = {maskForGroupWire_hi_hi_1, maskForGroupWire_hi_lo_1};
  wire [3:0]    _maskForGroupWire_T_261 = 4'h1 << maskCounterInGroup;
  wire [7:0]    maskForGroupWire_lo_lo_lo_lo_lo_2 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]    maskForGroupWire_lo_lo_lo_lo_hi_2 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]   maskForGroupWire_lo_lo_lo_lo_2 = {maskForGroupWire_lo_lo_lo_lo_hi_2, maskForGroupWire_lo_lo_lo_lo_lo_2};
  wire [7:0]    maskForGroupWire_lo_lo_lo_hi_lo_2 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]    maskForGroupWire_lo_lo_lo_hi_hi_2 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]   maskForGroupWire_lo_lo_lo_hi_2 = {maskForGroupWire_lo_lo_lo_hi_hi_2, maskForGroupWire_lo_lo_lo_hi_lo_2};
  wire [31:0]   maskForGroupWire_lo_lo_lo_2 = {maskForGroupWire_lo_lo_lo_hi_2, maskForGroupWire_lo_lo_lo_lo_2};
  wire [7:0]    maskForGroupWire_lo_lo_hi_lo_lo_2 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]    maskForGroupWire_lo_lo_hi_lo_hi_2 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]   maskForGroupWire_lo_lo_hi_lo_2 = {maskForGroupWire_lo_lo_hi_lo_hi_2, maskForGroupWire_lo_lo_hi_lo_lo_2};
  wire [7:0]    maskForGroupWire_lo_lo_hi_hi_lo_2 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]    maskForGroupWire_lo_lo_hi_hi_hi_2 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]   maskForGroupWire_lo_lo_hi_hi_2 = {maskForGroupWire_lo_lo_hi_hi_hi_2, maskForGroupWire_lo_lo_hi_hi_lo_2};
  wire [31:0]   maskForGroupWire_lo_lo_hi_2 = {maskForGroupWire_lo_lo_hi_hi_2, maskForGroupWire_lo_lo_hi_lo_2};
  wire [63:0]   maskForGroupWire_lo_lo_2 = {maskForGroupWire_lo_lo_hi_2, maskForGroupWire_lo_lo_lo_2};
  wire [7:0]    maskForGroupWire_lo_hi_lo_lo_lo_2 = {{4{maskWire[17]}}, {4{maskWire[16]}}};
  wire [7:0]    maskForGroupWire_lo_hi_lo_lo_hi_2 = {{4{maskWire[19]}}, {4{maskWire[18]}}};
  wire [15:0]   maskForGroupWire_lo_hi_lo_lo_2 = {maskForGroupWire_lo_hi_lo_lo_hi_2, maskForGroupWire_lo_hi_lo_lo_lo_2};
  wire [7:0]    maskForGroupWire_lo_hi_lo_hi_lo_2 = {{4{maskWire[21]}}, {4{maskWire[20]}}};
  wire [7:0]    maskForGroupWire_lo_hi_lo_hi_hi_2 = {{4{maskWire[23]}}, {4{maskWire[22]}}};
  wire [15:0]   maskForGroupWire_lo_hi_lo_hi_2 = {maskForGroupWire_lo_hi_lo_hi_hi_2, maskForGroupWire_lo_hi_lo_hi_lo_2};
  wire [31:0]   maskForGroupWire_lo_hi_lo_2 = {maskForGroupWire_lo_hi_lo_hi_2, maskForGroupWire_lo_hi_lo_lo_2};
  wire [7:0]    maskForGroupWire_lo_hi_hi_lo_lo_2 = {{4{maskWire[25]}}, {4{maskWire[24]}}};
  wire [7:0]    maskForGroupWire_lo_hi_hi_lo_hi_2 = {{4{maskWire[27]}}, {4{maskWire[26]}}};
  wire [15:0]   maskForGroupWire_lo_hi_hi_lo_2 = {maskForGroupWire_lo_hi_hi_lo_hi_2, maskForGroupWire_lo_hi_hi_lo_lo_2};
  wire [7:0]    maskForGroupWire_lo_hi_hi_hi_lo_2 = {{4{maskWire[29]}}, {4{maskWire[28]}}};
  wire [7:0]    maskForGroupWire_lo_hi_hi_hi_hi_2 = {{4{maskWire[31]}}, {4{maskWire[30]}}};
  wire [15:0]   maskForGroupWire_lo_hi_hi_hi_2 = {maskForGroupWire_lo_hi_hi_hi_hi_2, maskForGroupWire_lo_hi_hi_hi_lo_2};
  wire [31:0]   maskForGroupWire_lo_hi_hi_2 = {maskForGroupWire_lo_hi_hi_hi_2, maskForGroupWire_lo_hi_hi_lo_2};
  wire [63:0]   maskForGroupWire_lo_hi_2 = {maskForGroupWire_lo_hi_hi_2, maskForGroupWire_lo_hi_lo_2};
  wire [127:0]  maskForGroupWire_lo_2 = {maskForGroupWire_lo_hi_2, maskForGroupWire_lo_lo_2};
  wire [7:0]    maskForGroupWire_hi_lo_lo_lo_lo_2 = {{4{maskWire[33]}}, {4{maskWire[32]}}};
  wire [7:0]    maskForGroupWire_hi_lo_lo_lo_hi_2 = {{4{maskWire[35]}}, {4{maskWire[34]}}};
  wire [15:0]   maskForGroupWire_hi_lo_lo_lo_2 = {maskForGroupWire_hi_lo_lo_lo_hi_2, maskForGroupWire_hi_lo_lo_lo_lo_2};
  wire [7:0]    maskForGroupWire_hi_lo_lo_hi_lo_2 = {{4{maskWire[37]}}, {4{maskWire[36]}}};
  wire [7:0]    maskForGroupWire_hi_lo_lo_hi_hi_2 = {{4{maskWire[39]}}, {4{maskWire[38]}}};
  wire [15:0]   maskForGroupWire_hi_lo_lo_hi_2 = {maskForGroupWire_hi_lo_lo_hi_hi_2, maskForGroupWire_hi_lo_lo_hi_lo_2};
  wire [31:0]   maskForGroupWire_hi_lo_lo_2 = {maskForGroupWire_hi_lo_lo_hi_2, maskForGroupWire_hi_lo_lo_lo_2};
  wire [7:0]    maskForGroupWire_hi_lo_hi_lo_lo_2 = {{4{maskWire[41]}}, {4{maskWire[40]}}};
  wire [7:0]    maskForGroupWire_hi_lo_hi_lo_hi_2 = {{4{maskWire[43]}}, {4{maskWire[42]}}};
  wire [15:0]   maskForGroupWire_hi_lo_hi_lo_2 = {maskForGroupWire_hi_lo_hi_lo_hi_2, maskForGroupWire_hi_lo_hi_lo_lo_2};
  wire [7:0]    maskForGroupWire_hi_lo_hi_hi_lo_2 = {{4{maskWire[45]}}, {4{maskWire[44]}}};
  wire [7:0]    maskForGroupWire_hi_lo_hi_hi_hi_2 = {{4{maskWire[47]}}, {4{maskWire[46]}}};
  wire [15:0]   maskForGroupWire_hi_lo_hi_hi_2 = {maskForGroupWire_hi_lo_hi_hi_hi_2, maskForGroupWire_hi_lo_hi_hi_lo_2};
  wire [31:0]   maskForGroupWire_hi_lo_hi_2 = {maskForGroupWire_hi_lo_hi_hi_2, maskForGroupWire_hi_lo_hi_lo_2};
  wire [63:0]   maskForGroupWire_hi_lo_2 = {maskForGroupWire_hi_lo_hi_2, maskForGroupWire_hi_lo_lo_2};
  wire [7:0]    maskForGroupWire_hi_hi_lo_lo_lo_2 = {{4{maskWire[49]}}, {4{maskWire[48]}}};
  wire [7:0]    maskForGroupWire_hi_hi_lo_lo_hi_2 = {{4{maskWire[51]}}, {4{maskWire[50]}}};
  wire [15:0]   maskForGroupWire_hi_hi_lo_lo_2 = {maskForGroupWire_hi_hi_lo_lo_hi_2, maskForGroupWire_hi_hi_lo_lo_lo_2};
  wire [7:0]    maskForGroupWire_hi_hi_lo_hi_lo_2 = {{4{maskWire[53]}}, {4{maskWire[52]}}};
  wire [7:0]    maskForGroupWire_hi_hi_lo_hi_hi_2 = {{4{maskWire[55]}}, {4{maskWire[54]}}};
  wire [15:0]   maskForGroupWire_hi_hi_lo_hi_2 = {maskForGroupWire_hi_hi_lo_hi_hi_2, maskForGroupWire_hi_hi_lo_hi_lo_2};
  wire [31:0]   maskForGroupWire_hi_hi_lo_2 = {maskForGroupWire_hi_hi_lo_hi_2, maskForGroupWire_hi_hi_lo_lo_2};
  wire [7:0]    maskForGroupWire_hi_hi_hi_lo_lo_2 = {{4{maskWire[57]}}, {4{maskWire[56]}}};
  wire [7:0]    maskForGroupWire_hi_hi_hi_lo_hi_2 = {{4{maskWire[59]}}, {4{maskWire[58]}}};
  wire [15:0]   maskForGroupWire_hi_hi_hi_lo_2 = {maskForGroupWire_hi_hi_hi_lo_hi_2, maskForGroupWire_hi_hi_hi_lo_lo_2};
  wire [7:0]    maskForGroupWire_hi_hi_hi_hi_lo_2 = {{4{maskWire[61]}}, {4{maskWire[60]}}};
  wire [7:0]    maskForGroupWire_hi_hi_hi_hi_hi_2 = {{4{maskWire[63]}}, {4{maskWire[62]}}};
  wire [15:0]   maskForGroupWire_hi_hi_hi_hi_2 = {maskForGroupWire_hi_hi_hi_hi_hi_2, maskForGroupWire_hi_hi_hi_hi_lo_2};
  wire [31:0]   maskForGroupWire_hi_hi_hi_2 = {maskForGroupWire_hi_hi_hi_hi_2, maskForGroupWire_hi_hi_hi_lo_2};
  wire [63:0]   maskForGroupWire_hi_hi_2 = {maskForGroupWire_hi_hi_hi_2, maskForGroupWire_hi_hi_lo_2};
  wire [127:0]  maskForGroupWire_hi_2 = {maskForGroupWire_hi_hi_2, maskForGroupWire_hi_lo_2};
  wire [7:0]    maskForGroupWire_lo_lo_lo_lo_lo_3 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]    maskForGroupWire_lo_lo_lo_lo_hi_3 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]   maskForGroupWire_lo_lo_lo_lo_3 = {maskForGroupWire_lo_lo_lo_lo_hi_3, maskForGroupWire_lo_lo_lo_lo_lo_3};
  wire [7:0]    maskForGroupWire_lo_lo_lo_hi_lo_3 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]    maskForGroupWire_lo_lo_lo_hi_hi_3 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]   maskForGroupWire_lo_lo_lo_hi_3 = {maskForGroupWire_lo_lo_lo_hi_hi_3, maskForGroupWire_lo_lo_lo_hi_lo_3};
  wire [31:0]   maskForGroupWire_lo_lo_lo_3 = {maskForGroupWire_lo_lo_lo_hi_3, maskForGroupWire_lo_lo_lo_lo_3};
  wire [7:0]    maskForGroupWire_lo_lo_hi_lo_lo_3 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]    maskForGroupWire_lo_lo_hi_lo_hi_3 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]   maskForGroupWire_lo_lo_hi_lo_3 = {maskForGroupWire_lo_lo_hi_lo_hi_3, maskForGroupWire_lo_lo_hi_lo_lo_3};
  wire [7:0]    maskForGroupWire_lo_lo_hi_hi_lo_3 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]    maskForGroupWire_lo_lo_hi_hi_hi_3 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]   maskForGroupWire_lo_lo_hi_hi_3 = {maskForGroupWire_lo_lo_hi_hi_hi_3, maskForGroupWire_lo_lo_hi_hi_lo_3};
  wire [31:0]   maskForGroupWire_lo_lo_hi_3 = {maskForGroupWire_lo_lo_hi_hi_3, maskForGroupWire_lo_lo_hi_lo_3};
  wire [63:0]   maskForGroupWire_lo_lo_3 = {maskForGroupWire_lo_lo_hi_3, maskForGroupWire_lo_lo_lo_3};
  wire [7:0]    maskForGroupWire_lo_hi_lo_lo_lo_3 = {{4{maskWire[17]}}, {4{maskWire[16]}}};
  wire [7:0]    maskForGroupWire_lo_hi_lo_lo_hi_3 = {{4{maskWire[19]}}, {4{maskWire[18]}}};
  wire [15:0]   maskForGroupWire_lo_hi_lo_lo_3 = {maskForGroupWire_lo_hi_lo_lo_hi_3, maskForGroupWire_lo_hi_lo_lo_lo_3};
  wire [7:0]    maskForGroupWire_lo_hi_lo_hi_lo_3 = {{4{maskWire[21]}}, {4{maskWire[20]}}};
  wire [7:0]    maskForGroupWire_lo_hi_lo_hi_hi_3 = {{4{maskWire[23]}}, {4{maskWire[22]}}};
  wire [15:0]   maskForGroupWire_lo_hi_lo_hi_3 = {maskForGroupWire_lo_hi_lo_hi_hi_3, maskForGroupWire_lo_hi_lo_hi_lo_3};
  wire [31:0]   maskForGroupWire_lo_hi_lo_3 = {maskForGroupWire_lo_hi_lo_hi_3, maskForGroupWire_lo_hi_lo_lo_3};
  wire [7:0]    maskForGroupWire_lo_hi_hi_lo_lo_3 = {{4{maskWire[25]}}, {4{maskWire[24]}}};
  wire [7:0]    maskForGroupWire_lo_hi_hi_lo_hi_3 = {{4{maskWire[27]}}, {4{maskWire[26]}}};
  wire [15:0]   maskForGroupWire_lo_hi_hi_lo_3 = {maskForGroupWire_lo_hi_hi_lo_hi_3, maskForGroupWire_lo_hi_hi_lo_lo_3};
  wire [7:0]    maskForGroupWire_lo_hi_hi_hi_lo_3 = {{4{maskWire[29]}}, {4{maskWire[28]}}};
  wire [7:0]    maskForGroupWire_lo_hi_hi_hi_hi_3 = {{4{maskWire[31]}}, {4{maskWire[30]}}};
  wire [15:0]   maskForGroupWire_lo_hi_hi_hi_3 = {maskForGroupWire_lo_hi_hi_hi_hi_3, maskForGroupWire_lo_hi_hi_hi_lo_3};
  wire [31:0]   maskForGroupWire_lo_hi_hi_3 = {maskForGroupWire_lo_hi_hi_hi_3, maskForGroupWire_lo_hi_hi_lo_3};
  wire [63:0]   maskForGroupWire_lo_hi_3 = {maskForGroupWire_lo_hi_hi_3, maskForGroupWire_lo_hi_lo_3};
  wire [127:0]  maskForGroupWire_lo_3 = {maskForGroupWire_lo_hi_3, maskForGroupWire_lo_lo_3};
  wire [7:0]    maskForGroupWire_hi_lo_lo_lo_lo_3 = {{4{maskWire[33]}}, {4{maskWire[32]}}};
  wire [7:0]    maskForGroupWire_hi_lo_lo_lo_hi_3 = {{4{maskWire[35]}}, {4{maskWire[34]}}};
  wire [15:0]   maskForGroupWire_hi_lo_lo_lo_3 = {maskForGroupWire_hi_lo_lo_lo_hi_3, maskForGroupWire_hi_lo_lo_lo_lo_3};
  wire [7:0]    maskForGroupWire_hi_lo_lo_hi_lo_3 = {{4{maskWire[37]}}, {4{maskWire[36]}}};
  wire [7:0]    maskForGroupWire_hi_lo_lo_hi_hi_3 = {{4{maskWire[39]}}, {4{maskWire[38]}}};
  wire [15:0]   maskForGroupWire_hi_lo_lo_hi_3 = {maskForGroupWire_hi_lo_lo_hi_hi_3, maskForGroupWire_hi_lo_lo_hi_lo_3};
  wire [31:0]   maskForGroupWire_hi_lo_lo_3 = {maskForGroupWire_hi_lo_lo_hi_3, maskForGroupWire_hi_lo_lo_lo_3};
  wire [7:0]    maskForGroupWire_hi_lo_hi_lo_lo_3 = {{4{maskWire[41]}}, {4{maskWire[40]}}};
  wire [7:0]    maskForGroupWire_hi_lo_hi_lo_hi_3 = {{4{maskWire[43]}}, {4{maskWire[42]}}};
  wire [15:0]   maskForGroupWire_hi_lo_hi_lo_3 = {maskForGroupWire_hi_lo_hi_lo_hi_3, maskForGroupWire_hi_lo_hi_lo_lo_3};
  wire [7:0]    maskForGroupWire_hi_lo_hi_hi_lo_3 = {{4{maskWire[45]}}, {4{maskWire[44]}}};
  wire [7:0]    maskForGroupWire_hi_lo_hi_hi_hi_3 = {{4{maskWire[47]}}, {4{maskWire[46]}}};
  wire [15:0]   maskForGroupWire_hi_lo_hi_hi_3 = {maskForGroupWire_hi_lo_hi_hi_hi_3, maskForGroupWire_hi_lo_hi_hi_lo_3};
  wire [31:0]   maskForGroupWire_hi_lo_hi_3 = {maskForGroupWire_hi_lo_hi_hi_3, maskForGroupWire_hi_lo_hi_lo_3};
  wire [63:0]   maskForGroupWire_hi_lo_3 = {maskForGroupWire_hi_lo_hi_3, maskForGroupWire_hi_lo_lo_3};
  wire [7:0]    maskForGroupWire_hi_hi_lo_lo_lo_3 = {{4{maskWire[49]}}, {4{maskWire[48]}}};
  wire [7:0]    maskForGroupWire_hi_hi_lo_lo_hi_3 = {{4{maskWire[51]}}, {4{maskWire[50]}}};
  wire [15:0]   maskForGroupWire_hi_hi_lo_lo_3 = {maskForGroupWire_hi_hi_lo_lo_hi_3, maskForGroupWire_hi_hi_lo_lo_lo_3};
  wire [7:0]    maskForGroupWire_hi_hi_lo_hi_lo_3 = {{4{maskWire[53]}}, {4{maskWire[52]}}};
  wire [7:0]    maskForGroupWire_hi_hi_lo_hi_hi_3 = {{4{maskWire[55]}}, {4{maskWire[54]}}};
  wire [15:0]   maskForGroupWire_hi_hi_lo_hi_3 = {maskForGroupWire_hi_hi_lo_hi_hi_3, maskForGroupWire_hi_hi_lo_hi_lo_3};
  wire [31:0]   maskForGroupWire_hi_hi_lo_3 = {maskForGroupWire_hi_hi_lo_hi_3, maskForGroupWire_hi_hi_lo_lo_3};
  wire [7:0]    maskForGroupWire_hi_hi_hi_lo_lo_3 = {{4{maskWire[57]}}, {4{maskWire[56]}}};
  wire [7:0]    maskForGroupWire_hi_hi_hi_lo_hi_3 = {{4{maskWire[59]}}, {4{maskWire[58]}}};
  wire [15:0]   maskForGroupWire_hi_hi_hi_lo_3 = {maskForGroupWire_hi_hi_hi_lo_hi_3, maskForGroupWire_hi_hi_hi_lo_lo_3};
  wire [7:0]    maskForGroupWire_hi_hi_hi_hi_lo_3 = {{4{maskWire[61]}}, {4{maskWire[60]}}};
  wire [7:0]    maskForGroupWire_hi_hi_hi_hi_hi_3 = {{4{maskWire[63]}}, {4{maskWire[62]}}};
  wire [15:0]   maskForGroupWire_hi_hi_hi_hi_3 = {maskForGroupWire_hi_hi_hi_hi_hi_3, maskForGroupWire_hi_hi_hi_hi_lo_3};
  wire [31:0]   maskForGroupWire_hi_hi_hi_3 = {maskForGroupWire_hi_hi_hi_hi_3, maskForGroupWire_hi_hi_hi_lo_3};
  wire [63:0]   maskForGroupWire_hi_hi_3 = {maskForGroupWire_hi_hi_hi_3, maskForGroupWire_hi_hi_lo_3};
  wire [127:0]  maskForGroupWire_hi_3 = {maskForGroupWire_hi_hi_3, maskForGroupWire_hi_lo_3};
  wire [7:0]    maskForGroupWire_lo_lo_lo_lo_lo_4 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]    maskForGroupWire_lo_lo_lo_lo_hi_4 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]   maskForGroupWire_lo_lo_lo_lo_4 = {maskForGroupWire_lo_lo_lo_lo_hi_4, maskForGroupWire_lo_lo_lo_lo_lo_4};
  wire [7:0]    maskForGroupWire_lo_lo_lo_hi_lo_4 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]    maskForGroupWire_lo_lo_lo_hi_hi_4 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]   maskForGroupWire_lo_lo_lo_hi_4 = {maskForGroupWire_lo_lo_lo_hi_hi_4, maskForGroupWire_lo_lo_lo_hi_lo_4};
  wire [31:0]   maskForGroupWire_lo_lo_lo_4 = {maskForGroupWire_lo_lo_lo_hi_4, maskForGroupWire_lo_lo_lo_lo_4};
  wire [7:0]    maskForGroupWire_lo_lo_hi_lo_lo_4 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]    maskForGroupWire_lo_lo_hi_lo_hi_4 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]   maskForGroupWire_lo_lo_hi_lo_4 = {maskForGroupWire_lo_lo_hi_lo_hi_4, maskForGroupWire_lo_lo_hi_lo_lo_4};
  wire [7:0]    maskForGroupWire_lo_lo_hi_hi_lo_4 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]    maskForGroupWire_lo_lo_hi_hi_hi_4 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]   maskForGroupWire_lo_lo_hi_hi_4 = {maskForGroupWire_lo_lo_hi_hi_hi_4, maskForGroupWire_lo_lo_hi_hi_lo_4};
  wire [31:0]   maskForGroupWire_lo_lo_hi_4 = {maskForGroupWire_lo_lo_hi_hi_4, maskForGroupWire_lo_lo_hi_lo_4};
  wire [63:0]   maskForGroupWire_lo_lo_4 = {maskForGroupWire_lo_lo_hi_4, maskForGroupWire_lo_lo_lo_4};
  wire [7:0]    maskForGroupWire_lo_hi_lo_lo_lo_4 = {{4{maskWire[17]}}, {4{maskWire[16]}}};
  wire [7:0]    maskForGroupWire_lo_hi_lo_lo_hi_4 = {{4{maskWire[19]}}, {4{maskWire[18]}}};
  wire [15:0]   maskForGroupWire_lo_hi_lo_lo_4 = {maskForGroupWire_lo_hi_lo_lo_hi_4, maskForGroupWire_lo_hi_lo_lo_lo_4};
  wire [7:0]    maskForGroupWire_lo_hi_lo_hi_lo_4 = {{4{maskWire[21]}}, {4{maskWire[20]}}};
  wire [7:0]    maskForGroupWire_lo_hi_lo_hi_hi_4 = {{4{maskWire[23]}}, {4{maskWire[22]}}};
  wire [15:0]   maskForGroupWire_lo_hi_lo_hi_4 = {maskForGroupWire_lo_hi_lo_hi_hi_4, maskForGroupWire_lo_hi_lo_hi_lo_4};
  wire [31:0]   maskForGroupWire_lo_hi_lo_4 = {maskForGroupWire_lo_hi_lo_hi_4, maskForGroupWire_lo_hi_lo_lo_4};
  wire [7:0]    maskForGroupWire_lo_hi_hi_lo_lo_4 = {{4{maskWire[25]}}, {4{maskWire[24]}}};
  wire [7:0]    maskForGroupWire_lo_hi_hi_lo_hi_4 = {{4{maskWire[27]}}, {4{maskWire[26]}}};
  wire [15:0]   maskForGroupWire_lo_hi_hi_lo_4 = {maskForGroupWire_lo_hi_hi_lo_hi_4, maskForGroupWire_lo_hi_hi_lo_lo_4};
  wire [7:0]    maskForGroupWire_lo_hi_hi_hi_lo_4 = {{4{maskWire[29]}}, {4{maskWire[28]}}};
  wire [7:0]    maskForGroupWire_lo_hi_hi_hi_hi_4 = {{4{maskWire[31]}}, {4{maskWire[30]}}};
  wire [15:0]   maskForGroupWire_lo_hi_hi_hi_4 = {maskForGroupWire_lo_hi_hi_hi_hi_4, maskForGroupWire_lo_hi_hi_hi_lo_4};
  wire [31:0]   maskForGroupWire_lo_hi_hi_4 = {maskForGroupWire_lo_hi_hi_hi_4, maskForGroupWire_lo_hi_hi_lo_4};
  wire [63:0]   maskForGroupWire_lo_hi_4 = {maskForGroupWire_lo_hi_hi_4, maskForGroupWire_lo_hi_lo_4};
  wire [127:0]  maskForGroupWire_lo_4 = {maskForGroupWire_lo_hi_4, maskForGroupWire_lo_lo_4};
  wire [7:0]    maskForGroupWire_hi_lo_lo_lo_lo_4 = {{4{maskWire[33]}}, {4{maskWire[32]}}};
  wire [7:0]    maskForGroupWire_hi_lo_lo_lo_hi_4 = {{4{maskWire[35]}}, {4{maskWire[34]}}};
  wire [15:0]   maskForGroupWire_hi_lo_lo_lo_4 = {maskForGroupWire_hi_lo_lo_lo_hi_4, maskForGroupWire_hi_lo_lo_lo_lo_4};
  wire [7:0]    maskForGroupWire_hi_lo_lo_hi_lo_4 = {{4{maskWire[37]}}, {4{maskWire[36]}}};
  wire [7:0]    maskForGroupWire_hi_lo_lo_hi_hi_4 = {{4{maskWire[39]}}, {4{maskWire[38]}}};
  wire [15:0]   maskForGroupWire_hi_lo_lo_hi_4 = {maskForGroupWire_hi_lo_lo_hi_hi_4, maskForGroupWire_hi_lo_lo_hi_lo_4};
  wire [31:0]   maskForGroupWire_hi_lo_lo_4 = {maskForGroupWire_hi_lo_lo_hi_4, maskForGroupWire_hi_lo_lo_lo_4};
  wire [7:0]    maskForGroupWire_hi_lo_hi_lo_lo_4 = {{4{maskWire[41]}}, {4{maskWire[40]}}};
  wire [7:0]    maskForGroupWire_hi_lo_hi_lo_hi_4 = {{4{maskWire[43]}}, {4{maskWire[42]}}};
  wire [15:0]   maskForGroupWire_hi_lo_hi_lo_4 = {maskForGroupWire_hi_lo_hi_lo_hi_4, maskForGroupWire_hi_lo_hi_lo_lo_4};
  wire [7:0]    maskForGroupWire_hi_lo_hi_hi_lo_4 = {{4{maskWire[45]}}, {4{maskWire[44]}}};
  wire [7:0]    maskForGroupWire_hi_lo_hi_hi_hi_4 = {{4{maskWire[47]}}, {4{maskWire[46]}}};
  wire [15:0]   maskForGroupWire_hi_lo_hi_hi_4 = {maskForGroupWire_hi_lo_hi_hi_hi_4, maskForGroupWire_hi_lo_hi_hi_lo_4};
  wire [31:0]   maskForGroupWire_hi_lo_hi_4 = {maskForGroupWire_hi_lo_hi_hi_4, maskForGroupWire_hi_lo_hi_lo_4};
  wire [63:0]   maskForGroupWire_hi_lo_4 = {maskForGroupWire_hi_lo_hi_4, maskForGroupWire_hi_lo_lo_4};
  wire [7:0]    maskForGroupWire_hi_hi_lo_lo_lo_4 = {{4{maskWire[49]}}, {4{maskWire[48]}}};
  wire [7:0]    maskForGroupWire_hi_hi_lo_lo_hi_4 = {{4{maskWire[51]}}, {4{maskWire[50]}}};
  wire [15:0]   maskForGroupWire_hi_hi_lo_lo_4 = {maskForGroupWire_hi_hi_lo_lo_hi_4, maskForGroupWire_hi_hi_lo_lo_lo_4};
  wire [7:0]    maskForGroupWire_hi_hi_lo_hi_lo_4 = {{4{maskWire[53]}}, {4{maskWire[52]}}};
  wire [7:0]    maskForGroupWire_hi_hi_lo_hi_hi_4 = {{4{maskWire[55]}}, {4{maskWire[54]}}};
  wire [15:0]   maskForGroupWire_hi_hi_lo_hi_4 = {maskForGroupWire_hi_hi_lo_hi_hi_4, maskForGroupWire_hi_hi_lo_hi_lo_4};
  wire [31:0]   maskForGroupWire_hi_hi_lo_4 = {maskForGroupWire_hi_hi_lo_hi_4, maskForGroupWire_hi_hi_lo_lo_4};
  wire [7:0]    maskForGroupWire_hi_hi_hi_lo_lo_4 = {{4{maskWire[57]}}, {4{maskWire[56]}}};
  wire [7:0]    maskForGroupWire_hi_hi_hi_lo_hi_4 = {{4{maskWire[59]}}, {4{maskWire[58]}}};
  wire [15:0]   maskForGroupWire_hi_hi_hi_lo_4 = {maskForGroupWire_hi_hi_hi_lo_hi_4, maskForGroupWire_hi_hi_hi_lo_lo_4};
  wire [7:0]    maskForGroupWire_hi_hi_hi_hi_lo_4 = {{4{maskWire[61]}}, {4{maskWire[60]}}};
  wire [7:0]    maskForGroupWire_hi_hi_hi_hi_hi_4 = {{4{maskWire[63]}}, {4{maskWire[62]}}};
  wire [15:0]   maskForGroupWire_hi_hi_hi_hi_4 = {maskForGroupWire_hi_hi_hi_hi_hi_4, maskForGroupWire_hi_hi_hi_hi_lo_4};
  wire [31:0]   maskForGroupWire_hi_hi_hi_4 = {maskForGroupWire_hi_hi_hi_hi_4, maskForGroupWire_hi_hi_hi_lo_4};
  wire [63:0]   maskForGroupWire_hi_hi_4 = {maskForGroupWire_hi_hi_hi_4, maskForGroupWire_hi_hi_lo_4};
  wire [127:0]  maskForGroupWire_hi_4 = {maskForGroupWire_hi_hi_4, maskForGroupWire_hi_lo_4};
  wire [7:0]    maskForGroupWire_lo_lo_lo_lo_lo_5 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]    maskForGroupWire_lo_lo_lo_lo_hi_5 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]   maskForGroupWire_lo_lo_lo_lo_5 = {maskForGroupWire_lo_lo_lo_lo_hi_5, maskForGroupWire_lo_lo_lo_lo_lo_5};
  wire [7:0]    maskForGroupWire_lo_lo_lo_hi_lo_5 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]    maskForGroupWire_lo_lo_lo_hi_hi_5 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]   maskForGroupWire_lo_lo_lo_hi_5 = {maskForGroupWire_lo_lo_lo_hi_hi_5, maskForGroupWire_lo_lo_lo_hi_lo_5};
  wire [31:0]   maskForGroupWire_lo_lo_lo_5 = {maskForGroupWire_lo_lo_lo_hi_5, maskForGroupWire_lo_lo_lo_lo_5};
  wire [7:0]    maskForGroupWire_lo_lo_hi_lo_lo_5 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]    maskForGroupWire_lo_lo_hi_lo_hi_5 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]   maskForGroupWire_lo_lo_hi_lo_5 = {maskForGroupWire_lo_lo_hi_lo_hi_5, maskForGroupWire_lo_lo_hi_lo_lo_5};
  wire [7:0]    maskForGroupWire_lo_lo_hi_hi_lo_5 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]    maskForGroupWire_lo_lo_hi_hi_hi_5 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]   maskForGroupWire_lo_lo_hi_hi_5 = {maskForGroupWire_lo_lo_hi_hi_hi_5, maskForGroupWire_lo_lo_hi_hi_lo_5};
  wire [31:0]   maskForGroupWire_lo_lo_hi_5 = {maskForGroupWire_lo_lo_hi_hi_5, maskForGroupWire_lo_lo_hi_lo_5};
  wire [63:0]   maskForGroupWire_lo_lo_5 = {maskForGroupWire_lo_lo_hi_5, maskForGroupWire_lo_lo_lo_5};
  wire [7:0]    maskForGroupWire_lo_hi_lo_lo_lo_5 = {{4{maskWire[17]}}, {4{maskWire[16]}}};
  wire [7:0]    maskForGroupWire_lo_hi_lo_lo_hi_5 = {{4{maskWire[19]}}, {4{maskWire[18]}}};
  wire [15:0]   maskForGroupWire_lo_hi_lo_lo_5 = {maskForGroupWire_lo_hi_lo_lo_hi_5, maskForGroupWire_lo_hi_lo_lo_lo_5};
  wire [7:0]    maskForGroupWire_lo_hi_lo_hi_lo_5 = {{4{maskWire[21]}}, {4{maskWire[20]}}};
  wire [7:0]    maskForGroupWire_lo_hi_lo_hi_hi_5 = {{4{maskWire[23]}}, {4{maskWire[22]}}};
  wire [15:0]   maskForGroupWire_lo_hi_lo_hi_5 = {maskForGroupWire_lo_hi_lo_hi_hi_5, maskForGroupWire_lo_hi_lo_hi_lo_5};
  wire [31:0]   maskForGroupWire_lo_hi_lo_5 = {maskForGroupWire_lo_hi_lo_hi_5, maskForGroupWire_lo_hi_lo_lo_5};
  wire [7:0]    maskForGroupWire_lo_hi_hi_lo_lo_5 = {{4{maskWire[25]}}, {4{maskWire[24]}}};
  wire [7:0]    maskForGroupWire_lo_hi_hi_lo_hi_5 = {{4{maskWire[27]}}, {4{maskWire[26]}}};
  wire [15:0]   maskForGroupWire_lo_hi_hi_lo_5 = {maskForGroupWire_lo_hi_hi_lo_hi_5, maskForGroupWire_lo_hi_hi_lo_lo_5};
  wire [7:0]    maskForGroupWire_lo_hi_hi_hi_lo_5 = {{4{maskWire[29]}}, {4{maskWire[28]}}};
  wire [7:0]    maskForGroupWire_lo_hi_hi_hi_hi_5 = {{4{maskWire[31]}}, {4{maskWire[30]}}};
  wire [15:0]   maskForGroupWire_lo_hi_hi_hi_5 = {maskForGroupWire_lo_hi_hi_hi_hi_5, maskForGroupWire_lo_hi_hi_hi_lo_5};
  wire [31:0]   maskForGroupWire_lo_hi_hi_5 = {maskForGroupWire_lo_hi_hi_hi_5, maskForGroupWire_lo_hi_hi_lo_5};
  wire [63:0]   maskForGroupWire_lo_hi_5 = {maskForGroupWire_lo_hi_hi_5, maskForGroupWire_lo_hi_lo_5};
  wire [127:0]  maskForGroupWire_lo_5 = {maskForGroupWire_lo_hi_5, maskForGroupWire_lo_lo_5};
  wire [7:0]    maskForGroupWire_hi_lo_lo_lo_lo_5 = {{4{maskWire[33]}}, {4{maskWire[32]}}};
  wire [7:0]    maskForGroupWire_hi_lo_lo_lo_hi_5 = {{4{maskWire[35]}}, {4{maskWire[34]}}};
  wire [15:0]   maskForGroupWire_hi_lo_lo_lo_5 = {maskForGroupWire_hi_lo_lo_lo_hi_5, maskForGroupWire_hi_lo_lo_lo_lo_5};
  wire [7:0]    maskForGroupWire_hi_lo_lo_hi_lo_5 = {{4{maskWire[37]}}, {4{maskWire[36]}}};
  wire [7:0]    maskForGroupWire_hi_lo_lo_hi_hi_5 = {{4{maskWire[39]}}, {4{maskWire[38]}}};
  wire [15:0]   maskForGroupWire_hi_lo_lo_hi_5 = {maskForGroupWire_hi_lo_lo_hi_hi_5, maskForGroupWire_hi_lo_lo_hi_lo_5};
  wire [31:0]   maskForGroupWire_hi_lo_lo_5 = {maskForGroupWire_hi_lo_lo_hi_5, maskForGroupWire_hi_lo_lo_lo_5};
  wire [7:0]    maskForGroupWire_hi_lo_hi_lo_lo_5 = {{4{maskWire[41]}}, {4{maskWire[40]}}};
  wire [7:0]    maskForGroupWire_hi_lo_hi_lo_hi_5 = {{4{maskWire[43]}}, {4{maskWire[42]}}};
  wire [15:0]   maskForGroupWire_hi_lo_hi_lo_5 = {maskForGroupWire_hi_lo_hi_lo_hi_5, maskForGroupWire_hi_lo_hi_lo_lo_5};
  wire [7:0]    maskForGroupWire_hi_lo_hi_hi_lo_5 = {{4{maskWire[45]}}, {4{maskWire[44]}}};
  wire [7:0]    maskForGroupWire_hi_lo_hi_hi_hi_5 = {{4{maskWire[47]}}, {4{maskWire[46]}}};
  wire [15:0]   maskForGroupWire_hi_lo_hi_hi_5 = {maskForGroupWire_hi_lo_hi_hi_hi_5, maskForGroupWire_hi_lo_hi_hi_lo_5};
  wire [31:0]   maskForGroupWire_hi_lo_hi_5 = {maskForGroupWire_hi_lo_hi_hi_5, maskForGroupWire_hi_lo_hi_lo_5};
  wire [63:0]   maskForGroupWire_hi_lo_5 = {maskForGroupWire_hi_lo_hi_5, maskForGroupWire_hi_lo_lo_5};
  wire [7:0]    maskForGroupWire_hi_hi_lo_lo_lo_5 = {{4{maskWire[49]}}, {4{maskWire[48]}}};
  wire [7:0]    maskForGroupWire_hi_hi_lo_lo_hi_5 = {{4{maskWire[51]}}, {4{maskWire[50]}}};
  wire [15:0]   maskForGroupWire_hi_hi_lo_lo_5 = {maskForGroupWire_hi_hi_lo_lo_hi_5, maskForGroupWire_hi_hi_lo_lo_lo_5};
  wire [7:0]    maskForGroupWire_hi_hi_lo_hi_lo_5 = {{4{maskWire[53]}}, {4{maskWire[52]}}};
  wire [7:0]    maskForGroupWire_hi_hi_lo_hi_hi_5 = {{4{maskWire[55]}}, {4{maskWire[54]}}};
  wire [15:0]   maskForGroupWire_hi_hi_lo_hi_5 = {maskForGroupWire_hi_hi_lo_hi_hi_5, maskForGroupWire_hi_hi_lo_hi_lo_5};
  wire [31:0]   maskForGroupWire_hi_hi_lo_5 = {maskForGroupWire_hi_hi_lo_hi_5, maskForGroupWire_hi_hi_lo_lo_5};
  wire [7:0]    maskForGroupWire_hi_hi_hi_lo_lo_5 = {{4{maskWire[57]}}, {4{maskWire[56]}}};
  wire [7:0]    maskForGroupWire_hi_hi_hi_lo_hi_5 = {{4{maskWire[59]}}, {4{maskWire[58]}}};
  wire [15:0]   maskForGroupWire_hi_hi_hi_lo_5 = {maskForGroupWire_hi_hi_hi_lo_hi_5, maskForGroupWire_hi_hi_hi_lo_lo_5};
  wire [7:0]    maskForGroupWire_hi_hi_hi_hi_lo_5 = {{4{maskWire[61]}}, {4{maskWire[60]}}};
  wire [7:0]    maskForGroupWire_hi_hi_hi_hi_hi_5 = {{4{maskWire[63]}}, {4{maskWire[62]}}};
  wire [15:0]   maskForGroupWire_hi_hi_hi_hi_5 = {maskForGroupWire_hi_hi_hi_hi_hi_5, maskForGroupWire_hi_hi_hi_hi_lo_5};
  wire [31:0]   maskForGroupWire_hi_hi_hi_5 = {maskForGroupWire_hi_hi_hi_hi_5, maskForGroupWire_hi_hi_hi_lo_5};
  wire [63:0]   maskForGroupWire_hi_hi_5 = {maskForGroupWire_hi_hi_hi_5, maskForGroupWire_hi_hi_lo_5};
  wire [127:0]  maskForGroupWire_hi_5 = {maskForGroupWire_hi_hi_5, maskForGroupWire_hi_lo_5};
  wire [63:0]   maskForGroupWire =
    (dataEEWOH[0] ? maskWire : 64'h0) | (dataEEWOH[1] ? (maskCounterInGroup[0] ? maskForGroupWire_hi : maskForGroupWire_lo_1) : 64'h0)
    | (dataEEWOH[2]
         ? (_maskForGroupWire_T_261[0] ? maskForGroupWire_lo_2[63:0] : 64'h0) | (_maskForGroupWire_T_261[1] ? maskForGroupWire_lo_3[127:64] : 64'h0) | (_maskForGroupWire_T_261[2] ? maskForGroupWire_hi_4[63:0] : 64'h0)
           | (_maskForGroupWire_T_261[3] ? maskForGroupWire_hi_5[127:64] : 64'h0)
         : 64'h0);
  wire [1:0]    initSendState_lo = maskForGroupWire[1:0];
  wire [1:0]    initSendState_hi = maskForGroupWire[3:2];
  wire          initSendState_0 = |{initSendState_hi, initSendState_lo};
  wire [1:0]    initSendState_lo_1 = maskForGroupWire[5:4];
  wire [1:0]    initSendState_hi_1 = maskForGroupWire[7:6];
  wire          initSendState_1 = |{initSendState_hi_1, initSendState_lo_1};
  wire [1:0]    initSendState_lo_2 = maskForGroupWire[9:8];
  wire [1:0]    initSendState_hi_2 = maskForGroupWire[11:10];
  wire          initSendState_2 = |{initSendState_hi_2, initSendState_lo_2};
  wire [1:0]    initSendState_lo_3 = maskForGroupWire[13:12];
  wire [1:0]    initSendState_hi_3 = maskForGroupWire[15:14];
  wire          initSendState_3 = |{initSendState_hi_3, initSendState_lo_3};
  wire [1:0]    initSendState_lo_4 = maskForGroupWire[17:16];
  wire [1:0]    initSendState_hi_4 = maskForGroupWire[19:18];
  wire          initSendState_4 = |{initSendState_hi_4, initSendState_lo_4};
  wire [1:0]    initSendState_lo_5 = maskForGroupWire[21:20];
  wire [1:0]    initSendState_hi_5 = maskForGroupWire[23:22];
  wire          initSendState_5 = |{initSendState_hi_5, initSendState_lo_5};
  wire [1:0]    initSendState_lo_6 = maskForGroupWire[25:24];
  wire [1:0]    initSendState_hi_6 = maskForGroupWire[27:26];
  wire          initSendState_6 = |{initSendState_hi_6, initSendState_lo_6};
  wire [1:0]    initSendState_lo_7 = maskForGroupWire[29:28];
  wire [1:0]    initSendState_hi_7 = maskForGroupWire[31:30];
  wire          initSendState_7 = |{initSendState_hi_7, initSendState_lo_7};
  wire [1:0]    initSendState_lo_8 = maskForGroupWire[33:32];
  wire [1:0]    initSendState_hi_8 = maskForGroupWire[35:34];
  wire          initSendState_8 = |{initSendState_hi_8, initSendState_lo_8};
  wire [1:0]    initSendState_lo_9 = maskForGroupWire[37:36];
  wire [1:0]    initSendState_hi_9 = maskForGroupWire[39:38];
  wire          initSendState_9 = |{initSendState_hi_9, initSendState_lo_9};
  wire [1:0]    initSendState_lo_10 = maskForGroupWire[41:40];
  wire [1:0]    initSendState_hi_10 = maskForGroupWire[43:42];
  wire          initSendState_10 = |{initSendState_hi_10, initSendState_lo_10};
  wire [1:0]    initSendState_lo_11 = maskForGroupWire[45:44];
  wire [1:0]    initSendState_hi_11 = maskForGroupWire[47:46];
  wire          initSendState_11 = |{initSendState_hi_11, initSendState_lo_11};
  wire [1:0]    initSendState_lo_12 = maskForGroupWire[49:48];
  wire [1:0]    initSendState_hi_12 = maskForGroupWire[51:50];
  wire          initSendState_12 = |{initSendState_hi_12, initSendState_lo_12};
  wire [1:0]    initSendState_lo_13 = maskForGroupWire[53:52];
  wire [1:0]    initSendState_hi_13 = maskForGroupWire[55:54];
  wire          initSendState_13 = |{initSendState_hi_13, initSendState_lo_13};
  wire [1:0]    initSendState_lo_14 = maskForGroupWire[57:56];
  wire [1:0]    initSendState_hi_14 = maskForGroupWire[59:58];
  wire          initSendState_14 = |{initSendState_hi_14, initSendState_lo_14};
  wire [1:0]    initSendState_lo_15 = maskForGroupWire[61:60];
  wire [1:0]    initSendState_hi_15 = maskForGroupWire[63:62];
  wire          initSendState_15 = |{initSendState_hi_15, initSendState_lo_15};
  reg  [511:0]  accessData_0;
  reg  [511:0]  accessData_1;
  reg  [511:0]  accessData_2;
  reg  [511:0]  accessData_3;
  reg  [511:0]  accessData_4;
  reg  [511:0]  accessData_5;
  reg  [511:0]  accessData_6;
  reg  [511:0]  accessData_7;
  reg  [2:0]    accessPtr;
  reg           accessState_0;
  reg           accessState_1;
  reg           accessState_2;
  reg           accessState_3;
  reg           accessState_4;
  reg           accessState_5;
  reg           accessState_6;
  reg           accessState_7;
  reg           accessState_8;
  reg           accessState_9;
  reg           accessState_10;
  reg           accessState_11;
  reg           accessState_12;
  reg           accessState_13;
  reg           accessState_14;
  reg           accessState_15;
  wire          accessStateUpdate_0;
  wire          accessStateUpdate_1;
  wire [1:0]    accessStateCheck_lo_lo_lo = {accessStateUpdate_1, accessStateUpdate_0};
  wire          accessStateUpdate_2;
  wire          accessStateUpdate_3;
  wire [1:0]    accessStateCheck_lo_lo_hi = {accessStateUpdate_3, accessStateUpdate_2};
  wire [3:0]    accessStateCheck_lo_lo = {accessStateCheck_lo_lo_hi, accessStateCheck_lo_lo_lo};
  wire          accessStateUpdate_4;
  wire          accessStateUpdate_5;
  wire [1:0]    accessStateCheck_lo_hi_lo = {accessStateUpdate_5, accessStateUpdate_4};
  wire          accessStateUpdate_6;
  wire          accessStateUpdate_7;
  wire [1:0]    accessStateCheck_lo_hi_hi = {accessStateUpdate_7, accessStateUpdate_6};
  wire [3:0]    accessStateCheck_lo_hi = {accessStateCheck_lo_hi_hi, accessStateCheck_lo_hi_lo};
  wire [7:0]    accessStateCheck_lo = {accessStateCheck_lo_hi, accessStateCheck_lo_lo};
  wire          accessStateUpdate_8;
  wire          accessStateUpdate_9;
  wire [1:0]    accessStateCheck_hi_lo_lo = {accessStateUpdate_9, accessStateUpdate_8};
  wire          accessStateUpdate_10;
  wire          accessStateUpdate_11;
  wire [1:0]    accessStateCheck_hi_lo_hi = {accessStateUpdate_11, accessStateUpdate_10};
  wire [3:0]    accessStateCheck_hi_lo = {accessStateCheck_hi_lo_hi, accessStateCheck_hi_lo_lo};
  wire          accessStateUpdate_12;
  wire          accessStateUpdate_13;
  wire [1:0]    accessStateCheck_hi_hi_lo = {accessStateUpdate_13, accessStateUpdate_12};
  wire          accessStateUpdate_14;
  wire          accessStateUpdate_15;
  wire [1:0]    accessStateCheck_hi_hi_hi = {accessStateUpdate_15, accessStateUpdate_14};
  wire [3:0]    accessStateCheck_hi_hi = {accessStateCheck_hi_hi_hi, accessStateCheck_hi_hi_lo};
  wire [7:0]    accessStateCheck_hi = {accessStateCheck_hi_hi, accessStateCheck_hi_lo};
  wire          accessStateCheck = {accessStateCheck_hi, accessStateCheck_lo} == 16'h0;
  reg  [3:0]    dataGroup;
  reg  [511:0]  dataBuffer_0;
  reg  [511:0]  dataBuffer_1;
  reg  [511:0]  dataBuffer_2;
  reg  [511:0]  dataBuffer_3;
  reg  [511:0]  dataBuffer_4;
  reg  [511:0]  dataBuffer_5;
  reg  [511:0]  dataBuffer_6;
  reg  [511:0]  dataBuffer_7;
  reg  [4:0]    bufferBaseCacheLineIndex;
  reg  [2:0]    cacheLineIndexInBuffer;
  wire [5:0]    initOffset = lsuRequestReg_rs1Data[5:0];
  wire          invalidInstruction = csrInterface_vl == 11'h0;
  reg           invalidInstructionNext;
  wire          wholeType = lsuRequest_bits_instructionInformation_lumop[3];
  wire [2:0]    nfCorrection = wholeType ? 3'h0 : lsuRequest_bits_instructionInformation_nf;
  reg  [3:0]    segmentInstructionIndexInterval;
  wire [17:0]   bytePerInstruction = {3'h0, {11'h0, {1'h0, nfCorrection} + 4'h1} * {4'h0, csrInterface_vl}} << lsuRequest_bits_instructionInformation_eew;
  wire [17:0]   accessMemSize = bytePerInstruction + {12'h0, lsuRequest_bits_rs1Data[5:0]};
  wire [11:0]   lastCacheLineIndex = accessMemSize[17:6] - {11'h0, accessMemSize[5:0] == 6'h0};
  wire [11:0]   lastWriteVrfIndex = bytePerInstruction[17:6] - {11'h0, bytePerInstruction[5:0] == 6'h0};
  reg  [11:0]   lastWriteVrfIndexReg;
  reg           lastCacheNeedPush;
  reg  [11:0]   cacheLineNumberReg;
  wire          memRequest_valid_0;
  wire          _lastCacheRequest_T = memRequest_ready_0 & memRequest_valid_0;
  reg  [4:0]    cacheLineIndex;
  wire [4:0]    memRequest_bits_src_0 = cacheLineIndex;
  wire [4:0]    nextCacheLineIndex = cacheLineIndex + 5'h1;
  wire          validInstruction = ~invalidInstruction & lsuRequest_valid;
  wire          lastRequest = cacheLineNumberReg == {7'h0, cacheLineIndex};
  reg           sendRequest;
  assign requestAddress = {lsuRequestReg_rs1Data[31:6] + {21'h0, cacheLineIndex}, 6'h0};
  wire [31:0]   memRequest_bits_address_0 = requestAddress;
  reg           writeReadyReg;
  assign memRequest_valid_0 = sendRequest & ~addressConflict;
  wire          memResponse_ready_0;
  wire          unalignedEnqueueFire = memResponse_ready_0 & memResponse_valid_0;
  wire          anyLastCacheLineAck = unalignedEnqueueFire & {7'h0, memResponse_bits_index_0} == cacheLineNumberReg;
  wire          alignedDequeueValid;
  wire [511:0]  alignedDequeue_bits_data_lo_136;
  reg           unalignedCacheLine_valid;
  reg  [511:0]  unalignedCacheLine_bits_data;
  reg  [4:0]    unalignedCacheLine_bits_index;
  wire [4:0]    alignedDequeue_bits_index = unalignedCacheLine_bits_index;
  wire          alignedDequeue_ready;
  assign unalignedEnqueueReady = alignedDequeue_ready | ~unalignedCacheLine_valid;
  assign memResponse_ready_0 = unalignedEnqueueReady;
  wire [4:0]    nextIndex = unalignedCacheLine_valid ? unalignedCacheLine_bits_index + 5'h1 : 5'h0;
  assign alignedDequeueValid = unalignedCacheLine_valid & (memResponse_valid_0 | {7'h0, unalignedCacheLine_bits_index} == cacheLineNumberReg & lastCacheNeedPush);
  wire          alignedDequeue_valid = alignedDequeueValid;
  wire          _bufferTailFire_T = alignedDequeue_ready & alignedDequeue_valid;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_lo = {unalignedCacheLine_bits_data[8], unalignedCacheLine_bits_data[0]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_hi = {unalignedCacheLine_bits_data[24], unalignedCacheLine_bits_data[16]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo = {alignedDequeue_bits_data_lo_lo_lo_lo_lo_hi, alignedDequeue_bits_data_lo_lo_lo_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_lo = {unalignedCacheLine_bits_data[40], unalignedCacheLine_bits_data[32]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_hi = {unalignedCacheLine_bits_data[56], unalignedCacheLine_bits_data[48]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_hi, alignedDequeue_bits_data_lo_lo_lo_lo_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo_lo = {alignedDequeue_bits_data_lo_lo_lo_lo_hi, alignedDequeue_bits_data_lo_lo_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_lo = {unalignedCacheLine_bits_data[72], unalignedCacheLine_bits_data[64]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_hi = {unalignedCacheLine_bits_data[88], unalignedCacheLine_bits_data[80]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo = {alignedDequeue_bits_data_lo_lo_lo_hi_lo_hi, alignedDequeue_bits_data_lo_lo_lo_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_lo = {unalignedCacheLine_bits_data[104], unalignedCacheLine_bits_data[96]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_hi = {unalignedCacheLine_bits_data[120], unalignedCacheLine_bits_data[112]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_hi, alignedDequeue_bits_data_lo_lo_lo_hi_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo_hi = {alignedDequeue_bits_data_lo_lo_lo_hi_hi, alignedDequeue_bits_data_lo_lo_lo_hi_lo};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_lo = {alignedDequeue_bits_data_lo_lo_lo_hi, alignedDequeue_bits_data_lo_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_lo = {unalignedCacheLine_bits_data[136], unalignedCacheLine_bits_data[128]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_hi = {unalignedCacheLine_bits_data[152], unalignedCacheLine_bits_data[144]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo = {alignedDequeue_bits_data_lo_lo_hi_lo_lo_hi, alignedDequeue_bits_data_lo_lo_hi_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_lo = {unalignedCacheLine_bits_data[168], unalignedCacheLine_bits_data[160]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_hi = {unalignedCacheLine_bits_data[184], unalignedCacheLine_bits_data[176]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_hi, alignedDequeue_bits_data_lo_lo_hi_lo_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi_lo = {alignedDequeue_bits_data_lo_lo_hi_lo_hi, alignedDequeue_bits_data_lo_lo_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_lo = {unalignedCacheLine_bits_data[200], unalignedCacheLine_bits_data[192]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_hi = {unalignedCacheLine_bits_data[216], unalignedCacheLine_bits_data[208]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo = {alignedDequeue_bits_data_lo_lo_hi_hi_lo_hi, alignedDequeue_bits_data_lo_lo_hi_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_lo = {unalignedCacheLine_bits_data[232], unalignedCacheLine_bits_data[224]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_hi = {unalignedCacheLine_bits_data[248], unalignedCacheLine_bits_data[240]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_hi, alignedDequeue_bits_data_lo_lo_hi_hi_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi_hi = {alignedDequeue_bits_data_lo_lo_hi_hi_hi, alignedDequeue_bits_data_lo_lo_hi_hi_lo};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_hi = {alignedDequeue_bits_data_lo_lo_hi_hi, alignedDequeue_bits_data_lo_lo_hi_lo};
  wire [31:0]   alignedDequeue_bits_data_lo_lo = {alignedDequeue_bits_data_lo_lo_hi, alignedDequeue_bits_data_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_lo = {unalignedCacheLine_bits_data[264], unalignedCacheLine_bits_data[256]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_hi = {unalignedCacheLine_bits_data[280], unalignedCacheLine_bits_data[272]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo = {alignedDequeue_bits_data_lo_hi_lo_lo_lo_hi, alignedDequeue_bits_data_lo_hi_lo_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_lo = {unalignedCacheLine_bits_data[296], unalignedCacheLine_bits_data[288]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_hi = {unalignedCacheLine_bits_data[312], unalignedCacheLine_bits_data[304]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_hi, alignedDequeue_bits_data_lo_hi_lo_lo_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo_lo = {alignedDequeue_bits_data_lo_hi_lo_lo_hi, alignedDequeue_bits_data_lo_hi_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_lo = {unalignedCacheLine_bits_data[328], unalignedCacheLine_bits_data[320]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_hi = {unalignedCacheLine_bits_data[344], unalignedCacheLine_bits_data[336]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo = {alignedDequeue_bits_data_lo_hi_lo_hi_lo_hi, alignedDequeue_bits_data_lo_hi_lo_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_lo = {unalignedCacheLine_bits_data[360], unalignedCacheLine_bits_data[352]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_hi = {unalignedCacheLine_bits_data[376], unalignedCacheLine_bits_data[368]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_hi, alignedDequeue_bits_data_lo_hi_lo_hi_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo_hi = {alignedDequeue_bits_data_lo_hi_lo_hi_hi, alignedDequeue_bits_data_lo_hi_lo_hi_lo};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_lo = {alignedDequeue_bits_data_lo_hi_lo_hi, alignedDequeue_bits_data_lo_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_lo = {unalignedCacheLine_bits_data[392], unalignedCacheLine_bits_data[384]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_hi = {unalignedCacheLine_bits_data[408], unalignedCacheLine_bits_data[400]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo = {alignedDequeue_bits_data_lo_hi_hi_lo_lo_hi, alignedDequeue_bits_data_lo_hi_hi_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_lo = {unalignedCacheLine_bits_data[424], unalignedCacheLine_bits_data[416]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_hi = {unalignedCacheLine_bits_data[440], unalignedCacheLine_bits_data[432]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_hi, alignedDequeue_bits_data_lo_hi_hi_lo_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi_lo = {alignedDequeue_bits_data_lo_hi_hi_lo_hi, alignedDequeue_bits_data_lo_hi_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_lo = {unalignedCacheLine_bits_data[456], unalignedCacheLine_bits_data[448]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_hi = {unalignedCacheLine_bits_data[472], unalignedCacheLine_bits_data[464]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo = {alignedDequeue_bits_data_lo_hi_hi_hi_lo_hi, alignedDequeue_bits_data_lo_hi_hi_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_lo = {unalignedCacheLine_bits_data[488], unalignedCacheLine_bits_data[480]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_hi = {unalignedCacheLine_bits_data[504], unalignedCacheLine_bits_data[496]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_hi, alignedDequeue_bits_data_lo_hi_hi_hi_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi_hi = {alignedDequeue_bits_data_lo_hi_hi_hi_hi, alignedDequeue_bits_data_lo_hi_hi_hi_lo};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_hi = {alignedDequeue_bits_data_lo_hi_hi_hi, alignedDequeue_bits_data_lo_hi_hi_lo};
  wire [31:0]   alignedDequeue_bits_data_lo_hi = {alignedDequeue_bits_data_lo_hi_hi, alignedDequeue_bits_data_lo_hi_lo};
  wire [63:0]   alignedDequeue_bits_data_lo = {alignedDequeue_bits_data_lo_hi, alignedDequeue_bits_data_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_lo = {memResponse_bits_data_0[8], memResponse_bits_data_0[0]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_hi = {memResponse_bits_data_0[24], memResponse_bits_data_0[16]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo = {alignedDequeue_bits_data_hi_lo_lo_lo_lo_hi, alignedDequeue_bits_data_hi_lo_lo_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_lo = {memResponse_bits_data_0[40], memResponse_bits_data_0[32]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_hi = {memResponse_bits_data_0[56], memResponse_bits_data_0[48]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_hi, alignedDequeue_bits_data_hi_lo_lo_lo_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo_lo = {alignedDequeue_bits_data_hi_lo_lo_lo_hi, alignedDequeue_bits_data_hi_lo_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_lo = {memResponse_bits_data_0[72], memResponse_bits_data_0[64]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_hi = {memResponse_bits_data_0[88], memResponse_bits_data_0[80]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo = {alignedDequeue_bits_data_hi_lo_lo_hi_lo_hi, alignedDequeue_bits_data_hi_lo_lo_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_lo = {memResponse_bits_data_0[104], memResponse_bits_data_0[96]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_hi = {memResponse_bits_data_0[120], memResponse_bits_data_0[112]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_hi, alignedDequeue_bits_data_hi_lo_lo_hi_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo_hi = {alignedDequeue_bits_data_hi_lo_lo_hi_hi, alignedDequeue_bits_data_hi_lo_lo_hi_lo};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_lo = {alignedDequeue_bits_data_hi_lo_lo_hi, alignedDequeue_bits_data_hi_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_lo = {memResponse_bits_data_0[136], memResponse_bits_data_0[128]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_hi = {memResponse_bits_data_0[152], memResponse_bits_data_0[144]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo = {alignedDequeue_bits_data_hi_lo_hi_lo_lo_hi, alignedDequeue_bits_data_hi_lo_hi_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_lo = {memResponse_bits_data_0[168], memResponse_bits_data_0[160]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_hi = {memResponse_bits_data_0[184], memResponse_bits_data_0[176]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_hi, alignedDequeue_bits_data_hi_lo_hi_lo_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi_lo = {alignedDequeue_bits_data_hi_lo_hi_lo_hi, alignedDequeue_bits_data_hi_lo_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_lo = {memResponse_bits_data_0[200], memResponse_bits_data_0[192]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_hi = {memResponse_bits_data_0[216], memResponse_bits_data_0[208]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo = {alignedDequeue_bits_data_hi_lo_hi_hi_lo_hi, alignedDequeue_bits_data_hi_lo_hi_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_lo = {memResponse_bits_data_0[232], memResponse_bits_data_0[224]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_hi = {memResponse_bits_data_0[248], memResponse_bits_data_0[240]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_hi, alignedDequeue_bits_data_hi_lo_hi_hi_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi_hi = {alignedDequeue_bits_data_hi_lo_hi_hi_hi, alignedDequeue_bits_data_hi_lo_hi_hi_lo};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_hi = {alignedDequeue_bits_data_hi_lo_hi_hi, alignedDequeue_bits_data_hi_lo_hi_lo};
  wire [31:0]   alignedDequeue_bits_data_hi_lo = {alignedDequeue_bits_data_hi_lo_hi, alignedDequeue_bits_data_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_lo = {memResponse_bits_data_0[264], memResponse_bits_data_0[256]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_hi = {memResponse_bits_data_0[280], memResponse_bits_data_0[272]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo = {alignedDequeue_bits_data_hi_hi_lo_lo_lo_hi, alignedDequeue_bits_data_hi_hi_lo_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_lo = {memResponse_bits_data_0[296], memResponse_bits_data_0[288]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_hi = {memResponse_bits_data_0[312], memResponse_bits_data_0[304]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_hi, alignedDequeue_bits_data_hi_hi_lo_lo_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo_lo = {alignedDequeue_bits_data_hi_hi_lo_lo_hi, alignedDequeue_bits_data_hi_hi_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_lo = {memResponse_bits_data_0[328], memResponse_bits_data_0[320]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_hi = {memResponse_bits_data_0[344], memResponse_bits_data_0[336]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo = {alignedDequeue_bits_data_hi_hi_lo_hi_lo_hi, alignedDequeue_bits_data_hi_hi_lo_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_lo = {memResponse_bits_data_0[360], memResponse_bits_data_0[352]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_hi = {memResponse_bits_data_0[376], memResponse_bits_data_0[368]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_hi, alignedDequeue_bits_data_hi_hi_lo_hi_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo_hi = {alignedDequeue_bits_data_hi_hi_lo_hi_hi, alignedDequeue_bits_data_hi_hi_lo_hi_lo};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_lo = {alignedDequeue_bits_data_hi_hi_lo_hi, alignedDequeue_bits_data_hi_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_lo = {memResponse_bits_data_0[392], memResponse_bits_data_0[384]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_hi = {memResponse_bits_data_0[408], memResponse_bits_data_0[400]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo = {alignedDequeue_bits_data_hi_hi_hi_lo_lo_hi, alignedDequeue_bits_data_hi_hi_hi_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_lo = {memResponse_bits_data_0[424], memResponse_bits_data_0[416]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_hi = {memResponse_bits_data_0[440], memResponse_bits_data_0[432]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_hi, alignedDequeue_bits_data_hi_hi_hi_lo_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi_lo = {alignedDequeue_bits_data_hi_hi_hi_lo_hi, alignedDequeue_bits_data_hi_hi_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_lo = {memResponse_bits_data_0[456], memResponse_bits_data_0[448]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_hi = {memResponse_bits_data_0[472], memResponse_bits_data_0[464]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo = {alignedDequeue_bits_data_hi_hi_hi_hi_lo_hi, alignedDequeue_bits_data_hi_hi_hi_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_lo = {memResponse_bits_data_0[488], memResponse_bits_data_0[480]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_hi = {memResponse_bits_data_0[504], memResponse_bits_data_0[496]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_hi, alignedDequeue_bits_data_hi_hi_hi_hi_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi_hi = {alignedDequeue_bits_data_hi_hi_hi_hi_hi, alignedDequeue_bits_data_hi_hi_hi_hi_lo};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_hi = {alignedDequeue_bits_data_hi_hi_hi_hi, alignedDequeue_bits_data_hi_hi_hi_lo};
  wire [31:0]   alignedDequeue_bits_data_hi_hi = {alignedDequeue_bits_data_hi_hi_hi, alignedDequeue_bits_data_hi_hi_lo};
  wire [63:0]   alignedDequeue_bits_data_hi = {alignedDequeue_bits_data_hi_hi, alignedDequeue_bits_data_hi_lo};
  wire [127:0]  _GEN_4 = {122'h0, initOffset};
  wire [127:0]  _alignedDequeue_bits_data_T_1026 = {alignedDequeue_bits_data_hi, alignedDequeue_bits_data_lo} >> _GEN_4;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_lo_1 = {unalignedCacheLine_bits_data[9], unalignedCacheLine_bits_data[1]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_hi_1 = {unalignedCacheLine_bits_data[25], unalignedCacheLine_bits_data[17]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_1 = {alignedDequeue_bits_data_lo_lo_lo_lo_lo_hi_1, alignedDequeue_bits_data_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_lo_1 = {unalignedCacheLine_bits_data[41], unalignedCacheLine_bits_data[33]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_hi_1 = {unalignedCacheLine_bits_data[57], unalignedCacheLine_bits_data[49]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_1 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_hi_1, alignedDequeue_bits_data_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo_lo_1 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_1, alignedDequeue_bits_data_lo_lo_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_lo_1 = {unalignedCacheLine_bits_data[73], unalignedCacheLine_bits_data[65]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_hi_1 = {unalignedCacheLine_bits_data[89], unalignedCacheLine_bits_data[81]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_1 = {alignedDequeue_bits_data_lo_lo_lo_hi_lo_hi_1, alignedDequeue_bits_data_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_lo_1 = {unalignedCacheLine_bits_data[105], unalignedCacheLine_bits_data[97]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_hi_1 = {unalignedCacheLine_bits_data[121], unalignedCacheLine_bits_data[113]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_1 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_hi_1, alignedDequeue_bits_data_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo_hi_1 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_1, alignedDequeue_bits_data_lo_lo_lo_hi_lo_1};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_lo_1 = {alignedDequeue_bits_data_lo_lo_lo_hi_1, alignedDequeue_bits_data_lo_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_lo_1 = {unalignedCacheLine_bits_data[137], unalignedCacheLine_bits_data[129]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_hi_1 = {unalignedCacheLine_bits_data[153], unalignedCacheLine_bits_data[145]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_1 = {alignedDequeue_bits_data_lo_lo_hi_lo_lo_hi_1, alignedDequeue_bits_data_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_lo_1 = {unalignedCacheLine_bits_data[169], unalignedCacheLine_bits_data[161]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_hi_1 = {unalignedCacheLine_bits_data[185], unalignedCacheLine_bits_data[177]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_1 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_hi_1, alignedDequeue_bits_data_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi_lo_1 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_1, alignedDequeue_bits_data_lo_lo_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_lo_1 = {unalignedCacheLine_bits_data[201], unalignedCacheLine_bits_data[193]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_hi_1 = {unalignedCacheLine_bits_data[217], unalignedCacheLine_bits_data[209]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_1 = {alignedDequeue_bits_data_lo_lo_hi_hi_lo_hi_1, alignedDequeue_bits_data_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_lo_1 = {unalignedCacheLine_bits_data[233], unalignedCacheLine_bits_data[225]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_hi_1 = {unalignedCacheLine_bits_data[249], unalignedCacheLine_bits_data[241]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_1 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_hi_1, alignedDequeue_bits_data_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi_hi_1 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_1, alignedDequeue_bits_data_lo_lo_hi_hi_lo_1};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_hi_1 = {alignedDequeue_bits_data_lo_lo_hi_hi_1, alignedDequeue_bits_data_lo_lo_hi_lo_1};
  wire [31:0]   alignedDequeue_bits_data_lo_lo_1 = {alignedDequeue_bits_data_lo_lo_hi_1, alignedDequeue_bits_data_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_lo_1 = {unalignedCacheLine_bits_data[265], unalignedCacheLine_bits_data[257]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_hi_1 = {unalignedCacheLine_bits_data[281], unalignedCacheLine_bits_data[273]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_1 = {alignedDequeue_bits_data_lo_hi_lo_lo_lo_hi_1, alignedDequeue_bits_data_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_lo_1 = {unalignedCacheLine_bits_data[297], unalignedCacheLine_bits_data[289]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_hi_1 = {unalignedCacheLine_bits_data[313], unalignedCacheLine_bits_data[305]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_1 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_hi_1, alignedDequeue_bits_data_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo_lo_1 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_1, alignedDequeue_bits_data_lo_hi_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_lo_1 = {unalignedCacheLine_bits_data[329], unalignedCacheLine_bits_data[321]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_hi_1 = {unalignedCacheLine_bits_data[345], unalignedCacheLine_bits_data[337]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_1 = {alignedDequeue_bits_data_lo_hi_lo_hi_lo_hi_1, alignedDequeue_bits_data_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_lo_1 = {unalignedCacheLine_bits_data[361], unalignedCacheLine_bits_data[353]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_hi_1 = {unalignedCacheLine_bits_data[377], unalignedCacheLine_bits_data[369]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_1 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_hi_1, alignedDequeue_bits_data_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo_hi_1 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_1, alignedDequeue_bits_data_lo_hi_lo_hi_lo_1};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_lo_1 = {alignedDequeue_bits_data_lo_hi_lo_hi_1, alignedDequeue_bits_data_lo_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_lo_1 = {unalignedCacheLine_bits_data[393], unalignedCacheLine_bits_data[385]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_hi_1 = {unalignedCacheLine_bits_data[409], unalignedCacheLine_bits_data[401]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_1 = {alignedDequeue_bits_data_lo_hi_hi_lo_lo_hi_1, alignedDequeue_bits_data_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_lo_1 = {unalignedCacheLine_bits_data[425], unalignedCacheLine_bits_data[417]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_hi_1 = {unalignedCacheLine_bits_data[441], unalignedCacheLine_bits_data[433]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_1 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_hi_1, alignedDequeue_bits_data_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi_lo_1 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_1, alignedDequeue_bits_data_lo_hi_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_lo_1 = {unalignedCacheLine_bits_data[457], unalignedCacheLine_bits_data[449]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_hi_1 = {unalignedCacheLine_bits_data[473], unalignedCacheLine_bits_data[465]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_1 = {alignedDequeue_bits_data_lo_hi_hi_hi_lo_hi_1, alignedDequeue_bits_data_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_lo_1 = {unalignedCacheLine_bits_data[489], unalignedCacheLine_bits_data[481]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_hi_1 = {unalignedCacheLine_bits_data[505], unalignedCacheLine_bits_data[497]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_1 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_hi_1, alignedDequeue_bits_data_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi_hi_1 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_1, alignedDequeue_bits_data_lo_hi_hi_hi_lo_1};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_hi_1 = {alignedDequeue_bits_data_lo_hi_hi_hi_1, alignedDequeue_bits_data_lo_hi_hi_lo_1};
  wire [31:0]   alignedDequeue_bits_data_lo_hi_1 = {alignedDequeue_bits_data_lo_hi_hi_1, alignedDequeue_bits_data_lo_hi_lo_1};
  wire [63:0]   alignedDequeue_bits_data_lo_1 = {alignedDequeue_bits_data_lo_hi_1, alignedDequeue_bits_data_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_lo_1 = {memResponse_bits_data_0[9], memResponse_bits_data_0[1]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_hi_1 = {memResponse_bits_data_0[25], memResponse_bits_data_0[17]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_1 = {alignedDequeue_bits_data_hi_lo_lo_lo_lo_hi_1, alignedDequeue_bits_data_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_lo_1 = {memResponse_bits_data_0[41], memResponse_bits_data_0[33]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_hi_1 = {memResponse_bits_data_0[57], memResponse_bits_data_0[49]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_1 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_hi_1, alignedDequeue_bits_data_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo_lo_1 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_1, alignedDequeue_bits_data_hi_lo_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_lo_1 = {memResponse_bits_data_0[73], memResponse_bits_data_0[65]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_hi_1 = {memResponse_bits_data_0[89], memResponse_bits_data_0[81]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_1 = {alignedDequeue_bits_data_hi_lo_lo_hi_lo_hi_1, alignedDequeue_bits_data_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_lo_1 = {memResponse_bits_data_0[105], memResponse_bits_data_0[97]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_hi_1 = {memResponse_bits_data_0[121], memResponse_bits_data_0[113]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_1 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_hi_1, alignedDequeue_bits_data_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo_hi_1 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_1, alignedDequeue_bits_data_hi_lo_lo_hi_lo_1};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_lo_1 = {alignedDequeue_bits_data_hi_lo_lo_hi_1, alignedDequeue_bits_data_hi_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_lo_1 = {memResponse_bits_data_0[137], memResponse_bits_data_0[129]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_hi_1 = {memResponse_bits_data_0[153], memResponse_bits_data_0[145]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_1 = {alignedDequeue_bits_data_hi_lo_hi_lo_lo_hi_1, alignedDequeue_bits_data_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_lo_1 = {memResponse_bits_data_0[169], memResponse_bits_data_0[161]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_hi_1 = {memResponse_bits_data_0[185], memResponse_bits_data_0[177]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_1 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_hi_1, alignedDequeue_bits_data_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi_lo_1 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_1, alignedDequeue_bits_data_hi_lo_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_lo_1 = {memResponse_bits_data_0[201], memResponse_bits_data_0[193]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_hi_1 = {memResponse_bits_data_0[217], memResponse_bits_data_0[209]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_1 = {alignedDequeue_bits_data_hi_lo_hi_hi_lo_hi_1, alignedDequeue_bits_data_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_lo_1 = {memResponse_bits_data_0[233], memResponse_bits_data_0[225]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_hi_1 = {memResponse_bits_data_0[249], memResponse_bits_data_0[241]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_1 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_hi_1, alignedDequeue_bits_data_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi_hi_1 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_1, alignedDequeue_bits_data_hi_lo_hi_hi_lo_1};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_hi_1 = {alignedDequeue_bits_data_hi_lo_hi_hi_1, alignedDequeue_bits_data_hi_lo_hi_lo_1};
  wire [31:0]   alignedDequeue_bits_data_hi_lo_1 = {alignedDequeue_bits_data_hi_lo_hi_1, alignedDequeue_bits_data_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_lo_1 = {memResponse_bits_data_0[265], memResponse_bits_data_0[257]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_hi_1 = {memResponse_bits_data_0[281], memResponse_bits_data_0[273]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_1 = {alignedDequeue_bits_data_hi_hi_lo_lo_lo_hi_1, alignedDequeue_bits_data_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_lo_1 = {memResponse_bits_data_0[297], memResponse_bits_data_0[289]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_hi_1 = {memResponse_bits_data_0[313], memResponse_bits_data_0[305]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_1 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_hi_1, alignedDequeue_bits_data_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo_lo_1 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_1, alignedDequeue_bits_data_hi_hi_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_lo_1 = {memResponse_bits_data_0[329], memResponse_bits_data_0[321]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_hi_1 = {memResponse_bits_data_0[345], memResponse_bits_data_0[337]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_1 = {alignedDequeue_bits_data_hi_hi_lo_hi_lo_hi_1, alignedDequeue_bits_data_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_lo_1 = {memResponse_bits_data_0[361], memResponse_bits_data_0[353]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_hi_1 = {memResponse_bits_data_0[377], memResponse_bits_data_0[369]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_1 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_hi_1, alignedDequeue_bits_data_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo_hi_1 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_1, alignedDequeue_bits_data_hi_hi_lo_hi_lo_1};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_lo_1 = {alignedDequeue_bits_data_hi_hi_lo_hi_1, alignedDequeue_bits_data_hi_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_lo_1 = {memResponse_bits_data_0[393], memResponse_bits_data_0[385]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_hi_1 = {memResponse_bits_data_0[409], memResponse_bits_data_0[401]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_1 = {alignedDequeue_bits_data_hi_hi_hi_lo_lo_hi_1, alignedDequeue_bits_data_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_lo_1 = {memResponse_bits_data_0[425], memResponse_bits_data_0[417]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_hi_1 = {memResponse_bits_data_0[441], memResponse_bits_data_0[433]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_1 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_hi_1, alignedDequeue_bits_data_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi_lo_1 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_1, alignedDequeue_bits_data_hi_hi_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_lo_1 = {memResponse_bits_data_0[457], memResponse_bits_data_0[449]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_hi_1 = {memResponse_bits_data_0[473], memResponse_bits_data_0[465]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_1 = {alignedDequeue_bits_data_hi_hi_hi_hi_lo_hi_1, alignedDequeue_bits_data_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_lo_1 = {memResponse_bits_data_0[489], memResponse_bits_data_0[481]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_hi_1 = {memResponse_bits_data_0[505], memResponse_bits_data_0[497]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_1 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_hi_1, alignedDequeue_bits_data_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi_hi_1 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_1, alignedDequeue_bits_data_hi_hi_hi_hi_lo_1};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_hi_1 = {alignedDequeue_bits_data_hi_hi_hi_hi_1, alignedDequeue_bits_data_hi_hi_hi_lo_1};
  wire [31:0]   alignedDequeue_bits_data_hi_hi_1 = {alignedDequeue_bits_data_hi_hi_hi_1, alignedDequeue_bits_data_hi_hi_lo_1};
  wire [63:0]   alignedDequeue_bits_data_hi_1 = {alignedDequeue_bits_data_hi_hi_1, alignedDequeue_bits_data_hi_lo_1};
  wire [127:0]  _alignedDequeue_bits_data_T_1156 = {alignedDequeue_bits_data_hi_1, alignedDequeue_bits_data_lo_1} >> _GEN_4;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_lo_2 = {unalignedCacheLine_bits_data[10], unalignedCacheLine_bits_data[2]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_hi_2 = {unalignedCacheLine_bits_data[26], unalignedCacheLine_bits_data[18]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_2 = {alignedDequeue_bits_data_lo_lo_lo_lo_lo_hi_2, alignedDequeue_bits_data_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_lo_2 = {unalignedCacheLine_bits_data[42], unalignedCacheLine_bits_data[34]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_hi_2 = {unalignedCacheLine_bits_data[58], unalignedCacheLine_bits_data[50]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_2 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_hi_2, alignedDequeue_bits_data_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo_lo_2 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_2, alignedDequeue_bits_data_lo_lo_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_lo_2 = {unalignedCacheLine_bits_data[74], unalignedCacheLine_bits_data[66]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_hi_2 = {unalignedCacheLine_bits_data[90], unalignedCacheLine_bits_data[82]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_2 = {alignedDequeue_bits_data_lo_lo_lo_hi_lo_hi_2, alignedDequeue_bits_data_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_lo_2 = {unalignedCacheLine_bits_data[106], unalignedCacheLine_bits_data[98]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_hi_2 = {unalignedCacheLine_bits_data[122], unalignedCacheLine_bits_data[114]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_2 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_hi_2, alignedDequeue_bits_data_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo_hi_2 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_2, alignedDequeue_bits_data_lo_lo_lo_hi_lo_2};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_lo_2 = {alignedDequeue_bits_data_lo_lo_lo_hi_2, alignedDequeue_bits_data_lo_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_lo_2 = {unalignedCacheLine_bits_data[138], unalignedCacheLine_bits_data[130]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_hi_2 = {unalignedCacheLine_bits_data[154], unalignedCacheLine_bits_data[146]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_2 = {alignedDequeue_bits_data_lo_lo_hi_lo_lo_hi_2, alignedDequeue_bits_data_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_lo_2 = {unalignedCacheLine_bits_data[170], unalignedCacheLine_bits_data[162]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_hi_2 = {unalignedCacheLine_bits_data[186], unalignedCacheLine_bits_data[178]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_2 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_hi_2, alignedDequeue_bits_data_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi_lo_2 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_2, alignedDequeue_bits_data_lo_lo_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_lo_2 = {unalignedCacheLine_bits_data[202], unalignedCacheLine_bits_data[194]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_hi_2 = {unalignedCacheLine_bits_data[218], unalignedCacheLine_bits_data[210]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_2 = {alignedDequeue_bits_data_lo_lo_hi_hi_lo_hi_2, alignedDequeue_bits_data_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_lo_2 = {unalignedCacheLine_bits_data[234], unalignedCacheLine_bits_data[226]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_hi_2 = {unalignedCacheLine_bits_data[250], unalignedCacheLine_bits_data[242]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_2 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_hi_2, alignedDequeue_bits_data_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi_hi_2 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_2, alignedDequeue_bits_data_lo_lo_hi_hi_lo_2};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_hi_2 = {alignedDequeue_bits_data_lo_lo_hi_hi_2, alignedDequeue_bits_data_lo_lo_hi_lo_2};
  wire [31:0]   alignedDequeue_bits_data_lo_lo_2 = {alignedDequeue_bits_data_lo_lo_hi_2, alignedDequeue_bits_data_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_lo_2 = {unalignedCacheLine_bits_data[266], unalignedCacheLine_bits_data[258]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_hi_2 = {unalignedCacheLine_bits_data[282], unalignedCacheLine_bits_data[274]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_2 = {alignedDequeue_bits_data_lo_hi_lo_lo_lo_hi_2, alignedDequeue_bits_data_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_lo_2 = {unalignedCacheLine_bits_data[298], unalignedCacheLine_bits_data[290]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_hi_2 = {unalignedCacheLine_bits_data[314], unalignedCacheLine_bits_data[306]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_2 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_hi_2, alignedDequeue_bits_data_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo_lo_2 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_2, alignedDequeue_bits_data_lo_hi_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_lo_2 = {unalignedCacheLine_bits_data[330], unalignedCacheLine_bits_data[322]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_hi_2 = {unalignedCacheLine_bits_data[346], unalignedCacheLine_bits_data[338]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_2 = {alignedDequeue_bits_data_lo_hi_lo_hi_lo_hi_2, alignedDequeue_bits_data_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_lo_2 = {unalignedCacheLine_bits_data[362], unalignedCacheLine_bits_data[354]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_hi_2 = {unalignedCacheLine_bits_data[378], unalignedCacheLine_bits_data[370]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_2 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_hi_2, alignedDequeue_bits_data_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo_hi_2 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_2, alignedDequeue_bits_data_lo_hi_lo_hi_lo_2};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_lo_2 = {alignedDequeue_bits_data_lo_hi_lo_hi_2, alignedDequeue_bits_data_lo_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_lo_2 = {unalignedCacheLine_bits_data[394], unalignedCacheLine_bits_data[386]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_hi_2 = {unalignedCacheLine_bits_data[410], unalignedCacheLine_bits_data[402]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_2 = {alignedDequeue_bits_data_lo_hi_hi_lo_lo_hi_2, alignedDequeue_bits_data_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_lo_2 = {unalignedCacheLine_bits_data[426], unalignedCacheLine_bits_data[418]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_hi_2 = {unalignedCacheLine_bits_data[442], unalignedCacheLine_bits_data[434]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_2 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_hi_2, alignedDequeue_bits_data_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi_lo_2 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_2, alignedDequeue_bits_data_lo_hi_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_lo_2 = {unalignedCacheLine_bits_data[458], unalignedCacheLine_bits_data[450]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_hi_2 = {unalignedCacheLine_bits_data[474], unalignedCacheLine_bits_data[466]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_2 = {alignedDequeue_bits_data_lo_hi_hi_hi_lo_hi_2, alignedDequeue_bits_data_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_lo_2 = {unalignedCacheLine_bits_data[490], unalignedCacheLine_bits_data[482]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_hi_2 = {unalignedCacheLine_bits_data[506], unalignedCacheLine_bits_data[498]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_2 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_hi_2, alignedDequeue_bits_data_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi_hi_2 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_2, alignedDequeue_bits_data_lo_hi_hi_hi_lo_2};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_hi_2 = {alignedDequeue_bits_data_lo_hi_hi_hi_2, alignedDequeue_bits_data_lo_hi_hi_lo_2};
  wire [31:0]   alignedDequeue_bits_data_lo_hi_2 = {alignedDequeue_bits_data_lo_hi_hi_2, alignedDequeue_bits_data_lo_hi_lo_2};
  wire [63:0]   alignedDequeue_bits_data_lo_2 = {alignedDequeue_bits_data_lo_hi_2, alignedDequeue_bits_data_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_lo_2 = {memResponse_bits_data_0[10], memResponse_bits_data_0[2]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_hi_2 = {memResponse_bits_data_0[26], memResponse_bits_data_0[18]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_2 = {alignedDequeue_bits_data_hi_lo_lo_lo_lo_hi_2, alignedDequeue_bits_data_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_lo_2 = {memResponse_bits_data_0[42], memResponse_bits_data_0[34]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_hi_2 = {memResponse_bits_data_0[58], memResponse_bits_data_0[50]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_2 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_hi_2, alignedDequeue_bits_data_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo_lo_2 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_2, alignedDequeue_bits_data_hi_lo_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_lo_2 = {memResponse_bits_data_0[74], memResponse_bits_data_0[66]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_hi_2 = {memResponse_bits_data_0[90], memResponse_bits_data_0[82]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_2 = {alignedDequeue_bits_data_hi_lo_lo_hi_lo_hi_2, alignedDequeue_bits_data_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_lo_2 = {memResponse_bits_data_0[106], memResponse_bits_data_0[98]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_hi_2 = {memResponse_bits_data_0[122], memResponse_bits_data_0[114]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_2 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_hi_2, alignedDequeue_bits_data_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo_hi_2 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_2, alignedDequeue_bits_data_hi_lo_lo_hi_lo_2};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_lo_2 = {alignedDequeue_bits_data_hi_lo_lo_hi_2, alignedDequeue_bits_data_hi_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_lo_2 = {memResponse_bits_data_0[138], memResponse_bits_data_0[130]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_hi_2 = {memResponse_bits_data_0[154], memResponse_bits_data_0[146]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_2 = {alignedDequeue_bits_data_hi_lo_hi_lo_lo_hi_2, alignedDequeue_bits_data_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_lo_2 = {memResponse_bits_data_0[170], memResponse_bits_data_0[162]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_hi_2 = {memResponse_bits_data_0[186], memResponse_bits_data_0[178]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_2 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_hi_2, alignedDequeue_bits_data_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi_lo_2 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_2, alignedDequeue_bits_data_hi_lo_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_lo_2 = {memResponse_bits_data_0[202], memResponse_bits_data_0[194]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_hi_2 = {memResponse_bits_data_0[218], memResponse_bits_data_0[210]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_2 = {alignedDequeue_bits_data_hi_lo_hi_hi_lo_hi_2, alignedDequeue_bits_data_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_lo_2 = {memResponse_bits_data_0[234], memResponse_bits_data_0[226]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_hi_2 = {memResponse_bits_data_0[250], memResponse_bits_data_0[242]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_2 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_hi_2, alignedDequeue_bits_data_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi_hi_2 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_2, alignedDequeue_bits_data_hi_lo_hi_hi_lo_2};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_hi_2 = {alignedDequeue_bits_data_hi_lo_hi_hi_2, alignedDequeue_bits_data_hi_lo_hi_lo_2};
  wire [31:0]   alignedDequeue_bits_data_hi_lo_2 = {alignedDequeue_bits_data_hi_lo_hi_2, alignedDequeue_bits_data_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_lo_2 = {memResponse_bits_data_0[266], memResponse_bits_data_0[258]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_hi_2 = {memResponse_bits_data_0[282], memResponse_bits_data_0[274]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_2 = {alignedDequeue_bits_data_hi_hi_lo_lo_lo_hi_2, alignedDequeue_bits_data_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_lo_2 = {memResponse_bits_data_0[298], memResponse_bits_data_0[290]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_hi_2 = {memResponse_bits_data_0[314], memResponse_bits_data_0[306]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_2 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_hi_2, alignedDequeue_bits_data_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo_lo_2 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_2, alignedDequeue_bits_data_hi_hi_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_lo_2 = {memResponse_bits_data_0[330], memResponse_bits_data_0[322]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_hi_2 = {memResponse_bits_data_0[346], memResponse_bits_data_0[338]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_2 = {alignedDequeue_bits_data_hi_hi_lo_hi_lo_hi_2, alignedDequeue_bits_data_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_lo_2 = {memResponse_bits_data_0[362], memResponse_bits_data_0[354]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_hi_2 = {memResponse_bits_data_0[378], memResponse_bits_data_0[370]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_2 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_hi_2, alignedDequeue_bits_data_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo_hi_2 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_2, alignedDequeue_bits_data_hi_hi_lo_hi_lo_2};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_lo_2 = {alignedDequeue_bits_data_hi_hi_lo_hi_2, alignedDequeue_bits_data_hi_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_lo_2 = {memResponse_bits_data_0[394], memResponse_bits_data_0[386]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_hi_2 = {memResponse_bits_data_0[410], memResponse_bits_data_0[402]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_2 = {alignedDequeue_bits_data_hi_hi_hi_lo_lo_hi_2, alignedDequeue_bits_data_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_lo_2 = {memResponse_bits_data_0[426], memResponse_bits_data_0[418]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_hi_2 = {memResponse_bits_data_0[442], memResponse_bits_data_0[434]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_2 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_hi_2, alignedDequeue_bits_data_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi_lo_2 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_2, alignedDequeue_bits_data_hi_hi_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_lo_2 = {memResponse_bits_data_0[458], memResponse_bits_data_0[450]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_hi_2 = {memResponse_bits_data_0[474], memResponse_bits_data_0[466]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_2 = {alignedDequeue_bits_data_hi_hi_hi_hi_lo_hi_2, alignedDequeue_bits_data_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_lo_2 = {memResponse_bits_data_0[490], memResponse_bits_data_0[482]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_hi_2 = {memResponse_bits_data_0[506], memResponse_bits_data_0[498]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_2 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_hi_2, alignedDequeue_bits_data_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi_hi_2 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_2, alignedDequeue_bits_data_hi_hi_hi_hi_lo_2};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_hi_2 = {alignedDequeue_bits_data_hi_hi_hi_hi_2, alignedDequeue_bits_data_hi_hi_hi_lo_2};
  wire [31:0]   alignedDequeue_bits_data_hi_hi_2 = {alignedDequeue_bits_data_hi_hi_hi_2, alignedDequeue_bits_data_hi_hi_lo_2};
  wire [63:0]   alignedDequeue_bits_data_hi_2 = {alignedDequeue_bits_data_hi_hi_2, alignedDequeue_bits_data_hi_lo_2};
  wire [127:0]  _alignedDequeue_bits_data_T_1286 = {alignedDequeue_bits_data_hi_2, alignedDequeue_bits_data_lo_2} >> _GEN_4;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_lo_3 = {unalignedCacheLine_bits_data[11], unalignedCacheLine_bits_data[3]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_hi_3 = {unalignedCacheLine_bits_data[27], unalignedCacheLine_bits_data[19]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_3 = {alignedDequeue_bits_data_lo_lo_lo_lo_lo_hi_3, alignedDequeue_bits_data_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_lo_3 = {unalignedCacheLine_bits_data[43], unalignedCacheLine_bits_data[35]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_hi_3 = {unalignedCacheLine_bits_data[59], unalignedCacheLine_bits_data[51]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_3 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_hi_3, alignedDequeue_bits_data_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo_lo_3 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_3, alignedDequeue_bits_data_lo_lo_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_lo_3 = {unalignedCacheLine_bits_data[75], unalignedCacheLine_bits_data[67]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_hi_3 = {unalignedCacheLine_bits_data[91], unalignedCacheLine_bits_data[83]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_3 = {alignedDequeue_bits_data_lo_lo_lo_hi_lo_hi_3, alignedDequeue_bits_data_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_lo_3 = {unalignedCacheLine_bits_data[107], unalignedCacheLine_bits_data[99]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_hi_3 = {unalignedCacheLine_bits_data[123], unalignedCacheLine_bits_data[115]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_3 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_hi_3, alignedDequeue_bits_data_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo_hi_3 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_3, alignedDequeue_bits_data_lo_lo_lo_hi_lo_3};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_lo_3 = {alignedDequeue_bits_data_lo_lo_lo_hi_3, alignedDequeue_bits_data_lo_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_lo_3 = {unalignedCacheLine_bits_data[139], unalignedCacheLine_bits_data[131]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_hi_3 = {unalignedCacheLine_bits_data[155], unalignedCacheLine_bits_data[147]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_3 = {alignedDequeue_bits_data_lo_lo_hi_lo_lo_hi_3, alignedDequeue_bits_data_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_lo_3 = {unalignedCacheLine_bits_data[171], unalignedCacheLine_bits_data[163]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_hi_3 = {unalignedCacheLine_bits_data[187], unalignedCacheLine_bits_data[179]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_3 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_hi_3, alignedDequeue_bits_data_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi_lo_3 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_3, alignedDequeue_bits_data_lo_lo_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_lo_3 = {unalignedCacheLine_bits_data[203], unalignedCacheLine_bits_data[195]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_hi_3 = {unalignedCacheLine_bits_data[219], unalignedCacheLine_bits_data[211]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_3 = {alignedDequeue_bits_data_lo_lo_hi_hi_lo_hi_3, alignedDequeue_bits_data_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_lo_3 = {unalignedCacheLine_bits_data[235], unalignedCacheLine_bits_data[227]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_hi_3 = {unalignedCacheLine_bits_data[251], unalignedCacheLine_bits_data[243]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_3 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_hi_3, alignedDequeue_bits_data_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi_hi_3 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_3, alignedDequeue_bits_data_lo_lo_hi_hi_lo_3};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_hi_3 = {alignedDequeue_bits_data_lo_lo_hi_hi_3, alignedDequeue_bits_data_lo_lo_hi_lo_3};
  wire [31:0]   alignedDequeue_bits_data_lo_lo_3 = {alignedDequeue_bits_data_lo_lo_hi_3, alignedDequeue_bits_data_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_lo_3 = {unalignedCacheLine_bits_data[267], unalignedCacheLine_bits_data[259]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_hi_3 = {unalignedCacheLine_bits_data[283], unalignedCacheLine_bits_data[275]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_3 = {alignedDequeue_bits_data_lo_hi_lo_lo_lo_hi_3, alignedDequeue_bits_data_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_lo_3 = {unalignedCacheLine_bits_data[299], unalignedCacheLine_bits_data[291]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_hi_3 = {unalignedCacheLine_bits_data[315], unalignedCacheLine_bits_data[307]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_3 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_hi_3, alignedDequeue_bits_data_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo_lo_3 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_3, alignedDequeue_bits_data_lo_hi_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_lo_3 = {unalignedCacheLine_bits_data[331], unalignedCacheLine_bits_data[323]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_hi_3 = {unalignedCacheLine_bits_data[347], unalignedCacheLine_bits_data[339]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_3 = {alignedDequeue_bits_data_lo_hi_lo_hi_lo_hi_3, alignedDequeue_bits_data_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_lo_3 = {unalignedCacheLine_bits_data[363], unalignedCacheLine_bits_data[355]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_hi_3 = {unalignedCacheLine_bits_data[379], unalignedCacheLine_bits_data[371]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_3 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_hi_3, alignedDequeue_bits_data_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo_hi_3 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_3, alignedDequeue_bits_data_lo_hi_lo_hi_lo_3};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_lo_3 = {alignedDequeue_bits_data_lo_hi_lo_hi_3, alignedDequeue_bits_data_lo_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_lo_3 = {unalignedCacheLine_bits_data[395], unalignedCacheLine_bits_data[387]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_hi_3 = {unalignedCacheLine_bits_data[411], unalignedCacheLine_bits_data[403]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_3 = {alignedDequeue_bits_data_lo_hi_hi_lo_lo_hi_3, alignedDequeue_bits_data_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_lo_3 = {unalignedCacheLine_bits_data[427], unalignedCacheLine_bits_data[419]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_hi_3 = {unalignedCacheLine_bits_data[443], unalignedCacheLine_bits_data[435]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_3 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_hi_3, alignedDequeue_bits_data_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi_lo_3 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_3, alignedDequeue_bits_data_lo_hi_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_lo_3 = {unalignedCacheLine_bits_data[459], unalignedCacheLine_bits_data[451]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_hi_3 = {unalignedCacheLine_bits_data[475], unalignedCacheLine_bits_data[467]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_3 = {alignedDequeue_bits_data_lo_hi_hi_hi_lo_hi_3, alignedDequeue_bits_data_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_lo_3 = {unalignedCacheLine_bits_data[491], unalignedCacheLine_bits_data[483]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_hi_3 = {unalignedCacheLine_bits_data[507], unalignedCacheLine_bits_data[499]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_3 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_hi_3, alignedDequeue_bits_data_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi_hi_3 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_3, alignedDequeue_bits_data_lo_hi_hi_hi_lo_3};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_hi_3 = {alignedDequeue_bits_data_lo_hi_hi_hi_3, alignedDequeue_bits_data_lo_hi_hi_lo_3};
  wire [31:0]   alignedDequeue_bits_data_lo_hi_3 = {alignedDequeue_bits_data_lo_hi_hi_3, alignedDequeue_bits_data_lo_hi_lo_3};
  wire [63:0]   alignedDequeue_bits_data_lo_3 = {alignedDequeue_bits_data_lo_hi_3, alignedDequeue_bits_data_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_lo_3 = {memResponse_bits_data_0[11], memResponse_bits_data_0[3]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_hi_3 = {memResponse_bits_data_0[27], memResponse_bits_data_0[19]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_3 = {alignedDequeue_bits_data_hi_lo_lo_lo_lo_hi_3, alignedDequeue_bits_data_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_lo_3 = {memResponse_bits_data_0[43], memResponse_bits_data_0[35]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_hi_3 = {memResponse_bits_data_0[59], memResponse_bits_data_0[51]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_3 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_hi_3, alignedDequeue_bits_data_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo_lo_3 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_3, alignedDequeue_bits_data_hi_lo_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_lo_3 = {memResponse_bits_data_0[75], memResponse_bits_data_0[67]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_hi_3 = {memResponse_bits_data_0[91], memResponse_bits_data_0[83]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_3 = {alignedDequeue_bits_data_hi_lo_lo_hi_lo_hi_3, alignedDequeue_bits_data_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_lo_3 = {memResponse_bits_data_0[107], memResponse_bits_data_0[99]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_hi_3 = {memResponse_bits_data_0[123], memResponse_bits_data_0[115]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_3 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_hi_3, alignedDequeue_bits_data_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo_hi_3 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_3, alignedDequeue_bits_data_hi_lo_lo_hi_lo_3};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_lo_3 = {alignedDequeue_bits_data_hi_lo_lo_hi_3, alignedDequeue_bits_data_hi_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_lo_3 = {memResponse_bits_data_0[139], memResponse_bits_data_0[131]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_hi_3 = {memResponse_bits_data_0[155], memResponse_bits_data_0[147]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_3 = {alignedDequeue_bits_data_hi_lo_hi_lo_lo_hi_3, alignedDequeue_bits_data_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_lo_3 = {memResponse_bits_data_0[171], memResponse_bits_data_0[163]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_hi_3 = {memResponse_bits_data_0[187], memResponse_bits_data_0[179]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_3 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_hi_3, alignedDequeue_bits_data_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi_lo_3 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_3, alignedDequeue_bits_data_hi_lo_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_lo_3 = {memResponse_bits_data_0[203], memResponse_bits_data_0[195]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_hi_3 = {memResponse_bits_data_0[219], memResponse_bits_data_0[211]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_3 = {alignedDequeue_bits_data_hi_lo_hi_hi_lo_hi_3, alignedDequeue_bits_data_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_lo_3 = {memResponse_bits_data_0[235], memResponse_bits_data_0[227]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_hi_3 = {memResponse_bits_data_0[251], memResponse_bits_data_0[243]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_3 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_hi_3, alignedDequeue_bits_data_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi_hi_3 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_3, alignedDequeue_bits_data_hi_lo_hi_hi_lo_3};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_hi_3 = {alignedDequeue_bits_data_hi_lo_hi_hi_3, alignedDequeue_bits_data_hi_lo_hi_lo_3};
  wire [31:0]   alignedDequeue_bits_data_hi_lo_3 = {alignedDequeue_bits_data_hi_lo_hi_3, alignedDequeue_bits_data_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_lo_3 = {memResponse_bits_data_0[267], memResponse_bits_data_0[259]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_hi_3 = {memResponse_bits_data_0[283], memResponse_bits_data_0[275]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_3 = {alignedDequeue_bits_data_hi_hi_lo_lo_lo_hi_3, alignedDequeue_bits_data_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_lo_3 = {memResponse_bits_data_0[299], memResponse_bits_data_0[291]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_hi_3 = {memResponse_bits_data_0[315], memResponse_bits_data_0[307]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_3 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_hi_3, alignedDequeue_bits_data_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo_lo_3 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_3, alignedDequeue_bits_data_hi_hi_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_lo_3 = {memResponse_bits_data_0[331], memResponse_bits_data_0[323]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_hi_3 = {memResponse_bits_data_0[347], memResponse_bits_data_0[339]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_3 = {alignedDequeue_bits_data_hi_hi_lo_hi_lo_hi_3, alignedDequeue_bits_data_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_lo_3 = {memResponse_bits_data_0[363], memResponse_bits_data_0[355]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_hi_3 = {memResponse_bits_data_0[379], memResponse_bits_data_0[371]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_3 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_hi_3, alignedDequeue_bits_data_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo_hi_3 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_3, alignedDequeue_bits_data_hi_hi_lo_hi_lo_3};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_lo_3 = {alignedDequeue_bits_data_hi_hi_lo_hi_3, alignedDequeue_bits_data_hi_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_lo_3 = {memResponse_bits_data_0[395], memResponse_bits_data_0[387]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_hi_3 = {memResponse_bits_data_0[411], memResponse_bits_data_0[403]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_3 = {alignedDequeue_bits_data_hi_hi_hi_lo_lo_hi_3, alignedDequeue_bits_data_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_lo_3 = {memResponse_bits_data_0[427], memResponse_bits_data_0[419]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_hi_3 = {memResponse_bits_data_0[443], memResponse_bits_data_0[435]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_3 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_hi_3, alignedDequeue_bits_data_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi_lo_3 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_3, alignedDequeue_bits_data_hi_hi_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_lo_3 = {memResponse_bits_data_0[459], memResponse_bits_data_0[451]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_hi_3 = {memResponse_bits_data_0[475], memResponse_bits_data_0[467]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_3 = {alignedDequeue_bits_data_hi_hi_hi_hi_lo_hi_3, alignedDequeue_bits_data_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_lo_3 = {memResponse_bits_data_0[491], memResponse_bits_data_0[483]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_hi_3 = {memResponse_bits_data_0[507], memResponse_bits_data_0[499]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_3 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_hi_3, alignedDequeue_bits_data_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi_hi_3 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_3, alignedDequeue_bits_data_hi_hi_hi_hi_lo_3};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_hi_3 = {alignedDequeue_bits_data_hi_hi_hi_hi_3, alignedDequeue_bits_data_hi_hi_hi_lo_3};
  wire [31:0]   alignedDequeue_bits_data_hi_hi_3 = {alignedDequeue_bits_data_hi_hi_hi_3, alignedDequeue_bits_data_hi_hi_lo_3};
  wire [63:0]   alignedDequeue_bits_data_hi_3 = {alignedDequeue_bits_data_hi_hi_3, alignedDequeue_bits_data_hi_lo_3};
  wire [127:0]  _alignedDequeue_bits_data_T_1416 = {alignedDequeue_bits_data_hi_3, alignedDequeue_bits_data_lo_3} >> _GEN_4;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_lo_4 = {unalignedCacheLine_bits_data[12], unalignedCacheLine_bits_data[4]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_hi_4 = {unalignedCacheLine_bits_data[28], unalignedCacheLine_bits_data[20]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_4 = {alignedDequeue_bits_data_lo_lo_lo_lo_lo_hi_4, alignedDequeue_bits_data_lo_lo_lo_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_lo_4 = {unalignedCacheLine_bits_data[44], unalignedCacheLine_bits_data[36]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_hi_4 = {unalignedCacheLine_bits_data[60], unalignedCacheLine_bits_data[52]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_4 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_hi_4, alignedDequeue_bits_data_lo_lo_lo_lo_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo_lo_4 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_4, alignedDequeue_bits_data_lo_lo_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_lo_4 = {unalignedCacheLine_bits_data[76], unalignedCacheLine_bits_data[68]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_hi_4 = {unalignedCacheLine_bits_data[92], unalignedCacheLine_bits_data[84]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_4 = {alignedDequeue_bits_data_lo_lo_lo_hi_lo_hi_4, alignedDequeue_bits_data_lo_lo_lo_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_lo_4 = {unalignedCacheLine_bits_data[108], unalignedCacheLine_bits_data[100]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_hi_4 = {unalignedCacheLine_bits_data[124], unalignedCacheLine_bits_data[116]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_4 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_hi_4, alignedDequeue_bits_data_lo_lo_lo_hi_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo_hi_4 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_4, alignedDequeue_bits_data_lo_lo_lo_hi_lo_4};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_lo_4 = {alignedDequeue_bits_data_lo_lo_lo_hi_4, alignedDequeue_bits_data_lo_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_lo_4 = {unalignedCacheLine_bits_data[140], unalignedCacheLine_bits_data[132]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_hi_4 = {unalignedCacheLine_bits_data[156], unalignedCacheLine_bits_data[148]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_4 = {alignedDequeue_bits_data_lo_lo_hi_lo_lo_hi_4, alignedDequeue_bits_data_lo_lo_hi_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_lo_4 = {unalignedCacheLine_bits_data[172], unalignedCacheLine_bits_data[164]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_hi_4 = {unalignedCacheLine_bits_data[188], unalignedCacheLine_bits_data[180]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_4 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_hi_4, alignedDequeue_bits_data_lo_lo_hi_lo_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi_lo_4 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_4, alignedDequeue_bits_data_lo_lo_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_lo_4 = {unalignedCacheLine_bits_data[204], unalignedCacheLine_bits_data[196]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_hi_4 = {unalignedCacheLine_bits_data[220], unalignedCacheLine_bits_data[212]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_4 = {alignedDequeue_bits_data_lo_lo_hi_hi_lo_hi_4, alignedDequeue_bits_data_lo_lo_hi_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_lo_4 = {unalignedCacheLine_bits_data[236], unalignedCacheLine_bits_data[228]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_hi_4 = {unalignedCacheLine_bits_data[252], unalignedCacheLine_bits_data[244]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_4 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_hi_4, alignedDequeue_bits_data_lo_lo_hi_hi_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi_hi_4 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_4, alignedDequeue_bits_data_lo_lo_hi_hi_lo_4};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_hi_4 = {alignedDequeue_bits_data_lo_lo_hi_hi_4, alignedDequeue_bits_data_lo_lo_hi_lo_4};
  wire [31:0]   alignedDequeue_bits_data_lo_lo_4 = {alignedDequeue_bits_data_lo_lo_hi_4, alignedDequeue_bits_data_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_lo_4 = {unalignedCacheLine_bits_data[268], unalignedCacheLine_bits_data[260]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_hi_4 = {unalignedCacheLine_bits_data[284], unalignedCacheLine_bits_data[276]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_4 = {alignedDequeue_bits_data_lo_hi_lo_lo_lo_hi_4, alignedDequeue_bits_data_lo_hi_lo_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_lo_4 = {unalignedCacheLine_bits_data[300], unalignedCacheLine_bits_data[292]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_hi_4 = {unalignedCacheLine_bits_data[316], unalignedCacheLine_bits_data[308]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_4 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_hi_4, alignedDequeue_bits_data_lo_hi_lo_lo_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo_lo_4 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_4, alignedDequeue_bits_data_lo_hi_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_lo_4 = {unalignedCacheLine_bits_data[332], unalignedCacheLine_bits_data[324]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_hi_4 = {unalignedCacheLine_bits_data[348], unalignedCacheLine_bits_data[340]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_4 = {alignedDequeue_bits_data_lo_hi_lo_hi_lo_hi_4, alignedDequeue_bits_data_lo_hi_lo_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_lo_4 = {unalignedCacheLine_bits_data[364], unalignedCacheLine_bits_data[356]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_hi_4 = {unalignedCacheLine_bits_data[380], unalignedCacheLine_bits_data[372]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_4 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_hi_4, alignedDequeue_bits_data_lo_hi_lo_hi_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo_hi_4 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_4, alignedDequeue_bits_data_lo_hi_lo_hi_lo_4};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_lo_4 = {alignedDequeue_bits_data_lo_hi_lo_hi_4, alignedDequeue_bits_data_lo_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_lo_4 = {unalignedCacheLine_bits_data[396], unalignedCacheLine_bits_data[388]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_hi_4 = {unalignedCacheLine_bits_data[412], unalignedCacheLine_bits_data[404]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_4 = {alignedDequeue_bits_data_lo_hi_hi_lo_lo_hi_4, alignedDequeue_bits_data_lo_hi_hi_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_lo_4 = {unalignedCacheLine_bits_data[428], unalignedCacheLine_bits_data[420]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_hi_4 = {unalignedCacheLine_bits_data[444], unalignedCacheLine_bits_data[436]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_4 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_hi_4, alignedDequeue_bits_data_lo_hi_hi_lo_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi_lo_4 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_4, alignedDequeue_bits_data_lo_hi_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_lo_4 = {unalignedCacheLine_bits_data[460], unalignedCacheLine_bits_data[452]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_hi_4 = {unalignedCacheLine_bits_data[476], unalignedCacheLine_bits_data[468]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_4 = {alignedDequeue_bits_data_lo_hi_hi_hi_lo_hi_4, alignedDequeue_bits_data_lo_hi_hi_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_lo_4 = {unalignedCacheLine_bits_data[492], unalignedCacheLine_bits_data[484]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_hi_4 = {unalignedCacheLine_bits_data[508], unalignedCacheLine_bits_data[500]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_4 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_hi_4, alignedDequeue_bits_data_lo_hi_hi_hi_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi_hi_4 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_4, alignedDequeue_bits_data_lo_hi_hi_hi_lo_4};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_hi_4 = {alignedDequeue_bits_data_lo_hi_hi_hi_4, alignedDequeue_bits_data_lo_hi_hi_lo_4};
  wire [31:0]   alignedDequeue_bits_data_lo_hi_4 = {alignedDequeue_bits_data_lo_hi_hi_4, alignedDequeue_bits_data_lo_hi_lo_4};
  wire [63:0]   alignedDequeue_bits_data_lo_4 = {alignedDequeue_bits_data_lo_hi_4, alignedDequeue_bits_data_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_lo_4 = {memResponse_bits_data_0[12], memResponse_bits_data_0[4]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_hi_4 = {memResponse_bits_data_0[28], memResponse_bits_data_0[20]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_4 = {alignedDequeue_bits_data_hi_lo_lo_lo_lo_hi_4, alignedDequeue_bits_data_hi_lo_lo_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_lo_4 = {memResponse_bits_data_0[44], memResponse_bits_data_0[36]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_hi_4 = {memResponse_bits_data_0[60], memResponse_bits_data_0[52]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_4 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_hi_4, alignedDequeue_bits_data_hi_lo_lo_lo_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo_lo_4 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_4, alignedDequeue_bits_data_hi_lo_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_lo_4 = {memResponse_bits_data_0[76], memResponse_bits_data_0[68]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_hi_4 = {memResponse_bits_data_0[92], memResponse_bits_data_0[84]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_4 = {alignedDequeue_bits_data_hi_lo_lo_hi_lo_hi_4, alignedDequeue_bits_data_hi_lo_lo_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_lo_4 = {memResponse_bits_data_0[108], memResponse_bits_data_0[100]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_hi_4 = {memResponse_bits_data_0[124], memResponse_bits_data_0[116]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_4 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_hi_4, alignedDequeue_bits_data_hi_lo_lo_hi_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo_hi_4 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_4, alignedDequeue_bits_data_hi_lo_lo_hi_lo_4};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_lo_4 = {alignedDequeue_bits_data_hi_lo_lo_hi_4, alignedDequeue_bits_data_hi_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_lo_4 = {memResponse_bits_data_0[140], memResponse_bits_data_0[132]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_hi_4 = {memResponse_bits_data_0[156], memResponse_bits_data_0[148]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_4 = {alignedDequeue_bits_data_hi_lo_hi_lo_lo_hi_4, alignedDequeue_bits_data_hi_lo_hi_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_lo_4 = {memResponse_bits_data_0[172], memResponse_bits_data_0[164]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_hi_4 = {memResponse_bits_data_0[188], memResponse_bits_data_0[180]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_4 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_hi_4, alignedDequeue_bits_data_hi_lo_hi_lo_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi_lo_4 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_4, alignedDequeue_bits_data_hi_lo_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_lo_4 = {memResponse_bits_data_0[204], memResponse_bits_data_0[196]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_hi_4 = {memResponse_bits_data_0[220], memResponse_bits_data_0[212]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_4 = {alignedDequeue_bits_data_hi_lo_hi_hi_lo_hi_4, alignedDequeue_bits_data_hi_lo_hi_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_lo_4 = {memResponse_bits_data_0[236], memResponse_bits_data_0[228]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_hi_4 = {memResponse_bits_data_0[252], memResponse_bits_data_0[244]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_4 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_hi_4, alignedDequeue_bits_data_hi_lo_hi_hi_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi_hi_4 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_4, alignedDequeue_bits_data_hi_lo_hi_hi_lo_4};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_hi_4 = {alignedDequeue_bits_data_hi_lo_hi_hi_4, alignedDequeue_bits_data_hi_lo_hi_lo_4};
  wire [31:0]   alignedDequeue_bits_data_hi_lo_4 = {alignedDequeue_bits_data_hi_lo_hi_4, alignedDequeue_bits_data_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_lo_4 = {memResponse_bits_data_0[268], memResponse_bits_data_0[260]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_hi_4 = {memResponse_bits_data_0[284], memResponse_bits_data_0[276]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_4 = {alignedDequeue_bits_data_hi_hi_lo_lo_lo_hi_4, alignedDequeue_bits_data_hi_hi_lo_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_lo_4 = {memResponse_bits_data_0[300], memResponse_bits_data_0[292]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_hi_4 = {memResponse_bits_data_0[316], memResponse_bits_data_0[308]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_4 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_hi_4, alignedDequeue_bits_data_hi_hi_lo_lo_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo_lo_4 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_4, alignedDequeue_bits_data_hi_hi_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_lo_4 = {memResponse_bits_data_0[332], memResponse_bits_data_0[324]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_hi_4 = {memResponse_bits_data_0[348], memResponse_bits_data_0[340]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_4 = {alignedDequeue_bits_data_hi_hi_lo_hi_lo_hi_4, alignedDequeue_bits_data_hi_hi_lo_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_lo_4 = {memResponse_bits_data_0[364], memResponse_bits_data_0[356]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_hi_4 = {memResponse_bits_data_0[380], memResponse_bits_data_0[372]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_4 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_hi_4, alignedDequeue_bits_data_hi_hi_lo_hi_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo_hi_4 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_4, alignedDequeue_bits_data_hi_hi_lo_hi_lo_4};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_lo_4 = {alignedDequeue_bits_data_hi_hi_lo_hi_4, alignedDequeue_bits_data_hi_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_lo_4 = {memResponse_bits_data_0[396], memResponse_bits_data_0[388]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_hi_4 = {memResponse_bits_data_0[412], memResponse_bits_data_0[404]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_4 = {alignedDequeue_bits_data_hi_hi_hi_lo_lo_hi_4, alignedDequeue_bits_data_hi_hi_hi_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_lo_4 = {memResponse_bits_data_0[428], memResponse_bits_data_0[420]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_hi_4 = {memResponse_bits_data_0[444], memResponse_bits_data_0[436]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_4 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_hi_4, alignedDequeue_bits_data_hi_hi_hi_lo_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi_lo_4 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_4, alignedDequeue_bits_data_hi_hi_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_lo_4 = {memResponse_bits_data_0[460], memResponse_bits_data_0[452]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_hi_4 = {memResponse_bits_data_0[476], memResponse_bits_data_0[468]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_4 = {alignedDequeue_bits_data_hi_hi_hi_hi_lo_hi_4, alignedDequeue_bits_data_hi_hi_hi_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_lo_4 = {memResponse_bits_data_0[492], memResponse_bits_data_0[484]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_hi_4 = {memResponse_bits_data_0[508], memResponse_bits_data_0[500]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_4 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_hi_4, alignedDequeue_bits_data_hi_hi_hi_hi_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi_hi_4 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_4, alignedDequeue_bits_data_hi_hi_hi_hi_lo_4};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_hi_4 = {alignedDequeue_bits_data_hi_hi_hi_hi_4, alignedDequeue_bits_data_hi_hi_hi_lo_4};
  wire [31:0]   alignedDequeue_bits_data_hi_hi_4 = {alignedDequeue_bits_data_hi_hi_hi_4, alignedDequeue_bits_data_hi_hi_lo_4};
  wire [63:0]   alignedDequeue_bits_data_hi_4 = {alignedDequeue_bits_data_hi_hi_4, alignedDequeue_bits_data_hi_lo_4};
  wire [127:0]  _alignedDequeue_bits_data_T_1546 = {alignedDequeue_bits_data_hi_4, alignedDequeue_bits_data_lo_4} >> _GEN_4;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_lo_5 = {unalignedCacheLine_bits_data[13], unalignedCacheLine_bits_data[5]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_hi_5 = {unalignedCacheLine_bits_data[29], unalignedCacheLine_bits_data[21]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_5 = {alignedDequeue_bits_data_lo_lo_lo_lo_lo_hi_5, alignedDequeue_bits_data_lo_lo_lo_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_lo_5 = {unalignedCacheLine_bits_data[45], unalignedCacheLine_bits_data[37]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_hi_5 = {unalignedCacheLine_bits_data[61], unalignedCacheLine_bits_data[53]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_5 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_hi_5, alignedDequeue_bits_data_lo_lo_lo_lo_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo_lo_5 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_5, alignedDequeue_bits_data_lo_lo_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_lo_5 = {unalignedCacheLine_bits_data[77], unalignedCacheLine_bits_data[69]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_hi_5 = {unalignedCacheLine_bits_data[93], unalignedCacheLine_bits_data[85]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_5 = {alignedDequeue_bits_data_lo_lo_lo_hi_lo_hi_5, alignedDequeue_bits_data_lo_lo_lo_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_lo_5 = {unalignedCacheLine_bits_data[109], unalignedCacheLine_bits_data[101]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_hi_5 = {unalignedCacheLine_bits_data[125], unalignedCacheLine_bits_data[117]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_5 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_hi_5, alignedDequeue_bits_data_lo_lo_lo_hi_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo_hi_5 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_5, alignedDequeue_bits_data_lo_lo_lo_hi_lo_5};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_lo_5 = {alignedDequeue_bits_data_lo_lo_lo_hi_5, alignedDequeue_bits_data_lo_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_lo_5 = {unalignedCacheLine_bits_data[141], unalignedCacheLine_bits_data[133]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_hi_5 = {unalignedCacheLine_bits_data[157], unalignedCacheLine_bits_data[149]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_5 = {alignedDequeue_bits_data_lo_lo_hi_lo_lo_hi_5, alignedDequeue_bits_data_lo_lo_hi_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_lo_5 = {unalignedCacheLine_bits_data[173], unalignedCacheLine_bits_data[165]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_hi_5 = {unalignedCacheLine_bits_data[189], unalignedCacheLine_bits_data[181]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_5 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_hi_5, alignedDequeue_bits_data_lo_lo_hi_lo_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi_lo_5 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_5, alignedDequeue_bits_data_lo_lo_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_lo_5 = {unalignedCacheLine_bits_data[205], unalignedCacheLine_bits_data[197]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_hi_5 = {unalignedCacheLine_bits_data[221], unalignedCacheLine_bits_data[213]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_5 = {alignedDequeue_bits_data_lo_lo_hi_hi_lo_hi_5, alignedDequeue_bits_data_lo_lo_hi_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_lo_5 = {unalignedCacheLine_bits_data[237], unalignedCacheLine_bits_data[229]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_hi_5 = {unalignedCacheLine_bits_data[253], unalignedCacheLine_bits_data[245]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_5 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_hi_5, alignedDequeue_bits_data_lo_lo_hi_hi_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi_hi_5 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_5, alignedDequeue_bits_data_lo_lo_hi_hi_lo_5};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_hi_5 = {alignedDequeue_bits_data_lo_lo_hi_hi_5, alignedDequeue_bits_data_lo_lo_hi_lo_5};
  wire [31:0]   alignedDequeue_bits_data_lo_lo_5 = {alignedDequeue_bits_data_lo_lo_hi_5, alignedDequeue_bits_data_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_lo_5 = {unalignedCacheLine_bits_data[269], unalignedCacheLine_bits_data[261]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_hi_5 = {unalignedCacheLine_bits_data[285], unalignedCacheLine_bits_data[277]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_5 = {alignedDequeue_bits_data_lo_hi_lo_lo_lo_hi_5, alignedDequeue_bits_data_lo_hi_lo_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_lo_5 = {unalignedCacheLine_bits_data[301], unalignedCacheLine_bits_data[293]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_hi_5 = {unalignedCacheLine_bits_data[317], unalignedCacheLine_bits_data[309]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_5 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_hi_5, alignedDequeue_bits_data_lo_hi_lo_lo_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo_lo_5 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_5, alignedDequeue_bits_data_lo_hi_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_lo_5 = {unalignedCacheLine_bits_data[333], unalignedCacheLine_bits_data[325]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_hi_5 = {unalignedCacheLine_bits_data[349], unalignedCacheLine_bits_data[341]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_5 = {alignedDequeue_bits_data_lo_hi_lo_hi_lo_hi_5, alignedDequeue_bits_data_lo_hi_lo_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_lo_5 = {unalignedCacheLine_bits_data[365], unalignedCacheLine_bits_data[357]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_hi_5 = {unalignedCacheLine_bits_data[381], unalignedCacheLine_bits_data[373]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_5 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_hi_5, alignedDequeue_bits_data_lo_hi_lo_hi_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo_hi_5 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_5, alignedDequeue_bits_data_lo_hi_lo_hi_lo_5};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_lo_5 = {alignedDequeue_bits_data_lo_hi_lo_hi_5, alignedDequeue_bits_data_lo_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_lo_5 = {unalignedCacheLine_bits_data[397], unalignedCacheLine_bits_data[389]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_hi_5 = {unalignedCacheLine_bits_data[413], unalignedCacheLine_bits_data[405]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_5 = {alignedDequeue_bits_data_lo_hi_hi_lo_lo_hi_5, alignedDequeue_bits_data_lo_hi_hi_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_lo_5 = {unalignedCacheLine_bits_data[429], unalignedCacheLine_bits_data[421]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_hi_5 = {unalignedCacheLine_bits_data[445], unalignedCacheLine_bits_data[437]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_5 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_hi_5, alignedDequeue_bits_data_lo_hi_hi_lo_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi_lo_5 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_5, alignedDequeue_bits_data_lo_hi_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_lo_5 = {unalignedCacheLine_bits_data[461], unalignedCacheLine_bits_data[453]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_hi_5 = {unalignedCacheLine_bits_data[477], unalignedCacheLine_bits_data[469]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_5 = {alignedDequeue_bits_data_lo_hi_hi_hi_lo_hi_5, alignedDequeue_bits_data_lo_hi_hi_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_lo_5 = {unalignedCacheLine_bits_data[493], unalignedCacheLine_bits_data[485]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_hi_5 = {unalignedCacheLine_bits_data[509], unalignedCacheLine_bits_data[501]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_5 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_hi_5, alignedDequeue_bits_data_lo_hi_hi_hi_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi_hi_5 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_5, alignedDequeue_bits_data_lo_hi_hi_hi_lo_5};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_hi_5 = {alignedDequeue_bits_data_lo_hi_hi_hi_5, alignedDequeue_bits_data_lo_hi_hi_lo_5};
  wire [31:0]   alignedDequeue_bits_data_lo_hi_5 = {alignedDequeue_bits_data_lo_hi_hi_5, alignedDequeue_bits_data_lo_hi_lo_5};
  wire [63:0]   alignedDequeue_bits_data_lo_5 = {alignedDequeue_bits_data_lo_hi_5, alignedDequeue_bits_data_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_lo_5 = {memResponse_bits_data_0[13], memResponse_bits_data_0[5]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_hi_5 = {memResponse_bits_data_0[29], memResponse_bits_data_0[21]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_5 = {alignedDequeue_bits_data_hi_lo_lo_lo_lo_hi_5, alignedDequeue_bits_data_hi_lo_lo_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_lo_5 = {memResponse_bits_data_0[45], memResponse_bits_data_0[37]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_hi_5 = {memResponse_bits_data_0[61], memResponse_bits_data_0[53]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_5 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_hi_5, alignedDequeue_bits_data_hi_lo_lo_lo_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo_lo_5 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_5, alignedDequeue_bits_data_hi_lo_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_lo_5 = {memResponse_bits_data_0[77], memResponse_bits_data_0[69]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_hi_5 = {memResponse_bits_data_0[93], memResponse_bits_data_0[85]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_5 = {alignedDequeue_bits_data_hi_lo_lo_hi_lo_hi_5, alignedDequeue_bits_data_hi_lo_lo_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_lo_5 = {memResponse_bits_data_0[109], memResponse_bits_data_0[101]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_hi_5 = {memResponse_bits_data_0[125], memResponse_bits_data_0[117]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_5 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_hi_5, alignedDequeue_bits_data_hi_lo_lo_hi_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo_hi_5 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_5, alignedDequeue_bits_data_hi_lo_lo_hi_lo_5};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_lo_5 = {alignedDequeue_bits_data_hi_lo_lo_hi_5, alignedDequeue_bits_data_hi_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_lo_5 = {memResponse_bits_data_0[141], memResponse_bits_data_0[133]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_hi_5 = {memResponse_bits_data_0[157], memResponse_bits_data_0[149]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_5 = {alignedDequeue_bits_data_hi_lo_hi_lo_lo_hi_5, alignedDequeue_bits_data_hi_lo_hi_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_lo_5 = {memResponse_bits_data_0[173], memResponse_bits_data_0[165]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_hi_5 = {memResponse_bits_data_0[189], memResponse_bits_data_0[181]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_5 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_hi_5, alignedDequeue_bits_data_hi_lo_hi_lo_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi_lo_5 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_5, alignedDequeue_bits_data_hi_lo_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_lo_5 = {memResponse_bits_data_0[205], memResponse_bits_data_0[197]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_hi_5 = {memResponse_bits_data_0[221], memResponse_bits_data_0[213]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_5 = {alignedDequeue_bits_data_hi_lo_hi_hi_lo_hi_5, alignedDequeue_bits_data_hi_lo_hi_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_lo_5 = {memResponse_bits_data_0[237], memResponse_bits_data_0[229]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_hi_5 = {memResponse_bits_data_0[253], memResponse_bits_data_0[245]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_5 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_hi_5, alignedDequeue_bits_data_hi_lo_hi_hi_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi_hi_5 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_5, alignedDequeue_bits_data_hi_lo_hi_hi_lo_5};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_hi_5 = {alignedDequeue_bits_data_hi_lo_hi_hi_5, alignedDequeue_bits_data_hi_lo_hi_lo_5};
  wire [31:0]   alignedDequeue_bits_data_hi_lo_5 = {alignedDequeue_bits_data_hi_lo_hi_5, alignedDequeue_bits_data_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_lo_5 = {memResponse_bits_data_0[269], memResponse_bits_data_0[261]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_hi_5 = {memResponse_bits_data_0[285], memResponse_bits_data_0[277]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_5 = {alignedDequeue_bits_data_hi_hi_lo_lo_lo_hi_5, alignedDequeue_bits_data_hi_hi_lo_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_lo_5 = {memResponse_bits_data_0[301], memResponse_bits_data_0[293]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_hi_5 = {memResponse_bits_data_0[317], memResponse_bits_data_0[309]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_5 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_hi_5, alignedDequeue_bits_data_hi_hi_lo_lo_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo_lo_5 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_5, alignedDequeue_bits_data_hi_hi_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_lo_5 = {memResponse_bits_data_0[333], memResponse_bits_data_0[325]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_hi_5 = {memResponse_bits_data_0[349], memResponse_bits_data_0[341]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_5 = {alignedDequeue_bits_data_hi_hi_lo_hi_lo_hi_5, alignedDequeue_bits_data_hi_hi_lo_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_lo_5 = {memResponse_bits_data_0[365], memResponse_bits_data_0[357]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_hi_5 = {memResponse_bits_data_0[381], memResponse_bits_data_0[373]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_5 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_hi_5, alignedDequeue_bits_data_hi_hi_lo_hi_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo_hi_5 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_5, alignedDequeue_bits_data_hi_hi_lo_hi_lo_5};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_lo_5 = {alignedDequeue_bits_data_hi_hi_lo_hi_5, alignedDequeue_bits_data_hi_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_lo_5 = {memResponse_bits_data_0[397], memResponse_bits_data_0[389]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_hi_5 = {memResponse_bits_data_0[413], memResponse_bits_data_0[405]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_5 = {alignedDequeue_bits_data_hi_hi_hi_lo_lo_hi_5, alignedDequeue_bits_data_hi_hi_hi_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_lo_5 = {memResponse_bits_data_0[429], memResponse_bits_data_0[421]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_hi_5 = {memResponse_bits_data_0[445], memResponse_bits_data_0[437]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_5 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_hi_5, alignedDequeue_bits_data_hi_hi_hi_lo_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi_lo_5 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_5, alignedDequeue_bits_data_hi_hi_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_lo_5 = {memResponse_bits_data_0[461], memResponse_bits_data_0[453]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_hi_5 = {memResponse_bits_data_0[477], memResponse_bits_data_0[469]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_5 = {alignedDequeue_bits_data_hi_hi_hi_hi_lo_hi_5, alignedDequeue_bits_data_hi_hi_hi_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_lo_5 = {memResponse_bits_data_0[493], memResponse_bits_data_0[485]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_hi_5 = {memResponse_bits_data_0[509], memResponse_bits_data_0[501]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_5 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_hi_5, alignedDequeue_bits_data_hi_hi_hi_hi_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi_hi_5 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_5, alignedDequeue_bits_data_hi_hi_hi_hi_lo_5};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_hi_5 = {alignedDequeue_bits_data_hi_hi_hi_hi_5, alignedDequeue_bits_data_hi_hi_hi_lo_5};
  wire [31:0]   alignedDequeue_bits_data_hi_hi_5 = {alignedDequeue_bits_data_hi_hi_hi_5, alignedDequeue_bits_data_hi_hi_lo_5};
  wire [63:0]   alignedDequeue_bits_data_hi_5 = {alignedDequeue_bits_data_hi_hi_5, alignedDequeue_bits_data_hi_lo_5};
  wire [127:0]  _alignedDequeue_bits_data_T_1676 = {alignedDequeue_bits_data_hi_5, alignedDequeue_bits_data_lo_5} >> _GEN_4;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_lo_6 = {unalignedCacheLine_bits_data[14], unalignedCacheLine_bits_data[6]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_hi_6 = {unalignedCacheLine_bits_data[30], unalignedCacheLine_bits_data[22]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_6 = {alignedDequeue_bits_data_lo_lo_lo_lo_lo_hi_6, alignedDequeue_bits_data_lo_lo_lo_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_lo_6 = {unalignedCacheLine_bits_data[46], unalignedCacheLine_bits_data[38]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_hi_6 = {unalignedCacheLine_bits_data[62], unalignedCacheLine_bits_data[54]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_6 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_hi_6, alignedDequeue_bits_data_lo_lo_lo_lo_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo_lo_6 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_6, alignedDequeue_bits_data_lo_lo_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_lo_6 = {unalignedCacheLine_bits_data[78], unalignedCacheLine_bits_data[70]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_hi_6 = {unalignedCacheLine_bits_data[94], unalignedCacheLine_bits_data[86]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_6 = {alignedDequeue_bits_data_lo_lo_lo_hi_lo_hi_6, alignedDequeue_bits_data_lo_lo_lo_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_lo_6 = {unalignedCacheLine_bits_data[110], unalignedCacheLine_bits_data[102]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_hi_6 = {unalignedCacheLine_bits_data[126], unalignedCacheLine_bits_data[118]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_6 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_hi_6, alignedDequeue_bits_data_lo_lo_lo_hi_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo_hi_6 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_6, alignedDequeue_bits_data_lo_lo_lo_hi_lo_6};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_lo_6 = {alignedDequeue_bits_data_lo_lo_lo_hi_6, alignedDequeue_bits_data_lo_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_lo_6 = {unalignedCacheLine_bits_data[142], unalignedCacheLine_bits_data[134]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_hi_6 = {unalignedCacheLine_bits_data[158], unalignedCacheLine_bits_data[150]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_6 = {alignedDequeue_bits_data_lo_lo_hi_lo_lo_hi_6, alignedDequeue_bits_data_lo_lo_hi_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_lo_6 = {unalignedCacheLine_bits_data[174], unalignedCacheLine_bits_data[166]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_hi_6 = {unalignedCacheLine_bits_data[190], unalignedCacheLine_bits_data[182]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_6 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_hi_6, alignedDequeue_bits_data_lo_lo_hi_lo_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi_lo_6 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_6, alignedDequeue_bits_data_lo_lo_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_lo_6 = {unalignedCacheLine_bits_data[206], unalignedCacheLine_bits_data[198]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_hi_6 = {unalignedCacheLine_bits_data[222], unalignedCacheLine_bits_data[214]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_6 = {alignedDequeue_bits_data_lo_lo_hi_hi_lo_hi_6, alignedDequeue_bits_data_lo_lo_hi_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_lo_6 = {unalignedCacheLine_bits_data[238], unalignedCacheLine_bits_data[230]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_hi_6 = {unalignedCacheLine_bits_data[254], unalignedCacheLine_bits_data[246]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_6 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_hi_6, alignedDequeue_bits_data_lo_lo_hi_hi_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi_hi_6 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_6, alignedDequeue_bits_data_lo_lo_hi_hi_lo_6};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_hi_6 = {alignedDequeue_bits_data_lo_lo_hi_hi_6, alignedDequeue_bits_data_lo_lo_hi_lo_6};
  wire [31:0]   alignedDequeue_bits_data_lo_lo_6 = {alignedDequeue_bits_data_lo_lo_hi_6, alignedDequeue_bits_data_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_lo_6 = {unalignedCacheLine_bits_data[270], unalignedCacheLine_bits_data[262]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_hi_6 = {unalignedCacheLine_bits_data[286], unalignedCacheLine_bits_data[278]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_6 = {alignedDequeue_bits_data_lo_hi_lo_lo_lo_hi_6, alignedDequeue_bits_data_lo_hi_lo_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_lo_6 = {unalignedCacheLine_bits_data[302], unalignedCacheLine_bits_data[294]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_hi_6 = {unalignedCacheLine_bits_data[318], unalignedCacheLine_bits_data[310]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_6 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_hi_6, alignedDequeue_bits_data_lo_hi_lo_lo_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo_lo_6 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_6, alignedDequeue_bits_data_lo_hi_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_lo_6 = {unalignedCacheLine_bits_data[334], unalignedCacheLine_bits_data[326]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_hi_6 = {unalignedCacheLine_bits_data[350], unalignedCacheLine_bits_data[342]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_6 = {alignedDequeue_bits_data_lo_hi_lo_hi_lo_hi_6, alignedDequeue_bits_data_lo_hi_lo_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_lo_6 = {unalignedCacheLine_bits_data[366], unalignedCacheLine_bits_data[358]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_hi_6 = {unalignedCacheLine_bits_data[382], unalignedCacheLine_bits_data[374]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_6 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_hi_6, alignedDequeue_bits_data_lo_hi_lo_hi_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo_hi_6 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_6, alignedDequeue_bits_data_lo_hi_lo_hi_lo_6};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_lo_6 = {alignedDequeue_bits_data_lo_hi_lo_hi_6, alignedDequeue_bits_data_lo_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_lo_6 = {unalignedCacheLine_bits_data[398], unalignedCacheLine_bits_data[390]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_hi_6 = {unalignedCacheLine_bits_data[414], unalignedCacheLine_bits_data[406]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_6 = {alignedDequeue_bits_data_lo_hi_hi_lo_lo_hi_6, alignedDequeue_bits_data_lo_hi_hi_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_lo_6 = {unalignedCacheLine_bits_data[430], unalignedCacheLine_bits_data[422]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_hi_6 = {unalignedCacheLine_bits_data[446], unalignedCacheLine_bits_data[438]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_6 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_hi_6, alignedDequeue_bits_data_lo_hi_hi_lo_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi_lo_6 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_6, alignedDequeue_bits_data_lo_hi_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_lo_6 = {unalignedCacheLine_bits_data[462], unalignedCacheLine_bits_data[454]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_hi_6 = {unalignedCacheLine_bits_data[478], unalignedCacheLine_bits_data[470]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_6 = {alignedDequeue_bits_data_lo_hi_hi_hi_lo_hi_6, alignedDequeue_bits_data_lo_hi_hi_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_lo_6 = {unalignedCacheLine_bits_data[494], unalignedCacheLine_bits_data[486]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_hi_6 = {unalignedCacheLine_bits_data[510], unalignedCacheLine_bits_data[502]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_6 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_hi_6, alignedDequeue_bits_data_lo_hi_hi_hi_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi_hi_6 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_6, alignedDequeue_bits_data_lo_hi_hi_hi_lo_6};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_hi_6 = {alignedDequeue_bits_data_lo_hi_hi_hi_6, alignedDequeue_bits_data_lo_hi_hi_lo_6};
  wire [31:0]   alignedDequeue_bits_data_lo_hi_6 = {alignedDequeue_bits_data_lo_hi_hi_6, alignedDequeue_bits_data_lo_hi_lo_6};
  wire [63:0]   alignedDequeue_bits_data_lo_6 = {alignedDequeue_bits_data_lo_hi_6, alignedDequeue_bits_data_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_lo_6 = {memResponse_bits_data_0[14], memResponse_bits_data_0[6]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_hi_6 = {memResponse_bits_data_0[30], memResponse_bits_data_0[22]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_6 = {alignedDequeue_bits_data_hi_lo_lo_lo_lo_hi_6, alignedDequeue_bits_data_hi_lo_lo_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_lo_6 = {memResponse_bits_data_0[46], memResponse_bits_data_0[38]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_hi_6 = {memResponse_bits_data_0[62], memResponse_bits_data_0[54]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_6 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_hi_6, alignedDequeue_bits_data_hi_lo_lo_lo_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo_lo_6 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_6, alignedDequeue_bits_data_hi_lo_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_lo_6 = {memResponse_bits_data_0[78], memResponse_bits_data_0[70]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_hi_6 = {memResponse_bits_data_0[94], memResponse_bits_data_0[86]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_6 = {alignedDequeue_bits_data_hi_lo_lo_hi_lo_hi_6, alignedDequeue_bits_data_hi_lo_lo_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_lo_6 = {memResponse_bits_data_0[110], memResponse_bits_data_0[102]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_hi_6 = {memResponse_bits_data_0[126], memResponse_bits_data_0[118]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_6 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_hi_6, alignedDequeue_bits_data_hi_lo_lo_hi_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo_hi_6 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_6, alignedDequeue_bits_data_hi_lo_lo_hi_lo_6};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_lo_6 = {alignedDequeue_bits_data_hi_lo_lo_hi_6, alignedDequeue_bits_data_hi_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_lo_6 = {memResponse_bits_data_0[142], memResponse_bits_data_0[134]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_hi_6 = {memResponse_bits_data_0[158], memResponse_bits_data_0[150]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_6 = {alignedDequeue_bits_data_hi_lo_hi_lo_lo_hi_6, alignedDequeue_bits_data_hi_lo_hi_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_lo_6 = {memResponse_bits_data_0[174], memResponse_bits_data_0[166]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_hi_6 = {memResponse_bits_data_0[190], memResponse_bits_data_0[182]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_6 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_hi_6, alignedDequeue_bits_data_hi_lo_hi_lo_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi_lo_6 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_6, alignedDequeue_bits_data_hi_lo_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_lo_6 = {memResponse_bits_data_0[206], memResponse_bits_data_0[198]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_hi_6 = {memResponse_bits_data_0[222], memResponse_bits_data_0[214]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_6 = {alignedDequeue_bits_data_hi_lo_hi_hi_lo_hi_6, alignedDequeue_bits_data_hi_lo_hi_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_lo_6 = {memResponse_bits_data_0[238], memResponse_bits_data_0[230]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_hi_6 = {memResponse_bits_data_0[254], memResponse_bits_data_0[246]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_6 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_hi_6, alignedDequeue_bits_data_hi_lo_hi_hi_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi_hi_6 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_6, alignedDequeue_bits_data_hi_lo_hi_hi_lo_6};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_hi_6 = {alignedDequeue_bits_data_hi_lo_hi_hi_6, alignedDequeue_bits_data_hi_lo_hi_lo_6};
  wire [31:0]   alignedDequeue_bits_data_hi_lo_6 = {alignedDequeue_bits_data_hi_lo_hi_6, alignedDequeue_bits_data_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_lo_6 = {memResponse_bits_data_0[270], memResponse_bits_data_0[262]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_hi_6 = {memResponse_bits_data_0[286], memResponse_bits_data_0[278]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_6 = {alignedDequeue_bits_data_hi_hi_lo_lo_lo_hi_6, alignedDequeue_bits_data_hi_hi_lo_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_lo_6 = {memResponse_bits_data_0[302], memResponse_bits_data_0[294]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_hi_6 = {memResponse_bits_data_0[318], memResponse_bits_data_0[310]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_6 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_hi_6, alignedDequeue_bits_data_hi_hi_lo_lo_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo_lo_6 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_6, alignedDequeue_bits_data_hi_hi_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_lo_6 = {memResponse_bits_data_0[334], memResponse_bits_data_0[326]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_hi_6 = {memResponse_bits_data_0[350], memResponse_bits_data_0[342]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_6 = {alignedDequeue_bits_data_hi_hi_lo_hi_lo_hi_6, alignedDequeue_bits_data_hi_hi_lo_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_lo_6 = {memResponse_bits_data_0[366], memResponse_bits_data_0[358]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_hi_6 = {memResponse_bits_data_0[382], memResponse_bits_data_0[374]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_6 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_hi_6, alignedDequeue_bits_data_hi_hi_lo_hi_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo_hi_6 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_6, alignedDequeue_bits_data_hi_hi_lo_hi_lo_6};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_lo_6 = {alignedDequeue_bits_data_hi_hi_lo_hi_6, alignedDequeue_bits_data_hi_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_lo_6 = {memResponse_bits_data_0[398], memResponse_bits_data_0[390]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_hi_6 = {memResponse_bits_data_0[414], memResponse_bits_data_0[406]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_6 = {alignedDequeue_bits_data_hi_hi_hi_lo_lo_hi_6, alignedDequeue_bits_data_hi_hi_hi_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_lo_6 = {memResponse_bits_data_0[430], memResponse_bits_data_0[422]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_hi_6 = {memResponse_bits_data_0[446], memResponse_bits_data_0[438]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_6 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_hi_6, alignedDequeue_bits_data_hi_hi_hi_lo_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi_lo_6 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_6, alignedDequeue_bits_data_hi_hi_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_lo_6 = {memResponse_bits_data_0[462], memResponse_bits_data_0[454]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_hi_6 = {memResponse_bits_data_0[478], memResponse_bits_data_0[470]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_6 = {alignedDequeue_bits_data_hi_hi_hi_hi_lo_hi_6, alignedDequeue_bits_data_hi_hi_hi_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_lo_6 = {memResponse_bits_data_0[494], memResponse_bits_data_0[486]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_hi_6 = {memResponse_bits_data_0[510], memResponse_bits_data_0[502]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_6 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_hi_6, alignedDequeue_bits_data_hi_hi_hi_hi_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi_hi_6 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_6, alignedDequeue_bits_data_hi_hi_hi_hi_lo_6};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_hi_6 = {alignedDequeue_bits_data_hi_hi_hi_hi_6, alignedDequeue_bits_data_hi_hi_hi_lo_6};
  wire [31:0]   alignedDequeue_bits_data_hi_hi_6 = {alignedDequeue_bits_data_hi_hi_hi_6, alignedDequeue_bits_data_hi_hi_lo_6};
  wire [63:0]   alignedDequeue_bits_data_hi_6 = {alignedDequeue_bits_data_hi_hi_6, alignedDequeue_bits_data_hi_lo_6};
  wire [127:0]  _alignedDequeue_bits_data_T_1806 = {alignedDequeue_bits_data_hi_6, alignedDequeue_bits_data_lo_6} >> _GEN_4;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_lo_7 = {unalignedCacheLine_bits_data[15], unalignedCacheLine_bits_data[7]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_hi_7 = {unalignedCacheLine_bits_data[31], unalignedCacheLine_bits_data[23]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_7 = {alignedDequeue_bits_data_lo_lo_lo_lo_lo_hi_7, alignedDequeue_bits_data_lo_lo_lo_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_lo_7 = {unalignedCacheLine_bits_data[47], unalignedCacheLine_bits_data[39]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_hi_7 = {unalignedCacheLine_bits_data[63], unalignedCacheLine_bits_data[55]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_7 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_hi_7, alignedDequeue_bits_data_lo_lo_lo_lo_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo_lo_7 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_7, alignedDequeue_bits_data_lo_lo_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_lo_7 = {unalignedCacheLine_bits_data[79], unalignedCacheLine_bits_data[71]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_hi_7 = {unalignedCacheLine_bits_data[95], unalignedCacheLine_bits_data[87]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_7 = {alignedDequeue_bits_data_lo_lo_lo_hi_lo_hi_7, alignedDequeue_bits_data_lo_lo_lo_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_lo_7 = {unalignedCacheLine_bits_data[111], unalignedCacheLine_bits_data[103]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_hi_7 = {unalignedCacheLine_bits_data[127], unalignedCacheLine_bits_data[119]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_7 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_hi_7, alignedDequeue_bits_data_lo_lo_lo_hi_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo_hi_7 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_7, alignedDequeue_bits_data_lo_lo_lo_hi_lo_7};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_lo_7 = {alignedDequeue_bits_data_lo_lo_lo_hi_7, alignedDequeue_bits_data_lo_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_lo_7 = {unalignedCacheLine_bits_data[143], unalignedCacheLine_bits_data[135]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_hi_7 = {unalignedCacheLine_bits_data[159], unalignedCacheLine_bits_data[151]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_7 = {alignedDequeue_bits_data_lo_lo_hi_lo_lo_hi_7, alignedDequeue_bits_data_lo_lo_hi_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_lo_7 = {unalignedCacheLine_bits_data[175], unalignedCacheLine_bits_data[167]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_hi_7 = {unalignedCacheLine_bits_data[191], unalignedCacheLine_bits_data[183]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_7 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_hi_7, alignedDequeue_bits_data_lo_lo_hi_lo_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi_lo_7 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_7, alignedDequeue_bits_data_lo_lo_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_lo_7 = {unalignedCacheLine_bits_data[207], unalignedCacheLine_bits_data[199]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_hi_7 = {unalignedCacheLine_bits_data[223], unalignedCacheLine_bits_data[215]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_7 = {alignedDequeue_bits_data_lo_lo_hi_hi_lo_hi_7, alignedDequeue_bits_data_lo_lo_hi_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_lo_7 = {unalignedCacheLine_bits_data[239], unalignedCacheLine_bits_data[231]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_hi_7 = {unalignedCacheLine_bits_data[255], unalignedCacheLine_bits_data[247]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_7 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_hi_7, alignedDequeue_bits_data_lo_lo_hi_hi_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi_hi_7 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_7, alignedDequeue_bits_data_lo_lo_hi_hi_lo_7};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_hi_7 = {alignedDequeue_bits_data_lo_lo_hi_hi_7, alignedDequeue_bits_data_lo_lo_hi_lo_7};
  wire [31:0]   alignedDequeue_bits_data_lo_lo_7 = {alignedDequeue_bits_data_lo_lo_hi_7, alignedDequeue_bits_data_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_lo_7 = {unalignedCacheLine_bits_data[271], unalignedCacheLine_bits_data[263]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_hi_7 = {unalignedCacheLine_bits_data[287], unalignedCacheLine_bits_data[279]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_7 = {alignedDequeue_bits_data_lo_hi_lo_lo_lo_hi_7, alignedDequeue_bits_data_lo_hi_lo_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_lo_7 = {unalignedCacheLine_bits_data[303], unalignedCacheLine_bits_data[295]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_hi_7 = {unalignedCacheLine_bits_data[319], unalignedCacheLine_bits_data[311]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_7 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_hi_7, alignedDequeue_bits_data_lo_hi_lo_lo_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo_lo_7 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_7, alignedDequeue_bits_data_lo_hi_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_lo_7 = {unalignedCacheLine_bits_data[335], unalignedCacheLine_bits_data[327]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_hi_7 = {unalignedCacheLine_bits_data[351], unalignedCacheLine_bits_data[343]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_7 = {alignedDequeue_bits_data_lo_hi_lo_hi_lo_hi_7, alignedDequeue_bits_data_lo_hi_lo_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_lo_7 = {unalignedCacheLine_bits_data[367], unalignedCacheLine_bits_data[359]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_hi_7 = {unalignedCacheLine_bits_data[383], unalignedCacheLine_bits_data[375]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_7 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_hi_7, alignedDequeue_bits_data_lo_hi_lo_hi_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo_hi_7 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_7, alignedDequeue_bits_data_lo_hi_lo_hi_lo_7};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_lo_7 = {alignedDequeue_bits_data_lo_hi_lo_hi_7, alignedDequeue_bits_data_lo_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_lo_7 = {unalignedCacheLine_bits_data[399], unalignedCacheLine_bits_data[391]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_hi_7 = {unalignedCacheLine_bits_data[415], unalignedCacheLine_bits_data[407]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_7 = {alignedDequeue_bits_data_lo_hi_hi_lo_lo_hi_7, alignedDequeue_bits_data_lo_hi_hi_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_lo_7 = {unalignedCacheLine_bits_data[431], unalignedCacheLine_bits_data[423]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_hi_7 = {unalignedCacheLine_bits_data[447], unalignedCacheLine_bits_data[439]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_7 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_hi_7, alignedDequeue_bits_data_lo_hi_hi_lo_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi_lo_7 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_7, alignedDequeue_bits_data_lo_hi_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_lo_7 = {unalignedCacheLine_bits_data[463], unalignedCacheLine_bits_data[455]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_hi_7 = {unalignedCacheLine_bits_data[479], unalignedCacheLine_bits_data[471]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_7 = {alignedDequeue_bits_data_lo_hi_hi_hi_lo_hi_7, alignedDequeue_bits_data_lo_hi_hi_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_lo_7 = {unalignedCacheLine_bits_data[495], unalignedCacheLine_bits_data[487]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_hi_7 = {unalignedCacheLine_bits_data[511], unalignedCacheLine_bits_data[503]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_7 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_hi_7, alignedDequeue_bits_data_lo_hi_hi_hi_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi_hi_7 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_7, alignedDequeue_bits_data_lo_hi_hi_hi_lo_7};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_hi_7 = {alignedDequeue_bits_data_lo_hi_hi_hi_7, alignedDequeue_bits_data_lo_hi_hi_lo_7};
  wire [31:0]   alignedDequeue_bits_data_lo_hi_7 = {alignedDequeue_bits_data_lo_hi_hi_7, alignedDequeue_bits_data_lo_hi_lo_7};
  wire [63:0]   alignedDequeue_bits_data_lo_7 = {alignedDequeue_bits_data_lo_hi_7, alignedDequeue_bits_data_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_lo_7 = {memResponse_bits_data_0[15], memResponse_bits_data_0[7]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_hi_7 = {memResponse_bits_data_0[31], memResponse_bits_data_0[23]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_7 = {alignedDequeue_bits_data_hi_lo_lo_lo_lo_hi_7, alignedDequeue_bits_data_hi_lo_lo_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_lo_7 = {memResponse_bits_data_0[47], memResponse_bits_data_0[39]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_hi_7 = {memResponse_bits_data_0[63], memResponse_bits_data_0[55]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_7 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_hi_7, alignedDequeue_bits_data_hi_lo_lo_lo_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo_lo_7 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_7, alignedDequeue_bits_data_hi_lo_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_lo_7 = {memResponse_bits_data_0[79], memResponse_bits_data_0[71]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_hi_7 = {memResponse_bits_data_0[95], memResponse_bits_data_0[87]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_7 = {alignedDequeue_bits_data_hi_lo_lo_hi_lo_hi_7, alignedDequeue_bits_data_hi_lo_lo_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_lo_7 = {memResponse_bits_data_0[111], memResponse_bits_data_0[103]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_hi_7 = {memResponse_bits_data_0[127], memResponse_bits_data_0[119]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_7 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_hi_7, alignedDequeue_bits_data_hi_lo_lo_hi_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo_hi_7 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_7, alignedDequeue_bits_data_hi_lo_lo_hi_lo_7};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_lo_7 = {alignedDequeue_bits_data_hi_lo_lo_hi_7, alignedDequeue_bits_data_hi_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_lo_7 = {memResponse_bits_data_0[143], memResponse_bits_data_0[135]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_hi_7 = {memResponse_bits_data_0[159], memResponse_bits_data_0[151]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_7 = {alignedDequeue_bits_data_hi_lo_hi_lo_lo_hi_7, alignedDequeue_bits_data_hi_lo_hi_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_lo_7 = {memResponse_bits_data_0[175], memResponse_bits_data_0[167]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_hi_7 = {memResponse_bits_data_0[191], memResponse_bits_data_0[183]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_7 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_hi_7, alignedDequeue_bits_data_hi_lo_hi_lo_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi_lo_7 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_7, alignedDequeue_bits_data_hi_lo_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_lo_7 = {memResponse_bits_data_0[207], memResponse_bits_data_0[199]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_hi_7 = {memResponse_bits_data_0[223], memResponse_bits_data_0[215]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_7 = {alignedDequeue_bits_data_hi_lo_hi_hi_lo_hi_7, alignedDequeue_bits_data_hi_lo_hi_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_lo_7 = {memResponse_bits_data_0[239], memResponse_bits_data_0[231]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_hi_7 = {memResponse_bits_data_0[255], memResponse_bits_data_0[247]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_7 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_hi_7, alignedDequeue_bits_data_hi_lo_hi_hi_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi_hi_7 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_7, alignedDequeue_bits_data_hi_lo_hi_hi_lo_7};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_hi_7 = {alignedDequeue_bits_data_hi_lo_hi_hi_7, alignedDequeue_bits_data_hi_lo_hi_lo_7};
  wire [31:0]   alignedDequeue_bits_data_hi_lo_7 = {alignedDequeue_bits_data_hi_lo_hi_7, alignedDequeue_bits_data_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_lo_7 = {memResponse_bits_data_0[271], memResponse_bits_data_0[263]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_hi_7 = {memResponse_bits_data_0[287], memResponse_bits_data_0[279]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_7 = {alignedDequeue_bits_data_hi_hi_lo_lo_lo_hi_7, alignedDequeue_bits_data_hi_hi_lo_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_lo_7 = {memResponse_bits_data_0[303], memResponse_bits_data_0[295]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_hi_7 = {memResponse_bits_data_0[319], memResponse_bits_data_0[311]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_7 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_hi_7, alignedDequeue_bits_data_hi_hi_lo_lo_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo_lo_7 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_7, alignedDequeue_bits_data_hi_hi_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_lo_7 = {memResponse_bits_data_0[335], memResponse_bits_data_0[327]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_hi_7 = {memResponse_bits_data_0[351], memResponse_bits_data_0[343]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_7 = {alignedDequeue_bits_data_hi_hi_lo_hi_lo_hi_7, alignedDequeue_bits_data_hi_hi_lo_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_lo_7 = {memResponse_bits_data_0[367], memResponse_bits_data_0[359]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_hi_7 = {memResponse_bits_data_0[383], memResponse_bits_data_0[375]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_7 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_hi_7, alignedDequeue_bits_data_hi_hi_lo_hi_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo_hi_7 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_7, alignedDequeue_bits_data_hi_hi_lo_hi_lo_7};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_lo_7 = {alignedDequeue_bits_data_hi_hi_lo_hi_7, alignedDequeue_bits_data_hi_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_lo_7 = {memResponse_bits_data_0[399], memResponse_bits_data_0[391]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_hi_7 = {memResponse_bits_data_0[415], memResponse_bits_data_0[407]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_7 = {alignedDequeue_bits_data_hi_hi_hi_lo_lo_hi_7, alignedDequeue_bits_data_hi_hi_hi_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_lo_7 = {memResponse_bits_data_0[431], memResponse_bits_data_0[423]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_hi_7 = {memResponse_bits_data_0[447], memResponse_bits_data_0[439]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_7 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_hi_7, alignedDequeue_bits_data_hi_hi_hi_lo_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi_lo_7 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_7, alignedDequeue_bits_data_hi_hi_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_lo_7 = {memResponse_bits_data_0[463], memResponse_bits_data_0[455]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_hi_7 = {memResponse_bits_data_0[479], memResponse_bits_data_0[471]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_7 = {alignedDequeue_bits_data_hi_hi_hi_hi_lo_hi_7, alignedDequeue_bits_data_hi_hi_hi_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_lo_7 = {memResponse_bits_data_0[495], memResponse_bits_data_0[487]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_hi_7 = {memResponse_bits_data_0[511], memResponse_bits_data_0[503]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_7 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_hi_7, alignedDequeue_bits_data_hi_hi_hi_hi_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi_hi_7 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_7, alignedDequeue_bits_data_hi_hi_hi_hi_lo_7};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_hi_7 = {alignedDequeue_bits_data_hi_hi_hi_hi_7, alignedDequeue_bits_data_hi_hi_hi_lo_7};
  wire [31:0]   alignedDequeue_bits_data_hi_hi_7 = {alignedDequeue_bits_data_hi_hi_hi_7, alignedDequeue_bits_data_hi_hi_lo_7};
  wire [63:0]   alignedDequeue_bits_data_hi_7 = {alignedDequeue_bits_data_hi_hi_7, alignedDequeue_bits_data_hi_lo_7};
  wire [127:0]  _alignedDequeue_bits_data_T_1936 = {alignedDequeue_bits_data_hi_7, alignedDequeue_bits_data_lo_7} >> _GEN_4;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_8 = {_alignedDequeue_bits_data_T_1156[0], _alignedDequeue_bits_data_T_1026[0]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_8 = {_alignedDequeue_bits_data_T_1416[0], _alignedDequeue_bits_data_T_1286[0]};
  wire [3:0]    alignedDequeue_bits_data_lo_8 = {alignedDequeue_bits_data_lo_hi_8, alignedDequeue_bits_data_lo_lo_8};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_8 = {_alignedDequeue_bits_data_T_1676[0], _alignedDequeue_bits_data_T_1546[0]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_8 = {_alignedDequeue_bits_data_T_1936[0], _alignedDequeue_bits_data_T_1806[0]};
  wire [3:0]    alignedDequeue_bits_data_hi_8 = {alignedDequeue_bits_data_hi_hi_8, alignedDequeue_bits_data_hi_lo_8};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_9 = {_alignedDequeue_bits_data_T_1156[1], _alignedDequeue_bits_data_T_1026[1]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_9 = {_alignedDequeue_bits_data_T_1416[1], _alignedDequeue_bits_data_T_1286[1]};
  wire [3:0]    alignedDequeue_bits_data_lo_9 = {alignedDequeue_bits_data_lo_hi_9, alignedDequeue_bits_data_lo_lo_9};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_9 = {_alignedDequeue_bits_data_T_1676[1], _alignedDequeue_bits_data_T_1546[1]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_9 = {_alignedDequeue_bits_data_T_1936[1], _alignedDequeue_bits_data_T_1806[1]};
  wire [3:0]    alignedDequeue_bits_data_hi_9 = {alignedDequeue_bits_data_hi_hi_9, alignedDequeue_bits_data_hi_lo_9};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_10 = {_alignedDequeue_bits_data_T_1156[2], _alignedDequeue_bits_data_T_1026[2]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_10 = {_alignedDequeue_bits_data_T_1416[2], _alignedDequeue_bits_data_T_1286[2]};
  wire [3:0]    alignedDequeue_bits_data_lo_10 = {alignedDequeue_bits_data_lo_hi_10, alignedDequeue_bits_data_lo_lo_10};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_10 = {_alignedDequeue_bits_data_T_1676[2], _alignedDequeue_bits_data_T_1546[2]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_10 = {_alignedDequeue_bits_data_T_1936[2], _alignedDequeue_bits_data_T_1806[2]};
  wire [3:0]    alignedDequeue_bits_data_hi_10 = {alignedDequeue_bits_data_hi_hi_10, alignedDequeue_bits_data_hi_lo_10};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_11 = {_alignedDequeue_bits_data_T_1156[3], _alignedDequeue_bits_data_T_1026[3]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_11 = {_alignedDequeue_bits_data_T_1416[3], _alignedDequeue_bits_data_T_1286[3]};
  wire [3:0]    alignedDequeue_bits_data_lo_11 = {alignedDequeue_bits_data_lo_hi_11, alignedDequeue_bits_data_lo_lo_11};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_11 = {_alignedDequeue_bits_data_T_1676[3], _alignedDequeue_bits_data_T_1546[3]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_11 = {_alignedDequeue_bits_data_T_1936[3], _alignedDequeue_bits_data_T_1806[3]};
  wire [3:0]    alignedDequeue_bits_data_hi_11 = {alignedDequeue_bits_data_hi_hi_11, alignedDequeue_bits_data_hi_lo_11};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_12 = {_alignedDequeue_bits_data_T_1156[4], _alignedDequeue_bits_data_T_1026[4]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_12 = {_alignedDequeue_bits_data_T_1416[4], _alignedDequeue_bits_data_T_1286[4]};
  wire [3:0]    alignedDequeue_bits_data_lo_12 = {alignedDequeue_bits_data_lo_hi_12, alignedDequeue_bits_data_lo_lo_12};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_12 = {_alignedDequeue_bits_data_T_1676[4], _alignedDequeue_bits_data_T_1546[4]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_12 = {_alignedDequeue_bits_data_T_1936[4], _alignedDequeue_bits_data_T_1806[4]};
  wire [3:0]    alignedDequeue_bits_data_hi_12 = {alignedDequeue_bits_data_hi_hi_12, alignedDequeue_bits_data_hi_lo_12};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_13 = {_alignedDequeue_bits_data_T_1156[5], _alignedDequeue_bits_data_T_1026[5]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_13 = {_alignedDequeue_bits_data_T_1416[5], _alignedDequeue_bits_data_T_1286[5]};
  wire [3:0]    alignedDequeue_bits_data_lo_13 = {alignedDequeue_bits_data_lo_hi_13, alignedDequeue_bits_data_lo_lo_13};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_13 = {_alignedDequeue_bits_data_T_1676[5], _alignedDequeue_bits_data_T_1546[5]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_13 = {_alignedDequeue_bits_data_T_1936[5], _alignedDequeue_bits_data_T_1806[5]};
  wire [3:0]    alignedDequeue_bits_data_hi_13 = {alignedDequeue_bits_data_hi_hi_13, alignedDequeue_bits_data_hi_lo_13};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_14 = {_alignedDequeue_bits_data_T_1156[6], _alignedDequeue_bits_data_T_1026[6]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_14 = {_alignedDequeue_bits_data_T_1416[6], _alignedDequeue_bits_data_T_1286[6]};
  wire [3:0]    alignedDequeue_bits_data_lo_14 = {alignedDequeue_bits_data_lo_hi_14, alignedDequeue_bits_data_lo_lo_14};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_14 = {_alignedDequeue_bits_data_T_1676[6], _alignedDequeue_bits_data_T_1546[6]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_14 = {_alignedDequeue_bits_data_T_1936[6], _alignedDequeue_bits_data_T_1806[6]};
  wire [3:0]    alignedDequeue_bits_data_hi_14 = {alignedDequeue_bits_data_hi_hi_14, alignedDequeue_bits_data_hi_lo_14};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_15 = {_alignedDequeue_bits_data_T_1156[7], _alignedDequeue_bits_data_T_1026[7]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_15 = {_alignedDequeue_bits_data_T_1416[7], _alignedDequeue_bits_data_T_1286[7]};
  wire [3:0]    alignedDequeue_bits_data_lo_15 = {alignedDequeue_bits_data_lo_hi_15, alignedDequeue_bits_data_lo_lo_15};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_15 = {_alignedDequeue_bits_data_T_1676[7], _alignedDequeue_bits_data_T_1546[7]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_15 = {_alignedDequeue_bits_data_T_1936[7], _alignedDequeue_bits_data_T_1806[7]};
  wire [3:0]    alignedDequeue_bits_data_hi_15 = {alignedDequeue_bits_data_hi_hi_15, alignedDequeue_bits_data_hi_lo_15};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_16 = {_alignedDequeue_bits_data_T_1156[8], _alignedDequeue_bits_data_T_1026[8]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_16 = {_alignedDequeue_bits_data_T_1416[8], _alignedDequeue_bits_data_T_1286[8]};
  wire [3:0]    alignedDequeue_bits_data_lo_16 = {alignedDequeue_bits_data_lo_hi_16, alignedDequeue_bits_data_lo_lo_16};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_16 = {_alignedDequeue_bits_data_T_1676[8], _alignedDequeue_bits_data_T_1546[8]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_16 = {_alignedDequeue_bits_data_T_1936[8], _alignedDequeue_bits_data_T_1806[8]};
  wire [3:0]    alignedDequeue_bits_data_hi_16 = {alignedDequeue_bits_data_hi_hi_16, alignedDequeue_bits_data_hi_lo_16};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_17 = {_alignedDequeue_bits_data_T_1156[9], _alignedDequeue_bits_data_T_1026[9]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_17 = {_alignedDequeue_bits_data_T_1416[9], _alignedDequeue_bits_data_T_1286[9]};
  wire [3:0]    alignedDequeue_bits_data_lo_17 = {alignedDequeue_bits_data_lo_hi_17, alignedDequeue_bits_data_lo_lo_17};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_17 = {_alignedDequeue_bits_data_T_1676[9], _alignedDequeue_bits_data_T_1546[9]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_17 = {_alignedDequeue_bits_data_T_1936[9], _alignedDequeue_bits_data_T_1806[9]};
  wire [3:0]    alignedDequeue_bits_data_hi_17 = {alignedDequeue_bits_data_hi_hi_17, alignedDequeue_bits_data_hi_lo_17};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_18 = {_alignedDequeue_bits_data_T_1156[10], _alignedDequeue_bits_data_T_1026[10]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_18 = {_alignedDequeue_bits_data_T_1416[10], _alignedDequeue_bits_data_T_1286[10]};
  wire [3:0]    alignedDequeue_bits_data_lo_18 = {alignedDequeue_bits_data_lo_hi_18, alignedDequeue_bits_data_lo_lo_18};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_18 = {_alignedDequeue_bits_data_T_1676[10], _alignedDequeue_bits_data_T_1546[10]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_18 = {_alignedDequeue_bits_data_T_1936[10], _alignedDequeue_bits_data_T_1806[10]};
  wire [3:0]    alignedDequeue_bits_data_hi_18 = {alignedDequeue_bits_data_hi_hi_18, alignedDequeue_bits_data_hi_lo_18};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_19 = {_alignedDequeue_bits_data_T_1156[11], _alignedDequeue_bits_data_T_1026[11]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_19 = {_alignedDequeue_bits_data_T_1416[11], _alignedDequeue_bits_data_T_1286[11]};
  wire [3:0]    alignedDequeue_bits_data_lo_19 = {alignedDequeue_bits_data_lo_hi_19, alignedDequeue_bits_data_lo_lo_19};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_19 = {_alignedDequeue_bits_data_T_1676[11], _alignedDequeue_bits_data_T_1546[11]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_19 = {_alignedDequeue_bits_data_T_1936[11], _alignedDequeue_bits_data_T_1806[11]};
  wire [3:0]    alignedDequeue_bits_data_hi_19 = {alignedDequeue_bits_data_hi_hi_19, alignedDequeue_bits_data_hi_lo_19};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_20 = {_alignedDequeue_bits_data_T_1156[12], _alignedDequeue_bits_data_T_1026[12]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_20 = {_alignedDequeue_bits_data_T_1416[12], _alignedDequeue_bits_data_T_1286[12]};
  wire [3:0]    alignedDequeue_bits_data_lo_20 = {alignedDequeue_bits_data_lo_hi_20, alignedDequeue_bits_data_lo_lo_20};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_20 = {_alignedDequeue_bits_data_T_1676[12], _alignedDequeue_bits_data_T_1546[12]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_20 = {_alignedDequeue_bits_data_T_1936[12], _alignedDequeue_bits_data_T_1806[12]};
  wire [3:0]    alignedDequeue_bits_data_hi_20 = {alignedDequeue_bits_data_hi_hi_20, alignedDequeue_bits_data_hi_lo_20};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_21 = {_alignedDequeue_bits_data_T_1156[13], _alignedDequeue_bits_data_T_1026[13]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_21 = {_alignedDequeue_bits_data_T_1416[13], _alignedDequeue_bits_data_T_1286[13]};
  wire [3:0]    alignedDequeue_bits_data_lo_21 = {alignedDequeue_bits_data_lo_hi_21, alignedDequeue_bits_data_lo_lo_21};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_21 = {_alignedDequeue_bits_data_T_1676[13], _alignedDequeue_bits_data_T_1546[13]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_21 = {_alignedDequeue_bits_data_T_1936[13], _alignedDequeue_bits_data_T_1806[13]};
  wire [3:0]    alignedDequeue_bits_data_hi_21 = {alignedDequeue_bits_data_hi_hi_21, alignedDequeue_bits_data_hi_lo_21};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_22 = {_alignedDequeue_bits_data_T_1156[14], _alignedDequeue_bits_data_T_1026[14]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_22 = {_alignedDequeue_bits_data_T_1416[14], _alignedDequeue_bits_data_T_1286[14]};
  wire [3:0]    alignedDequeue_bits_data_lo_22 = {alignedDequeue_bits_data_lo_hi_22, alignedDequeue_bits_data_lo_lo_22};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_22 = {_alignedDequeue_bits_data_T_1676[14], _alignedDequeue_bits_data_T_1546[14]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_22 = {_alignedDequeue_bits_data_T_1936[14], _alignedDequeue_bits_data_T_1806[14]};
  wire [3:0]    alignedDequeue_bits_data_hi_22 = {alignedDequeue_bits_data_hi_hi_22, alignedDequeue_bits_data_hi_lo_22};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_23 = {_alignedDequeue_bits_data_T_1156[15], _alignedDequeue_bits_data_T_1026[15]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_23 = {_alignedDequeue_bits_data_T_1416[15], _alignedDequeue_bits_data_T_1286[15]};
  wire [3:0]    alignedDequeue_bits_data_lo_23 = {alignedDequeue_bits_data_lo_hi_23, alignedDequeue_bits_data_lo_lo_23};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_23 = {_alignedDequeue_bits_data_T_1676[15], _alignedDequeue_bits_data_T_1546[15]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_23 = {_alignedDequeue_bits_data_T_1936[15], _alignedDequeue_bits_data_T_1806[15]};
  wire [3:0]    alignedDequeue_bits_data_hi_23 = {alignedDequeue_bits_data_hi_hi_23, alignedDequeue_bits_data_hi_lo_23};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_24 = {_alignedDequeue_bits_data_T_1156[16], _alignedDequeue_bits_data_T_1026[16]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_24 = {_alignedDequeue_bits_data_T_1416[16], _alignedDequeue_bits_data_T_1286[16]};
  wire [3:0]    alignedDequeue_bits_data_lo_24 = {alignedDequeue_bits_data_lo_hi_24, alignedDequeue_bits_data_lo_lo_24};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_24 = {_alignedDequeue_bits_data_T_1676[16], _alignedDequeue_bits_data_T_1546[16]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_24 = {_alignedDequeue_bits_data_T_1936[16], _alignedDequeue_bits_data_T_1806[16]};
  wire [3:0]    alignedDequeue_bits_data_hi_24 = {alignedDequeue_bits_data_hi_hi_24, alignedDequeue_bits_data_hi_lo_24};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_25 = {_alignedDequeue_bits_data_T_1156[17], _alignedDequeue_bits_data_T_1026[17]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_25 = {_alignedDequeue_bits_data_T_1416[17], _alignedDequeue_bits_data_T_1286[17]};
  wire [3:0]    alignedDequeue_bits_data_lo_25 = {alignedDequeue_bits_data_lo_hi_25, alignedDequeue_bits_data_lo_lo_25};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_25 = {_alignedDequeue_bits_data_T_1676[17], _alignedDequeue_bits_data_T_1546[17]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_25 = {_alignedDequeue_bits_data_T_1936[17], _alignedDequeue_bits_data_T_1806[17]};
  wire [3:0]    alignedDequeue_bits_data_hi_25 = {alignedDequeue_bits_data_hi_hi_25, alignedDequeue_bits_data_hi_lo_25};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_26 = {_alignedDequeue_bits_data_T_1156[18], _alignedDequeue_bits_data_T_1026[18]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_26 = {_alignedDequeue_bits_data_T_1416[18], _alignedDequeue_bits_data_T_1286[18]};
  wire [3:0]    alignedDequeue_bits_data_lo_26 = {alignedDequeue_bits_data_lo_hi_26, alignedDequeue_bits_data_lo_lo_26};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_26 = {_alignedDequeue_bits_data_T_1676[18], _alignedDequeue_bits_data_T_1546[18]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_26 = {_alignedDequeue_bits_data_T_1936[18], _alignedDequeue_bits_data_T_1806[18]};
  wire [3:0]    alignedDequeue_bits_data_hi_26 = {alignedDequeue_bits_data_hi_hi_26, alignedDequeue_bits_data_hi_lo_26};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_27 = {_alignedDequeue_bits_data_T_1156[19], _alignedDequeue_bits_data_T_1026[19]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_27 = {_alignedDequeue_bits_data_T_1416[19], _alignedDequeue_bits_data_T_1286[19]};
  wire [3:0]    alignedDequeue_bits_data_lo_27 = {alignedDequeue_bits_data_lo_hi_27, alignedDequeue_bits_data_lo_lo_27};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_27 = {_alignedDequeue_bits_data_T_1676[19], _alignedDequeue_bits_data_T_1546[19]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_27 = {_alignedDequeue_bits_data_T_1936[19], _alignedDequeue_bits_data_T_1806[19]};
  wire [3:0]    alignedDequeue_bits_data_hi_27 = {alignedDequeue_bits_data_hi_hi_27, alignedDequeue_bits_data_hi_lo_27};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_28 = {_alignedDequeue_bits_data_T_1156[20], _alignedDequeue_bits_data_T_1026[20]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_28 = {_alignedDequeue_bits_data_T_1416[20], _alignedDequeue_bits_data_T_1286[20]};
  wire [3:0]    alignedDequeue_bits_data_lo_28 = {alignedDequeue_bits_data_lo_hi_28, alignedDequeue_bits_data_lo_lo_28};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_28 = {_alignedDequeue_bits_data_T_1676[20], _alignedDequeue_bits_data_T_1546[20]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_28 = {_alignedDequeue_bits_data_T_1936[20], _alignedDequeue_bits_data_T_1806[20]};
  wire [3:0]    alignedDequeue_bits_data_hi_28 = {alignedDequeue_bits_data_hi_hi_28, alignedDequeue_bits_data_hi_lo_28};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_29 = {_alignedDequeue_bits_data_T_1156[21], _alignedDequeue_bits_data_T_1026[21]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_29 = {_alignedDequeue_bits_data_T_1416[21], _alignedDequeue_bits_data_T_1286[21]};
  wire [3:0]    alignedDequeue_bits_data_lo_29 = {alignedDequeue_bits_data_lo_hi_29, alignedDequeue_bits_data_lo_lo_29};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_29 = {_alignedDequeue_bits_data_T_1676[21], _alignedDequeue_bits_data_T_1546[21]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_29 = {_alignedDequeue_bits_data_T_1936[21], _alignedDequeue_bits_data_T_1806[21]};
  wire [3:0]    alignedDequeue_bits_data_hi_29 = {alignedDequeue_bits_data_hi_hi_29, alignedDequeue_bits_data_hi_lo_29};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_30 = {_alignedDequeue_bits_data_T_1156[22], _alignedDequeue_bits_data_T_1026[22]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_30 = {_alignedDequeue_bits_data_T_1416[22], _alignedDequeue_bits_data_T_1286[22]};
  wire [3:0]    alignedDequeue_bits_data_lo_30 = {alignedDequeue_bits_data_lo_hi_30, alignedDequeue_bits_data_lo_lo_30};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_30 = {_alignedDequeue_bits_data_T_1676[22], _alignedDequeue_bits_data_T_1546[22]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_30 = {_alignedDequeue_bits_data_T_1936[22], _alignedDequeue_bits_data_T_1806[22]};
  wire [3:0]    alignedDequeue_bits_data_hi_30 = {alignedDequeue_bits_data_hi_hi_30, alignedDequeue_bits_data_hi_lo_30};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_31 = {_alignedDequeue_bits_data_T_1156[23], _alignedDequeue_bits_data_T_1026[23]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_31 = {_alignedDequeue_bits_data_T_1416[23], _alignedDequeue_bits_data_T_1286[23]};
  wire [3:0]    alignedDequeue_bits_data_lo_31 = {alignedDequeue_bits_data_lo_hi_31, alignedDequeue_bits_data_lo_lo_31};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_31 = {_alignedDequeue_bits_data_T_1676[23], _alignedDequeue_bits_data_T_1546[23]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_31 = {_alignedDequeue_bits_data_T_1936[23], _alignedDequeue_bits_data_T_1806[23]};
  wire [3:0]    alignedDequeue_bits_data_hi_31 = {alignedDequeue_bits_data_hi_hi_31, alignedDequeue_bits_data_hi_lo_31};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_32 = {_alignedDequeue_bits_data_T_1156[24], _alignedDequeue_bits_data_T_1026[24]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_32 = {_alignedDequeue_bits_data_T_1416[24], _alignedDequeue_bits_data_T_1286[24]};
  wire [3:0]    alignedDequeue_bits_data_lo_32 = {alignedDequeue_bits_data_lo_hi_32, alignedDequeue_bits_data_lo_lo_32};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_32 = {_alignedDequeue_bits_data_T_1676[24], _alignedDequeue_bits_data_T_1546[24]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_32 = {_alignedDequeue_bits_data_T_1936[24], _alignedDequeue_bits_data_T_1806[24]};
  wire [3:0]    alignedDequeue_bits_data_hi_32 = {alignedDequeue_bits_data_hi_hi_32, alignedDequeue_bits_data_hi_lo_32};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_33 = {_alignedDequeue_bits_data_T_1156[25], _alignedDequeue_bits_data_T_1026[25]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_33 = {_alignedDequeue_bits_data_T_1416[25], _alignedDequeue_bits_data_T_1286[25]};
  wire [3:0]    alignedDequeue_bits_data_lo_33 = {alignedDequeue_bits_data_lo_hi_33, alignedDequeue_bits_data_lo_lo_33};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_33 = {_alignedDequeue_bits_data_T_1676[25], _alignedDequeue_bits_data_T_1546[25]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_33 = {_alignedDequeue_bits_data_T_1936[25], _alignedDequeue_bits_data_T_1806[25]};
  wire [3:0]    alignedDequeue_bits_data_hi_33 = {alignedDequeue_bits_data_hi_hi_33, alignedDequeue_bits_data_hi_lo_33};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_34 = {_alignedDequeue_bits_data_T_1156[26], _alignedDequeue_bits_data_T_1026[26]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_34 = {_alignedDequeue_bits_data_T_1416[26], _alignedDequeue_bits_data_T_1286[26]};
  wire [3:0]    alignedDequeue_bits_data_lo_34 = {alignedDequeue_bits_data_lo_hi_34, alignedDequeue_bits_data_lo_lo_34};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_34 = {_alignedDequeue_bits_data_T_1676[26], _alignedDequeue_bits_data_T_1546[26]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_34 = {_alignedDequeue_bits_data_T_1936[26], _alignedDequeue_bits_data_T_1806[26]};
  wire [3:0]    alignedDequeue_bits_data_hi_34 = {alignedDequeue_bits_data_hi_hi_34, alignedDequeue_bits_data_hi_lo_34};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_35 = {_alignedDequeue_bits_data_T_1156[27], _alignedDequeue_bits_data_T_1026[27]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_35 = {_alignedDequeue_bits_data_T_1416[27], _alignedDequeue_bits_data_T_1286[27]};
  wire [3:0]    alignedDequeue_bits_data_lo_35 = {alignedDequeue_bits_data_lo_hi_35, alignedDequeue_bits_data_lo_lo_35};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_35 = {_alignedDequeue_bits_data_T_1676[27], _alignedDequeue_bits_data_T_1546[27]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_35 = {_alignedDequeue_bits_data_T_1936[27], _alignedDequeue_bits_data_T_1806[27]};
  wire [3:0]    alignedDequeue_bits_data_hi_35 = {alignedDequeue_bits_data_hi_hi_35, alignedDequeue_bits_data_hi_lo_35};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_36 = {_alignedDequeue_bits_data_T_1156[28], _alignedDequeue_bits_data_T_1026[28]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_36 = {_alignedDequeue_bits_data_T_1416[28], _alignedDequeue_bits_data_T_1286[28]};
  wire [3:0]    alignedDequeue_bits_data_lo_36 = {alignedDequeue_bits_data_lo_hi_36, alignedDequeue_bits_data_lo_lo_36};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_36 = {_alignedDequeue_bits_data_T_1676[28], _alignedDequeue_bits_data_T_1546[28]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_36 = {_alignedDequeue_bits_data_T_1936[28], _alignedDequeue_bits_data_T_1806[28]};
  wire [3:0]    alignedDequeue_bits_data_hi_36 = {alignedDequeue_bits_data_hi_hi_36, alignedDequeue_bits_data_hi_lo_36};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_37 = {_alignedDequeue_bits_data_T_1156[29], _alignedDequeue_bits_data_T_1026[29]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_37 = {_alignedDequeue_bits_data_T_1416[29], _alignedDequeue_bits_data_T_1286[29]};
  wire [3:0]    alignedDequeue_bits_data_lo_37 = {alignedDequeue_bits_data_lo_hi_37, alignedDequeue_bits_data_lo_lo_37};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_37 = {_alignedDequeue_bits_data_T_1676[29], _alignedDequeue_bits_data_T_1546[29]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_37 = {_alignedDequeue_bits_data_T_1936[29], _alignedDequeue_bits_data_T_1806[29]};
  wire [3:0]    alignedDequeue_bits_data_hi_37 = {alignedDequeue_bits_data_hi_hi_37, alignedDequeue_bits_data_hi_lo_37};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_38 = {_alignedDequeue_bits_data_T_1156[30], _alignedDequeue_bits_data_T_1026[30]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_38 = {_alignedDequeue_bits_data_T_1416[30], _alignedDequeue_bits_data_T_1286[30]};
  wire [3:0]    alignedDequeue_bits_data_lo_38 = {alignedDequeue_bits_data_lo_hi_38, alignedDequeue_bits_data_lo_lo_38};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_38 = {_alignedDequeue_bits_data_T_1676[30], _alignedDequeue_bits_data_T_1546[30]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_38 = {_alignedDequeue_bits_data_T_1936[30], _alignedDequeue_bits_data_T_1806[30]};
  wire [3:0]    alignedDequeue_bits_data_hi_38 = {alignedDequeue_bits_data_hi_hi_38, alignedDequeue_bits_data_hi_lo_38};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_39 = {_alignedDequeue_bits_data_T_1156[31], _alignedDequeue_bits_data_T_1026[31]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_39 = {_alignedDequeue_bits_data_T_1416[31], _alignedDequeue_bits_data_T_1286[31]};
  wire [3:0]    alignedDequeue_bits_data_lo_39 = {alignedDequeue_bits_data_lo_hi_39, alignedDequeue_bits_data_lo_lo_39};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_39 = {_alignedDequeue_bits_data_T_1676[31], _alignedDequeue_bits_data_T_1546[31]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_39 = {_alignedDequeue_bits_data_T_1936[31], _alignedDequeue_bits_data_T_1806[31]};
  wire [3:0]    alignedDequeue_bits_data_hi_39 = {alignedDequeue_bits_data_hi_hi_39, alignedDequeue_bits_data_hi_lo_39};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_40 = {_alignedDequeue_bits_data_T_1156[32], _alignedDequeue_bits_data_T_1026[32]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_40 = {_alignedDequeue_bits_data_T_1416[32], _alignedDequeue_bits_data_T_1286[32]};
  wire [3:0]    alignedDequeue_bits_data_lo_40 = {alignedDequeue_bits_data_lo_hi_40, alignedDequeue_bits_data_lo_lo_40};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_40 = {_alignedDequeue_bits_data_T_1676[32], _alignedDequeue_bits_data_T_1546[32]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_40 = {_alignedDequeue_bits_data_T_1936[32], _alignedDequeue_bits_data_T_1806[32]};
  wire [3:0]    alignedDequeue_bits_data_hi_40 = {alignedDequeue_bits_data_hi_hi_40, alignedDequeue_bits_data_hi_lo_40};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_41 = {_alignedDequeue_bits_data_T_1156[33], _alignedDequeue_bits_data_T_1026[33]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_41 = {_alignedDequeue_bits_data_T_1416[33], _alignedDequeue_bits_data_T_1286[33]};
  wire [3:0]    alignedDequeue_bits_data_lo_41 = {alignedDequeue_bits_data_lo_hi_41, alignedDequeue_bits_data_lo_lo_41};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_41 = {_alignedDequeue_bits_data_T_1676[33], _alignedDequeue_bits_data_T_1546[33]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_41 = {_alignedDequeue_bits_data_T_1936[33], _alignedDequeue_bits_data_T_1806[33]};
  wire [3:0]    alignedDequeue_bits_data_hi_41 = {alignedDequeue_bits_data_hi_hi_41, alignedDequeue_bits_data_hi_lo_41};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_42 = {_alignedDequeue_bits_data_T_1156[34], _alignedDequeue_bits_data_T_1026[34]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_42 = {_alignedDequeue_bits_data_T_1416[34], _alignedDequeue_bits_data_T_1286[34]};
  wire [3:0]    alignedDequeue_bits_data_lo_42 = {alignedDequeue_bits_data_lo_hi_42, alignedDequeue_bits_data_lo_lo_42};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_42 = {_alignedDequeue_bits_data_T_1676[34], _alignedDequeue_bits_data_T_1546[34]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_42 = {_alignedDequeue_bits_data_T_1936[34], _alignedDequeue_bits_data_T_1806[34]};
  wire [3:0]    alignedDequeue_bits_data_hi_42 = {alignedDequeue_bits_data_hi_hi_42, alignedDequeue_bits_data_hi_lo_42};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_43 = {_alignedDequeue_bits_data_T_1156[35], _alignedDequeue_bits_data_T_1026[35]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_43 = {_alignedDequeue_bits_data_T_1416[35], _alignedDequeue_bits_data_T_1286[35]};
  wire [3:0]    alignedDequeue_bits_data_lo_43 = {alignedDequeue_bits_data_lo_hi_43, alignedDequeue_bits_data_lo_lo_43};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_43 = {_alignedDequeue_bits_data_T_1676[35], _alignedDequeue_bits_data_T_1546[35]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_43 = {_alignedDequeue_bits_data_T_1936[35], _alignedDequeue_bits_data_T_1806[35]};
  wire [3:0]    alignedDequeue_bits_data_hi_43 = {alignedDequeue_bits_data_hi_hi_43, alignedDequeue_bits_data_hi_lo_43};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_44 = {_alignedDequeue_bits_data_T_1156[36], _alignedDequeue_bits_data_T_1026[36]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_44 = {_alignedDequeue_bits_data_T_1416[36], _alignedDequeue_bits_data_T_1286[36]};
  wire [3:0]    alignedDequeue_bits_data_lo_44 = {alignedDequeue_bits_data_lo_hi_44, alignedDequeue_bits_data_lo_lo_44};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_44 = {_alignedDequeue_bits_data_T_1676[36], _alignedDequeue_bits_data_T_1546[36]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_44 = {_alignedDequeue_bits_data_T_1936[36], _alignedDequeue_bits_data_T_1806[36]};
  wire [3:0]    alignedDequeue_bits_data_hi_44 = {alignedDequeue_bits_data_hi_hi_44, alignedDequeue_bits_data_hi_lo_44};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_45 = {_alignedDequeue_bits_data_T_1156[37], _alignedDequeue_bits_data_T_1026[37]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_45 = {_alignedDequeue_bits_data_T_1416[37], _alignedDequeue_bits_data_T_1286[37]};
  wire [3:0]    alignedDequeue_bits_data_lo_45 = {alignedDequeue_bits_data_lo_hi_45, alignedDequeue_bits_data_lo_lo_45};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_45 = {_alignedDequeue_bits_data_T_1676[37], _alignedDequeue_bits_data_T_1546[37]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_45 = {_alignedDequeue_bits_data_T_1936[37], _alignedDequeue_bits_data_T_1806[37]};
  wire [3:0]    alignedDequeue_bits_data_hi_45 = {alignedDequeue_bits_data_hi_hi_45, alignedDequeue_bits_data_hi_lo_45};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_46 = {_alignedDequeue_bits_data_T_1156[38], _alignedDequeue_bits_data_T_1026[38]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_46 = {_alignedDequeue_bits_data_T_1416[38], _alignedDequeue_bits_data_T_1286[38]};
  wire [3:0]    alignedDequeue_bits_data_lo_46 = {alignedDequeue_bits_data_lo_hi_46, alignedDequeue_bits_data_lo_lo_46};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_46 = {_alignedDequeue_bits_data_T_1676[38], _alignedDequeue_bits_data_T_1546[38]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_46 = {_alignedDequeue_bits_data_T_1936[38], _alignedDequeue_bits_data_T_1806[38]};
  wire [3:0]    alignedDequeue_bits_data_hi_46 = {alignedDequeue_bits_data_hi_hi_46, alignedDequeue_bits_data_hi_lo_46};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_47 = {_alignedDequeue_bits_data_T_1156[39], _alignedDequeue_bits_data_T_1026[39]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_47 = {_alignedDequeue_bits_data_T_1416[39], _alignedDequeue_bits_data_T_1286[39]};
  wire [3:0]    alignedDequeue_bits_data_lo_47 = {alignedDequeue_bits_data_lo_hi_47, alignedDequeue_bits_data_lo_lo_47};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_47 = {_alignedDequeue_bits_data_T_1676[39], _alignedDequeue_bits_data_T_1546[39]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_47 = {_alignedDequeue_bits_data_T_1936[39], _alignedDequeue_bits_data_T_1806[39]};
  wire [3:0]    alignedDequeue_bits_data_hi_47 = {alignedDequeue_bits_data_hi_hi_47, alignedDequeue_bits_data_hi_lo_47};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_48 = {_alignedDequeue_bits_data_T_1156[40], _alignedDequeue_bits_data_T_1026[40]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_48 = {_alignedDequeue_bits_data_T_1416[40], _alignedDequeue_bits_data_T_1286[40]};
  wire [3:0]    alignedDequeue_bits_data_lo_48 = {alignedDequeue_bits_data_lo_hi_48, alignedDequeue_bits_data_lo_lo_48};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_48 = {_alignedDequeue_bits_data_T_1676[40], _alignedDequeue_bits_data_T_1546[40]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_48 = {_alignedDequeue_bits_data_T_1936[40], _alignedDequeue_bits_data_T_1806[40]};
  wire [3:0]    alignedDequeue_bits_data_hi_48 = {alignedDequeue_bits_data_hi_hi_48, alignedDequeue_bits_data_hi_lo_48};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_49 = {_alignedDequeue_bits_data_T_1156[41], _alignedDequeue_bits_data_T_1026[41]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_49 = {_alignedDequeue_bits_data_T_1416[41], _alignedDequeue_bits_data_T_1286[41]};
  wire [3:0]    alignedDequeue_bits_data_lo_49 = {alignedDequeue_bits_data_lo_hi_49, alignedDequeue_bits_data_lo_lo_49};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_49 = {_alignedDequeue_bits_data_T_1676[41], _alignedDequeue_bits_data_T_1546[41]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_49 = {_alignedDequeue_bits_data_T_1936[41], _alignedDequeue_bits_data_T_1806[41]};
  wire [3:0]    alignedDequeue_bits_data_hi_49 = {alignedDequeue_bits_data_hi_hi_49, alignedDequeue_bits_data_hi_lo_49};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_50 = {_alignedDequeue_bits_data_T_1156[42], _alignedDequeue_bits_data_T_1026[42]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_50 = {_alignedDequeue_bits_data_T_1416[42], _alignedDequeue_bits_data_T_1286[42]};
  wire [3:0]    alignedDequeue_bits_data_lo_50 = {alignedDequeue_bits_data_lo_hi_50, alignedDequeue_bits_data_lo_lo_50};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_50 = {_alignedDequeue_bits_data_T_1676[42], _alignedDequeue_bits_data_T_1546[42]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_50 = {_alignedDequeue_bits_data_T_1936[42], _alignedDequeue_bits_data_T_1806[42]};
  wire [3:0]    alignedDequeue_bits_data_hi_50 = {alignedDequeue_bits_data_hi_hi_50, alignedDequeue_bits_data_hi_lo_50};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_51 = {_alignedDequeue_bits_data_T_1156[43], _alignedDequeue_bits_data_T_1026[43]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_51 = {_alignedDequeue_bits_data_T_1416[43], _alignedDequeue_bits_data_T_1286[43]};
  wire [3:0]    alignedDequeue_bits_data_lo_51 = {alignedDequeue_bits_data_lo_hi_51, alignedDequeue_bits_data_lo_lo_51};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_51 = {_alignedDequeue_bits_data_T_1676[43], _alignedDequeue_bits_data_T_1546[43]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_51 = {_alignedDequeue_bits_data_T_1936[43], _alignedDequeue_bits_data_T_1806[43]};
  wire [3:0]    alignedDequeue_bits_data_hi_51 = {alignedDequeue_bits_data_hi_hi_51, alignedDequeue_bits_data_hi_lo_51};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_52 = {_alignedDequeue_bits_data_T_1156[44], _alignedDequeue_bits_data_T_1026[44]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_52 = {_alignedDequeue_bits_data_T_1416[44], _alignedDequeue_bits_data_T_1286[44]};
  wire [3:0]    alignedDequeue_bits_data_lo_52 = {alignedDequeue_bits_data_lo_hi_52, alignedDequeue_bits_data_lo_lo_52};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_52 = {_alignedDequeue_bits_data_T_1676[44], _alignedDequeue_bits_data_T_1546[44]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_52 = {_alignedDequeue_bits_data_T_1936[44], _alignedDequeue_bits_data_T_1806[44]};
  wire [3:0]    alignedDequeue_bits_data_hi_52 = {alignedDequeue_bits_data_hi_hi_52, alignedDequeue_bits_data_hi_lo_52};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_53 = {_alignedDequeue_bits_data_T_1156[45], _alignedDequeue_bits_data_T_1026[45]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_53 = {_alignedDequeue_bits_data_T_1416[45], _alignedDequeue_bits_data_T_1286[45]};
  wire [3:0]    alignedDequeue_bits_data_lo_53 = {alignedDequeue_bits_data_lo_hi_53, alignedDequeue_bits_data_lo_lo_53};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_53 = {_alignedDequeue_bits_data_T_1676[45], _alignedDequeue_bits_data_T_1546[45]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_53 = {_alignedDequeue_bits_data_T_1936[45], _alignedDequeue_bits_data_T_1806[45]};
  wire [3:0]    alignedDequeue_bits_data_hi_53 = {alignedDequeue_bits_data_hi_hi_53, alignedDequeue_bits_data_hi_lo_53};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_54 = {_alignedDequeue_bits_data_T_1156[46], _alignedDequeue_bits_data_T_1026[46]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_54 = {_alignedDequeue_bits_data_T_1416[46], _alignedDequeue_bits_data_T_1286[46]};
  wire [3:0]    alignedDequeue_bits_data_lo_54 = {alignedDequeue_bits_data_lo_hi_54, alignedDequeue_bits_data_lo_lo_54};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_54 = {_alignedDequeue_bits_data_T_1676[46], _alignedDequeue_bits_data_T_1546[46]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_54 = {_alignedDequeue_bits_data_T_1936[46], _alignedDequeue_bits_data_T_1806[46]};
  wire [3:0]    alignedDequeue_bits_data_hi_54 = {alignedDequeue_bits_data_hi_hi_54, alignedDequeue_bits_data_hi_lo_54};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_55 = {_alignedDequeue_bits_data_T_1156[47], _alignedDequeue_bits_data_T_1026[47]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_55 = {_alignedDequeue_bits_data_T_1416[47], _alignedDequeue_bits_data_T_1286[47]};
  wire [3:0]    alignedDequeue_bits_data_lo_55 = {alignedDequeue_bits_data_lo_hi_55, alignedDequeue_bits_data_lo_lo_55};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_55 = {_alignedDequeue_bits_data_T_1676[47], _alignedDequeue_bits_data_T_1546[47]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_55 = {_alignedDequeue_bits_data_T_1936[47], _alignedDequeue_bits_data_T_1806[47]};
  wire [3:0]    alignedDequeue_bits_data_hi_55 = {alignedDequeue_bits_data_hi_hi_55, alignedDequeue_bits_data_hi_lo_55};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_56 = {_alignedDequeue_bits_data_T_1156[48], _alignedDequeue_bits_data_T_1026[48]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_56 = {_alignedDequeue_bits_data_T_1416[48], _alignedDequeue_bits_data_T_1286[48]};
  wire [3:0]    alignedDequeue_bits_data_lo_56 = {alignedDequeue_bits_data_lo_hi_56, alignedDequeue_bits_data_lo_lo_56};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_56 = {_alignedDequeue_bits_data_T_1676[48], _alignedDequeue_bits_data_T_1546[48]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_56 = {_alignedDequeue_bits_data_T_1936[48], _alignedDequeue_bits_data_T_1806[48]};
  wire [3:0]    alignedDequeue_bits_data_hi_56 = {alignedDequeue_bits_data_hi_hi_56, alignedDequeue_bits_data_hi_lo_56};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_57 = {_alignedDequeue_bits_data_T_1156[49], _alignedDequeue_bits_data_T_1026[49]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_57 = {_alignedDequeue_bits_data_T_1416[49], _alignedDequeue_bits_data_T_1286[49]};
  wire [3:0]    alignedDequeue_bits_data_lo_57 = {alignedDequeue_bits_data_lo_hi_57, alignedDequeue_bits_data_lo_lo_57};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_57 = {_alignedDequeue_bits_data_T_1676[49], _alignedDequeue_bits_data_T_1546[49]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_57 = {_alignedDequeue_bits_data_T_1936[49], _alignedDequeue_bits_data_T_1806[49]};
  wire [3:0]    alignedDequeue_bits_data_hi_57 = {alignedDequeue_bits_data_hi_hi_57, alignedDequeue_bits_data_hi_lo_57};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_58 = {_alignedDequeue_bits_data_T_1156[50], _alignedDequeue_bits_data_T_1026[50]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_58 = {_alignedDequeue_bits_data_T_1416[50], _alignedDequeue_bits_data_T_1286[50]};
  wire [3:0]    alignedDequeue_bits_data_lo_58 = {alignedDequeue_bits_data_lo_hi_58, alignedDequeue_bits_data_lo_lo_58};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_58 = {_alignedDequeue_bits_data_T_1676[50], _alignedDequeue_bits_data_T_1546[50]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_58 = {_alignedDequeue_bits_data_T_1936[50], _alignedDequeue_bits_data_T_1806[50]};
  wire [3:0]    alignedDequeue_bits_data_hi_58 = {alignedDequeue_bits_data_hi_hi_58, alignedDequeue_bits_data_hi_lo_58};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_59 = {_alignedDequeue_bits_data_T_1156[51], _alignedDequeue_bits_data_T_1026[51]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_59 = {_alignedDequeue_bits_data_T_1416[51], _alignedDequeue_bits_data_T_1286[51]};
  wire [3:0]    alignedDequeue_bits_data_lo_59 = {alignedDequeue_bits_data_lo_hi_59, alignedDequeue_bits_data_lo_lo_59};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_59 = {_alignedDequeue_bits_data_T_1676[51], _alignedDequeue_bits_data_T_1546[51]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_59 = {_alignedDequeue_bits_data_T_1936[51], _alignedDequeue_bits_data_T_1806[51]};
  wire [3:0]    alignedDequeue_bits_data_hi_59 = {alignedDequeue_bits_data_hi_hi_59, alignedDequeue_bits_data_hi_lo_59};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_60 = {_alignedDequeue_bits_data_T_1156[52], _alignedDequeue_bits_data_T_1026[52]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_60 = {_alignedDequeue_bits_data_T_1416[52], _alignedDequeue_bits_data_T_1286[52]};
  wire [3:0]    alignedDequeue_bits_data_lo_60 = {alignedDequeue_bits_data_lo_hi_60, alignedDequeue_bits_data_lo_lo_60};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_60 = {_alignedDequeue_bits_data_T_1676[52], _alignedDequeue_bits_data_T_1546[52]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_60 = {_alignedDequeue_bits_data_T_1936[52], _alignedDequeue_bits_data_T_1806[52]};
  wire [3:0]    alignedDequeue_bits_data_hi_60 = {alignedDequeue_bits_data_hi_hi_60, alignedDequeue_bits_data_hi_lo_60};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_61 = {_alignedDequeue_bits_data_T_1156[53], _alignedDequeue_bits_data_T_1026[53]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_61 = {_alignedDequeue_bits_data_T_1416[53], _alignedDequeue_bits_data_T_1286[53]};
  wire [3:0]    alignedDequeue_bits_data_lo_61 = {alignedDequeue_bits_data_lo_hi_61, alignedDequeue_bits_data_lo_lo_61};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_61 = {_alignedDequeue_bits_data_T_1676[53], _alignedDequeue_bits_data_T_1546[53]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_61 = {_alignedDequeue_bits_data_T_1936[53], _alignedDequeue_bits_data_T_1806[53]};
  wire [3:0]    alignedDequeue_bits_data_hi_61 = {alignedDequeue_bits_data_hi_hi_61, alignedDequeue_bits_data_hi_lo_61};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_62 = {_alignedDequeue_bits_data_T_1156[54], _alignedDequeue_bits_data_T_1026[54]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_62 = {_alignedDequeue_bits_data_T_1416[54], _alignedDequeue_bits_data_T_1286[54]};
  wire [3:0]    alignedDequeue_bits_data_lo_62 = {alignedDequeue_bits_data_lo_hi_62, alignedDequeue_bits_data_lo_lo_62};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_62 = {_alignedDequeue_bits_data_T_1676[54], _alignedDequeue_bits_data_T_1546[54]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_62 = {_alignedDequeue_bits_data_T_1936[54], _alignedDequeue_bits_data_T_1806[54]};
  wire [3:0]    alignedDequeue_bits_data_hi_62 = {alignedDequeue_bits_data_hi_hi_62, alignedDequeue_bits_data_hi_lo_62};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_63 = {_alignedDequeue_bits_data_T_1156[55], _alignedDequeue_bits_data_T_1026[55]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_63 = {_alignedDequeue_bits_data_T_1416[55], _alignedDequeue_bits_data_T_1286[55]};
  wire [3:0]    alignedDequeue_bits_data_lo_63 = {alignedDequeue_bits_data_lo_hi_63, alignedDequeue_bits_data_lo_lo_63};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_63 = {_alignedDequeue_bits_data_T_1676[55], _alignedDequeue_bits_data_T_1546[55]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_63 = {_alignedDequeue_bits_data_T_1936[55], _alignedDequeue_bits_data_T_1806[55]};
  wire [3:0]    alignedDequeue_bits_data_hi_63 = {alignedDequeue_bits_data_hi_hi_63, alignedDequeue_bits_data_hi_lo_63};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_64 = {_alignedDequeue_bits_data_T_1156[56], _alignedDequeue_bits_data_T_1026[56]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_64 = {_alignedDequeue_bits_data_T_1416[56], _alignedDequeue_bits_data_T_1286[56]};
  wire [3:0]    alignedDequeue_bits_data_lo_64 = {alignedDequeue_bits_data_lo_hi_64, alignedDequeue_bits_data_lo_lo_64};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_64 = {_alignedDequeue_bits_data_T_1676[56], _alignedDequeue_bits_data_T_1546[56]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_64 = {_alignedDequeue_bits_data_T_1936[56], _alignedDequeue_bits_data_T_1806[56]};
  wire [3:0]    alignedDequeue_bits_data_hi_64 = {alignedDequeue_bits_data_hi_hi_64, alignedDequeue_bits_data_hi_lo_64};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_65 = {_alignedDequeue_bits_data_T_1156[57], _alignedDequeue_bits_data_T_1026[57]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_65 = {_alignedDequeue_bits_data_T_1416[57], _alignedDequeue_bits_data_T_1286[57]};
  wire [3:0]    alignedDequeue_bits_data_lo_65 = {alignedDequeue_bits_data_lo_hi_65, alignedDequeue_bits_data_lo_lo_65};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_65 = {_alignedDequeue_bits_data_T_1676[57], _alignedDequeue_bits_data_T_1546[57]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_65 = {_alignedDequeue_bits_data_T_1936[57], _alignedDequeue_bits_data_T_1806[57]};
  wire [3:0]    alignedDequeue_bits_data_hi_65 = {alignedDequeue_bits_data_hi_hi_65, alignedDequeue_bits_data_hi_lo_65};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_66 = {_alignedDequeue_bits_data_T_1156[58], _alignedDequeue_bits_data_T_1026[58]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_66 = {_alignedDequeue_bits_data_T_1416[58], _alignedDequeue_bits_data_T_1286[58]};
  wire [3:0]    alignedDequeue_bits_data_lo_66 = {alignedDequeue_bits_data_lo_hi_66, alignedDequeue_bits_data_lo_lo_66};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_66 = {_alignedDequeue_bits_data_T_1676[58], _alignedDequeue_bits_data_T_1546[58]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_66 = {_alignedDequeue_bits_data_T_1936[58], _alignedDequeue_bits_data_T_1806[58]};
  wire [3:0]    alignedDequeue_bits_data_hi_66 = {alignedDequeue_bits_data_hi_hi_66, alignedDequeue_bits_data_hi_lo_66};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_67 = {_alignedDequeue_bits_data_T_1156[59], _alignedDequeue_bits_data_T_1026[59]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_67 = {_alignedDequeue_bits_data_T_1416[59], _alignedDequeue_bits_data_T_1286[59]};
  wire [3:0]    alignedDequeue_bits_data_lo_67 = {alignedDequeue_bits_data_lo_hi_67, alignedDequeue_bits_data_lo_lo_67};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_67 = {_alignedDequeue_bits_data_T_1676[59], _alignedDequeue_bits_data_T_1546[59]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_67 = {_alignedDequeue_bits_data_T_1936[59], _alignedDequeue_bits_data_T_1806[59]};
  wire [3:0]    alignedDequeue_bits_data_hi_67 = {alignedDequeue_bits_data_hi_hi_67, alignedDequeue_bits_data_hi_lo_67};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_68 = {_alignedDequeue_bits_data_T_1156[60], _alignedDequeue_bits_data_T_1026[60]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_68 = {_alignedDequeue_bits_data_T_1416[60], _alignedDequeue_bits_data_T_1286[60]};
  wire [3:0]    alignedDequeue_bits_data_lo_68 = {alignedDequeue_bits_data_lo_hi_68, alignedDequeue_bits_data_lo_lo_68};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_68 = {_alignedDequeue_bits_data_T_1676[60], _alignedDequeue_bits_data_T_1546[60]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_68 = {_alignedDequeue_bits_data_T_1936[60], _alignedDequeue_bits_data_T_1806[60]};
  wire [3:0]    alignedDequeue_bits_data_hi_68 = {alignedDequeue_bits_data_hi_hi_68, alignedDequeue_bits_data_hi_lo_68};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_69 = {_alignedDequeue_bits_data_T_1156[61], _alignedDequeue_bits_data_T_1026[61]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_69 = {_alignedDequeue_bits_data_T_1416[61], _alignedDequeue_bits_data_T_1286[61]};
  wire [3:0]    alignedDequeue_bits_data_lo_69 = {alignedDequeue_bits_data_lo_hi_69, alignedDequeue_bits_data_lo_lo_69};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_69 = {_alignedDequeue_bits_data_T_1676[61], _alignedDequeue_bits_data_T_1546[61]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_69 = {_alignedDequeue_bits_data_T_1936[61], _alignedDequeue_bits_data_T_1806[61]};
  wire [3:0]    alignedDequeue_bits_data_hi_69 = {alignedDequeue_bits_data_hi_hi_69, alignedDequeue_bits_data_hi_lo_69};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_70 = {_alignedDequeue_bits_data_T_1156[62], _alignedDequeue_bits_data_T_1026[62]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_70 = {_alignedDequeue_bits_data_T_1416[62], _alignedDequeue_bits_data_T_1286[62]};
  wire [3:0]    alignedDequeue_bits_data_lo_70 = {alignedDequeue_bits_data_lo_hi_70, alignedDequeue_bits_data_lo_lo_70};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_70 = {_alignedDequeue_bits_data_T_1676[62], _alignedDequeue_bits_data_T_1546[62]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_70 = {_alignedDequeue_bits_data_T_1936[62], _alignedDequeue_bits_data_T_1806[62]};
  wire [3:0]    alignedDequeue_bits_data_hi_70 = {alignedDequeue_bits_data_hi_hi_70, alignedDequeue_bits_data_hi_lo_70};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_71 = {_alignedDequeue_bits_data_T_1156[63], _alignedDequeue_bits_data_T_1026[63]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_71 = {_alignedDequeue_bits_data_T_1416[63], _alignedDequeue_bits_data_T_1286[63]};
  wire [3:0]    alignedDequeue_bits_data_lo_71 = {alignedDequeue_bits_data_lo_hi_71, alignedDequeue_bits_data_lo_lo_71};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_71 = {_alignedDequeue_bits_data_T_1676[63], _alignedDequeue_bits_data_T_1546[63]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_71 = {_alignedDequeue_bits_data_T_1936[63], _alignedDequeue_bits_data_T_1806[63]};
  wire [3:0]    alignedDequeue_bits_data_hi_71 = {alignedDequeue_bits_data_hi_hi_71, alignedDequeue_bits_data_hi_lo_71};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_72 = {_alignedDequeue_bits_data_T_1156[64], _alignedDequeue_bits_data_T_1026[64]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_72 = {_alignedDequeue_bits_data_T_1416[64], _alignedDequeue_bits_data_T_1286[64]};
  wire [3:0]    alignedDequeue_bits_data_lo_72 = {alignedDequeue_bits_data_lo_hi_72, alignedDequeue_bits_data_lo_lo_72};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_72 = {_alignedDequeue_bits_data_T_1676[64], _alignedDequeue_bits_data_T_1546[64]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_72 = {_alignedDequeue_bits_data_T_1936[64], _alignedDequeue_bits_data_T_1806[64]};
  wire [3:0]    alignedDequeue_bits_data_hi_72 = {alignedDequeue_bits_data_hi_hi_72, alignedDequeue_bits_data_hi_lo_72};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_73 = {_alignedDequeue_bits_data_T_1156[65], _alignedDequeue_bits_data_T_1026[65]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_73 = {_alignedDequeue_bits_data_T_1416[65], _alignedDequeue_bits_data_T_1286[65]};
  wire [3:0]    alignedDequeue_bits_data_lo_73 = {alignedDequeue_bits_data_lo_hi_73, alignedDequeue_bits_data_lo_lo_73};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_73 = {_alignedDequeue_bits_data_T_1676[65], _alignedDequeue_bits_data_T_1546[65]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_73 = {_alignedDequeue_bits_data_T_1936[65], _alignedDequeue_bits_data_T_1806[65]};
  wire [3:0]    alignedDequeue_bits_data_hi_73 = {alignedDequeue_bits_data_hi_hi_73, alignedDequeue_bits_data_hi_lo_73};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_74 = {_alignedDequeue_bits_data_T_1156[66], _alignedDequeue_bits_data_T_1026[66]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_74 = {_alignedDequeue_bits_data_T_1416[66], _alignedDequeue_bits_data_T_1286[66]};
  wire [3:0]    alignedDequeue_bits_data_lo_74 = {alignedDequeue_bits_data_lo_hi_74, alignedDequeue_bits_data_lo_lo_74};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_74 = {_alignedDequeue_bits_data_T_1676[66], _alignedDequeue_bits_data_T_1546[66]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_74 = {_alignedDequeue_bits_data_T_1936[66], _alignedDequeue_bits_data_T_1806[66]};
  wire [3:0]    alignedDequeue_bits_data_hi_74 = {alignedDequeue_bits_data_hi_hi_74, alignedDequeue_bits_data_hi_lo_74};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_75 = {_alignedDequeue_bits_data_T_1156[67], _alignedDequeue_bits_data_T_1026[67]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_75 = {_alignedDequeue_bits_data_T_1416[67], _alignedDequeue_bits_data_T_1286[67]};
  wire [3:0]    alignedDequeue_bits_data_lo_75 = {alignedDequeue_bits_data_lo_hi_75, alignedDequeue_bits_data_lo_lo_75};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_75 = {_alignedDequeue_bits_data_T_1676[67], _alignedDequeue_bits_data_T_1546[67]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_75 = {_alignedDequeue_bits_data_T_1936[67], _alignedDequeue_bits_data_T_1806[67]};
  wire [3:0]    alignedDequeue_bits_data_hi_75 = {alignedDequeue_bits_data_hi_hi_75, alignedDequeue_bits_data_hi_lo_75};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_76 = {_alignedDequeue_bits_data_T_1156[68], _alignedDequeue_bits_data_T_1026[68]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_76 = {_alignedDequeue_bits_data_T_1416[68], _alignedDequeue_bits_data_T_1286[68]};
  wire [3:0]    alignedDequeue_bits_data_lo_76 = {alignedDequeue_bits_data_lo_hi_76, alignedDequeue_bits_data_lo_lo_76};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_76 = {_alignedDequeue_bits_data_T_1676[68], _alignedDequeue_bits_data_T_1546[68]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_76 = {_alignedDequeue_bits_data_T_1936[68], _alignedDequeue_bits_data_T_1806[68]};
  wire [3:0]    alignedDequeue_bits_data_hi_76 = {alignedDequeue_bits_data_hi_hi_76, alignedDequeue_bits_data_hi_lo_76};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_77 = {_alignedDequeue_bits_data_T_1156[69], _alignedDequeue_bits_data_T_1026[69]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_77 = {_alignedDequeue_bits_data_T_1416[69], _alignedDequeue_bits_data_T_1286[69]};
  wire [3:0]    alignedDequeue_bits_data_lo_77 = {alignedDequeue_bits_data_lo_hi_77, alignedDequeue_bits_data_lo_lo_77};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_77 = {_alignedDequeue_bits_data_T_1676[69], _alignedDequeue_bits_data_T_1546[69]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_77 = {_alignedDequeue_bits_data_T_1936[69], _alignedDequeue_bits_data_T_1806[69]};
  wire [3:0]    alignedDequeue_bits_data_hi_77 = {alignedDequeue_bits_data_hi_hi_77, alignedDequeue_bits_data_hi_lo_77};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_78 = {_alignedDequeue_bits_data_T_1156[70], _alignedDequeue_bits_data_T_1026[70]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_78 = {_alignedDequeue_bits_data_T_1416[70], _alignedDequeue_bits_data_T_1286[70]};
  wire [3:0]    alignedDequeue_bits_data_lo_78 = {alignedDequeue_bits_data_lo_hi_78, alignedDequeue_bits_data_lo_lo_78};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_78 = {_alignedDequeue_bits_data_T_1676[70], _alignedDequeue_bits_data_T_1546[70]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_78 = {_alignedDequeue_bits_data_T_1936[70], _alignedDequeue_bits_data_T_1806[70]};
  wire [3:0]    alignedDequeue_bits_data_hi_78 = {alignedDequeue_bits_data_hi_hi_78, alignedDequeue_bits_data_hi_lo_78};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_79 = {_alignedDequeue_bits_data_T_1156[71], _alignedDequeue_bits_data_T_1026[71]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_79 = {_alignedDequeue_bits_data_T_1416[71], _alignedDequeue_bits_data_T_1286[71]};
  wire [3:0]    alignedDequeue_bits_data_lo_79 = {alignedDequeue_bits_data_lo_hi_79, alignedDequeue_bits_data_lo_lo_79};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_79 = {_alignedDequeue_bits_data_T_1676[71], _alignedDequeue_bits_data_T_1546[71]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_79 = {_alignedDequeue_bits_data_T_1936[71], _alignedDequeue_bits_data_T_1806[71]};
  wire [3:0]    alignedDequeue_bits_data_hi_79 = {alignedDequeue_bits_data_hi_hi_79, alignedDequeue_bits_data_hi_lo_79};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_80 = {_alignedDequeue_bits_data_T_1156[72], _alignedDequeue_bits_data_T_1026[72]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_80 = {_alignedDequeue_bits_data_T_1416[72], _alignedDequeue_bits_data_T_1286[72]};
  wire [3:0]    alignedDequeue_bits_data_lo_80 = {alignedDequeue_bits_data_lo_hi_80, alignedDequeue_bits_data_lo_lo_80};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_80 = {_alignedDequeue_bits_data_T_1676[72], _alignedDequeue_bits_data_T_1546[72]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_80 = {_alignedDequeue_bits_data_T_1936[72], _alignedDequeue_bits_data_T_1806[72]};
  wire [3:0]    alignedDequeue_bits_data_hi_80 = {alignedDequeue_bits_data_hi_hi_80, alignedDequeue_bits_data_hi_lo_80};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_81 = {_alignedDequeue_bits_data_T_1156[73], _alignedDequeue_bits_data_T_1026[73]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_81 = {_alignedDequeue_bits_data_T_1416[73], _alignedDequeue_bits_data_T_1286[73]};
  wire [3:0]    alignedDequeue_bits_data_lo_81 = {alignedDequeue_bits_data_lo_hi_81, alignedDequeue_bits_data_lo_lo_81};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_81 = {_alignedDequeue_bits_data_T_1676[73], _alignedDequeue_bits_data_T_1546[73]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_81 = {_alignedDequeue_bits_data_T_1936[73], _alignedDequeue_bits_data_T_1806[73]};
  wire [3:0]    alignedDequeue_bits_data_hi_81 = {alignedDequeue_bits_data_hi_hi_81, alignedDequeue_bits_data_hi_lo_81};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_82 = {_alignedDequeue_bits_data_T_1156[74], _alignedDequeue_bits_data_T_1026[74]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_82 = {_alignedDequeue_bits_data_T_1416[74], _alignedDequeue_bits_data_T_1286[74]};
  wire [3:0]    alignedDequeue_bits_data_lo_82 = {alignedDequeue_bits_data_lo_hi_82, alignedDequeue_bits_data_lo_lo_82};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_82 = {_alignedDequeue_bits_data_T_1676[74], _alignedDequeue_bits_data_T_1546[74]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_82 = {_alignedDequeue_bits_data_T_1936[74], _alignedDequeue_bits_data_T_1806[74]};
  wire [3:0]    alignedDequeue_bits_data_hi_82 = {alignedDequeue_bits_data_hi_hi_82, alignedDequeue_bits_data_hi_lo_82};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_83 = {_alignedDequeue_bits_data_T_1156[75], _alignedDequeue_bits_data_T_1026[75]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_83 = {_alignedDequeue_bits_data_T_1416[75], _alignedDequeue_bits_data_T_1286[75]};
  wire [3:0]    alignedDequeue_bits_data_lo_83 = {alignedDequeue_bits_data_lo_hi_83, alignedDequeue_bits_data_lo_lo_83};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_83 = {_alignedDequeue_bits_data_T_1676[75], _alignedDequeue_bits_data_T_1546[75]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_83 = {_alignedDequeue_bits_data_T_1936[75], _alignedDequeue_bits_data_T_1806[75]};
  wire [3:0]    alignedDequeue_bits_data_hi_83 = {alignedDequeue_bits_data_hi_hi_83, alignedDequeue_bits_data_hi_lo_83};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_84 = {_alignedDequeue_bits_data_T_1156[76], _alignedDequeue_bits_data_T_1026[76]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_84 = {_alignedDequeue_bits_data_T_1416[76], _alignedDequeue_bits_data_T_1286[76]};
  wire [3:0]    alignedDequeue_bits_data_lo_84 = {alignedDequeue_bits_data_lo_hi_84, alignedDequeue_bits_data_lo_lo_84};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_84 = {_alignedDequeue_bits_data_T_1676[76], _alignedDequeue_bits_data_T_1546[76]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_84 = {_alignedDequeue_bits_data_T_1936[76], _alignedDequeue_bits_data_T_1806[76]};
  wire [3:0]    alignedDequeue_bits_data_hi_84 = {alignedDequeue_bits_data_hi_hi_84, alignedDequeue_bits_data_hi_lo_84};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_85 = {_alignedDequeue_bits_data_T_1156[77], _alignedDequeue_bits_data_T_1026[77]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_85 = {_alignedDequeue_bits_data_T_1416[77], _alignedDequeue_bits_data_T_1286[77]};
  wire [3:0]    alignedDequeue_bits_data_lo_85 = {alignedDequeue_bits_data_lo_hi_85, alignedDequeue_bits_data_lo_lo_85};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_85 = {_alignedDequeue_bits_data_T_1676[77], _alignedDequeue_bits_data_T_1546[77]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_85 = {_alignedDequeue_bits_data_T_1936[77], _alignedDequeue_bits_data_T_1806[77]};
  wire [3:0]    alignedDequeue_bits_data_hi_85 = {alignedDequeue_bits_data_hi_hi_85, alignedDequeue_bits_data_hi_lo_85};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_86 = {_alignedDequeue_bits_data_T_1156[78], _alignedDequeue_bits_data_T_1026[78]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_86 = {_alignedDequeue_bits_data_T_1416[78], _alignedDequeue_bits_data_T_1286[78]};
  wire [3:0]    alignedDequeue_bits_data_lo_86 = {alignedDequeue_bits_data_lo_hi_86, alignedDequeue_bits_data_lo_lo_86};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_86 = {_alignedDequeue_bits_data_T_1676[78], _alignedDequeue_bits_data_T_1546[78]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_86 = {_alignedDequeue_bits_data_T_1936[78], _alignedDequeue_bits_data_T_1806[78]};
  wire [3:0]    alignedDequeue_bits_data_hi_86 = {alignedDequeue_bits_data_hi_hi_86, alignedDequeue_bits_data_hi_lo_86};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_87 = {_alignedDequeue_bits_data_T_1156[79], _alignedDequeue_bits_data_T_1026[79]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_87 = {_alignedDequeue_bits_data_T_1416[79], _alignedDequeue_bits_data_T_1286[79]};
  wire [3:0]    alignedDequeue_bits_data_lo_87 = {alignedDequeue_bits_data_lo_hi_87, alignedDequeue_bits_data_lo_lo_87};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_87 = {_alignedDequeue_bits_data_T_1676[79], _alignedDequeue_bits_data_T_1546[79]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_87 = {_alignedDequeue_bits_data_T_1936[79], _alignedDequeue_bits_data_T_1806[79]};
  wire [3:0]    alignedDequeue_bits_data_hi_87 = {alignedDequeue_bits_data_hi_hi_87, alignedDequeue_bits_data_hi_lo_87};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_88 = {_alignedDequeue_bits_data_T_1156[80], _alignedDequeue_bits_data_T_1026[80]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_88 = {_alignedDequeue_bits_data_T_1416[80], _alignedDequeue_bits_data_T_1286[80]};
  wire [3:0]    alignedDequeue_bits_data_lo_88 = {alignedDequeue_bits_data_lo_hi_88, alignedDequeue_bits_data_lo_lo_88};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_88 = {_alignedDequeue_bits_data_T_1676[80], _alignedDequeue_bits_data_T_1546[80]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_88 = {_alignedDequeue_bits_data_T_1936[80], _alignedDequeue_bits_data_T_1806[80]};
  wire [3:0]    alignedDequeue_bits_data_hi_88 = {alignedDequeue_bits_data_hi_hi_88, alignedDequeue_bits_data_hi_lo_88};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_89 = {_alignedDequeue_bits_data_T_1156[81], _alignedDequeue_bits_data_T_1026[81]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_89 = {_alignedDequeue_bits_data_T_1416[81], _alignedDequeue_bits_data_T_1286[81]};
  wire [3:0]    alignedDequeue_bits_data_lo_89 = {alignedDequeue_bits_data_lo_hi_89, alignedDequeue_bits_data_lo_lo_89};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_89 = {_alignedDequeue_bits_data_T_1676[81], _alignedDequeue_bits_data_T_1546[81]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_89 = {_alignedDequeue_bits_data_T_1936[81], _alignedDequeue_bits_data_T_1806[81]};
  wire [3:0]    alignedDequeue_bits_data_hi_89 = {alignedDequeue_bits_data_hi_hi_89, alignedDequeue_bits_data_hi_lo_89};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_90 = {_alignedDequeue_bits_data_T_1156[82], _alignedDequeue_bits_data_T_1026[82]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_90 = {_alignedDequeue_bits_data_T_1416[82], _alignedDequeue_bits_data_T_1286[82]};
  wire [3:0]    alignedDequeue_bits_data_lo_90 = {alignedDequeue_bits_data_lo_hi_90, alignedDequeue_bits_data_lo_lo_90};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_90 = {_alignedDequeue_bits_data_T_1676[82], _alignedDequeue_bits_data_T_1546[82]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_90 = {_alignedDequeue_bits_data_T_1936[82], _alignedDequeue_bits_data_T_1806[82]};
  wire [3:0]    alignedDequeue_bits_data_hi_90 = {alignedDequeue_bits_data_hi_hi_90, alignedDequeue_bits_data_hi_lo_90};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_91 = {_alignedDequeue_bits_data_T_1156[83], _alignedDequeue_bits_data_T_1026[83]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_91 = {_alignedDequeue_bits_data_T_1416[83], _alignedDequeue_bits_data_T_1286[83]};
  wire [3:0]    alignedDequeue_bits_data_lo_91 = {alignedDequeue_bits_data_lo_hi_91, alignedDequeue_bits_data_lo_lo_91};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_91 = {_alignedDequeue_bits_data_T_1676[83], _alignedDequeue_bits_data_T_1546[83]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_91 = {_alignedDequeue_bits_data_T_1936[83], _alignedDequeue_bits_data_T_1806[83]};
  wire [3:0]    alignedDequeue_bits_data_hi_91 = {alignedDequeue_bits_data_hi_hi_91, alignedDequeue_bits_data_hi_lo_91};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_92 = {_alignedDequeue_bits_data_T_1156[84], _alignedDequeue_bits_data_T_1026[84]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_92 = {_alignedDequeue_bits_data_T_1416[84], _alignedDequeue_bits_data_T_1286[84]};
  wire [3:0]    alignedDequeue_bits_data_lo_92 = {alignedDequeue_bits_data_lo_hi_92, alignedDequeue_bits_data_lo_lo_92};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_92 = {_alignedDequeue_bits_data_T_1676[84], _alignedDequeue_bits_data_T_1546[84]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_92 = {_alignedDequeue_bits_data_T_1936[84], _alignedDequeue_bits_data_T_1806[84]};
  wire [3:0]    alignedDequeue_bits_data_hi_92 = {alignedDequeue_bits_data_hi_hi_92, alignedDequeue_bits_data_hi_lo_92};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_93 = {_alignedDequeue_bits_data_T_1156[85], _alignedDequeue_bits_data_T_1026[85]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_93 = {_alignedDequeue_bits_data_T_1416[85], _alignedDequeue_bits_data_T_1286[85]};
  wire [3:0]    alignedDequeue_bits_data_lo_93 = {alignedDequeue_bits_data_lo_hi_93, alignedDequeue_bits_data_lo_lo_93};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_93 = {_alignedDequeue_bits_data_T_1676[85], _alignedDequeue_bits_data_T_1546[85]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_93 = {_alignedDequeue_bits_data_T_1936[85], _alignedDequeue_bits_data_T_1806[85]};
  wire [3:0]    alignedDequeue_bits_data_hi_93 = {alignedDequeue_bits_data_hi_hi_93, alignedDequeue_bits_data_hi_lo_93};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_94 = {_alignedDequeue_bits_data_T_1156[86], _alignedDequeue_bits_data_T_1026[86]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_94 = {_alignedDequeue_bits_data_T_1416[86], _alignedDequeue_bits_data_T_1286[86]};
  wire [3:0]    alignedDequeue_bits_data_lo_94 = {alignedDequeue_bits_data_lo_hi_94, alignedDequeue_bits_data_lo_lo_94};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_94 = {_alignedDequeue_bits_data_T_1676[86], _alignedDequeue_bits_data_T_1546[86]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_94 = {_alignedDequeue_bits_data_T_1936[86], _alignedDequeue_bits_data_T_1806[86]};
  wire [3:0]    alignedDequeue_bits_data_hi_94 = {alignedDequeue_bits_data_hi_hi_94, alignedDequeue_bits_data_hi_lo_94};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_95 = {_alignedDequeue_bits_data_T_1156[87], _alignedDequeue_bits_data_T_1026[87]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_95 = {_alignedDequeue_bits_data_T_1416[87], _alignedDequeue_bits_data_T_1286[87]};
  wire [3:0]    alignedDequeue_bits_data_lo_95 = {alignedDequeue_bits_data_lo_hi_95, alignedDequeue_bits_data_lo_lo_95};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_95 = {_alignedDequeue_bits_data_T_1676[87], _alignedDequeue_bits_data_T_1546[87]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_95 = {_alignedDequeue_bits_data_T_1936[87], _alignedDequeue_bits_data_T_1806[87]};
  wire [3:0]    alignedDequeue_bits_data_hi_95 = {alignedDequeue_bits_data_hi_hi_95, alignedDequeue_bits_data_hi_lo_95};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_96 = {_alignedDequeue_bits_data_T_1156[88], _alignedDequeue_bits_data_T_1026[88]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_96 = {_alignedDequeue_bits_data_T_1416[88], _alignedDequeue_bits_data_T_1286[88]};
  wire [3:0]    alignedDequeue_bits_data_lo_96 = {alignedDequeue_bits_data_lo_hi_96, alignedDequeue_bits_data_lo_lo_96};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_96 = {_alignedDequeue_bits_data_T_1676[88], _alignedDequeue_bits_data_T_1546[88]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_96 = {_alignedDequeue_bits_data_T_1936[88], _alignedDequeue_bits_data_T_1806[88]};
  wire [3:0]    alignedDequeue_bits_data_hi_96 = {alignedDequeue_bits_data_hi_hi_96, alignedDequeue_bits_data_hi_lo_96};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_97 = {_alignedDequeue_bits_data_T_1156[89], _alignedDequeue_bits_data_T_1026[89]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_97 = {_alignedDequeue_bits_data_T_1416[89], _alignedDequeue_bits_data_T_1286[89]};
  wire [3:0]    alignedDequeue_bits_data_lo_97 = {alignedDequeue_bits_data_lo_hi_97, alignedDequeue_bits_data_lo_lo_97};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_97 = {_alignedDequeue_bits_data_T_1676[89], _alignedDequeue_bits_data_T_1546[89]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_97 = {_alignedDequeue_bits_data_T_1936[89], _alignedDequeue_bits_data_T_1806[89]};
  wire [3:0]    alignedDequeue_bits_data_hi_97 = {alignedDequeue_bits_data_hi_hi_97, alignedDequeue_bits_data_hi_lo_97};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_98 = {_alignedDequeue_bits_data_T_1156[90], _alignedDequeue_bits_data_T_1026[90]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_98 = {_alignedDequeue_bits_data_T_1416[90], _alignedDequeue_bits_data_T_1286[90]};
  wire [3:0]    alignedDequeue_bits_data_lo_98 = {alignedDequeue_bits_data_lo_hi_98, alignedDequeue_bits_data_lo_lo_98};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_98 = {_alignedDequeue_bits_data_T_1676[90], _alignedDequeue_bits_data_T_1546[90]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_98 = {_alignedDequeue_bits_data_T_1936[90], _alignedDequeue_bits_data_T_1806[90]};
  wire [3:0]    alignedDequeue_bits_data_hi_98 = {alignedDequeue_bits_data_hi_hi_98, alignedDequeue_bits_data_hi_lo_98};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_99 = {_alignedDequeue_bits_data_T_1156[91], _alignedDequeue_bits_data_T_1026[91]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_99 = {_alignedDequeue_bits_data_T_1416[91], _alignedDequeue_bits_data_T_1286[91]};
  wire [3:0]    alignedDequeue_bits_data_lo_99 = {alignedDequeue_bits_data_lo_hi_99, alignedDequeue_bits_data_lo_lo_99};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_99 = {_alignedDequeue_bits_data_T_1676[91], _alignedDequeue_bits_data_T_1546[91]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_99 = {_alignedDequeue_bits_data_T_1936[91], _alignedDequeue_bits_data_T_1806[91]};
  wire [3:0]    alignedDequeue_bits_data_hi_99 = {alignedDequeue_bits_data_hi_hi_99, alignedDequeue_bits_data_hi_lo_99};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_100 = {_alignedDequeue_bits_data_T_1156[92], _alignedDequeue_bits_data_T_1026[92]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_100 = {_alignedDequeue_bits_data_T_1416[92], _alignedDequeue_bits_data_T_1286[92]};
  wire [3:0]    alignedDequeue_bits_data_lo_100 = {alignedDequeue_bits_data_lo_hi_100, alignedDequeue_bits_data_lo_lo_100};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_100 = {_alignedDequeue_bits_data_T_1676[92], _alignedDequeue_bits_data_T_1546[92]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_100 = {_alignedDequeue_bits_data_T_1936[92], _alignedDequeue_bits_data_T_1806[92]};
  wire [3:0]    alignedDequeue_bits_data_hi_100 = {alignedDequeue_bits_data_hi_hi_100, alignedDequeue_bits_data_hi_lo_100};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_101 = {_alignedDequeue_bits_data_T_1156[93], _alignedDequeue_bits_data_T_1026[93]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_101 = {_alignedDequeue_bits_data_T_1416[93], _alignedDequeue_bits_data_T_1286[93]};
  wire [3:0]    alignedDequeue_bits_data_lo_101 = {alignedDequeue_bits_data_lo_hi_101, alignedDequeue_bits_data_lo_lo_101};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_101 = {_alignedDequeue_bits_data_T_1676[93], _alignedDequeue_bits_data_T_1546[93]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_101 = {_alignedDequeue_bits_data_T_1936[93], _alignedDequeue_bits_data_T_1806[93]};
  wire [3:0]    alignedDequeue_bits_data_hi_101 = {alignedDequeue_bits_data_hi_hi_101, alignedDequeue_bits_data_hi_lo_101};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_102 = {_alignedDequeue_bits_data_T_1156[94], _alignedDequeue_bits_data_T_1026[94]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_102 = {_alignedDequeue_bits_data_T_1416[94], _alignedDequeue_bits_data_T_1286[94]};
  wire [3:0]    alignedDequeue_bits_data_lo_102 = {alignedDequeue_bits_data_lo_hi_102, alignedDequeue_bits_data_lo_lo_102};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_102 = {_alignedDequeue_bits_data_T_1676[94], _alignedDequeue_bits_data_T_1546[94]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_102 = {_alignedDequeue_bits_data_T_1936[94], _alignedDequeue_bits_data_T_1806[94]};
  wire [3:0]    alignedDequeue_bits_data_hi_102 = {alignedDequeue_bits_data_hi_hi_102, alignedDequeue_bits_data_hi_lo_102};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_103 = {_alignedDequeue_bits_data_T_1156[95], _alignedDequeue_bits_data_T_1026[95]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_103 = {_alignedDequeue_bits_data_T_1416[95], _alignedDequeue_bits_data_T_1286[95]};
  wire [3:0]    alignedDequeue_bits_data_lo_103 = {alignedDequeue_bits_data_lo_hi_103, alignedDequeue_bits_data_lo_lo_103};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_103 = {_alignedDequeue_bits_data_T_1676[95], _alignedDequeue_bits_data_T_1546[95]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_103 = {_alignedDequeue_bits_data_T_1936[95], _alignedDequeue_bits_data_T_1806[95]};
  wire [3:0]    alignedDequeue_bits_data_hi_103 = {alignedDequeue_bits_data_hi_hi_103, alignedDequeue_bits_data_hi_lo_103};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_104 = {_alignedDequeue_bits_data_T_1156[96], _alignedDequeue_bits_data_T_1026[96]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_104 = {_alignedDequeue_bits_data_T_1416[96], _alignedDequeue_bits_data_T_1286[96]};
  wire [3:0]    alignedDequeue_bits_data_lo_104 = {alignedDequeue_bits_data_lo_hi_104, alignedDequeue_bits_data_lo_lo_104};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_104 = {_alignedDequeue_bits_data_T_1676[96], _alignedDequeue_bits_data_T_1546[96]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_104 = {_alignedDequeue_bits_data_T_1936[96], _alignedDequeue_bits_data_T_1806[96]};
  wire [3:0]    alignedDequeue_bits_data_hi_104 = {alignedDequeue_bits_data_hi_hi_104, alignedDequeue_bits_data_hi_lo_104};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_105 = {_alignedDequeue_bits_data_T_1156[97], _alignedDequeue_bits_data_T_1026[97]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_105 = {_alignedDequeue_bits_data_T_1416[97], _alignedDequeue_bits_data_T_1286[97]};
  wire [3:0]    alignedDequeue_bits_data_lo_105 = {alignedDequeue_bits_data_lo_hi_105, alignedDequeue_bits_data_lo_lo_105};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_105 = {_alignedDequeue_bits_data_T_1676[97], _alignedDequeue_bits_data_T_1546[97]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_105 = {_alignedDequeue_bits_data_T_1936[97], _alignedDequeue_bits_data_T_1806[97]};
  wire [3:0]    alignedDequeue_bits_data_hi_105 = {alignedDequeue_bits_data_hi_hi_105, alignedDequeue_bits_data_hi_lo_105};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_106 = {_alignedDequeue_bits_data_T_1156[98], _alignedDequeue_bits_data_T_1026[98]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_106 = {_alignedDequeue_bits_data_T_1416[98], _alignedDequeue_bits_data_T_1286[98]};
  wire [3:0]    alignedDequeue_bits_data_lo_106 = {alignedDequeue_bits_data_lo_hi_106, alignedDequeue_bits_data_lo_lo_106};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_106 = {_alignedDequeue_bits_data_T_1676[98], _alignedDequeue_bits_data_T_1546[98]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_106 = {_alignedDequeue_bits_data_T_1936[98], _alignedDequeue_bits_data_T_1806[98]};
  wire [3:0]    alignedDequeue_bits_data_hi_106 = {alignedDequeue_bits_data_hi_hi_106, alignedDequeue_bits_data_hi_lo_106};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_107 = {_alignedDequeue_bits_data_T_1156[99], _alignedDequeue_bits_data_T_1026[99]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_107 = {_alignedDequeue_bits_data_T_1416[99], _alignedDequeue_bits_data_T_1286[99]};
  wire [3:0]    alignedDequeue_bits_data_lo_107 = {alignedDequeue_bits_data_lo_hi_107, alignedDequeue_bits_data_lo_lo_107};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_107 = {_alignedDequeue_bits_data_T_1676[99], _alignedDequeue_bits_data_T_1546[99]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_107 = {_alignedDequeue_bits_data_T_1936[99], _alignedDequeue_bits_data_T_1806[99]};
  wire [3:0]    alignedDequeue_bits_data_hi_107 = {alignedDequeue_bits_data_hi_hi_107, alignedDequeue_bits_data_hi_lo_107};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_108 = {_alignedDequeue_bits_data_T_1156[100], _alignedDequeue_bits_data_T_1026[100]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_108 = {_alignedDequeue_bits_data_T_1416[100], _alignedDequeue_bits_data_T_1286[100]};
  wire [3:0]    alignedDequeue_bits_data_lo_108 = {alignedDequeue_bits_data_lo_hi_108, alignedDequeue_bits_data_lo_lo_108};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_108 = {_alignedDequeue_bits_data_T_1676[100], _alignedDequeue_bits_data_T_1546[100]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_108 = {_alignedDequeue_bits_data_T_1936[100], _alignedDequeue_bits_data_T_1806[100]};
  wire [3:0]    alignedDequeue_bits_data_hi_108 = {alignedDequeue_bits_data_hi_hi_108, alignedDequeue_bits_data_hi_lo_108};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_109 = {_alignedDequeue_bits_data_T_1156[101], _alignedDequeue_bits_data_T_1026[101]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_109 = {_alignedDequeue_bits_data_T_1416[101], _alignedDequeue_bits_data_T_1286[101]};
  wire [3:0]    alignedDequeue_bits_data_lo_109 = {alignedDequeue_bits_data_lo_hi_109, alignedDequeue_bits_data_lo_lo_109};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_109 = {_alignedDequeue_bits_data_T_1676[101], _alignedDequeue_bits_data_T_1546[101]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_109 = {_alignedDequeue_bits_data_T_1936[101], _alignedDequeue_bits_data_T_1806[101]};
  wire [3:0]    alignedDequeue_bits_data_hi_109 = {alignedDequeue_bits_data_hi_hi_109, alignedDequeue_bits_data_hi_lo_109};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_110 = {_alignedDequeue_bits_data_T_1156[102], _alignedDequeue_bits_data_T_1026[102]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_110 = {_alignedDequeue_bits_data_T_1416[102], _alignedDequeue_bits_data_T_1286[102]};
  wire [3:0]    alignedDequeue_bits_data_lo_110 = {alignedDequeue_bits_data_lo_hi_110, alignedDequeue_bits_data_lo_lo_110};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_110 = {_alignedDequeue_bits_data_T_1676[102], _alignedDequeue_bits_data_T_1546[102]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_110 = {_alignedDequeue_bits_data_T_1936[102], _alignedDequeue_bits_data_T_1806[102]};
  wire [3:0]    alignedDequeue_bits_data_hi_110 = {alignedDequeue_bits_data_hi_hi_110, alignedDequeue_bits_data_hi_lo_110};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_111 = {_alignedDequeue_bits_data_T_1156[103], _alignedDequeue_bits_data_T_1026[103]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_111 = {_alignedDequeue_bits_data_T_1416[103], _alignedDequeue_bits_data_T_1286[103]};
  wire [3:0]    alignedDequeue_bits_data_lo_111 = {alignedDequeue_bits_data_lo_hi_111, alignedDequeue_bits_data_lo_lo_111};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_111 = {_alignedDequeue_bits_data_T_1676[103], _alignedDequeue_bits_data_T_1546[103]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_111 = {_alignedDequeue_bits_data_T_1936[103], _alignedDequeue_bits_data_T_1806[103]};
  wire [3:0]    alignedDequeue_bits_data_hi_111 = {alignedDequeue_bits_data_hi_hi_111, alignedDequeue_bits_data_hi_lo_111};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_112 = {_alignedDequeue_bits_data_T_1156[104], _alignedDequeue_bits_data_T_1026[104]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_112 = {_alignedDequeue_bits_data_T_1416[104], _alignedDequeue_bits_data_T_1286[104]};
  wire [3:0]    alignedDequeue_bits_data_lo_112 = {alignedDequeue_bits_data_lo_hi_112, alignedDequeue_bits_data_lo_lo_112};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_112 = {_alignedDequeue_bits_data_T_1676[104], _alignedDequeue_bits_data_T_1546[104]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_112 = {_alignedDequeue_bits_data_T_1936[104], _alignedDequeue_bits_data_T_1806[104]};
  wire [3:0]    alignedDequeue_bits_data_hi_112 = {alignedDequeue_bits_data_hi_hi_112, alignedDequeue_bits_data_hi_lo_112};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_113 = {_alignedDequeue_bits_data_T_1156[105], _alignedDequeue_bits_data_T_1026[105]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_113 = {_alignedDequeue_bits_data_T_1416[105], _alignedDequeue_bits_data_T_1286[105]};
  wire [3:0]    alignedDequeue_bits_data_lo_113 = {alignedDequeue_bits_data_lo_hi_113, alignedDequeue_bits_data_lo_lo_113};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_113 = {_alignedDequeue_bits_data_T_1676[105], _alignedDequeue_bits_data_T_1546[105]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_113 = {_alignedDequeue_bits_data_T_1936[105], _alignedDequeue_bits_data_T_1806[105]};
  wire [3:0]    alignedDequeue_bits_data_hi_113 = {alignedDequeue_bits_data_hi_hi_113, alignedDequeue_bits_data_hi_lo_113};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_114 = {_alignedDequeue_bits_data_T_1156[106], _alignedDequeue_bits_data_T_1026[106]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_114 = {_alignedDequeue_bits_data_T_1416[106], _alignedDequeue_bits_data_T_1286[106]};
  wire [3:0]    alignedDequeue_bits_data_lo_114 = {alignedDequeue_bits_data_lo_hi_114, alignedDequeue_bits_data_lo_lo_114};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_114 = {_alignedDequeue_bits_data_T_1676[106], _alignedDequeue_bits_data_T_1546[106]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_114 = {_alignedDequeue_bits_data_T_1936[106], _alignedDequeue_bits_data_T_1806[106]};
  wire [3:0]    alignedDequeue_bits_data_hi_114 = {alignedDequeue_bits_data_hi_hi_114, alignedDequeue_bits_data_hi_lo_114};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_115 = {_alignedDequeue_bits_data_T_1156[107], _alignedDequeue_bits_data_T_1026[107]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_115 = {_alignedDequeue_bits_data_T_1416[107], _alignedDequeue_bits_data_T_1286[107]};
  wire [3:0]    alignedDequeue_bits_data_lo_115 = {alignedDequeue_bits_data_lo_hi_115, alignedDequeue_bits_data_lo_lo_115};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_115 = {_alignedDequeue_bits_data_T_1676[107], _alignedDequeue_bits_data_T_1546[107]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_115 = {_alignedDequeue_bits_data_T_1936[107], _alignedDequeue_bits_data_T_1806[107]};
  wire [3:0]    alignedDequeue_bits_data_hi_115 = {alignedDequeue_bits_data_hi_hi_115, alignedDequeue_bits_data_hi_lo_115};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_116 = {_alignedDequeue_bits_data_T_1156[108], _alignedDequeue_bits_data_T_1026[108]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_116 = {_alignedDequeue_bits_data_T_1416[108], _alignedDequeue_bits_data_T_1286[108]};
  wire [3:0]    alignedDequeue_bits_data_lo_116 = {alignedDequeue_bits_data_lo_hi_116, alignedDequeue_bits_data_lo_lo_116};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_116 = {_alignedDequeue_bits_data_T_1676[108], _alignedDequeue_bits_data_T_1546[108]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_116 = {_alignedDequeue_bits_data_T_1936[108], _alignedDequeue_bits_data_T_1806[108]};
  wire [3:0]    alignedDequeue_bits_data_hi_116 = {alignedDequeue_bits_data_hi_hi_116, alignedDequeue_bits_data_hi_lo_116};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_117 = {_alignedDequeue_bits_data_T_1156[109], _alignedDequeue_bits_data_T_1026[109]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_117 = {_alignedDequeue_bits_data_T_1416[109], _alignedDequeue_bits_data_T_1286[109]};
  wire [3:0]    alignedDequeue_bits_data_lo_117 = {alignedDequeue_bits_data_lo_hi_117, alignedDequeue_bits_data_lo_lo_117};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_117 = {_alignedDequeue_bits_data_T_1676[109], _alignedDequeue_bits_data_T_1546[109]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_117 = {_alignedDequeue_bits_data_T_1936[109], _alignedDequeue_bits_data_T_1806[109]};
  wire [3:0]    alignedDequeue_bits_data_hi_117 = {alignedDequeue_bits_data_hi_hi_117, alignedDequeue_bits_data_hi_lo_117};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_118 = {_alignedDequeue_bits_data_T_1156[110], _alignedDequeue_bits_data_T_1026[110]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_118 = {_alignedDequeue_bits_data_T_1416[110], _alignedDequeue_bits_data_T_1286[110]};
  wire [3:0]    alignedDequeue_bits_data_lo_118 = {alignedDequeue_bits_data_lo_hi_118, alignedDequeue_bits_data_lo_lo_118};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_118 = {_alignedDequeue_bits_data_T_1676[110], _alignedDequeue_bits_data_T_1546[110]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_118 = {_alignedDequeue_bits_data_T_1936[110], _alignedDequeue_bits_data_T_1806[110]};
  wire [3:0]    alignedDequeue_bits_data_hi_118 = {alignedDequeue_bits_data_hi_hi_118, alignedDequeue_bits_data_hi_lo_118};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_119 = {_alignedDequeue_bits_data_T_1156[111], _alignedDequeue_bits_data_T_1026[111]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_119 = {_alignedDequeue_bits_data_T_1416[111], _alignedDequeue_bits_data_T_1286[111]};
  wire [3:0]    alignedDequeue_bits_data_lo_119 = {alignedDequeue_bits_data_lo_hi_119, alignedDequeue_bits_data_lo_lo_119};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_119 = {_alignedDequeue_bits_data_T_1676[111], _alignedDequeue_bits_data_T_1546[111]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_119 = {_alignedDequeue_bits_data_T_1936[111], _alignedDequeue_bits_data_T_1806[111]};
  wire [3:0]    alignedDequeue_bits_data_hi_119 = {alignedDequeue_bits_data_hi_hi_119, alignedDequeue_bits_data_hi_lo_119};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_120 = {_alignedDequeue_bits_data_T_1156[112], _alignedDequeue_bits_data_T_1026[112]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_120 = {_alignedDequeue_bits_data_T_1416[112], _alignedDequeue_bits_data_T_1286[112]};
  wire [3:0]    alignedDequeue_bits_data_lo_120 = {alignedDequeue_bits_data_lo_hi_120, alignedDequeue_bits_data_lo_lo_120};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_120 = {_alignedDequeue_bits_data_T_1676[112], _alignedDequeue_bits_data_T_1546[112]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_120 = {_alignedDequeue_bits_data_T_1936[112], _alignedDequeue_bits_data_T_1806[112]};
  wire [3:0]    alignedDequeue_bits_data_hi_120 = {alignedDequeue_bits_data_hi_hi_120, alignedDequeue_bits_data_hi_lo_120};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_121 = {_alignedDequeue_bits_data_T_1156[113], _alignedDequeue_bits_data_T_1026[113]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_121 = {_alignedDequeue_bits_data_T_1416[113], _alignedDequeue_bits_data_T_1286[113]};
  wire [3:0]    alignedDequeue_bits_data_lo_121 = {alignedDequeue_bits_data_lo_hi_121, alignedDequeue_bits_data_lo_lo_121};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_121 = {_alignedDequeue_bits_data_T_1676[113], _alignedDequeue_bits_data_T_1546[113]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_121 = {_alignedDequeue_bits_data_T_1936[113], _alignedDequeue_bits_data_T_1806[113]};
  wire [3:0]    alignedDequeue_bits_data_hi_121 = {alignedDequeue_bits_data_hi_hi_121, alignedDequeue_bits_data_hi_lo_121};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_122 = {_alignedDequeue_bits_data_T_1156[114], _alignedDequeue_bits_data_T_1026[114]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_122 = {_alignedDequeue_bits_data_T_1416[114], _alignedDequeue_bits_data_T_1286[114]};
  wire [3:0]    alignedDequeue_bits_data_lo_122 = {alignedDequeue_bits_data_lo_hi_122, alignedDequeue_bits_data_lo_lo_122};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_122 = {_alignedDequeue_bits_data_T_1676[114], _alignedDequeue_bits_data_T_1546[114]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_122 = {_alignedDequeue_bits_data_T_1936[114], _alignedDequeue_bits_data_T_1806[114]};
  wire [3:0]    alignedDequeue_bits_data_hi_122 = {alignedDequeue_bits_data_hi_hi_122, alignedDequeue_bits_data_hi_lo_122};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_123 = {_alignedDequeue_bits_data_T_1156[115], _alignedDequeue_bits_data_T_1026[115]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_123 = {_alignedDequeue_bits_data_T_1416[115], _alignedDequeue_bits_data_T_1286[115]};
  wire [3:0]    alignedDequeue_bits_data_lo_123 = {alignedDequeue_bits_data_lo_hi_123, alignedDequeue_bits_data_lo_lo_123};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_123 = {_alignedDequeue_bits_data_T_1676[115], _alignedDequeue_bits_data_T_1546[115]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_123 = {_alignedDequeue_bits_data_T_1936[115], _alignedDequeue_bits_data_T_1806[115]};
  wire [3:0]    alignedDequeue_bits_data_hi_123 = {alignedDequeue_bits_data_hi_hi_123, alignedDequeue_bits_data_hi_lo_123};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_124 = {_alignedDequeue_bits_data_T_1156[116], _alignedDequeue_bits_data_T_1026[116]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_124 = {_alignedDequeue_bits_data_T_1416[116], _alignedDequeue_bits_data_T_1286[116]};
  wire [3:0]    alignedDequeue_bits_data_lo_124 = {alignedDequeue_bits_data_lo_hi_124, alignedDequeue_bits_data_lo_lo_124};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_124 = {_alignedDequeue_bits_data_T_1676[116], _alignedDequeue_bits_data_T_1546[116]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_124 = {_alignedDequeue_bits_data_T_1936[116], _alignedDequeue_bits_data_T_1806[116]};
  wire [3:0]    alignedDequeue_bits_data_hi_124 = {alignedDequeue_bits_data_hi_hi_124, alignedDequeue_bits_data_hi_lo_124};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_125 = {_alignedDequeue_bits_data_T_1156[117], _alignedDequeue_bits_data_T_1026[117]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_125 = {_alignedDequeue_bits_data_T_1416[117], _alignedDequeue_bits_data_T_1286[117]};
  wire [3:0]    alignedDequeue_bits_data_lo_125 = {alignedDequeue_bits_data_lo_hi_125, alignedDequeue_bits_data_lo_lo_125};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_125 = {_alignedDequeue_bits_data_T_1676[117], _alignedDequeue_bits_data_T_1546[117]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_125 = {_alignedDequeue_bits_data_T_1936[117], _alignedDequeue_bits_data_T_1806[117]};
  wire [3:0]    alignedDequeue_bits_data_hi_125 = {alignedDequeue_bits_data_hi_hi_125, alignedDequeue_bits_data_hi_lo_125};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_126 = {_alignedDequeue_bits_data_T_1156[118], _alignedDequeue_bits_data_T_1026[118]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_126 = {_alignedDequeue_bits_data_T_1416[118], _alignedDequeue_bits_data_T_1286[118]};
  wire [3:0]    alignedDequeue_bits_data_lo_126 = {alignedDequeue_bits_data_lo_hi_126, alignedDequeue_bits_data_lo_lo_126};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_126 = {_alignedDequeue_bits_data_T_1676[118], _alignedDequeue_bits_data_T_1546[118]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_126 = {_alignedDequeue_bits_data_T_1936[118], _alignedDequeue_bits_data_T_1806[118]};
  wire [3:0]    alignedDequeue_bits_data_hi_126 = {alignedDequeue_bits_data_hi_hi_126, alignedDequeue_bits_data_hi_lo_126};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_127 = {_alignedDequeue_bits_data_T_1156[119], _alignedDequeue_bits_data_T_1026[119]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_127 = {_alignedDequeue_bits_data_T_1416[119], _alignedDequeue_bits_data_T_1286[119]};
  wire [3:0]    alignedDequeue_bits_data_lo_127 = {alignedDequeue_bits_data_lo_hi_127, alignedDequeue_bits_data_lo_lo_127};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_127 = {_alignedDequeue_bits_data_T_1676[119], _alignedDequeue_bits_data_T_1546[119]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_127 = {_alignedDequeue_bits_data_T_1936[119], _alignedDequeue_bits_data_T_1806[119]};
  wire [3:0]    alignedDequeue_bits_data_hi_127 = {alignedDequeue_bits_data_hi_hi_127, alignedDequeue_bits_data_hi_lo_127};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_128 = {_alignedDequeue_bits_data_T_1156[120], _alignedDequeue_bits_data_T_1026[120]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_128 = {_alignedDequeue_bits_data_T_1416[120], _alignedDequeue_bits_data_T_1286[120]};
  wire [3:0]    alignedDequeue_bits_data_lo_128 = {alignedDequeue_bits_data_lo_hi_128, alignedDequeue_bits_data_lo_lo_128};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_128 = {_alignedDequeue_bits_data_T_1676[120], _alignedDequeue_bits_data_T_1546[120]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_128 = {_alignedDequeue_bits_data_T_1936[120], _alignedDequeue_bits_data_T_1806[120]};
  wire [3:0]    alignedDequeue_bits_data_hi_128 = {alignedDequeue_bits_data_hi_hi_128, alignedDequeue_bits_data_hi_lo_128};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_129 = {_alignedDequeue_bits_data_T_1156[121], _alignedDequeue_bits_data_T_1026[121]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_129 = {_alignedDequeue_bits_data_T_1416[121], _alignedDequeue_bits_data_T_1286[121]};
  wire [3:0]    alignedDequeue_bits_data_lo_129 = {alignedDequeue_bits_data_lo_hi_129, alignedDequeue_bits_data_lo_lo_129};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_129 = {_alignedDequeue_bits_data_T_1676[121], _alignedDequeue_bits_data_T_1546[121]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_129 = {_alignedDequeue_bits_data_T_1936[121], _alignedDequeue_bits_data_T_1806[121]};
  wire [3:0]    alignedDequeue_bits_data_hi_129 = {alignedDequeue_bits_data_hi_hi_129, alignedDequeue_bits_data_hi_lo_129};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_130 = {_alignedDequeue_bits_data_T_1156[122], _alignedDequeue_bits_data_T_1026[122]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_130 = {_alignedDequeue_bits_data_T_1416[122], _alignedDequeue_bits_data_T_1286[122]};
  wire [3:0]    alignedDequeue_bits_data_lo_130 = {alignedDequeue_bits_data_lo_hi_130, alignedDequeue_bits_data_lo_lo_130};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_130 = {_alignedDequeue_bits_data_T_1676[122], _alignedDequeue_bits_data_T_1546[122]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_130 = {_alignedDequeue_bits_data_T_1936[122], _alignedDequeue_bits_data_T_1806[122]};
  wire [3:0]    alignedDequeue_bits_data_hi_130 = {alignedDequeue_bits_data_hi_hi_130, alignedDequeue_bits_data_hi_lo_130};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_131 = {_alignedDequeue_bits_data_T_1156[123], _alignedDequeue_bits_data_T_1026[123]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_131 = {_alignedDequeue_bits_data_T_1416[123], _alignedDequeue_bits_data_T_1286[123]};
  wire [3:0]    alignedDequeue_bits_data_lo_131 = {alignedDequeue_bits_data_lo_hi_131, alignedDequeue_bits_data_lo_lo_131};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_131 = {_alignedDequeue_bits_data_T_1676[123], _alignedDequeue_bits_data_T_1546[123]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_131 = {_alignedDequeue_bits_data_T_1936[123], _alignedDequeue_bits_data_T_1806[123]};
  wire [3:0]    alignedDequeue_bits_data_hi_131 = {alignedDequeue_bits_data_hi_hi_131, alignedDequeue_bits_data_hi_lo_131};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_132 = {_alignedDequeue_bits_data_T_1156[124], _alignedDequeue_bits_data_T_1026[124]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_132 = {_alignedDequeue_bits_data_T_1416[124], _alignedDequeue_bits_data_T_1286[124]};
  wire [3:0]    alignedDequeue_bits_data_lo_132 = {alignedDequeue_bits_data_lo_hi_132, alignedDequeue_bits_data_lo_lo_132};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_132 = {_alignedDequeue_bits_data_T_1676[124], _alignedDequeue_bits_data_T_1546[124]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_132 = {_alignedDequeue_bits_data_T_1936[124], _alignedDequeue_bits_data_T_1806[124]};
  wire [3:0]    alignedDequeue_bits_data_hi_132 = {alignedDequeue_bits_data_hi_hi_132, alignedDequeue_bits_data_hi_lo_132};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_133 = {_alignedDequeue_bits_data_T_1156[125], _alignedDequeue_bits_data_T_1026[125]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_133 = {_alignedDequeue_bits_data_T_1416[125], _alignedDequeue_bits_data_T_1286[125]};
  wire [3:0]    alignedDequeue_bits_data_lo_133 = {alignedDequeue_bits_data_lo_hi_133, alignedDequeue_bits_data_lo_lo_133};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_133 = {_alignedDequeue_bits_data_T_1676[125], _alignedDequeue_bits_data_T_1546[125]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_133 = {_alignedDequeue_bits_data_T_1936[125], _alignedDequeue_bits_data_T_1806[125]};
  wire [3:0]    alignedDequeue_bits_data_hi_133 = {alignedDequeue_bits_data_hi_hi_133, alignedDequeue_bits_data_hi_lo_133};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_134 = {_alignedDequeue_bits_data_T_1156[126], _alignedDequeue_bits_data_T_1026[126]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_134 = {_alignedDequeue_bits_data_T_1416[126], _alignedDequeue_bits_data_T_1286[126]};
  wire [3:0]    alignedDequeue_bits_data_lo_134 = {alignedDequeue_bits_data_lo_hi_134, alignedDequeue_bits_data_lo_lo_134};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_134 = {_alignedDequeue_bits_data_T_1676[126], _alignedDequeue_bits_data_T_1546[126]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_134 = {_alignedDequeue_bits_data_T_1936[126], _alignedDequeue_bits_data_T_1806[126]};
  wire [3:0]    alignedDequeue_bits_data_hi_134 = {alignedDequeue_bits_data_hi_hi_134, alignedDequeue_bits_data_hi_lo_134};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_135 = {_alignedDequeue_bits_data_T_1156[127], _alignedDequeue_bits_data_T_1026[127]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_135 = {_alignedDequeue_bits_data_T_1416[127], _alignedDequeue_bits_data_T_1286[127]};
  wire [3:0]    alignedDequeue_bits_data_lo_135 = {alignedDequeue_bits_data_lo_hi_135, alignedDequeue_bits_data_lo_lo_135};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_135 = {_alignedDequeue_bits_data_T_1676[127], _alignedDequeue_bits_data_T_1546[127]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_135 = {_alignedDequeue_bits_data_T_1936[127], _alignedDequeue_bits_data_T_1806[127]};
  wire [3:0]    alignedDequeue_bits_data_hi_135 = {alignedDequeue_bits_data_hi_hi_135, alignedDequeue_bits_data_hi_lo_135};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_lo_lo_lo_lo_8 = {alignedDequeue_bits_data_hi_9, alignedDequeue_bits_data_lo_9, alignedDequeue_bits_data_hi_8, alignedDequeue_bits_data_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_lo_lo_lo_hi_8 = {alignedDequeue_bits_data_hi_11, alignedDequeue_bits_data_lo_11, alignedDequeue_bits_data_hi_10, alignedDequeue_bits_data_lo_10};
  wire [31:0]   alignedDequeue_bits_data_lo_lo_lo_lo_lo_8 = {alignedDequeue_bits_data_lo_lo_lo_lo_lo_hi_8, alignedDequeue_bits_data_lo_lo_lo_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_lo_lo_hi_lo_8 = {alignedDequeue_bits_data_hi_13, alignedDequeue_bits_data_lo_13, alignedDequeue_bits_data_hi_12, alignedDequeue_bits_data_lo_12};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_lo_lo_hi_hi_8 = {alignedDequeue_bits_data_hi_15, alignedDequeue_bits_data_lo_15, alignedDequeue_bits_data_hi_14, alignedDequeue_bits_data_lo_14};
  wire [31:0]   alignedDequeue_bits_data_lo_lo_lo_lo_hi_8 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_hi_8, alignedDequeue_bits_data_lo_lo_lo_lo_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_lo_lo_lo_lo_8 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_8, alignedDequeue_bits_data_lo_lo_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_lo_hi_lo_lo_8 = {alignedDequeue_bits_data_hi_17, alignedDequeue_bits_data_lo_17, alignedDequeue_bits_data_hi_16, alignedDequeue_bits_data_lo_16};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_lo_hi_lo_hi_8 = {alignedDequeue_bits_data_hi_19, alignedDequeue_bits_data_lo_19, alignedDequeue_bits_data_hi_18, alignedDequeue_bits_data_lo_18};
  wire [31:0]   alignedDequeue_bits_data_lo_lo_lo_hi_lo_8 = {alignedDequeue_bits_data_lo_lo_lo_hi_lo_hi_8, alignedDequeue_bits_data_lo_lo_lo_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_lo_hi_hi_lo_8 = {alignedDequeue_bits_data_hi_21, alignedDequeue_bits_data_lo_21, alignedDequeue_bits_data_hi_20, alignedDequeue_bits_data_lo_20};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_lo_hi_hi_hi_8 = {alignedDequeue_bits_data_hi_23, alignedDequeue_bits_data_lo_23, alignedDequeue_bits_data_hi_22, alignedDequeue_bits_data_lo_22};
  wire [31:0]   alignedDequeue_bits_data_lo_lo_lo_hi_hi_8 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_hi_8, alignedDequeue_bits_data_lo_lo_lo_hi_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_lo_lo_lo_hi_8 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_8, alignedDequeue_bits_data_lo_lo_lo_hi_lo_8};
  wire [127:0]  alignedDequeue_bits_data_lo_lo_lo_8 = {alignedDequeue_bits_data_lo_lo_lo_hi_8, alignedDequeue_bits_data_lo_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_hi_lo_lo_lo_8 = {alignedDequeue_bits_data_hi_25, alignedDequeue_bits_data_lo_25, alignedDequeue_bits_data_hi_24, alignedDequeue_bits_data_lo_24};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_hi_lo_lo_hi_8 = {alignedDequeue_bits_data_hi_27, alignedDequeue_bits_data_lo_27, alignedDequeue_bits_data_hi_26, alignedDequeue_bits_data_lo_26};
  wire [31:0]   alignedDequeue_bits_data_lo_lo_hi_lo_lo_8 = {alignedDequeue_bits_data_lo_lo_hi_lo_lo_hi_8, alignedDequeue_bits_data_lo_lo_hi_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_hi_lo_hi_lo_8 = {alignedDequeue_bits_data_hi_29, alignedDequeue_bits_data_lo_29, alignedDequeue_bits_data_hi_28, alignedDequeue_bits_data_lo_28};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_hi_lo_hi_hi_8 = {alignedDequeue_bits_data_hi_31, alignedDequeue_bits_data_lo_31, alignedDequeue_bits_data_hi_30, alignedDequeue_bits_data_lo_30};
  wire [31:0]   alignedDequeue_bits_data_lo_lo_hi_lo_hi_8 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_hi_8, alignedDequeue_bits_data_lo_lo_hi_lo_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_lo_lo_hi_lo_8 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_8, alignedDequeue_bits_data_lo_lo_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_hi_hi_lo_lo_8 = {alignedDequeue_bits_data_hi_33, alignedDequeue_bits_data_lo_33, alignedDequeue_bits_data_hi_32, alignedDequeue_bits_data_lo_32};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_hi_hi_lo_hi_8 = {alignedDequeue_bits_data_hi_35, alignedDequeue_bits_data_lo_35, alignedDequeue_bits_data_hi_34, alignedDequeue_bits_data_lo_34};
  wire [31:0]   alignedDequeue_bits_data_lo_lo_hi_hi_lo_8 = {alignedDequeue_bits_data_lo_lo_hi_hi_lo_hi_8, alignedDequeue_bits_data_lo_lo_hi_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_hi_hi_hi_lo_8 = {alignedDequeue_bits_data_hi_37, alignedDequeue_bits_data_lo_37, alignedDequeue_bits_data_hi_36, alignedDequeue_bits_data_lo_36};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_hi_hi_hi_hi_8 = {alignedDequeue_bits_data_hi_39, alignedDequeue_bits_data_lo_39, alignedDequeue_bits_data_hi_38, alignedDequeue_bits_data_lo_38};
  wire [31:0]   alignedDequeue_bits_data_lo_lo_hi_hi_hi_8 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_hi_8, alignedDequeue_bits_data_lo_lo_hi_hi_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_lo_lo_hi_hi_8 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_8, alignedDequeue_bits_data_lo_lo_hi_hi_lo_8};
  wire [127:0]  alignedDequeue_bits_data_lo_lo_hi_8 = {alignedDequeue_bits_data_lo_lo_hi_hi_8, alignedDequeue_bits_data_lo_lo_hi_lo_8};
  wire [255:0]  alignedDequeue_bits_data_lo_lo_136 = {alignedDequeue_bits_data_lo_lo_hi_8, alignedDequeue_bits_data_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_lo_lo_lo_lo_8 = {alignedDequeue_bits_data_hi_41, alignedDequeue_bits_data_lo_41, alignedDequeue_bits_data_hi_40, alignedDequeue_bits_data_lo_40};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_lo_lo_lo_hi_8 = {alignedDequeue_bits_data_hi_43, alignedDequeue_bits_data_lo_43, alignedDequeue_bits_data_hi_42, alignedDequeue_bits_data_lo_42};
  wire [31:0]   alignedDequeue_bits_data_lo_hi_lo_lo_lo_8 = {alignedDequeue_bits_data_lo_hi_lo_lo_lo_hi_8, alignedDequeue_bits_data_lo_hi_lo_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_lo_lo_hi_lo_8 = {alignedDequeue_bits_data_hi_45, alignedDequeue_bits_data_lo_45, alignedDequeue_bits_data_hi_44, alignedDequeue_bits_data_lo_44};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_lo_lo_hi_hi_8 = {alignedDequeue_bits_data_hi_47, alignedDequeue_bits_data_lo_47, alignedDequeue_bits_data_hi_46, alignedDequeue_bits_data_lo_46};
  wire [31:0]   alignedDequeue_bits_data_lo_hi_lo_lo_hi_8 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_hi_8, alignedDequeue_bits_data_lo_hi_lo_lo_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_lo_hi_lo_lo_8 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_8, alignedDequeue_bits_data_lo_hi_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_lo_hi_lo_lo_8 = {alignedDequeue_bits_data_hi_49, alignedDequeue_bits_data_lo_49, alignedDequeue_bits_data_hi_48, alignedDequeue_bits_data_lo_48};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_lo_hi_lo_hi_8 = {alignedDequeue_bits_data_hi_51, alignedDequeue_bits_data_lo_51, alignedDequeue_bits_data_hi_50, alignedDequeue_bits_data_lo_50};
  wire [31:0]   alignedDequeue_bits_data_lo_hi_lo_hi_lo_8 = {alignedDequeue_bits_data_lo_hi_lo_hi_lo_hi_8, alignedDequeue_bits_data_lo_hi_lo_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_lo_hi_hi_lo_8 = {alignedDequeue_bits_data_hi_53, alignedDequeue_bits_data_lo_53, alignedDequeue_bits_data_hi_52, alignedDequeue_bits_data_lo_52};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_lo_hi_hi_hi_8 = {alignedDequeue_bits_data_hi_55, alignedDequeue_bits_data_lo_55, alignedDequeue_bits_data_hi_54, alignedDequeue_bits_data_lo_54};
  wire [31:0]   alignedDequeue_bits_data_lo_hi_lo_hi_hi_8 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_hi_8, alignedDequeue_bits_data_lo_hi_lo_hi_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_lo_hi_lo_hi_8 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_8, alignedDequeue_bits_data_lo_hi_lo_hi_lo_8};
  wire [127:0]  alignedDequeue_bits_data_lo_hi_lo_8 = {alignedDequeue_bits_data_lo_hi_lo_hi_8, alignedDequeue_bits_data_lo_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_hi_lo_lo_lo_8 = {alignedDequeue_bits_data_hi_57, alignedDequeue_bits_data_lo_57, alignedDequeue_bits_data_hi_56, alignedDequeue_bits_data_lo_56};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_hi_lo_lo_hi_8 = {alignedDequeue_bits_data_hi_59, alignedDequeue_bits_data_lo_59, alignedDequeue_bits_data_hi_58, alignedDequeue_bits_data_lo_58};
  wire [31:0]   alignedDequeue_bits_data_lo_hi_hi_lo_lo_8 = {alignedDequeue_bits_data_lo_hi_hi_lo_lo_hi_8, alignedDequeue_bits_data_lo_hi_hi_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_hi_lo_hi_lo_8 = {alignedDequeue_bits_data_hi_61, alignedDequeue_bits_data_lo_61, alignedDequeue_bits_data_hi_60, alignedDequeue_bits_data_lo_60};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_hi_lo_hi_hi_8 = {alignedDequeue_bits_data_hi_63, alignedDequeue_bits_data_lo_63, alignedDequeue_bits_data_hi_62, alignedDequeue_bits_data_lo_62};
  wire [31:0]   alignedDequeue_bits_data_lo_hi_hi_lo_hi_8 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_hi_8, alignedDequeue_bits_data_lo_hi_hi_lo_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_lo_hi_hi_lo_8 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_8, alignedDequeue_bits_data_lo_hi_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_hi_hi_lo_lo_8 = {alignedDequeue_bits_data_hi_65, alignedDequeue_bits_data_lo_65, alignedDequeue_bits_data_hi_64, alignedDequeue_bits_data_lo_64};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_hi_hi_lo_hi_8 = {alignedDequeue_bits_data_hi_67, alignedDequeue_bits_data_lo_67, alignedDequeue_bits_data_hi_66, alignedDequeue_bits_data_lo_66};
  wire [31:0]   alignedDequeue_bits_data_lo_hi_hi_hi_lo_8 = {alignedDequeue_bits_data_lo_hi_hi_hi_lo_hi_8, alignedDequeue_bits_data_lo_hi_hi_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_hi_hi_hi_lo_8 = {alignedDequeue_bits_data_hi_69, alignedDequeue_bits_data_lo_69, alignedDequeue_bits_data_hi_68, alignedDequeue_bits_data_lo_68};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_hi_hi_hi_hi_8 = {alignedDequeue_bits_data_hi_71, alignedDequeue_bits_data_lo_71, alignedDequeue_bits_data_hi_70, alignedDequeue_bits_data_lo_70};
  wire [31:0]   alignedDequeue_bits_data_lo_hi_hi_hi_hi_8 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_hi_8, alignedDequeue_bits_data_lo_hi_hi_hi_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_lo_hi_hi_hi_8 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_8, alignedDequeue_bits_data_lo_hi_hi_hi_lo_8};
  wire [127:0]  alignedDequeue_bits_data_lo_hi_hi_8 = {alignedDequeue_bits_data_lo_hi_hi_hi_8, alignedDequeue_bits_data_lo_hi_hi_lo_8};
  wire [255:0]  alignedDequeue_bits_data_lo_hi_136 = {alignedDequeue_bits_data_lo_hi_hi_8, alignedDequeue_bits_data_lo_hi_lo_8};
  assign alignedDequeue_bits_data_lo_136 = {alignedDequeue_bits_data_lo_hi_136, alignedDequeue_bits_data_lo_lo_136};
  wire [511:0]  alignedDequeue_bits_data = alignedDequeue_bits_data_lo_136;
  wire [15:0]   alignedDequeue_bits_data_hi_lo_lo_lo_lo_lo_8 = {alignedDequeue_bits_data_hi_73, alignedDequeue_bits_data_lo_73, alignedDequeue_bits_data_hi_72, alignedDequeue_bits_data_lo_72};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_lo_lo_lo_hi_8 = {alignedDequeue_bits_data_hi_75, alignedDequeue_bits_data_lo_75, alignedDequeue_bits_data_hi_74, alignedDequeue_bits_data_lo_74};
  wire [31:0]   alignedDequeue_bits_data_hi_lo_lo_lo_lo_8 = {alignedDequeue_bits_data_hi_lo_lo_lo_lo_hi_8, alignedDequeue_bits_data_hi_lo_lo_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_lo_lo_hi_lo_8 = {alignedDequeue_bits_data_hi_77, alignedDequeue_bits_data_lo_77, alignedDequeue_bits_data_hi_76, alignedDequeue_bits_data_lo_76};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_lo_lo_hi_hi_8 = {alignedDequeue_bits_data_hi_79, alignedDequeue_bits_data_lo_79, alignedDequeue_bits_data_hi_78, alignedDequeue_bits_data_lo_78};
  wire [31:0]   alignedDequeue_bits_data_hi_lo_lo_lo_hi_8 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_hi_8, alignedDequeue_bits_data_hi_lo_lo_lo_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_hi_lo_lo_lo_8 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_8, alignedDequeue_bits_data_hi_lo_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_lo_hi_lo_lo_8 = {alignedDequeue_bits_data_hi_81, alignedDequeue_bits_data_lo_81, alignedDequeue_bits_data_hi_80, alignedDequeue_bits_data_lo_80};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_lo_hi_lo_hi_8 = {alignedDequeue_bits_data_hi_83, alignedDequeue_bits_data_lo_83, alignedDequeue_bits_data_hi_82, alignedDequeue_bits_data_lo_82};
  wire [31:0]   alignedDequeue_bits_data_hi_lo_lo_hi_lo_8 = {alignedDequeue_bits_data_hi_lo_lo_hi_lo_hi_8, alignedDequeue_bits_data_hi_lo_lo_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_lo_hi_hi_lo_8 = {alignedDequeue_bits_data_hi_85, alignedDequeue_bits_data_lo_85, alignedDequeue_bits_data_hi_84, alignedDequeue_bits_data_lo_84};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_lo_hi_hi_hi_8 = {alignedDequeue_bits_data_hi_87, alignedDequeue_bits_data_lo_87, alignedDequeue_bits_data_hi_86, alignedDequeue_bits_data_lo_86};
  wire [31:0]   alignedDequeue_bits_data_hi_lo_lo_hi_hi_8 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_hi_8, alignedDequeue_bits_data_hi_lo_lo_hi_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_hi_lo_lo_hi_8 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_8, alignedDequeue_bits_data_hi_lo_lo_hi_lo_8};
  wire [127:0]  alignedDequeue_bits_data_hi_lo_lo_8 = {alignedDequeue_bits_data_hi_lo_lo_hi_8, alignedDequeue_bits_data_hi_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_hi_lo_lo_lo_8 = {alignedDequeue_bits_data_hi_89, alignedDequeue_bits_data_lo_89, alignedDequeue_bits_data_hi_88, alignedDequeue_bits_data_lo_88};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_hi_lo_lo_hi_8 = {alignedDequeue_bits_data_hi_91, alignedDequeue_bits_data_lo_91, alignedDequeue_bits_data_hi_90, alignedDequeue_bits_data_lo_90};
  wire [31:0]   alignedDequeue_bits_data_hi_lo_hi_lo_lo_8 = {alignedDequeue_bits_data_hi_lo_hi_lo_lo_hi_8, alignedDequeue_bits_data_hi_lo_hi_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_hi_lo_hi_lo_8 = {alignedDequeue_bits_data_hi_93, alignedDequeue_bits_data_lo_93, alignedDequeue_bits_data_hi_92, alignedDequeue_bits_data_lo_92};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_hi_lo_hi_hi_8 = {alignedDequeue_bits_data_hi_95, alignedDequeue_bits_data_lo_95, alignedDequeue_bits_data_hi_94, alignedDequeue_bits_data_lo_94};
  wire [31:0]   alignedDequeue_bits_data_hi_lo_hi_lo_hi_8 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_hi_8, alignedDequeue_bits_data_hi_lo_hi_lo_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_hi_lo_hi_lo_8 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_8, alignedDequeue_bits_data_hi_lo_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_hi_hi_lo_lo_8 = {alignedDequeue_bits_data_hi_97, alignedDequeue_bits_data_lo_97, alignedDequeue_bits_data_hi_96, alignedDequeue_bits_data_lo_96};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_hi_hi_lo_hi_8 = {alignedDequeue_bits_data_hi_99, alignedDequeue_bits_data_lo_99, alignedDequeue_bits_data_hi_98, alignedDequeue_bits_data_lo_98};
  wire [31:0]   alignedDequeue_bits_data_hi_lo_hi_hi_lo_8 = {alignedDequeue_bits_data_hi_lo_hi_hi_lo_hi_8, alignedDequeue_bits_data_hi_lo_hi_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_hi_hi_hi_lo_8 = {alignedDequeue_bits_data_hi_101, alignedDequeue_bits_data_lo_101, alignedDequeue_bits_data_hi_100, alignedDequeue_bits_data_lo_100};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_hi_hi_hi_hi_8 = {alignedDequeue_bits_data_hi_103, alignedDequeue_bits_data_lo_103, alignedDequeue_bits_data_hi_102, alignedDequeue_bits_data_lo_102};
  wire [31:0]   alignedDequeue_bits_data_hi_lo_hi_hi_hi_8 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_hi_8, alignedDequeue_bits_data_hi_lo_hi_hi_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_hi_lo_hi_hi_8 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_8, alignedDequeue_bits_data_hi_lo_hi_hi_lo_8};
  wire [127:0]  alignedDequeue_bits_data_hi_lo_hi_8 = {alignedDequeue_bits_data_hi_lo_hi_hi_8, alignedDequeue_bits_data_hi_lo_hi_lo_8};
  wire [255:0]  alignedDequeue_bits_data_hi_lo_136 = {alignedDequeue_bits_data_hi_lo_hi_8, alignedDequeue_bits_data_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_lo_lo_lo_lo_8 = {alignedDequeue_bits_data_hi_105, alignedDequeue_bits_data_lo_105, alignedDequeue_bits_data_hi_104, alignedDequeue_bits_data_lo_104};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_lo_lo_lo_hi_8 = {alignedDequeue_bits_data_hi_107, alignedDequeue_bits_data_lo_107, alignedDequeue_bits_data_hi_106, alignedDequeue_bits_data_lo_106};
  wire [31:0]   alignedDequeue_bits_data_hi_hi_lo_lo_lo_8 = {alignedDequeue_bits_data_hi_hi_lo_lo_lo_hi_8, alignedDequeue_bits_data_hi_hi_lo_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_lo_lo_hi_lo_8 = {alignedDequeue_bits_data_hi_109, alignedDequeue_bits_data_lo_109, alignedDequeue_bits_data_hi_108, alignedDequeue_bits_data_lo_108};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_lo_lo_hi_hi_8 = {alignedDequeue_bits_data_hi_111, alignedDequeue_bits_data_lo_111, alignedDequeue_bits_data_hi_110, alignedDequeue_bits_data_lo_110};
  wire [31:0]   alignedDequeue_bits_data_hi_hi_lo_lo_hi_8 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_hi_8, alignedDequeue_bits_data_hi_hi_lo_lo_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_hi_hi_lo_lo_8 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_8, alignedDequeue_bits_data_hi_hi_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_lo_hi_lo_lo_8 = {alignedDequeue_bits_data_hi_113, alignedDequeue_bits_data_lo_113, alignedDequeue_bits_data_hi_112, alignedDequeue_bits_data_lo_112};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_lo_hi_lo_hi_8 = {alignedDequeue_bits_data_hi_115, alignedDequeue_bits_data_lo_115, alignedDequeue_bits_data_hi_114, alignedDequeue_bits_data_lo_114};
  wire [31:0]   alignedDequeue_bits_data_hi_hi_lo_hi_lo_8 = {alignedDequeue_bits_data_hi_hi_lo_hi_lo_hi_8, alignedDequeue_bits_data_hi_hi_lo_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_lo_hi_hi_lo_8 = {alignedDequeue_bits_data_hi_117, alignedDequeue_bits_data_lo_117, alignedDequeue_bits_data_hi_116, alignedDequeue_bits_data_lo_116};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_lo_hi_hi_hi_8 = {alignedDequeue_bits_data_hi_119, alignedDequeue_bits_data_lo_119, alignedDequeue_bits_data_hi_118, alignedDequeue_bits_data_lo_118};
  wire [31:0]   alignedDequeue_bits_data_hi_hi_lo_hi_hi_8 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_hi_8, alignedDequeue_bits_data_hi_hi_lo_hi_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_hi_hi_lo_hi_8 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_8, alignedDequeue_bits_data_hi_hi_lo_hi_lo_8};
  wire [127:0]  alignedDequeue_bits_data_hi_hi_lo_8 = {alignedDequeue_bits_data_hi_hi_lo_hi_8, alignedDequeue_bits_data_hi_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_hi_lo_lo_lo_8 = {alignedDequeue_bits_data_hi_121, alignedDequeue_bits_data_lo_121, alignedDequeue_bits_data_hi_120, alignedDequeue_bits_data_lo_120};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_hi_lo_lo_hi_8 = {alignedDequeue_bits_data_hi_123, alignedDequeue_bits_data_lo_123, alignedDequeue_bits_data_hi_122, alignedDequeue_bits_data_lo_122};
  wire [31:0]   alignedDequeue_bits_data_hi_hi_hi_lo_lo_8 = {alignedDequeue_bits_data_hi_hi_hi_lo_lo_hi_8, alignedDequeue_bits_data_hi_hi_hi_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_hi_lo_hi_lo_8 = {alignedDequeue_bits_data_hi_125, alignedDequeue_bits_data_lo_125, alignedDequeue_bits_data_hi_124, alignedDequeue_bits_data_lo_124};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_hi_lo_hi_hi_8 = {alignedDequeue_bits_data_hi_127, alignedDequeue_bits_data_lo_127, alignedDequeue_bits_data_hi_126, alignedDequeue_bits_data_lo_126};
  wire [31:0]   alignedDequeue_bits_data_hi_hi_hi_lo_hi_8 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_hi_8, alignedDequeue_bits_data_hi_hi_hi_lo_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_hi_hi_hi_lo_8 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_8, alignedDequeue_bits_data_hi_hi_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_hi_hi_lo_lo_8 = {alignedDequeue_bits_data_hi_129, alignedDequeue_bits_data_lo_129, alignedDequeue_bits_data_hi_128, alignedDequeue_bits_data_lo_128};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_hi_hi_lo_hi_8 = {alignedDequeue_bits_data_hi_131, alignedDequeue_bits_data_lo_131, alignedDequeue_bits_data_hi_130, alignedDequeue_bits_data_lo_130};
  wire [31:0]   alignedDequeue_bits_data_hi_hi_hi_hi_lo_8 = {alignedDequeue_bits_data_hi_hi_hi_hi_lo_hi_8, alignedDequeue_bits_data_hi_hi_hi_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_hi_hi_hi_lo_8 = {alignedDequeue_bits_data_hi_133, alignedDequeue_bits_data_lo_133, alignedDequeue_bits_data_hi_132, alignedDequeue_bits_data_lo_132};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_hi_hi_hi_hi_8 = {alignedDequeue_bits_data_hi_135, alignedDequeue_bits_data_lo_135, alignedDequeue_bits_data_hi_134, alignedDequeue_bits_data_lo_134};
  wire [31:0]   alignedDequeue_bits_data_hi_hi_hi_hi_hi_8 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_hi_8, alignedDequeue_bits_data_hi_hi_hi_hi_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_hi_hi_hi_hi_8 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_8, alignedDequeue_bits_data_hi_hi_hi_hi_lo_8};
  wire [127:0]  alignedDequeue_bits_data_hi_hi_hi_8 = {alignedDequeue_bits_data_hi_hi_hi_hi_8, alignedDequeue_bits_data_hi_hi_hi_lo_8};
  wire [255:0]  alignedDequeue_bits_data_hi_hi_136 = {alignedDequeue_bits_data_hi_hi_hi_8, alignedDequeue_bits_data_hi_hi_lo_8};
  wire [511:0]  alignedDequeue_bits_data_hi_136 = {alignedDequeue_bits_data_hi_hi_136, alignedDequeue_bits_data_hi_lo_136};
  reg           bufferFull;
  wire          bufferTailFire;
  wire          bufferDequeueValid = bufferFull | bufferTailFire;
  wire          writeStageReady;
  wire          bufferDequeueReady;
  wire          bufferDequeueFire = bufferDequeueReady & bufferDequeueValid;
  assign alignedDequeue_ready = ~bufferFull;
  wire [7:0]    bufferEnqueueSelect = _bufferTailFire_T ? 8'h1 << cacheLineIndexInBuffer : 8'h0;
  wire [511:0]  dataBufferUpdate_0 = bufferEnqueueSelect[0] ? alignedDequeue_bits_data : dataBuffer_0;
  wire [511:0]  dataBufferUpdate_1 = bufferEnqueueSelect[1] ? alignedDequeue_bits_data : dataBuffer_1;
  wire [511:0]  dataBufferUpdate_2 = bufferEnqueueSelect[2] ? alignedDequeue_bits_data : dataBuffer_2;
  wire [511:0]  dataBufferUpdate_3 = bufferEnqueueSelect[3] ? alignedDequeue_bits_data : dataBuffer_3;
  wire [511:0]  dataBufferUpdate_4 = bufferEnqueueSelect[4] ? alignedDequeue_bits_data : dataBuffer_4;
  wire [511:0]  dataBufferUpdate_5 = bufferEnqueueSelect[5] ? alignedDequeue_bits_data : dataBuffer_5;
  wire [511:0]  dataBufferUpdate_6 = bufferEnqueueSelect[6] ? alignedDequeue_bits_data : dataBuffer_6;
  wire [511:0]  dataBufferUpdate_7 = bufferEnqueueSelect[7] ? alignedDequeue_bits_data : dataBuffer_7;
  wire [511:0]  dataSelect_0 = bufferFull ? dataBuffer_0 : dataBufferUpdate_0;
  wire [511:0]  dataSelect_1 = bufferFull ? dataBuffer_1 : dataBufferUpdate_1;
  wire [511:0]  dataSelect_2 = bufferFull ? dataBuffer_2 : dataBufferUpdate_2;
  wire [511:0]  dataSelect_3 = bufferFull ? dataBuffer_3 : dataBufferUpdate_3;
  wire [511:0]  dataSelect_4 = bufferFull ? dataBuffer_4 : dataBufferUpdate_4;
  wire [511:0]  dataSelect_5 = bufferFull ? dataBuffer_5 : dataBufferUpdate_5;
  wire [511:0]  dataSelect_6 = bufferFull ? dataBuffer_6 : dataBufferUpdate_6;
  wire [511:0]  dataSelect_7 = bufferFull ? dataBuffer_7 : dataBufferUpdate_7;
  wire          lastCacheLineForThisGroup = cacheLineIndexInBuffer == lsuRequestReg_instructionInformation_nf;
  wire          lastCacheLineForInst = {7'h0, alignedDequeue_bits_index} == lastWriteVrfIndexReg;
  assign bufferTailFire = _bufferTailFire_T & (lastCacheLineForThisGroup | lastCacheLineForInst);
  reg           waitForFirstDataGroup;
  wire          lastPtr = accessPtr == 3'h0;
  assign writeStageReady = lastPtr & accessStateCheck;
  assign bufferDequeueReady = writeStageReady;
  wire          _maskSelect_valid_output = bufferDequeueFire & isLastDataGroup;
  wire [1023:0] _GEN_5 = {dataSelect_1, dataSelect_0};
  wire [1023:0] dataGroup_lo_lo;
  assign dataGroup_lo_lo = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1;
  assign dataGroup_lo_lo_1 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2;
  assign dataGroup_lo_lo_2 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3;
  assign dataGroup_lo_lo_3 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4;
  assign dataGroup_lo_lo_4 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_5;
  assign dataGroup_lo_lo_5 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_6;
  assign dataGroup_lo_lo_6 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_7;
  assign dataGroup_lo_lo_7 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_8;
  assign dataGroup_lo_lo_8 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_9;
  assign dataGroup_lo_lo_9 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_10;
  assign dataGroup_lo_lo_10 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_11;
  assign dataGroup_lo_lo_11 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_12;
  assign dataGroup_lo_lo_12 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_13;
  assign dataGroup_lo_lo_13 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_14;
  assign dataGroup_lo_lo_14 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_15;
  assign dataGroup_lo_lo_15 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_16;
  assign dataGroup_lo_lo_16 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_17;
  assign dataGroup_lo_lo_17 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_18;
  assign dataGroup_lo_lo_18 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_19;
  assign dataGroup_lo_lo_19 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_20;
  assign dataGroup_lo_lo_20 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_21;
  assign dataGroup_lo_lo_21 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_22;
  assign dataGroup_lo_lo_22 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_23;
  assign dataGroup_lo_lo_23 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_24;
  assign dataGroup_lo_lo_24 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_25;
  assign dataGroup_lo_lo_25 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_26;
  assign dataGroup_lo_lo_26 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_27;
  assign dataGroup_lo_lo_27 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_28;
  assign dataGroup_lo_lo_28 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_29;
  assign dataGroup_lo_lo_29 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_30;
  assign dataGroup_lo_lo_30 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_31;
  assign dataGroup_lo_lo_31 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_32;
  assign dataGroup_lo_lo_32 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_33;
  assign dataGroup_lo_lo_33 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_34;
  assign dataGroup_lo_lo_34 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_35;
  assign dataGroup_lo_lo_35 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_36;
  assign dataGroup_lo_lo_36 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_37;
  assign dataGroup_lo_lo_37 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_38;
  assign dataGroup_lo_lo_38 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_39;
  assign dataGroup_lo_lo_39 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_40;
  assign dataGroup_lo_lo_40 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_41;
  assign dataGroup_lo_lo_41 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_42;
  assign dataGroup_lo_lo_42 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_43;
  assign dataGroup_lo_lo_43 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_44;
  assign dataGroup_lo_lo_44 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_45;
  assign dataGroup_lo_lo_45 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_46;
  assign dataGroup_lo_lo_46 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_47;
  assign dataGroup_lo_lo_47 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_48;
  assign dataGroup_lo_lo_48 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_49;
  assign dataGroup_lo_lo_49 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_50;
  assign dataGroup_lo_lo_50 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_51;
  assign dataGroup_lo_lo_51 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_52;
  assign dataGroup_lo_lo_52 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_53;
  assign dataGroup_lo_lo_53 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_54;
  assign dataGroup_lo_lo_54 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_55;
  assign dataGroup_lo_lo_55 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_56;
  assign dataGroup_lo_lo_56 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_57;
  assign dataGroup_lo_lo_57 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_58;
  assign dataGroup_lo_lo_58 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_59;
  assign dataGroup_lo_lo_59 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_60;
  assign dataGroup_lo_lo_60 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_61;
  assign dataGroup_lo_lo_61 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_62;
  assign dataGroup_lo_lo_62 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_63;
  assign dataGroup_lo_lo_63 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_64;
  assign dataGroup_lo_lo_64 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_65;
  assign dataGroup_lo_lo_65 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_66;
  assign dataGroup_lo_lo_66 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_67;
  assign dataGroup_lo_lo_67 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_68;
  assign dataGroup_lo_lo_68 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_69;
  assign dataGroup_lo_lo_69 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_70;
  assign dataGroup_lo_lo_70 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_71;
  assign dataGroup_lo_lo_71 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_72;
  assign dataGroup_lo_lo_72 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_73;
  assign dataGroup_lo_lo_73 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_74;
  assign dataGroup_lo_lo_74 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_75;
  assign dataGroup_lo_lo_75 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_76;
  assign dataGroup_lo_lo_76 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_77;
  assign dataGroup_lo_lo_77 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_78;
  assign dataGroup_lo_lo_78 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_79;
  assign dataGroup_lo_lo_79 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_80;
  assign dataGroup_lo_lo_80 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_81;
  assign dataGroup_lo_lo_81 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_82;
  assign dataGroup_lo_lo_82 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_83;
  assign dataGroup_lo_lo_83 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_84;
  assign dataGroup_lo_lo_84 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_85;
  assign dataGroup_lo_lo_85 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_86;
  assign dataGroup_lo_lo_86 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_87;
  assign dataGroup_lo_lo_87 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_88;
  assign dataGroup_lo_lo_88 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_89;
  assign dataGroup_lo_lo_89 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_90;
  assign dataGroup_lo_lo_90 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_91;
  assign dataGroup_lo_lo_91 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_92;
  assign dataGroup_lo_lo_92 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_93;
  assign dataGroup_lo_lo_93 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_94;
  assign dataGroup_lo_lo_94 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_95;
  assign dataGroup_lo_lo_95 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_96;
  assign dataGroup_lo_lo_96 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_97;
  assign dataGroup_lo_lo_97 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_98;
  assign dataGroup_lo_lo_98 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_99;
  assign dataGroup_lo_lo_99 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_100;
  assign dataGroup_lo_lo_100 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_101;
  assign dataGroup_lo_lo_101 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_102;
  assign dataGroup_lo_lo_102 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_103;
  assign dataGroup_lo_lo_103 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_104;
  assign dataGroup_lo_lo_104 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_105;
  assign dataGroup_lo_lo_105 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_106;
  assign dataGroup_lo_lo_106 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_107;
  assign dataGroup_lo_lo_107 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_108;
  assign dataGroup_lo_lo_108 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_109;
  assign dataGroup_lo_lo_109 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_110;
  assign dataGroup_lo_lo_110 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_111;
  assign dataGroup_lo_lo_111 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_112;
  assign dataGroup_lo_lo_112 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_113;
  assign dataGroup_lo_lo_113 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_114;
  assign dataGroup_lo_lo_114 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_115;
  assign dataGroup_lo_lo_115 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_116;
  assign dataGroup_lo_lo_116 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_117;
  assign dataGroup_lo_lo_117 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_118;
  assign dataGroup_lo_lo_118 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_119;
  assign dataGroup_lo_lo_119 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_120;
  assign dataGroup_lo_lo_120 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_121;
  assign dataGroup_lo_lo_121 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_122;
  assign dataGroup_lo_lo_122 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_123;
  assign dataGroup_lo_lo_123 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_124;
  assign dataGroup_lo_lo_124 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_125;
  assign dataGroup_lo_lo_125 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_126;
  assign dataGroup_lo_lo_126 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_127;
  assign dataGroup_lo_lo_127 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_128;
  assign dataGroup_lo_lo_128 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_129;
  assign dataGroup_lo_lo_129 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_130;
  assign dataGroup_lo_lo_130 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_131;
  assign dataGroup_lo_lo_131 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_132;
  assign dataGroup_lo_lo_132 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_133;
  assign dataGroup_lo_lo_133 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_134;
  assign dataGroup_lo_lo_134 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_135;
  assign dataGroup_lo_lo_135 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_136;
  assign dataGroup_lo_lo_136 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_137;
  assign dataGroup_lo_lo_137 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_138;
  assign dataGroup_lo_lo_138 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_139;
  assign dataGroup_lo_lo_139 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_140;
  assign dataGroup_lo_lo_140 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_141;
  assign dataGroup_lo_lo_141 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_142;
  assign dataGroup_lo_lo_142 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_143;
  assign dataGroup_lo_lo_143 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_144;
  assign dataGroup_lo_lo_144 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_145;
  assign dataGroup_lo_lo_145 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_146;
  assign dataGroup_lo_lo_146 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_147;
  assign dataGroup_lo_lo_147 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_148;
  assign dataGroup_lo_lo_148 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_149;
  assign dataGroup_lo_lo_149 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_150;
  assign dataGroup_lo_lo_150 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_151;
  assign dataGroup_lo_lo_151 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_152;
  assign dataGroup_lo_lo_152 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_153;
  assign dataGroup_lo_lo_153 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_154;
  assign dataGroup_lo_lo_154 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_155;
  assign dataGroup_lo_lo_155 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_156;
  assign dataGroup_lo_lo_156 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_157;
  assign dataGroup_lo_lo_157 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_158;
  assign dataGroup_lo_lo_158 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_159;
  assign dataGroup_lo_lo_159 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_160;
  assign dataGroup_lo_lo_160 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_161;
  assign dataGroup_lo_lo_161 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_162;
  assign dataGroup_lo_lo_162 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_163;
  assign dataGroup_lo_lo_163 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_164;
  assign dataGroup_lo_lo_164 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_165;
  assign dataGroup_lo_lo_165 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_166;
  assign dataGroup_lo_lo_166 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_167;
  assign dataGroup_lo_lo_167 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_168;
  assign dataGroup_lo_lo_168 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_169;
  assign dataGroup_lo_lo_169 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_170;
  assign dataGroup_lo_lo_170 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_171;
  assign dataGroup_lo_lo_171 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_172;
  assign dataGroup_lo_lo_172 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_173;
  assign dataGroup_lo_lo_173 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_174;
  assign dataGroup_lo_lo_174 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_175;
  assign dataGroup_lo_lo_175 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_176;
  assign dataGroup_lo_lo_176 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_177;
  assign dataGroup_lo_lo_177 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_178;
  assign dataGroup_lo_lo_178 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_179;
  assign dataGroup_lo_lo_179 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_180;
  assign dataGroup_lo_lo_180 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_181;
  assign dataGroup_lo_lo_181 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_182;
  assign dataGroup_lo_lo_182 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_183;
  assign dataGroup_lo_lo_183 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_184;
  assign dataGroup_lo_lo_184 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_185;
  assign dataGroup_lo_lo_185 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_186;
  assign dataGroup_lo_lo_186 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_187;
  assign dataGroup_lo_lo_187 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_188;
  assign dataGroup_lo_lo_188 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_189;
  assign dataGroup_lo_lo_189 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_190;
  assign dataGroup_lo_lo_190 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_191;
  assign dataGroup_lo_lo_191 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_192;
  assign dataGroup_lo_lo_192 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_193;
  assign dataGroup_lo_lo_193 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_194;
  assign dataGroup_lo_lo_194 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_195;
  assign dataGroup_lo_lo_195 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_196;
  assign dataGroup_lo_lo_196 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_197;
  assign dataGroup_lo_lo_197 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_198;
  assign dataGroup_lo_lo_198 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_199;
  assign dataGroup_lo_lo_199 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_200;
  assign dataGroup_lo_lo_200 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_201;
  assign dataGroup_lo_lo_201 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_202;
  assign dataGroup_lo_lo_202 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_203;
  assign dataGroup_lo_lo_203 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_204;
  assign dataGroup_lo_lo_204 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_205;
  assign dataGroup_lo_lo_205 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_206;
  assign dataGroup_lo_lo_206 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_207;
  assign dataGroup_lo_lo_207 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_208;
  assign dataGroup_lo_lo_208 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_209;
  assign dataGroup_lo_lo_209 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_210;
  assign dataGroup_lo_lo_210 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_211;
  assign dataGroup_lo_lo_211 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_212;
  assign dataGroup_lo_lo_212 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_213;
  assign dataGroup_lo_lo_213 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_214;
  assign dataGroup_lo_lo_214 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_215;
  assign dataGroup_lo_lo_215 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_216;
  assign dataGroup_lo_lo_216 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_217;
  assign dataGroup_lo_lo_217 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_218;
  assign dataGroup_lo_lo_218 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_219;
  assign dataGroup_lo_lo_219 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_220;
  assign dataGroup_lo_lo_220 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_221;
  assign dataGroup_lo_lo_221 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_222;
  assign dataGroup_lo_lo_222 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_223;
  assign dataGroup_lo_lo_223 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_224;
  assign dataGroup_lo_lo_224 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_225;
  assign dataGroup_lo_lo_225 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_226;
  assign dataGroup_lo_lo_226 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_227;
  assign dataGroup_lo_lo_227 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_228;
  assign dataGroup_lo_lo_228 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_229;
  assign dataGroup_lo_lo_229 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_230;
  assign dataGroup_lo_lo_230 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_231;
  assign dataGroup_lo_lo_231 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_232;
  assign dataGroup_lo_lo_232 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_233;
  assign dataGroup_lo_lo_233 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_234;
  assign dataGroup_lo_lo_234 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_235;
  assign dataGroup_lo_lo_235 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_236;
  assign dataGroup_lo_lo_236 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_237;
  assign dataGroup_lo_lo_237 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_238;
  assign dataGroup_lo_lo_238 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_239;
  assign dataGroup_lo_lo_239 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_240;
  assign dataGroup_lo_lo_240 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_241;
  assign dataGroup_lo_lo_241 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_242;
  assign dataGroup_lo_lo_242 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_243;
  assign dataGroup_lo_lo_243 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_244;
  assign dataGroup_lo_lo_244 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_245;
  assign dataGroup_lo_lo_245 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_246;
  assign dataGroup_lo_lo_246 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_247;
  assign dataGroup_lo_lo_247 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_248;
  assign dataGroup_lo_lo_248 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_249;
  assign dataGroup_lo_lo_249 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_250;
  assign dataGroup_lo_lo_250 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_251;
  assign dataGroup_lo_lo_251 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_252;
  assign dataGroup_lo_lo_252 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_253;
  assign dataGroup_lo_lo_253 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_254;
  assign dataGroup_lo_lo_254 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_255;
  assign dataGroup_lo_lo_255 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_256;
  assign dataGroup_lo_lo_256 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_257;
  assign dataGroup_lo_lo_257 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_258;
  assign dataGroup_lo_lo_258 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_259;
  assign dataGroup_lo_lo_259 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_260;
  assign dataGroup_lo_lo_260 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_261;
  assign dataGroup_lo_lo_261 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_262;
  assign dataGroup_lo_lo_262 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_263;
  assign dataGroup_lo_lo_263 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_264;
  assign dataGroup_lo_lo_264 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_265;
  assign dataGroup_lo_lo_265 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_266;
  assign dataGroup_lo_lo_266 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_267;
  assign dataGroup_lo_lo_267 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_268;
  assign dataGroup_lo_lo_268 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_269;
  assign dataGroup_lo_lo_269 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_270;
  assign dataGroup_lo_lo_270 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_271;
  assign dataGroup_lo_lo_271 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_272;
  assign dataGroup_lo_lo_272 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_273;
  assign dataGroup_lo_lo_273 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_274;
  assign dataGroup_lo_lo_274 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_275;
  assign dataGroup_lo_lo_275 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_276;
  assign dataGroup_lo_lo_276 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_277;
  assign dataGroup_lo_lo_277 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_278;
  assign dataGroup_lo_lo_278 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_279;
  assign dataGroup_lo_lo_279 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_280;
  assign dataGroup_lo_lo_280 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_281;
  assign dataGroup_lo_lo_281 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_282;
  assign dataGroup_lo_lo_282 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_283;
  assign dataGroup_lo_lo_283 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_284;
  assign dataGroup_lo_lo_284 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_285;
  assign dataGroup_lo_lo_285 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_286;
  assign dataGroup_lo_lo_286 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_287;
  assign dataGroup_lo_lo_287 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_288;
  assign dataGroup_lo_lo_288 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_289;
  assign dataGroup_lo_lo_289 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_290;
  assign dataGroup_lo_lo_290 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_291;
  assign dataGroup_lo_lo_291 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_292;
  assign dataGroup_lo_lo_292 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_293;
  assign dataGroup_lo_lo_293 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_294;
  assign dataGroup_lo_lo_294 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_295;
  assign dataGroup_lo_lo_295 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_296;
  assign dataGroup_lo_lo_296 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_297;
  assign dataGroup_lo_lo_297 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_298;
  assign dataGroup_lo_lo_298 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_299;
  assign dataGroup_lo_lo_299 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_300;
  assign dataGroup_lo_lo_300 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_301;
  assign dataGroup_lo_lo_301 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_302;
  assign dataGroup_lo_lo_302 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_303;
  assign dataGroup_lo_lo_303 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_304;
  assign dataGroup_lo_lo_304 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_305;
  assign dataGroup_lo_lo_305 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_306;
  assign dataGroup_lo_lo_306 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_307;
  assign dataGroup_lo_lo_307 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_308;
  assign dataGroup_lo_lo_308 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_309;
  assign dataGroup_lo_lo_309 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_310;
  assign dataGroup_lo_lo_310 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_311;
  assign dataGroup_lo_lo_311 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_312;
  assign dataGroup_lo_lo_312 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_313;
  assign dataGroup_lo_lo_313 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_314;
  assign dataGroup_lo_lo_314 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_315;
  assign dataGroup_lo_lo_315 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_316;
  assign dataGroup_lo_lo_316 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_317;
  assign dataGroup_lo_lo_317 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_318;
  assign dataGroup_lo_lo_318 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_319;
  assign dataGroup_lo_lo_319 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_320;
  assign dataGroup_lo_lo_320 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_321;
  assign dataGroup_lo_lo_321 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_322;
  assign dataGroup_lo_lo_322 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_323;
  assign dataGroup_lo_lo_323 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_324;
  assign dataGroup_lo_lo_324 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_325;
  assign dataGroup_lo_lo_325 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_326;
  assign dataGroup_lo_lo_326 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_327;
  assign dataGroup_lo_lo_327 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_328;
  assign dataGroup_lo_lo_328 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_329;
  assign dataGroup_lo_lo_329 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_330;
  assign dataGroup_lo_lo_330 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_331;
  assign dataGroup_lo_lo_331 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_332;
  assign dataGroup_lo_lo_332 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_333;
  assign dataGroup_lo_lo_333 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_334;
  assign dataGroup_lo_lo_334 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_335;
  assign dataGroup_lo_lo_335 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_336;
  assign dataGroup_lo_lo_336 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_337;
  assign dataGroup_lo_lo_337 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_338;
  assign dataGroup_lo_lo_338 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_339;
  assign dataGroup_lo_lo_339 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_340;
  assign dataGroup_lo_lo_340 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_341;
  assign dataGroup_lo_lo_341 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_342;
  assign dataGroup_lo_lo_342 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_343;
  assign dataGroup_lo_lo_343 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_344;
  assign dataGroup_lo_lo_344 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_345;
  assign dataGroup_lo_lo_345 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_346;
  assign dataGroup_lo_lo_346 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_347;
  assign dataGroup_lo_lo_347 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_348;
  assign dataGroup_lo_lo_348 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_349;
  assign dataGroup_lo_lo_349 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_350;
  assign dataGroup_lo_lo_350 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_351;
  assign dataGroup_lo_lo_351 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_352;
  assign dataGroup_lo_lo_352 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_353;
  assign dataGroup_lo_lo_353 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_354;
  assign dataGroup_lo_lo_354 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_355;
  assign dataGroup_lo_lo_355 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_356;
  assign dataGroup_lo_lo_356 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_357;
  assign dataGroup_lo_lo_357 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_358;
  assign dataGroup_lo_lo_358 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_359;
  assign dataGroup_lo_lo_359 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_360;
  assign dataGroup_lo_lo_360 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_361;
  assign dataGroup_lo_lo_361 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_362;
  assign dataGroup_lo_lo_362 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_363;
  assign dataGroup_lo_lo_363 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_364;
  assign dataGroup_lo_lo_364 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_365;
  assign dataGroup_lo_lo_365 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_366;
  assign dataGroup_lo_lo_366 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_367;
  assign dataGroup_lo_lo_367 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_368;
  assign dataGroup_lo_lo_368 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_369;
  assign dataGroup_lo_lo_369 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_370;
  assign dataGroup_lo_lo_370 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_371;
  assign dataGroup_lo_lo_371 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_372;
  assign dataGroup_lo_lo_372 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_373;
  assign dataGroup_lo_lo_373 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_374;
  assign dataGroup_lo_lo_374 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_375;
  assign dataGroup_lo_lo_375 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_376;
  assign dataGroup_lo_lo_376 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_377;
  assign dataGroup_lo_lo_377 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_378;
  assign dataGroup_lo_lo_378 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_379;
  assign dataGroup_lo_lo_379 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_380;
  assign dataGroup_lo_lo_380 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_381;
  assign dataGroup_lo_lo_381 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_382;
  assign dataGroup_lo_lo_382 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_383;
  assign dataGroup_lo_lo_383 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_384;
  assign dataGroup_lo_lo_384 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_385;
  assign dataGroup_lo_lo_385 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_386;
  assign dataGroup_lo_lo_386 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_387;
  assign dataGroup_lo_lo_387 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_388;
  assign dataGroup_lo_lo_388 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_389;
  assign dataGroup_lo_lo_389 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_390;
  assign dataGroup_lo_lo_390 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_391;
  assign dataGroup_lo_lo_391 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_392;
  assign dataGroup_lo_lo_392 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_393;
  assign dataGroup_lo_lo_393 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_394;
  assign dataGroup_lo_lo_394 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_395;
  assign dataGroup_lo_lo_395 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_396;
  assign dataGroup_lo_lo_396 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_397;
  assign dataGroup_lo_lo_397 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_398;
  assign dataGroup_lo_lo_398 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_399;
  assign dataGroup_lo_lo_399 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_400;
  assign dataGroup_lo_lo_400 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_401;
  assign dataGroup_lo_lo_401 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_402;
  assign dataGroup_lo_lo_402 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_403;
  assign dataGroup_lo_lo_403 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_404;
  assign dataGroup_lo_lo_404 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_405;
  assign dataGroup_lo_lo_405 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_406;
  assign dataGroup_lo_lo_406 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_407;
  assign dataGroup_lo_lo_407 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_408;
  assign dataGroup_lo_lo_408 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_409;
  assign dataGroup_lo_lo_409 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_410;
  assign dataGroup_lo_lo_410 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_411;
  assign dataGroup_lo_lo_411 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_412;
  assign dataGroup_lo_lo_412 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_413;
  assign dataGroup_lo_lo_413 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_414;
  assign dataGroup_lo_lo_414 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_415;
  assign dataGroup_lo_lo_415 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_416;
  assign dataGroup_lo_lo_416 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_417;
  assign dataGroup_lo_lo_417 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_418;
  assign dataGroup_lo_lo_418 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_419;
  assign dataGroup_lo_lo_419 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_420;
  assign dataGroup_lo_lo_420 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_421;
  assign dataGroup_lo_lo_421 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_422;
  assign dataGroup_lo_lo_422 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_423;
  assign dataGroup_lo_lo_423 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_424;
  assign dataGroup_lo_lo_424 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_425;
  assign dataGroup_lo_lo_425 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_426;
  assign dataGroup_lo_lo_426 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_427;
  assign dataGroup_lo_lo_427 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_428;
  assign dataGroup_lo_lo_428 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_429;
  assign dataGroup_lo_lo_429 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_430;
  assign dataGroup_lo_lo_430 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_431;
  assign dataGroup_lo_lo_431 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_432;
  assign dataGroup_lo_lo_432 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_433;
  assign dataGroup_lo_lo_433 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_434;
  assign dataGroup_lo_lo_434 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_435;
  assign dataGroup_lo_lo_435 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_436;
  assign dataGroup_lo_lo_436 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_437;
  assign dataGroup_lo_lo_437 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_438;
  assign dataGroup_lo_lo_438 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_439;
  assign dataGroup_lo_lo_439 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_440;
  assign dataGroup_lo_lo_440 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_441;
  assign dataGroup_lo_lo_441 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_442;
  assign dataGroup_lo_lo_442 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_443;
  assign dataGroup_lo_lo_443 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_444;
  assign dataGroup_lo_lo_444 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_445;
  assign dataGroup_lo_lo_445 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_446;
  assign dataGroup_lo_lo_446 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_447;
  assign dataGroup_lo_lo_447 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_448;
  assign dataGroup_lo_lo_448 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_449;
  assign dataGroup_lo_lo_449 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_450;
  assign dataGroup_lo_lo_450 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_451;
  assign dataGroup_lo_lo_451 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_452;
  assign dataGroup_lo_lo_452 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_453;
  assign dataGroup_lo_lo_453 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_454;
  assign dataGroup_lo_lo_454 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_455;
  assign dataGroup_lo_lo_455 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_456;
  assign dataGroup_lo_lo_456 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_457;
  assign dataGroup_lo_lo_457 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_458;
  assign dataGroup_lo_lo_458 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_459;
  assign dataGroup_lo_lo_459 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_460;
  assign dataGroup_lo_lo_460 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_461;
  assign dataGroup_lo_lo_461 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_462;
  assign dataGroup_lo_lo_462 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_463;
  assign dataGroup_lo_lo_463 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_464;
  assign dataGroup_lo_lo_464 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_465;
  assign dataGroup_lo_lo_465 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_466;
  assign dataGroup_lo_lo_466 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_467;
  assign dataGroup_lo_lo_467 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_468;
  assign dataGroup_lo_lo_468 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_469;
  assign dataGroup_lo_lo_469 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_470;
  assign dataGroup_lo_lo_470 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_471;
  assign dataGroup_lo_lo_471 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_472;
  assign dataGroup_lo_lo_472 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_473;
  assign dataGroup_lo_lo_473 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_474;
  assign dataGroup_lo_lo_474 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_475;
  assign dataGroup_lo_lo_475 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_476;
  assign dataGroup_lo_lo_476 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_477;
  assign dataGroup_lo_lo_477 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_478;
  assign dataGroup_lo_lo_478 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_479;
  assign dataGroup_lo_lo_479 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_480;
  assign dataGroup_lo_lo_480 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_481;
  assign dataGroup_lo_lo_481 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_482;
  assign dataGroup_lo_lo_482 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_483;
  assign dataGroup_lo_lo_483 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_484;
  assign dataGroup_lo_lo_484 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_485;
  assign dataGroup_lo_lo_485 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_486;
  assign dataGroup_lo_lo_486 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_487;
  assign dataGroup_lo_lo_487 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_488;
  assign dataGroup_lo_lo_488 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_489;
  assign dataGroup_lo_lo_489 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_490;
  assign dataGroup_lo_lo_490 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_491;
  assign dataGroup_lo_lo_491 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_492;
  assign dataGroup_lo_lo_492 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_493;
  assign dataGroup_lo_lo_493 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_494;
  assign dataGroup_lo_lo_494 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_495;
  assign dataGroup_lo_lo_495 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_496;
  assign dataGroup_lo_lo_496 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_497;
  assign dataGroup_lo_lo_497 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_498;
  assign dataGroup_lo_lo_498 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_499;
  assign dataGroup_lo_lo_499 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_500;
  assign dataGroup_lo_lo_500 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_501;
  assign dataGroup_lo_lo_501 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_502;
  assign dataGroup_lo_lo_502 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_503;
  assign dataGroup_lo_lo_503 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_504;
  assign dataGroup_lo_lo_504 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_505;
  assign dataGroup_lo_lo_505 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_506;
  assign dataGroup_lo_lo_506 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_507;
  assign dataGroup_lo_lo_507 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_508;
  assign dataGroup_lo_lo_508 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_509;
  assign dataGroup_lo_lo_509 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_510;
  assign dataGroup_lo_lo_510 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_511;
  assign dataGroup_lo_lo_511 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_512;
  assign dataGroup_lo_lo_512 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_513;
  assign dataGroup_lo_lo_513 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_514;
  assign dataGroup_lo_lo_514 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_515;
  assign dataGroup_lo_lo_515 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_516;
  assign dataGroup_lo_lo_516 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_517;
  assign dataGroup_lo_lo_517 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_518;
  assign dataGroup_lo_lo_518 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_519;
  assign dataGroup_lo_lo_519 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_520;
  assign dataGroup_lo_lo_520 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_521;
  assign dataGroup_lo_lo_521 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_522;
  assign dataGroup_lo_lo_522 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_523;
  assign dataGroup_lo_lo_523 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_524;
  assign dataGroup_lo_lo_524 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_525;
  assign dataGroup_lo_lo_525 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_526;
  assign dataGroup_lo_lo_526 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_527;
  assign dataGroup_lo_lo_527 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_528;
  assign dataGroup_lo_lo_528 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_529;
  assign dataGroup_lo_lo_529 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_530;
  assign dataGroup_lo_lo_530 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_531;
  assign dataGroup_lo_lo_531 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_532;
  assign dataGroup_lo_lo_532 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_533;
  assign dataGroup_lo_lo_533 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_534;
  assign dataGroup_lo_lo_534 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_535;
  assign dataGroup_lo_lo_535 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_536;
  assign dataGroup_lo_lo_536 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_537;
  assign dataGroup_lo_lo_537 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_538;
  assign dataGroup_lo_lo_538 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_539;
  assign dataGroup_lo_lo_539 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_540;
  assign dataGroup_lo_lo_540 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_541;
  assign dataGroup_lo_lo_541 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_542;
  assign dataGroup_lo_lo_542 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_543;
  assign dataGroup_lo_lo_543 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_544;
  assign dataGroup_lo_lo_544 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_545;
  assign dataGroup_lo_lo_545 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_546;
  assign dataGroup_lo_lo_546 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_547;
  assign dataGroup_lo_lo_547 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_548;
  assign dataGroup_lo_lo_548 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_549;
  assign dataGroup_lo_lo_549 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_550;
  assign dataGroup_lo_lo_550 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_551;
  assign dataGroup_lo_lo_551 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_552;
  assign dataGroup_lo_lo_552 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_553;
  assign dataGroup_lo_lo_553 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_554;
  assign dataGroup_lo_lo_554 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_555;
  assign dataGroup_lo_lo_555 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_556;
  assign dataGroup_lo_lo_556 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_557;
  assign dataGroup_lo_lo_557 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_558;
  assign dataGroup_lo_lo_558 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_559;
  assign dataGroup_lo_lo_559 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_560;
  assign dataGroup_lo_lo_560 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_561;
  assign dataGroup_lo_lo_561 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_562;
  assign dataGroup_lo_lo_562 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_563;
  assign dataGroup_lo_lo_563 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_564;
  assign dataGroup_lo_lo_564 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_565;
  assign dataGroup_lo_lo_565 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_566;
  assign dataGroup_lo_lo_566 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_567;
  assign dataGroup_lo_lo_567 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_568;
  assign dataGroup_lo_lo_568 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_569;
  assign dataGroup_lo_lo_569 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_570;
  assign dataGroup_lo_lo_570 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_571;
  assign dataGroup_lo_lo_571 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_572;
  assign dataGroup_lo_lo_572 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_573;
  assign dataGroup_lo_lo_573 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_574;
  assign dataGroup_lo_lo_574 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_575;
  assign dataGroup_lo_lo_575 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_576;
  assign dataGroup_lo_lo_576 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_577;
  assign dataGroup_lo_lo_577 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_578;
  assign dataGroup_lo_lo_578 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_579;
  assign dataGroup_lo_lo_579 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_580;
  assign dataGroup_lo_lo_580 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_581;
  assign dataGroup_lo_lo_581 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_582;
  assign dataGroup_lo_lo_582 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_583;
  assign dataGroup_lo_lo_583 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_584;
  assign dataGroup_lo_lo_584 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_585;
  assign dataGroup_lo_lo_585 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_586;
  assign dataGroup_lo_lo_586 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_587;
  assign dataGroup_lo_lo_587 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_588;
  assign dataGroup_lo_lo_588 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_589;
  assign dataGroup_lo_lo_589 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_590;
  assign dataGroup_lo_lo_590 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_591;
  assign dataGroup_lo_lo_591 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_592;
  assign dataGroup_lo_lo_592 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_593;
  assign dataGroup_lo_lo_593 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_594;
  assign dataGroup_lo_lo_594 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_595;
  assign dataGroup_lo_lo_595 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_596;
  assign dataGroup_lo_lo_596 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_597;
  assign dataGroup_lo_lo_597 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_598;
  assign dataGroup_lo_lo_598 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_599;
  assign dataGroup_lo_lo_599 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_600;
  assign dataGroup_lo_lo_600 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_601;
  assign dataGroup_lo_lo_601 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_602;
  assign dataGroup_lo_lo_602 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_603;
  assign dataGroup_lo_lo_603 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_604;
  assign dataGroup_lo_lo_604 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_605;
  assign dataGroup_lo_lo_605 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_606;
  assign dataGroup_lo_lo_606 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_607;
  assign dataGroup_lo_lo_607 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_608;
  assign dataGroup_lo_lo_608 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_609;
  assign dataGroup_lo_lo_609 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_610;
  assign dataGroup_lo_lo_610 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_611;
  assign dataGroup_lo_lo_611 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_612;
  assign dataGroup_lo_lo_612 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_613;
  assign dataGroup_lo_lo_613 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_614;
  assign dataGroup_lo_lo_614 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_615;
  assign dataGroup_lo_lo_615 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_616;
  assign dataGroup_lo_lo_616 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_617;
  assign dataGroup_lo_lo_617 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_618;
  assign dataGroup_lo_lo_618 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_619;
  assign dataGroup_lo_lo_619 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_620;
  assign dataGroup_lo_lo_620 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_621;
  assign dataGroup_lo_lo_621 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_622;
  assign dataGroup_lo_lo_622 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_623;
  assign dataGroup_lo_lo_623 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_624;
  assign dataGroup_lo_lo_624 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_625;
  assign dataGroup_lo_lo_625 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_626;
  assign dataGroup_lo_lo_626 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_627;
  assign dataGroup_lo_lo_627 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_628;
  assign dataGroup_lo_lo_628 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_629;
  assign dataGroup_lo_lo_629 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_630;
  assign dataGroup_lo_lo_630 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_631;
  assign dataGroup_lo_lo_631 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_632;
  assign dataGroup_lo_lo_632 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_633;
  assign dataGroup_lo_lo_633 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_634;
  assign dataGroup_lo_lo_634 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_635;
  assign dataGroup_lo_lo_635 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_636;
  assign dataGroup_lo_lo_636 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_637;
  assign dataGroup_lo_lo_637 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_638;
  assign dataGroup_lo_lo_638 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_639;
  assign dataGroup_lo_lo_639 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_640;
  assign dataGroup_lo_lo_640 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_641;
  assign dataGroup_lo_lo_641 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_642;
  assign dataGroup_lo_lo_642 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_643;
  assign dataGroup_lo_lo_643 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_644;
  assign dataGroup_lo_lo_644 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_645;
  assign dataGroup_lo_lo_645 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_646;
  assign dataGroup_lo_lo_646 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_647;
  assign dataGroup_lo_lo_647 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_648;
  assign dataGroup_lo_lo_648 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_649;
  assign dataGroup_lo_lo_649 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_650;
  assign dataGroup_lo_lo_650 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_651;
  assign dataGroup_lo_lo_651 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_652;
  assign dataGroup_lo_lo_652 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_653;
  assign dataGroup_lo_lo_653 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_654;
  assign dataGroup_lo_lo_654 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_655;
  assign dataGroup_lo_lo_655 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_656;
  assign dataGroup_lo_lo_656 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_657;
  assign dataGroup_lo_lo_657 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_658;
  assign dataGroup_lo_lo_658 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_659;
  assign dataGroup_lo_lo_659 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_660;
  assign dataGroup_lo_lo_660 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_661;
  assign dataGroup_lo_lo_661 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_662;
  assign dataGroup_lo_lo_662 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_663;
  assign dataGroup_lo_lo_663 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_664;
  assign dataGroup_lo_lo_664 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_665;
  assign dataGroup_lo_lo_665 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_666;
  assign dataGroup_lo_lo_666 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_667;
  assign dataGroup_lo_lo_667 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_668;
  assign dataGroup_lo_lo_668 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_669;
  assign dataGroup_lo_lo_669 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_670;
  assign dataGroup_lo_lo_670 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_671;
  assign dataGroup_lo_lo_671 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_672;
  assign dataGroup_lo_lo_672 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_673;
  assign dataGroup_lo_lo_673 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_674;
  assign dataGroup_lo_lo_674 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_675;
  assign dataGroup_lo_lo_675 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_676;
  assign dataGroup_lo_lo_676 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_677;
  assign dataGroup_lo_lo_677 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_678;
  assign dataGroup_lo_lo_678 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_679;
  assign dataGroup_lo_lo_679 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_680;
  assign dataGroup_lo_lo_680 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_681;
  assign dataGroup_lo_lo_681 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_682;
  assign dataGroup_lo_lo_682 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_683;
  assign dataGroup_lo_lo_683 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_684;
  assign dataGroup_lo_lo_684 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_685;
  assign dataGroup_lo_lo_685 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_686;
  assign dataGroup_lo_lo_686 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_687;
  assign dataGroup_lo_lo_687 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_688;
  assign dataGroup_lo_lo_688 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_689;
  assign dataGroup_lo_lo_689 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_690;
  assign dataGroup_lo_lo_690 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_691;
  assign dataGroup_lo_lo_691 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_692;
  assign dataGroup_lo_lo_692 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_693;
  assign dataGroup_lo_lo_693 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_694;
  assign dataGroup_lo_lo_694 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_695;
  assign dataGroup_lo_lo_695 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_696;
  assign dataGroup_lo_lo_696 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_697;
  assign dataGroup_lo_lo_697 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_698;
  assign dataGroup_lo_lo_698 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_699;
  assign dataGroup_lo_lo_699 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_700;
  assign dataGroup_lo_lo_700 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_701;
  assign dataGroup_lo_lo_701 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_702;
  assign dataGroup_lo_lo_702 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_703;
  assign dataGroup_lo_lo_703 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_704;
  assign dataGroup_lo_lo_704 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_705;
  assign dataGroup_lo_lo_705 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_706;
  assign dataGroup_lo_lo_706 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_707;
  assign dataGroup_lo_lo_707 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_708;
  assign dataGroup_lo_lo_708 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_709;
  assign dataGroup_lo_lo_709 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_710;
  assign dataGroup_lo_lo_710 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_711;
  assign dataGroup_lo_lo_711 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_712;
  assign dataGroup_lo_lo_712 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_713;
  assign dataGroup_lo_lo_713 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_714;
  assign dataGroup_lo_lo_714 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_715;
  assign dataGroup_lo_lo_715 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_716;
  assign dataGroup_lo_lo_716 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_717;
  assign dataGroup_lo_lo_717 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_718;
  assign dataGroup_lo_lo_718 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_719;
  assign dataGroup_lo_lo_719 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_720;
  assign dataGroup_lo_lo_720 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_721;
  assign dataGroup_lo_lo_721 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_722;
  assign dataGroup_lo_lo_722 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_723;
  assign dataGroup_lo_lo_723 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_724;
  assign dataGroup_lo_lo_724 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_725;
  assign dataGroup_lo_lo_725 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_726;
  assign dataGroup_lo_lo_726 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_727;
  assign dataGroup_lo_lo_727 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_728;
  assign dataGroup_lo_lo_728 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_729;
  assign dataGroup_lo_lo_729 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_730;
  assign dataGroup_lo_lo_730 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_731;
  assign dataGroup_lo_lo_731 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_732;
  assign dataGroup_lo_lo_732 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_733;
  assign dataGroup_lo_lo_733 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_734;
  assign dataGroup_lo_lo_734 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_735;
  assign dataGroup_lo_lo_735 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_736;
  assign dataGroup_lo_lo_736 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_737;
  assign dataGroup_lo_lo_737 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_738;
  assign dataGroup_lo_lo_738 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_739;
  assign dataGroup_lo_lo_739 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_740;
  assign dataGroup_lo_lo_740 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_741;
  assign dataGroup_lo_lo_741 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_742;
  assign dataGroup_lo_lo_742 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_743;
  assign dataGroup_lo_lo_743 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_744;
  assign dataGroup_lo_lo_744 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_745;
  assign dataGroup_lo_lo_745 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_746;
  assign dataGroup_lo_lo_746 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_747;
  assign dataGroup_lo_lo_747 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_748;
  assign dataGroup_lo_lo_748 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_749;
  assign dataGroup_lo_lo_749 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_750;
  assign dataGroup_lo_lo_750 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_751;
  assign dataGroup_lo_lo_751 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_752;
  assign dataGroup_lo_lo_752 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_753;
  assign dataGroup_lo_lo_753 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_754;
  assign dataGroup_lo_lo_754 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_755;
  assign dataGroup_lo_lo_755 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_756;
  assign dataGroup_lo_lo_756 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_757;
  assign dataGroup_lo_lo_757 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_758;
  assign dataGroup_lo_lo_758 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_759;
  assign dataGroup_lo_lo_759 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_760;
  assign dataGroup_lo_lo_760 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_761;
  assign dataGroup_lo_lo_761 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_762;
  assign dataGroup_lo_lo_762 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_763;
  assign dataGroup_lo_lo_763 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_764;
  assign dataGroup_lo_lo_764 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_765;
  assign dataGroup_lo_lo_765 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_766;
  assign dataGroup_lo_lo_766 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_767;
  assign dataGroup_lo_lo_767 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_768;
  assign dataGroup_lo_lo_768 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_769;
  assign dataGroup_lo_lo_769 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_770;
  assign dataGroup_lo_lo_770 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_771;
  assign dataGroup_lo_lo_771 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_772;
  assign dataGroup_lo_lo_772 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_773;
  assign dataGroup_lo_lo_773 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_774;
  assign dataGroup_lo_lo_774 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_775;
  assign dataGroup_lo_lo_775 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_776;
  assign dataGroup_lo_lo_776 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_777;
  assign dataGroup_lo_lo_777 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_778;
  assign dataGroup_lo_lo_778 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_779;
  assign dataGroup_lo_lo_779 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_780;
  assign dataGroup_lo_lo_780 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_781;
  assign dataGroup_lo_lo_781 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_782;
  assign dataGroup_lo_lo_782 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_783;
  assign dataGroup_lo_lo_783 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_784;
  assign dataGroup_lo_lo_784 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_785;
  assign dataGroup_lo_lo_785 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_786;
  assign dataGroup_lo_lo_786 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_787;
  assign dataGroup_lo_lo_787 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_788;
  assign dataGroup_lo_lo_788 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_789;
  assign dataGroup_lo_lo_789 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_790;
  assign dataGroup_lo_lo_790 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_791;
  assign dataGroup_lo_lo_791 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_792;
  assign dataGroup_lo_lo_792 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_793;
  assign dataGroup_lo_lo_793 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_794;
  assign dataGroup_lo_lo_794 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_795;
  assign dataGroup_lo_lo_795 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_796;
  assign dataGroup_lo_lo_796 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_797;
  assign dataGroup_lo_lo_797 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_798;
  assign dataGroup_lo_lo_798 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_799;
  assign dataGroup_lo_lo_799 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_800;
  assign dataGroup_lo_lo_800 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_801;
  assign dataGroup_lo_lo_801 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_802;
  assign dataGroup_lo_lo_802 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_803;
  assign dataGroup_lo_lo_803 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_804;
  assign dataGroup_lo_lo_804 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_805;
  assign dataGroup_lo_lo_805 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_806;
  assign dataGroup_lo_lo_806 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_807;
  assign dataGroup_lo_lo_807 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_808;
  assign dataGroup_lo_lo_808 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_809;
  assign dataGroup_lo_lo_809 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_810;
  assign dataGroup_lo_lo_810 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_811;
  assign dataGroup_lo_lo_811 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_812;
  assign dataGroup_lo_lo_812 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_813;
  assign dataGroup_lo_lo_813 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_814;
  assign dataGroup_lo_lo_814 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_815;
  assign dataGroup_lo_lo_815 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_816;
  assign dataGroup_lo_lo_816 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_817;
  assign dataGroup_lo_lo_817 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_818;
  assign dataGroup_lo_lo_818 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_819;
  assign dataGroup_lo_lo_819 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_820;
  assign dataGroup_lo_lo_820 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_821;
  assign dataGroup_lo_lo_821 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_822;
  assign dataGroup_lo_lo_822 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_823;
  assign dataGroup_lo_lo_823 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_824;
  assign dataGroup_lo_lo_824 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_825;
  assign dataGroup_lo_lo_825 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_826;
  assign dataGroup_lo_lo_826 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_827;
  assign dataGroup_lo_lo_827 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_828;
  assign dataGroup_lo_lo_828 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_829;
  assign dataGroup_lo_lo_829 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_830;
  assign dataGroup_lo_lo_830 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_831;
  assign dataGroup_lo_lo_831 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_832;
  assign dataGroup_lo_lo_832 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_833;
  assign dataGroup_lo_lo_833 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_834;
  assign dataGroup_lo_lo_834 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_835;
  assign dataGroup_lo_lo_835 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_836;
  assign dataGroup_lo_lo_836 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_837;
  assign dataGroup_lo_lo_837 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_838;
  assign dataGroup_lo_lo_838 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_839;
  assign dataGroup_lo_lo_839 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_840;
  assign dataGroup_lo_lo_840 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_841;
  assign dataGroup_lo_lo_841 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_842;
  assign dataGroup_lo_lo_842 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_843;
  assign dataGroup_lo_lo_843 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_844;
  assign dataGroup_lo_lo_844 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_845;
  assign dataGroup_lo_lo_845 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_846;
  assign dataGroup_lo_lo_846 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_847;
  assign dataGroup_lo_lo_847 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_848;
  assign dataGroup_lo_lo_848 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_849;
  assign dataGroup_lo_lo_849 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_850;
  assign dataGroup_lo_lo_850 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_851;
  assign dataGroup_lo_lo_851 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_852;
  assign dataGroup_lo_lo_852 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_853;
  assign dataGroup_lo_lo_853 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_854;
  assign dataGroup_lo_lo_854 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_855;
  assign dataGroup_lo_lo_855 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_856;
  assign dataGroup_lo_lo_856 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_857;
  assign dataGroup_lo_lo_857 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_858;
  assign dataGroup_lo_lo_858 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_859;
  assign dataGroup_lo_lo_859 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_860;
  assign dataGroup_lo_lo_860 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_861;
  assign dataGroup_lo_lo_861 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_862;
  assign dataGroup_lo_lo_862 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_863;
  assign dataGroup_lo_lo_863 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_864;
  assign dataGroup_lo_lo_864 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_865;
  assign dataGroup_lo_lo_865 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_866;
  assign dataGroup_lo_lo_866 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_867;
  assign dataGroup_lo_lo_867 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_868;
  assign dataGroup_lo_lo_868 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_869;
  assign dataGroup_lo_lo_869 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_870;
  assign dataGroup_lo_lo_870 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_871;
  assign dataGroup_lo_lo_871 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_872;
  assign dataGroup_lo_lo_872 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_873;
  assign dataGroup_lo_lo_873 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_874;
  assign dataGroup_lo_lo_874 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_875;
  assign dataGroup_lo_lo_875 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_876;
  assign dataGroup_lo_lo_876 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_877;
  assign dataGroup_lo_lo_877 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_878;
  assign dataGroup_lo_lo_878 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_879;
  assign dataGroup_lo_lo_879 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_880;
  assign dataGroup_lo_lo_880 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_881;
  assign dataGroup_lo_lo_881 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_882;
  assign dataGroup_lo_lo_882 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_883;
  assign dataGroup_lo_lo_883 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_884;
  assign dataGroup_lo_lo_884 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_885;
  assign dataGroup_lo_lo_885 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_886;
  assign dataGroup_lo_lo_886 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_887;
  assign dataGroup_lo_lo_887 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_888;
  assign dataGroup_lo_lo_888 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_889;
  assign dataGroup_lo_lo_889 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_890;
  assign dataGroup_lo_lo_890 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_891;
  assign dataGroup_lo_lo_891 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_892;
  assign dataGroup_lo_lo_892 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_893;
  assign dataGroup_lo_lo_893 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_894;
  assign dataGroup_lo_lo_894 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_895;
  assign dataGroup_lo_lo_895 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_896;
  assign dataGroup_lo_lo_896 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_897;
  assign dataGroup_lo_lo_897 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_898;
  assign dataGroup_lo_lo_898 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_899;
  assign dataGroup_lo_lo_899 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_900;
  assign dataGroup_lo_lo_900 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_901;
  assign dataGroup_lo_lo_901 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_902;
  assign dataGroup_lo_lo_902 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_903;
  assign dataGroup_lo_lo_903 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_904;
  assign dataGroup_lo_lo_904 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_905;
  assign dataGroup_lo_lo_905 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_906;
  assign dataGroup_lo_lo_906 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_907;
  assign dataGroup_lo_lo_907 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_908;
  assign dataGroup_lo_lo_908 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_909;
  assign dataGroup_lo_lo_909 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_910;
  assign dataGroup_lo_lo_910 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_911;
  assign dataGroup_lo_lo_911 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_912;
  assign dataGroup_lo_lo_912 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_913;
  assign dataGroup_lo_lo_913 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_914;
  assign dataGroup_lo_lo_914 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_915;
  assign dataGroup_lo_lo_915 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_916;
  assign dataGroup_lo_lo_916 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_917;
  assign dataGroup_lo_lo_917 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_918;
  assign dataGroup_lo_lo_918 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_919;
  assign dataGroup_lo_lo_919 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_920;
  assign dataGroup_lo_lo_920 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_921;
  assign dataGroup_lo_lo_921 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_922;
  assign dataGroup_lo_lo_922 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_923;
  assign dataGroup_lo_lo_923 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_924;
  assign dataGroup_lo_lo_924 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_925;
  assign dataGroup_lo_lo_925 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_926;
  assign dataGroup_lo_lo_926 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_927;
  assign dataGroup_lo_lo_927 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_928;
  assign dataGroup_lo_lo_928 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_929;
  assign dataGroup_lo_lo_929 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_930;
  assign dataGroup_lo_lo_930 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_931;
  assign dataGroup_lo_lo_931 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_932;
  assign dataGroup_lo_lo_932 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_933;
  assign dataGroup_lo_lo_933 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_934;
  assign dataGroup_lo_lo_934 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_935;
  assign dataGroup_lo_lo_935 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_936;
  assign dataGroup_lo_lo_936 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_937;
  assign dataGroup_lo_lo_937 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_938;
  assign dataGroup_lo_lo_938 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_939;
  assign dataGroup_lo_lo_939 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_940;
  assign dataGroup_lo_lo_940 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_941;
  assign dataGroup_lo_lo_941 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_942;
  assign dataGroup_lo_lo_942 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_943;
  assign dataGroup_lo_lo_943 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_944;
  assign dataGroup_lo_lo_944 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_945;
  assign dataGroup_lo_lo_945 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_946;
  assign dataGroup_lo_lo_946 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_947;
  assign dataGroup_lo_lo_947 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_948;
  assign dataGroup_lo_lo_948 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_949;
  assign dataGroup_lo_lo_949 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_950;
  assign dataGroup_lo_lo_950 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_951;
  assign dataGroup_lo_lo_951 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_952;
  assign dataGroup_lo_lo_952 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_953;
  assign dataGroup_lo_lo_953 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_954;
  assign dataGroup_lo_lo_954 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_955;
  assign dataGroup_lo_lo_955 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_956;
  assign dataGroup_lo_lo_956 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_957;
  assign dataGroup_lo_lo_957 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_958;
  assign dataGroup_lo_lo_958 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_959;
  assign dataGroup_lo_lo_959 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_960;
  assign dataGroup_lo_lo_960 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_961;
  assign dataGroup_lo_lo_961 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_962;
  assign dataGroup_lo_lo_962 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_963;
  assign dataGroup_lo_lo_963 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_964;
  assign dataGroup_lo_lo_964 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_965;
  assign dataGroup_lo_lo_965 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_966;
  assign dataGroup_lo_lo_966 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_967;
  assign dataGroup_lo_lo_967 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_968;
  assign dataGroup_lo_lo_968 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_969;
  assign dataGroup_lo_lo_969 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_970;
  assign dataGroup_lo_lo_970 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_971;
  assign dataGroup_lo_lo_971 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_972;
  assign dataGroup_lo_lo_972 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_973;
  assign dataGroup_lo_lo_973 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_974;
  assign dataGroup_lo_lo_974 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_975;
  assign dataGroup_lo_lo_975 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_976;
  assign dataGroup_lo_lo_976 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_977;
  assign dataGroup_lo_lo_977 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_978;
  assign dataGroup_lo_lo_978 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_979;
  assign dataGroup_lo_lo_979 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_980;
  assign dataGroup_lo_lo_980 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_981;
  assign dataGroup_lo_lo_981 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_982;
  assign dataGroup_lo_lo_982 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_983;
  assign dataGroup_lo_lo_983 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_984;
  assign dataGroup_lo_lo_984 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_985;
  assign dataGroup_lo_lo_985 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_986;
  assign dataGroup_lo_lo_986 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_987;
  assign dataGroup_lo_lo_987 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_988;
  assign dataGroup_lo_lo_988 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_989;
  assign dataGroup_lo_lo_989 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_990;
  assign dataGroup_lo_lo_990 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_991;
  assign dataGroup_lo_lo_991 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_992;
  assign dataGroup_lo_lo_992 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_993;
  assign dataGroup_lo_lo_993 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_994;
  assign dataGroup_lo_lo_994 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_995;
  assign dataGroup_lo_lo_995 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_996;
  assign dataGroup_lo_lo_996 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_997;
  assign dataGroup_lo_lo_997 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_998;
  assign dataGroup_lo_lo_998 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_999;
  assign dataGroup_lo_lo_999 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1000;
  assign dataGroup_lo_lo_1000 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1001;
  assign dataGroup_lo_lo_1001 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1002;
  assign dataGroup_lo_lo_1002 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1003;
  assign dataGroup_lo_lo_1003 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1004;
  assign dataGroup_lo_lo_1004 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1005;
  assign dataGroup_lo_lo_1005 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1006;
  assign dataGroup_lo_lo_1006 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1007;
  assign dataGroup_lo_lo_1007 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1008;
  assign dataGroup_lo_lo_1008 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1009;
  assign dataGroup_lo_lo_1009 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1010;
  assign dataGroup_lo_lo_1010 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1011;
  assign dataGroup_lo_lo_1011 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1012;
  assign dataGroup_lo_lo_1012 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1013;
  assign dataGroup_lo_lo_1013 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1014;
  assign dataGroup_lo_lo_1014 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1015;
  assign dataGroup_lo_lo_1015 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1016;
  assign dataGroup_lo_lo_1016 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1017;
  assign dataGroup_lo_lo_1017 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1018;
  assign dataGroup_lo_lo_1018 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1019;
  assign dataGroup_lo_lo_1019 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1020;
  assign dataGroup_lo_lo_1020 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1021;
  assign dataGroup_lo_lo_1021 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1022;
  assign dataGroup_lo_lo_1022 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1023;
  assign dataGroup_lo_lo_1023 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1024;
  assign dataGroup_lo_lo_1024 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1025;
  assign dataGroup_lo_lo_1025 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1026;
  assign dataGroup_lo_lo_1026 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1027;
  assign dataGroup_lo_lo_1027 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1028;
  assign dataGroup_lo_lo_1028 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1029;
  assign dataGroup_lo_lo_1029 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1030;
  assign dataGroup_lo_lo_1030 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1031;
  assign dataGroup_lo_lo_1031 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1032;
  assign dataGroup_lo_lo_1032 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1033;
  assign dataGroup_lo_lo_1033 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1034;
  assign dataGroup_lo_lo_1034 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1035;
  assign dataGroup_lo_lo_1035 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1036;
  assign dataGroup_lo_lo_1036 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1037;
  assign dataGroup_lo_lo_1037 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1038;
  assign dataGroup_lo_lo_1038 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1039;
  assign dataGroup_lo_lo_1039 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1040;
  assign dataGroup_lo_lo_1040 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1041;
  assign dataGroup_lo_lo_1041 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1042;
  assign dataGroup_lo_lo_1042 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1043;
  assign dataGroup_lo_lo_1043 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1044;
  assign dataGroup_lo_lo_1044 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1045;
  assign dataGroup_lo_lo_1045 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1046;
  assign dataGroup_lo_lo_1046 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1047;
  assign dataGroup_lo_lo_1047 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1048;
  assign dataGroup_lo_lo_1048 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1049;
  assign dataGroup_lo_lo_1049 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1050;
  assign dataGroup_lo_lo_1050 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1051;
  assign dataGroup_lo_lo_1051 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1052;
  assign dataGroup_lo_lo_1052 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1053;
  assign dataGroup_lo_lo_1053 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1054;
  assign dataGroup_lo_lo_1054 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1055;
  assign dataGroup_lo_lo_1055 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1056;
  assign dataGroup_lo_lo_1056 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1057;
  assign dataGroup_lo_lo_1057 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1058;
  assign dataGroup_lo_lo_1058 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1059;
  assign dataGroup_lo_lo_1059 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1060;
  assign dataGroup_lo_lo_1060 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1061;
  assign dataGroup_lo_lo_1061 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1062;
  assign dataGroup_lo_lo_1062 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1063;
  assign dataGroup_lo_lo_1063 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1064;
  assign dataGroup_lo_lo_1064 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1065;
  assign dataGroup_lo_lo_1065 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1066;
  assign dataGroup_lo_lo_1066 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1067;
  assign dataGroup_lo_lo_1067 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1068;
  assign dataGroup_lo_lo_1068 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1069;
  assign dataGroup_lo_lo_1069 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1070;
  assign dataGroup_lo_lo_1070 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1071;
  assign dataGroup_lo_lo_1071 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1072;
  assign dataGroup_lo_lo_1072 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1073;
  assign dataGroup_lo_lo_1073 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1074;
  assign dataGroup_lo_lo_1074 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1075;
  assign dataGroup_lo_lo_1075 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1076;
  assign dataGroup_lo_lo_1076 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1077;
  assign dataGroup_lo_lo_1077 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1078;
  assign dataGroup_lo_lo_1078 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1079;
  assign dataGroup_lo_lo_1079 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1080;
  assign dataGroup_lo_lo_1080 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1081;
  assign dataGroup_lo_lo_1081 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1082;
  assign dataGroup_lo_lo_1082 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1083;
  assign dataGroup_lo_lo_1083 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1084;
  assign dataGroup_lo_lo_1084 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1085;
  assign dataGroup_lo_lo_1085 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1086;
  assign dataGroup_lo_lo_1086 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1087;
  assign dataGroup_lo_lo_1087 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1088;
  assign dataGroup_lo_lo_1088 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1089;
  assign dataGroup_lo_lo_1089 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1090;
  assign dataGroup_lo_lo_1090 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1091;
  assign dataGroup_lo_lo_1091 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1092;
  assign dataGroup_lo_lo_1092 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1093;
  assign dataGroup_lo_lo_1093 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1094;
  assign dataGroup_lo_lo_1094 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1095;
  assign dataGroup_lo_lo_1095 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1096;
  assign dataGroup_lo_lo_1096 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1097;
  assign dataGroup_lo_lo_1097 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1098;
  assign dataGroup_lo_lo_1098 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1099;
  assign dataGroup_lo_lo_1099 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1100;
  assign dataGroup_lo_lo_1100 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1101;
  assign dataGroup_lo_lo_1101 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1102;
  assign dataGroup_lo_lo_1102 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1103;
  assign dataGroup_lo_lo_1103 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1104;
  assign dataGroup_lo_lo_1104 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1105;
  assign dataGroup_lo_lo_1105 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1106;
  assign dataGroup_lo_lo_1106 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1107;
  assign dataGroup_lo_lo_1107 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1108;
  assign dataGroup_lo_lo_1108 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1109;
  assign dataGroup_lo_lo_1109 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1110;
  assign dataGroup_lo_lo_1110 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1111;
  assign dataGroup_lo_lo_1111 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1112;
  assign dataGroup_lo_lo_1112 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1113;
  assign dataGroup_lo_lo_1113 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1114;
  assign dataGroup_lo_lo_1114 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1115;
  assign dataGroup_lo_lo_1115 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1116;
  assign dataGroup_lo_lo_1116 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1117;
  assign dataGroup_lo_lo_1117 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1118;
  assign dataGroup_lo_lo_1118 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1119;
  assign dataGroup_lo_lo_1119 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1120;
  assign dataGroup_lo_lo_1120 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1121;
  assign dataGroup_lo_lo_1121 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1122;
  assign dataGroup_lo_lo_1122 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1123;
  assign dataGroup_lo_lo_1123 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1124;
  assign dataGroup_lo_lo_1124 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1125;
  assign dataGroup_lo_lo_1125 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1126;
  assign dataGroup_lo_lo_1126 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1127;
  assign dataGroup_lo_lo_1127 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1128;
  assign dataGroup_lo_lo_1128 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1129;
  assign dataGroup_lo_lo_1129 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1130;
  assign dataGroup_lo_lo_1130 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1131;
  assign dataGroup_lo_lo_1131 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1132;
  assign dataGroup_lo_lo_1132 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1133;
  assign dataGroup_lo_lo_1133 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1134;
  assign dataGroup_lo_lo_1134 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1135;
  assign dataGroup_lo_lo_1135 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1136;
  assign dataGroup_lo_lo_1136 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1137;
  assign dataGroup_lo_lo_1137 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1138;
  assign dataGroup_lo_lo_1138 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1139;
  assign dataGroup_lo_lo_1139 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1140;
  assign dataGroup_lo_lo_1140 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1141;
  assign dataGroup_lo_lo_1141 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1142;
  assign dataGroup_lo_lo_1142 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1143;
  assign dataGroup_lo_lo_1143 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1144;
  assign dataGroup_lo_lo_1144 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1145;
  assign dataGroup_lo_lo_1145 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1146;
  assign dataGroup_lo_lo_1146 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1147;
  assign dataGroup_lo_lo_1147 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1148;
  assign dataGroup_lo_lo_1148 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1149;
  assign dataGroup_lo_lo_1149 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1150;
  assign dataGroup_lo_lo_1150 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1151;
  assign dataGroup_lo_lo_1151 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1152;
  assign dataGroup_lo_lo_1152 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1153;
  assign dataGroup_lo_lo_1153 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1154;
  assign dataGroup_lo_lo_1154 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1155;
  assign dataGroup_lo_lo_1155 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1156;
  assign dataGroup_lo_lo_1156 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1157;
  assign dataGroup_lo_lo_1157 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1158;
  assign dataGroup_lo_lo_1158 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1159;
  assign dataGroup_lo_lo_1159 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1160;
  assign dataGroup_lo_lo_1160 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1161;
  assign dataGroup_lo_lo_1161 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1162;
  assign dataGroup_lo_lo_1162 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1163;
  assign dataGroup_lo_lo_1163 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1164;
  assign dataGroup_lo_lo_1164 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1165;
  assign dataGroup_lo_lo_1165 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1166;
  assign dataGroup_lo_lo_1166 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1167;
  assign dataGroup_lo_lo_1167 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1168;
  assign dataGroup_lo_lo_1168 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1169;
  assign dataGroup_lo_lo_1169 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1170;
  assign dataGroup_lo_lo_1170 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1171;
  assign dataGroup_lo_lo_1171 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1172;
  assign dataGroup_lo_lo_1172 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1173;
  assign dataGroup_lo_lo_1173 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1174;
  assign dataGroup_lo_lo_1174 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1175;
  assign dataGroup_lo_lo_1175 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1176;
  assign dataGroup_lo_lo_1176 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1177;
  assign dataGroup_lo_lo_1177 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1178;
  assign dataGroup_lo_lo_1178 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1179;
  assign dataGroup_lo_lo_1179 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1180;
  assign dataGroup_lo_lo_1180 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1181;
  assign dataGroup_lo_lo_1181 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1182;
  assign dataGroup_lo_lo_1182 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1183;
  assign dataGroup_lo_lo_1183 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1184;
  assign dataGroup_lo_lo_1184 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1185;
  assign dataGroup_lo_lo_1185 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1186;
  assign dataGroup_lo_lo_1186 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1187;
  assign dataGroup_lo_lo_1187 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1188;
  assign dataGroup_lo_lo_1188 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1189;
  assign dataGroup_lo_lo_1189 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1190;
  assign dataGroup_lo_lo_1190 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1191;
  assign dataGroup_lo_lo_1191 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1192;
  assign dataGroup_lo_lo_1192 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1193;
  assign dataGroup_lo_lo_1193 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1194;
  assign dataGroup_lo_lo_1194 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1195;
  assign dataGroup_lo_lo_1195 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1196;
  assign dataGroup_lo_lo_1196 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1197;
  assign dataGroup_lo_lo_1197 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1198;
  assign dataGroup_lo_lo_1198 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1199;
  assign dataGroup_lo_lo_1199 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1200;
  assign dataGroup_lo_lo_1200 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1201;
  assign dataGroup_lo_lo_1201 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1202;
  assign dataGroup_lo_lo_1202 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1203;
  assign dataGroup_lo_lo_1203 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1204;
  assign dataGroup_lo_lo_1204 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1205;
  assign dataGroup_lo_lo_1205 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1206;
  assign dataGroup_lo_lo_1206 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1207;
  assign dataGroup_lo_lo_1207 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1208;
  assign dataGroup_lo_lo_1208 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1209;
  assign dataGroup_lo_lo_1209 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1210;
  assign dataGroup_lo_lo_1210 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1211;
  assign dataGroup_lo_lo_1211 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1212;
  assign dataGroup_lo_lo_1212 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1213;
  assign dataGroup_lo_lo_1213 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1214;
  assign dataGroup_lo_lo_1214 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1215;
  assign dataGroup_lo_lo_1215 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1216;
  assign dataGroup_lo_lo_1216 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1217;
  assign dataGroup_lo_lo_1217 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1218;
  assign dataGroup_lo_lo_1218 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1219;
  assign dataGroup_lo_lo_1219 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1220;
  assign dataGroup_lo_lo_1220 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1221;
  assign dataGroup_lo_lo_1221 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1222;
  assign dataGroup_lo_lo_1222 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1223;
  assign dataGroup_lo_lo_1223 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1224;
  assign dataGroup_lo_lo_1224 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1225;
  assign dataGroup_lo_lo_1225 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1226;
  assign dataGroup_lo_lo_1226 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1227;
  assign dataGroup_lo_lo_1227 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1228;
  assign dataGroup_lo_lo_1228 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1229;
  assign dataGroup_lo_lo_1229 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1230;
  assign dataGroup_lo_lo_1230 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1231;
  assign dataGroup_lo_lo_1231 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1232;
  assign dataGroup_lo_lo_1232 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1233;
  assign dataGroup_lo_lo_1233 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1234;
  assign dataGroup_lo_lo_1234 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1235;
  assign dataGroup_lo_lo_1235 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1236;
  assign dataGroup_lo_lo_1236 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1237;
  assign dataGroup_lo_lo_1237 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1238;
  assign dataGroup_lo_lo_1238 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1239;
  assign dataGroup_lo_lo_1239 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1240;
  assign dataGroup_lo_lo_1240 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1241;
  assign dataGroup_lo_lo_1241 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1242;
  assign dataGroup_lo_lo_1242 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1243;
  assign dataGroup_lo_lo_1243 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1244;
  assign dataGroup_lo_lo_1244 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1245;
  assign dataGroup_lo_lo_1245 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1246;
  assign dataGroup_lo_lo_1246 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1247;
  assign dataGroup_lo_lo_1247 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1248;
  assign dataGroup_lo_lo_1248 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1249;
  assign dataGroup_lo_lo_1249 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1250;
  assign dataGroup_lo_lo_1250 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1251;
  assign dataGroup_lo_lo_1251 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1252;
  assign dataGroup_lo_lo_1252 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1253;
  assign dataGroup_lo_lo_1253 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1254;
  assign dataGroup_lo_lo_1254 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1255;
  assign dataGroup_lo_lo_1255 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1256;
  assign dataGroup_lo_lo_1256 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1257;
  assign dataGroup_lo_lo_1257 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1258;
  assign dataGroup_lo_lo_1258 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1259;
  assign dataGroup_lo_lo_1259 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1260;
  assign dataGroup_lo_lo_1260 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1261;
  assign dataGroup_lo_lo_1261 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1262;
  assign dataGroup_lo_lo_1262 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1263;
  assign dataGroup_lo_lo_1263 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1264;
  assign dataGroup_lo_lo_1264 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1265;
  assign dataGroup_lo_lo_1265 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1266;
  assign dataGroup_lo_lo_1266 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1267;
  assign dataGroup_lo_lo_1267 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1268;
  assign dataGroup_lo_lo_1268 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1269;
  assign dataGroup_lo_lo_1269 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1270;
  assign dataGroup_lo_lo_1270 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1271;
  assign dataGroup_lo_lo_1271 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1272;
  assign dataGroup_lo_lo_1272 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1273;
  assign dataGroup_lo_lo_1273 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1274;
  assign dataGroup_lo_lo_1274 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1275;
  assign dataGroup_lo_lo_1275 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1276;
  assign dataGroup_lo_lo_1276 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1277;
  assign dataGroup_lo_lo_1277 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1278;
  assign dataGroup_lo_lo_1278 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1279;
  assign dataGroup_lo_lo_1279 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1280;
  assign dataGroup_lo_lo_1280 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1281;
  assign dataGroup_lo_lo_1281 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1282;
  assign dataGroup_lo_lo_1282 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1283;
  assign dataGroup_lo_lo_1283 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1284;
  assign dataGroup_lo_lo_1284 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1285;
  assign dataGroup_lo_lo_1285 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1286;
  assign dataGroup_lo_lo_1286 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1287;
  assign dataGroup_lo_lo_1287 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1288;
  assign dataGroup_lo_lo_1288 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1289;
  assign dataGroup_lo_lo_1289 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1290;
  assign dataGroup_lo_lo_1290 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1291;
  assign dataGroup_lo_lo_1291 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1292;
  assign dataGroup_lo_lo_1292 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1293;
  assign dataGroup_lo_lo_1293 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1294;
  assign dataGroup_lo_lo_1294 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1295;
  assign dataGroup_lo_lo_1295 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1296;
  assign dataGroup_lo_lo_1296 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1297;
  assign dataGroup_lo_lo_1297 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1298;
  assign dataGroup_lo_lo_1298 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1299;
  assign dataGroup_lo_lo_1299 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1300;
  assign dataGroup_lo_lo_1300 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1301;
  assign dataGroup_lo_lo_1301 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1302;
  assign dataGroup_lo_lo_1302 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1303;
  assign dataGroup_lo_lo_1303 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1304;
  assign dataGroup_lo_lo_1304 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1305;
  assign dataGroup_lo_lo_1305 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1306;
  assign dataGroup_lo_lo_1306 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1307;
  assign dataGroup_lo_lo_1307 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1308;
  assign dataGroup_lo_lo_1308 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1309;
  assign dataGroup_lo_lo_1309 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1310;
  assign dataGroup_lo_lo_1310 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1311;
  assign dataGroup_lo_lo_1311 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1312;
  assign dataGroup_lo_lo_1312 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1313;
  assign dataGroup_lo_lo_1313 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1314;
  assign dataGroup_lo_lo_1314 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1315;
  assign dataGroup_lo_lo_1315 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1316;
  assign dataGroup_lo_lo_1316 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1317;
  assign dataGroup_lo_lo_1317 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1318;
  assign dataGroup_lo_lo_1318 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1319;
  assign dataGroup_lo_lo_1319 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1320;
  assign dataGroup_lo_lo_1320 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1321;
  assign dataGroup_lo_lo_1321 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1322;
  assign dataGroup_lo_lo_1322 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1323;
  assign dataGroup_lo_lo_1323 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1324;
  assign dataGroup_lo_lo_1324 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1325;
  assign dataGroup_lo_lo_1325 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1326;
  assign dataGroup_lo_lo_1326 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1327;
  assign dataGroup_lo_lo_1327 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1328;
  assign dataGroup_lo_lo_1328 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1329;
  assign dataGroup_lo_lo_1329 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1330;
  assign dataGroup_lo_lo_1330 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1331;
  assign dataGroup_lo_lo_1331 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1332;
  assign dataGroup_lo_lo_1332 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1333;
  assign dataGroup_lo_lo_1333 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1334;
  assign dataGroup_lo_lo_1334 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1335;
  assign dataGroup_lo_lo_1335 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1336;
  assign dataGroup_lo_lo_1336 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1337;
  assign dataGroup_lo_lo_1337 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1338;
  assign dataGroup_lo_lo_1338 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1339;
  assign dataGroup_lo_lo_1339 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1340;
  assign dataGroup_lo_lo_1340 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1341;
  assign dataGroup_lo_lo_1341 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1342;
  assign dataGroup_lo_lo_1342 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1343;
  assign dataGroup_lo_lo_1343 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1344;
  assign dataGroup_lo_lo_1344 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1345;
  assign dataGroup_lo_lo_1345 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1346;
  assign dataGroup_lo_lo_1346 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1347;
  assign dataGroup_lo_lo_1347 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1348;
  assign dataGroup_lo_lo_1348 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1349;
  assign dataGroup_lo_lo_1349 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1350;
  assign dataGroup_lo_lo_1350 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1351;
  assign dataGroup_lo_lo_1351 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1352;
  assign dataGroup_lo_lo_1352 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1353;
  assign dataGroup_lo_lo_1353 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1354;
  assign dataGroup_lo_lo_1354 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1355;
  assign dataGroup_lo_lo_1355 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1356;
  assign dataGroup_lo_lo_1356 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1357;
  assign dataGroup_lo_lo_1357 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1358;
  assign dataGroup_lo_lo_1358 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1359;
  assign dataGroup_lo_lo_1359 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1360;
  assign dataGroup_lo_lo_1360 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1361;
  assign dataGroup_lo_lo_1361 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1362;
  assign dataGroup_lo_lo_1362 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1363;
  assign dataGroup_lo_lo_1363 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1364;
  assign dataGroup_lo_lo_1364 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1365;
  assign dataGroup_lo_lo_1365 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1366;
  assign dataGroup_lo_lo_1366 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1367;
  assign dataGroup_lo_lo_1367 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1368;
  assign dataGroup_lo_lo_1368 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1369;
  assign dataGroup_lo_lo_1369 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1370;
  assign dataGroup_lo_lo_1370 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1371;
  assign dataGroup_lo_lo_1371 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1372;
  assign dataGroup_lo_lo_1372 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1373;
  assign dataGroup_lo_lo_1373 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1374;
  assign dataGroup_lo_lo_1374 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1375;
  assign dataGroup_lo_lo_1375 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1376;
  assign dataGroup_lo_lo_1376 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1377;
  assign dataGroup_lo_lo_1377 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1378;
  assign dataGroup_lo_lo_1378 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1379;
  assign dataGroup_lo_lo_1379 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1380;
  assign dataGroup_lo_lo_1380 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1381;
  assign dataGroup_lo_lo_1381 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1382;
  assign dataGroup_lo_lo_1382 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1383;
  assign dataGroup_lo_lo_1383 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1384;
  assign dataGroup_lo_lo_1384 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1385;
  assign dataGroup_lo_lo_1385 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1386;
  assign dataGroup_lo_lo_1386 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1387;
  assign dataGroup_lo_lo_1387 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1388;
  assign dataGroup_lo_lo_1388 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1389;
  assign dataGroup_lo_lo_1389 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1390;
  assign dataGroup_lo_lo_1390 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1391;
  assign dataGroup_lo_lo_1391 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1392;
  assign dataGroup_lo_lo_1392 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1393;
  assign dataGroup_lo_lo_1393 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1394;
  assign dataGroup_lo_lo_1394 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1395;
  assign dataGroup_lo_lo_1395 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1396;
  assign dataGroup_lo_lo_1396 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1397;
  assign dataGroup_lo_lo_1397 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1398;
  assign dataGroup_lo_lo_1398 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1399;
  assign dataGroup_lo_lo_1399 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1400;
  assign dataGroup_lo_lo_1400 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1401;
  assign dataGroup_lo_lo_1401 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1402;
  assign dataGroup_lo_lo_1402 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1403;
  assign dataGroup_lo_lo_1403 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1404;
  assign dataGroup_lo_lo_1404 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1405;
  assign dataGroup_lo_lo_1405 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1406;
  assign dataGroup_lo_lo_1406 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1407;
  assign dataGroup_lo_lo_1407 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1408;
  assign dataGroup_lo_lo_1408 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1409;
  assign dataGroup_lo_lo_1409 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1410;
  assign dataGroup_lo_lo_1410 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1411;
  assign dataGroup_lo_lo_1411 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1412;
  assign dataGroup_lo_lo_1412 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1413;
  assign dataGroup_lo_lo_1413 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1414;
  assign dataGroup_lo_lo_1414 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1415;
  assign dataGroup_lo_lo_1415 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1416;
  assign dataGroup_lo_lo_1416 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1417;
  assign dataGroup_lo_lo_1417 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1418;
  assign dataGroup_lo_lo_1418 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1419;
  assign dataGroup_lo_lo_1419 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1420;
  assign dataGroup_lo_lo_1420 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1421;
  assign dataGroup_lo_lo_1421 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1422;
  assign dataGroup_lo_lo_1422 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1423;
  assign dataGroup_lo_lo_1423 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1424;
  assign dataGroup_lo_lo_1424 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1425;
  assign dataGroup_lo_lo_1425 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1426;
  assign dataGroup_lo_lo_1426 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1427;
  assign dataGroup_lo_lo_1427 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1428;
  assign dataGroup_lo_lo_1428 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1429;
  assign dataGroup_lo_lo_1429 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1430;
  assign dataGroup_lo_lo_1430 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1431;
  assign dataGroup_lo_lo_1431 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1432;
  assign dataGroup_lo_lo_1432 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1433;
  assign dataGroup_lo_lo_1433 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1434;
  assign dataGroup_lo_lo_1434 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1435;
  assign dataGroup_lo_lo_1435 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1436;
  assign dataGroup_lo_lo_1436 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1437;
  assign dataGroup_lo_lo_1437 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1438;
  assign dataGroup_lo_lo_1438 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1439;
  assign dataGroup_lo_lo_1439 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1440;
  assign dataGroup_lo_lo_1440 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1441;
  assign dataGroup_lo_lo_1441 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1442;
  assign dataGroup_lo_lo_1442 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1443;
  assign dataGroup_lo_lo_1443 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1444;
  assign dataGroup_lo_lo_1444 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1445;
  assign dataGroup_lo_lo_1445 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1446;
  assign dataGroup_lo_lo_1446 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1447;
  assign dataGroup_lo_lo_1447 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1448;
  assign dataGroup_lo_lo_1448 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1449;
  assign dataGroup_lo_lo_1449 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1450;
  assign dataGroup_lo_lo_1450 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1451;
  assign dataGroup_lo_lo_1451 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1452;
  assign dataGroup_lo_lo_1452 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1453;
  assign dataGroup_lo_lo_1453 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1454;
  assign dataGroup_lo_lo_1454 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1455;
  assign dataGroup_lo_lo_1455 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1456;
  assign dataGroup_lo_lo_1456 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1457;
  assign dataGroup_lo_lo_1457 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1458;
  assign dataGroup_lo_lo_1458 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1459;
  assign dataGroup_lo_lo_1459 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1460;
  assign dataGroup_lo_lo_1460 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1461;
  assign dataGroup_lo_lo_1461 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1462;
  assign dataGroup_lo_lo_1462 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1463;
  assign dataGroup_lo_lo_1463 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1464;
  assign dataGroup_lo_lo_1464 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1465;
  assign dataGroup_lo_lo_1465 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1466;
  assign dataGroup_lo_lo_1466 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1467;
  assign dataGroup_lo_lo_1467 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1468;
  assign dataGroup_lo_lo_1468 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1469;
  assign dataGroup_lo_lo_1469 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1470;
  assign dataGroup_lo_lo_1470 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1471;
  assign dataGroup_lo_lo_1471 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1472;
  assign dataGroup_lo_lo_1472 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1473;
  assign dataGroup_lo_lo_1473 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1474;
  assign dataGroup_lo_lo_1474 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1475;
  assign dataGroup_lo_lo_1475 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1476;
  assign dataGroup_lo_lo_1476 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1477;
  assign dataGroup_lo_lo_1477 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1478;
  assign dataGroup_lo_lo_1478 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1479;
  assign dataGroup_lo_lo_1479 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1480;
  assign dataGroup_lo_lo_1480 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1481;
  assign dataGroup_lo_lo_1481 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1482;
  assign dataGroup_lo_lo_1482 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1483;
  assign dataGroup_lo_lo_1483 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1484;
  assign dataGroup_lo_lo_1484 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1485;
  assign dataGroup_lo_lo_1485 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1486;
  assign dataGroup_lo_lo_1486 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1487;
  assign dataGroup_lo_lo_1487 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1488;
  assign dataGroup_lo_lo_1488 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1489;
  assign dataGroup_lo_lo_1489 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1490;
  assign dataGroup_lo_lo_1490 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1491;
  assign dataGroup_lo_lo_1491 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1492;
  assign dataGroup_lo_lo_1492 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1493;
  assign dataGroup_lo_lo_1493 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1494;
  assign dataGroup_lo_lo_1494 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1495;
  assign dataGroup_lo_lo_1495 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1496;
  assign dataGroup_lo_lo_1496 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1497;
  assign dataGroup_lo_lo_1497 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1498;
  assign dataGroup_lo_lo_1498 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1499;
  assign dataGroup_lo_lo_1499 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1500;
  assign dataGroup_lo_lo_1500 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1501;
  assign dataGroup_lo_lo_1501 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1502;
  assign dataGroup_lo_lo_1502 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1503;
  assign dataGroup_lo_lo_1503 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1504;
  assign dataGroup_lo_lo_1504 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1505;
  assign dataGroup_lo_lo_1505 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1506;
  assign dataGroup_lo_lo_1506 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1507;
  assign dataGroup_lo_lo_1507 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1508;
  assign dataGroup_lo_lo_1508 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1509;
  assign dataGroup_lo_lo_1509 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1510;
  assign dataGroup_lo_lo_1510 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1511;
  assign dataGroup_lo_lo_1511 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1512;
  assign dataGroup_lo_lo_1512 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1513;
  assign dataGroup_lo_lo_1513 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1514;
  assign dataGroup_lo_lo_1514 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1515;
  assign dataGroup_lo_lo_1515 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1516;
  assign dataGroup_lo_lo_1516 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1517;
  assign dataGroup_lo_lo_1517 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1518;
  assign dataGroup_lo_lo_1518 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1519;
  assign dataGroup_lo_lo_1519 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1520;
  assign dataGroup_lo_lo_1520 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1521;
  assign dataGroup_lo_lo_1521 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1522;
  assign dataGroup_lo_lo_1522 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1523;
  assign dataGroup_lo_lo_1523 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1524;
  assign dataGroup_lo_lo_1524 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1525;
  assign dataGroup_lo_lo_1525 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1526;
  assign dataGroup_lo_lo_1526 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1527;
  assign dataGroup_lo_lo_1527 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1528;
  assign dataGroup_lo_lo_1528 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1529;
  assign dataGroup_lo_lo_1529 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1530;
  assign dataGroup_lo_lo_1530 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1531;
  assign dataGroup_lo_lo_1531 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1532;
  assign dataGroup_lo_lo_1532 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1533;
  assign dataGroup_lo_lo_1533 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1534;
  assign dataGroup_lo_lo_1534 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1535;
  assign dataGroup_lo_lo_1535 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1536;
  assign dataGroup_lo_lo_1536 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1537;
  assign dataGroup_lo_lo_1537 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1538;
  assign dataGroup_lo_lo_1538 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1539;
  assign dataGroup_lo_lo_1539 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1540;
  assign dataGroup_lo_lo_1540 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1541;
  assign dataGroup_lo_lo_1541 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1542;
  assign dataGroup_lo_lo_1542 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1543;
  assign dataGroup_lo_lo_1543 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1544;
  assign dataGroup_lo_lo_1544 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1545;
  assign dataGroup_lo_lo_1545 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1546;
  assign dataGroup_lo_lo_1546 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1547;
  assign dataGroup_lo_lo_1547 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1548;
  assign dataGroup_lo_lo_1548 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1549;
  assign dataGroup_lo_lo_1549 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1550;
  assign dataGroup_lo_lo_1550 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1551;
  assign dataGroup_lo_lo_1551 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1552;
  assign dataGroup_lo_lo_1552 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1553;
  assign dataGroup_lo_lo_1553 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1554;
  assign dataGroup_lo_lo_1554 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1555;
  assign dataGroup_lo_lo_1555 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1556;
  assign dataGroup_lo_lo_1556 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1557;
  assign dataGroup_lo_lo_1557 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1558;
  assign dataGroup_lo_lo_1558 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1559;
  assign dataGroup_lo_lo_1559 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1560;
  assign dataGroup_lo_lo_1560 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1561;
  assign dataGroup_lo_lo_1561 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1562;
  assign dataGroup_lo_lo_1562 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1563;
  assign dataGroup_lo_lo_1563 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1564;
  assign dataGroup_lo_lo_1564 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1565;
  assign dataGroup_lo_lo_1565 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1566;
  assign dataGroup_lo_lo_1566 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1567;
  assign dataGroup_lo_lo_1567 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1568;
  assign dataGroup_lo_lo_1568 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1569;
  assign dataGroup_lo_lo_1569 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1570;
  assign dataGroup_lo_lo_1570 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1571;
  assign dataGroup_lo_lo_1571 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1572;
  assign dataGroup_lo_lo_1572 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1573;
  assign dataGroup_lo_lo_1573 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1574;
  assign dataGroup_lo_lo_1574 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1575;
  assign dataGroup_lo_lo_1575 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1576;
  assign dataGroup_lo_lo_1576 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1577;
  assign dataGroup_lo_lo_1577 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1578;
  assign dataGroup_lo_lo_1578 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1579;
  assign dataGroup_lo_lo_1579 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1580;
  assign dataGroup_lo_lo_1580 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1581;
  assign dataGroup_lo_lo_1581 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1582;
  assign dataGroup_lo_lo_1582 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1583;
  assign dataGroup_lo_lo_1583 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1584;
  assign dataGroup_lo_lo_1584 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1585;
  assign dataGroup_lo_lo_1585 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1586;
  assign dataGroup_lo_lo_1586 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1587;
  assign dataGroup_lo_lo_1587 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1588;
  assign dataGroup_lo_lo_1588 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1589;
  assign dataGroup_lo_lo_1589 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1590;
  assign dataGroup_lo_lo_1590 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1591;
  assign dataGroup_lo_lo_1591 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1592;
  assign dataGroup_lo_lo_1592 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1593;
  assign dataGroup_lo_lo_1593 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1594;
  assign dataGroup_lo_lo_1594 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1595;
  assign dataGroup_lo_lo_1595 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1596;
  assign dataGroup_lo_lo_1596 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1597;
  assign dataGroup_lo_lo_1597 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1598;
  assign dataGroup_lo_lo_1598 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1599;
  assign dataGroup_lo_lo_1599 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1600;
  assign dataGroup_lo_lo_1600 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1601;
  assign dataGroup_lo_lo_1601 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1602;
  assign dataGroup_lo_lo_1602 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1603;
  assign dataGroup_lo_lo_1603 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1604;
  assign dataGroup_lo_lo_1604 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1605;
  assign dataGroup_lo_lo_1605 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1606;
  assign dataGroup_lo_lo_1606 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1607;
  assign dataGroup_lo_lo_1607 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1608;
  assign dataGroup_lo_lo_1608 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1609;
  assign dataGroup_lo_lo_1609 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1610;
  assign dataGroup_lo_lo_1610 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1611;
  assign dataGroup_lo_lo_1611 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1612;
  assign dataGroup_lo_lo_1612 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1613;
  assign dataGroup_lo_lo_1613 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1614;
  assign dataGroup_lo_lo_1614 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1615;
  assign dataGroup_lo_lo_1615 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1616;
  assign dataGroup_lo_lo_1616 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1617;
  assign dataGroup_lo_lo_1617 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1618;
  assign dataGroup_lo_lo_1618 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1619;
  assign dataGroup_lo_lo_1619 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1620;
  assign dataGroup_lo_lo_1620 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1621;
  assign dataGroup_lo_lo_1621 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1622;
  assign dataGroup_lo_lo_1622 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1623;
  assign dataGroup_lo_lo_1623 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1624;
  assign dataGroup_lo_lo_1624 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1625;
  assign dataGroup_lo_lo_1625 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1626;
  assign dataGroup_lo_lo_1626 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1627;
  assign dataGroup_lo_lo_1627 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1628;
  assign dataGroup_lo_lo_1628 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1629;
  assign dataGroup_lo_lo_1629 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1630;
  assign dataGroup_lo_lo_1630 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1631;
  assign dataGroup_lo_lo_1631 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1632;
  assign dataGroup_lo_lo_1632 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1633;
  assign dataGroup_lo_lo_1633 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1634;
  assign dataGroup_lo_lo_1634 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1635;
  assign dataGroup_lo_lo_1635 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1636;
  assign dataGroup_lo_lo_1636 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1637;
  assign dataGroup_lo_lo_1637 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1638;
  assign dataGroup_lo_lo_1638 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1639;
  assign dataGroup_lo_lo_1639 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1640;
  assign dataGroup_lo_lo_1640 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1641;
  assign dataGroup_lo_lo_1641 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1642;
  assign dataGroup_lo_lo_1642 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1643;
  assign dataGroup_lo_lo_1643 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1644;
  assign dataGroup_lo_lo_1644 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1645;
  assign dataGroup_lo_lo_1645 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1646;
  assign dataGroup_lo_lo_1646 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1647;
  assign dataGroup_lo_lo_1647 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1648;
  assign dataGroup_lo_lo_1648 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1649;
  assign dataGroup_lo_lo_1649 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1650;
  assign dataGroup_lo_lo_1650 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1651;
  assign dataGroup_lo_lo_1651 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1652;
  assign dataGroup_lo_lo_1652 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1653;
  assign dataGroup_lo_lo_1653 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1654;
  assign dataGroup_lo_lo_1654 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1655;
  assign dataGroup_lo_lo_1655 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1656;
  assign dataGroup_lo_lo_1656 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1657;
  assign dataGroup_lo_lo_1657 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1658;
  assign dataGroup_lo_lo_1658 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1659;
  assign dataGroup_lo_lo_1659 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1660;
  assign dataGroup_lo_lo_1660 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1661;
  assign dataGroup_lo_lo_1661 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1662;
  assign dataGroup_lo_lo_1662 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1663;
  assign dataGroup_lo_lo_1663 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1664;
  assign dataGroup_lo_lo_1664 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1665;
  assign dataGroup_lo_lo_1665 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1666;
  assign dataGroup_lo_lo_1666 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1667;
  assign dataGroup_lo_lo_1667 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1668;
  assign dataGroup_lo_lo_1668 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1669;
  assign dataGroup_lo_lo_1669 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1670;
  assign dataGroup_lo_lo_1670 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1671;
  assign dataGroup_lo_lo_1671 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1672;
  assign dataGroup_lo_lo_1672 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1673;
  assign dataGroup_lo_lo_1673 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1674;
  assign dataGroup_lo_lo_1674 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1675;
  assign dataGroup_lo_lo_1675 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1676;
  assign dataGroup_lo_lo_1676 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1677;
  assign dataGroup_lo_lo_1677 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1678;
  assign dataGroup_lo_lo_1678 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1679;
  assign dataGroup_lo_lo_1679 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1680;
  assign dataGroup_lo_lo_1680 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1681;
  assign dataGroup_lo_lo_1681 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1682;
  assign dataGroup_lo_lo_1682 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1683;
  assign dataGroup_lo_lo_1683 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1684;
  assign dataGroup_lo_lo_1684 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1685;
  assign dataGroup_lo_lo_1685 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1686;
  assign dataGroup_lo_lo_1686 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1687;
  assign dataGroup_lo_lo_1687 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1688;
  assign dataGroup_lo_lo_1688 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1689;
  assign dataGroup_lo_lo_1689 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1690;
  assign dataGroup_lo_lo_1690 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1691;
  assign dataGroup_lo_lo_1691 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1692;
  assign dataGroup_lo_lo_1692 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1693;
  assign dataGroup_lo_lo_1693 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1694;
  assign dataGroup_lo_lo_1694 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1695;
  assign dataGroup_lo_lo_1695 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1696;
  assign dataGroup_lo_lo_1696 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1697;
  assign dataGroup_lo_lo_1697 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1698;
  assign dataGroup_lo_lo_1698 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1699;
  assign dataGroup_lo_lo_1699 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1700;
  assign dataGroup_lo_lo_1700 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1701;
  assign dataGroup_lo_lo_1701 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1702;
  assign dataGroup_lo_lo_1702 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1703;
  assign dataGroup_lo_lo_1703 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1704;
  assign dataGroup_lo_lo_1704 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1705;
  assign dataGroup_lo_lo_1705 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1706;
  assign dataGroup_lo_lo_1706 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1707;
  assign dataGroup_lo_lo_1707 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1708;
  assign dataGroup_lo_lo_1708 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1709;
  assign dataGroup_lo_lo_1709 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1710;
  assign dataGroup_lo_lo_1710 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1711;
  assign dataGroup_lo_lo_1711 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1712;
  assign dataGroup_lo_lo_1712 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1713;
  assign dataGroup_lo_lo_1713 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1714;
  assign dataGroup_lo_lo_1714 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1715;
  assign dataGroup_lo_lo_1715 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1716;
  assign dataGroup_lo_lo_1716 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1717;
  assign dataGroup_lo_lo_1717 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1718;
  assign dataGroup_lo_lo_1718 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1719;
  assign dataGroup_lo_lo_1719 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1720;
  assign dataGroup_lo_lo_1720 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1721;
  assign dataGroup_lo_lo_1721 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1722;
  assign dataGroup_lo_lo_1722 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1723;
  assign dataGroup_lo_lo_1723 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1724;
  assign dataGroup_lo_lo_1724 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1725;
  assign dataGroup_lo_lo_1725 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1726;
  assign dataGroup_lo_lo_1726 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1727;
  assign dataGroup_lo_lo_1727 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1728;
  assign dataGroup_lo_lo_1728 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1729;
  assign dataGroup_lo_lo_1729 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1730;
  assign dataGroup_lo_lo_1730 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1731;
  assign dataGroup_lo_lo_1731 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1732;
  assign dataGroup_lo_lo_1732 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1733;
  assign dataGroup_lo_lo_1733 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1734;
  assign dataGroup_lo_lo_1734 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1735;
  assign dataGroup_lo_lo_1735 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1736;
  assign dataGroup_lo_lo_1736 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1737;
  assign dataGroup_lo_lo_1737 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1738;
  assign dataGroup_lo_lo_1738 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1739;
  assign dataGroup_lo_lo_1739 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1740;
  assign dataGroup_lo_lo_1740 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1741;
  assign dataGroup_lo_lo_1741 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1742;
  assign dataGroup_lo_lo_1742 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1743;
  assign dataGroup_lo_lo_1743 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1744;
  assign dataGroup_lo_lo_1744 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1745;
  assign dataGroup_lo_lo_1745 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1746;
  assign dataGroup_lo_lo_1746 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1747;
  assign dataGroup_lo_lo_1747 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1748;
  assign dataGroup_lo_lo_1748 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1749;
  assign dataGroup_lo_lo_1749 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1750;
  assign dataGroup_lo_lo_1750 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1751;
  assign dataGroup_lo_lo_1751 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1752;
  assign dataGroup_lo_lo_1752 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1753;
  assign dataGroup_lo_lo_1753 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1754;
  assign dataGroup_lo_lo_1754 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1755;
  assign dataGroup_lo_lo_1755 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1756;
  assign dataGroup_lo_lo_1756 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1757;
  assign dataGroup_lo_lo_1757 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1758;
  assign dataGroup_lo_lo_1758 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1759;
  assign dataGroup_lo_lo_1759 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1760;
  assign dataGroup_lo_lo_1760 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1761;
  assign dataGroup_lo_lo_1761 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1762;
  assign dataGroup_lo_lo_1762 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1763;
  assign dataGroup_lo_lo_1763 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1764;
  assign dataGroup_lo_lo_1764 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1765;
  assign dataGroup_lo_lo_1765 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1766;
  assign dataGroup_lo_lo_1766 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1767;
  assign dataGroup_lo_lo_1767 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1768;
  assign dataGroup_lo_lo_1768 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1769;
  assign dataGroup_lo_lo_1769 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1770;
  assign dataGroup_lo_lo_1770 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1771;
  assign dataGroup_lo_lo_1771 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1772;
  assign dataGroup_lo_lo_1772 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1773;
  assign dataGroup_lo_lo_1773 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1774;
  assign dataGroup_lo_lo_1774 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1775;
  assign dataGroup_lo_lo_1775 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1776;
  assign dataGroup_lo_lo_1776 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1777;
  assign dataGroup_lo_lo_1777 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1778;
  assign dataGroup_lo_lo_1778 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1779;
  assign dataGroup_lo_lo_1779 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1780;
  assign dataGroup_lo_lo_1780 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1781;
  assign dataGroup_lo_lo_1781 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1782;
  assign dataGroup_lo_lo_1782 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1783;
  assign dataGroup_lo_lo_1783 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1784;
  assign dataGroup_lo_lo_1784 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1785;
  assign dataGroup_lo_lo_1785 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1786;
  assign dataGroup_lo_lo_1786 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1787;
  assign dataGroup_lo_lo_1787 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1788;
  assign dataGroup_lo_lo_1788 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1789;
  assign dataGroup_lo_lo_1789 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1790;
  assign dataGroup_lo_lo_1790 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1791;
  assign dataGroup_lo_lo_1791 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1792;
  assign dataGroup_lo_lo_1792 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1793;
  assign dataGroup_lo_lo_1793 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1794;
  assign dataGroup_lo_lo_1794 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1795;
  assign dataGroup_lo_lo_1795 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1796;
  assign dataGroup_lo_lo_1796 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1797;
  assign dataGroup_lo_lo_1797 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1798;
  assign dataGroup_lo_lo_1798 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1799;
  assign dataGroup_lo_lo_1799 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1800;
  assign dataGroup_lo_lo_1800 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1801;
  assign dataGroup_lo_lo_1801 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1802;
  assign dataGroup_lo_lo_1802 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1803;
  assign dataGroup_lo_lo_1803 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1804;
  assign dataGroup_lo_lo_1804 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1805;
  assign dataGroup_lo_lo_1805 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1806;
  assign dataGroup_lo_lo_1806 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1807;
  assign dataGroup_lo_lo_1807 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1808;
  assign dataGroup_lo_lo_1808 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1809;
  assign dataGroup_lo_lo_1809 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1810;
  assign dataGroup_lo_lo_1810 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1811;
  assign dataGroup_lo_lo_1811 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1812;
  assign dataGroup_lo_lo_1812 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1813;
  assign dataGroup_lo_lo_1813 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1814;
  assign dataGroup_lo_lo_1814 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1815;
  assign dataGroup_lo_lo_1815 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1816;
  assign dataGroup_lo_lo_1816 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1817;
  assign dataGroup_lo_lo_1817 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1818;
  assign dataGroup_lo_lo_1818 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1819;
  assign dataGroup_lo_lo_1819 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1820;
  assign dataGroup_lo_lo_1820 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1821;
  assign dataGroup_lo_lo_1821 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1822;
  assign dataGroup_lo_lo_1822 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1823;
  assign dataGroup_lo_lo_1823 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1824;
  assign dataGroup_lo_lo_1824 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1825;
  assign dataGroup_lo_lo_1825 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1826;
  assign dataGroup_lo_lo_1826 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1827;
  assign dataGroup_lo_lo_1827 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1828;
  assign dataGroup_lo_lo_1828 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1829;
  assign dataGroup_lo_lo_1829 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1830;
  assign dataGroup_lo_lo_1830 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1831;
  assign dataGroup_lo_lo_1831 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1832;
  assign dataGroup_lo_lo_1832 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1833;
  assign dataGroup_lo_lo_1833 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1834;
  assign dataGroup_lo_lo_1834 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1835;
  assign dataGroup_lo_lo_1835 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1836;
  assign dataGroup_lo_lo_1836 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1837;
  assign dataGroup_lo_lo_1837 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1838;
  assign dataGroup_lo_lo_1838 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1839;
  assign dataGroup_lo_lo_1839 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1840;
  assign dataGroup_lo_lo_1840 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1841;
  assign dataGroup_lo_lo_1841 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1842;
  assign dataGroup_lo_lo_1842 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1843;
  assign dataGroup_lo_lo_1843 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1844;
  assign dataGroup_lo_lo_1844 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1845;
  assign dataGroup_lo_lo_1845 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1846;
  assign dataGroup_lo_lo_1846 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1847;
  assign dataGroup_lo_lo_1847 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1848;
  assign dataGroup_lo_lo_1848 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1849;
  assign dataGroup_lo_lo_1849 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1850;
  assign dataGroup_lo_lo_1850 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1851;
  assign dataGroup_lo_lo_1851 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1852;
  assign dataGroup_lo_lo_1852 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1853;
  assign dataGroup_lo_lo_1853 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1854;
  assign dataGroup_lo_lo_1854 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1855;
  assign dataGroup_lo_lo_1855 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1856;
  assign dataGroup_lo_lo_1856 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1857;
  assign dataGroup_lo_lo_1857 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1858;
  assign dataGroup_lo_lo_1858 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1859;
  assign dataGroup_lo_lo_1859 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1860;
  assign dataGroup_lo_lo_1860 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1861;
  assign dataGroup_lo_lo_1861 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1862;
  assign dataGroup_lo_lo_1862 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1863;
  assign dataGroup_lo_lo_1863 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1864;
  assign dataGroup_lo_lo_1864 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1865;
  assign dataGroup_lo_lo_1865 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1866;
  assign dataGroup_lo_lo_1866 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1867;
  assign dataGroup_lo_lo_1867 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1868;
  assign dataGroup_lo_lo_1868 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1869;
  assign dataGroup_lo_lo_1869 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1870;
  assign dataGroup_lo_lo_1870 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1871;
  assign dataGroup_lo_lo_1871 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1872;
  assign dataGroup_lo_lo_1872 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1873;
  assign dataGroup_lo_lo_1873 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1874;
  assign dataGroup_lo_lo_1874 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1875;
  assign dataGroup_lo_lo_1875 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1876;
  assign dataGroup_lo_lo_1876 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1877;
  assign dataGroup_lo_lo_1877 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1878;
  assign dataGroup_lo_lo_1878 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1879;
  assign dataGroup_lo_lo_1879 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1880;
  assign dataGroup_lo_lo_1880 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1881;
  assign dataGroup_lo_lo_1881 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1882;
  assign dataGroup_lo_lo_1882 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1883;
  assign dataGroup_lo_lo_1883 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1884;
  assign dataGroup_lo_lo_1884 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1885;
  assign dataGroup_lo_lo_1885 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1886;
  assign dataGroup_lo_lo_1886 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1887;
  assign dataGroup_lo_lo_1887 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1888;
  assign dataGroup_lo_lo_1888 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1889;
  assign dataGroup_lo_lo_1889 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1890;
  assign dataGroup_lo_lo_1890 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1891;
  assign dataGroup_lo_lo_1891 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1892;
  assign dataGroup_lo_lo_1892 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1893;
  assign dataGroup_lo_lo_1893 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1894;
  assign dataGroup_lo_lo_1894 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1895;
  assign dataGroup_lo_lo_1895 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1896;
  assign dataGroup_lo_lo_1896 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1897;
  assign dataGroup_lo_lo_1897 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1898;
  assign dataGroup_lo_lo_1898 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1899;
  assign dataGroup_lo_lo_1899 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1900;
  assign dataGroup_lo_lo_1900 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1901;
  assign dataGroup_lo_lo_1901 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1902;
  assign dataGroup_lo_lo_1902 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1903;
  assign dataGroup_lo_lo_1903 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1904;
  assign dataGroup_lo_lo_1904 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1905;
  assign dataGroup_lo_lo_1905 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1906;
  assign dataGroup_lo_lo_1906 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1907;
  assign dataGroup_lo_lo_1907 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1908;
  assign dataGroup_lo_lo_1908 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1909;
  assign dataGroup_lo_lo_1909 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1910;
  assign dataGroup_lo_lo_1910 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1911;
  assign dataGroup_lo_lo_1911 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1912;
  assign dataGroup_lo_lo_1912 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1913;
  assign dataGroup_lo_lo_1913 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1914;
  assign dataGroup_lo_lo_1914 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1915;
  assign dataGroup_lo_lo_1915 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1916;
  assign dataGroup_lo_lo_1916 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1917;
  assign dataGroup_lo_lo_1917 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1918;
  assign dataGroup_lo_lo_1918 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1919;
  assign dataGroup_lo_lo_1919 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1920;
  assign dataGroup_lo_lo_1920 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1921;
  assign dataGroup_lo_lo_1921 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1922;
  assign dataGroup_lo_lo_1922 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1923;
  assign dataGroup_lo_lo_1923 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1924;
  assign dataGroup_lo_lo_1924 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1925;
  assign dataGroup_lo_lo_1925 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1926;
  assign dataGroup_lo_lo_1926 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1927;
  assign dataGroup_lo_lo_1927 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1928;
  assign dataGroup_lo_lo_1928 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1929;
  assign dataGroup_lo_lo_1929 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1930;
  assign dataGroup_lo_lo_1930 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1931;
  assign dataGroup_lo_lo_1931 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1932;
  assign dataGroup_lo_lo_1932 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1933;
  assign dataGroup_lo_lo_1933 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1934;
  assign dataGroup_lo_lo_1934 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1935;
  assign dataGroup_lo_lo_1935 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1936;
  assign dataGroup_lo_lo_1936 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1937;
  assign dataGroup_lo_lo_1937 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1938;
  assign dataGroup_lo_lo_1938 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1939;
  assign dataGroup_lo_lo_1939 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1940;
  assign dataGroup_lo_lo_1940 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1941;
  assign dataGroup_lo_lo_1941 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1942;
  assign dataGroup_lo_lo_1942 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1943;
  assign dataGroup_lo_lo_1943 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1944;
  assign dataGroup_lo_lo_1944 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1945;
  assign dataGroup_lo_lo_1945 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1946;
  assign dataGroup_lo_lo_1946 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1947;
  assign dataGroup_lo_lo_1947 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1948;
  assign dataGroup_lo_lo_1948 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1949;
  assign dataGroup_lo_lo_1949 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1950;
  assign dataGroup_lo_lo_1950 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1951;
  assign dataGroup_lo_lo_1951 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1952;
  assign dataGroup_lo_lo_1952 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1953;
  assign dataGroup_lo_lo_1953 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1954;
  assign dataGroup_lo_lo_1954 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1955;
  assign dataGroup_lo_lo_1955 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1956;
  assign dataGroup_lo_lo_1956 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1957;
  assign dataGroup_lo_lo_1957 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1958;
  assign dataGroup_lo_lo_1958 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1959;
  assign dataGroup_lo_lo_1959 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1960;
  assign dataGroup_lo_lo_1960 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1961;
  assign dataGroup_lo_lo_1961 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1962;
  assign dataGroup_lo_lo_1962 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1963;
  assign dataGroup_lo_lo_1963 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1964;
  assign dataGroup_lo_lo_1964 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1965;
  assign dataGroup_lo_lo_1965 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1966;
  assign dataGroup_lo_lo_1966 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1967;
  assign dataGroup_lo_lo_1967 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1968;
  assign dataGroup_lo_lo_1968 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1969;
  assign dataGroup_lo_lo_1969 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1970;
  assign dataGroup_lo_lo_1970 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1971;
  assign dataGroup_lo_lo_1971 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1972;
  assign dataGroup_lo_lo_1972 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1973;
  assign dataGroup_lo_lo_1973 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1974;
  assign dataGroup_lo_lo_1974 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1975;
  assign dataGroup_lo_lo_1975 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1976;
  assign dataGroup_lo_lo_1976 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1977;
  assign dataGroup_lo_lo_1977 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1978;
  assign dataGroup_lo_lo_1978 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1979;
  assign dataGroup_lo_lo_1979 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1980;
  assign dataGroup_lo_lo_1980 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1981;
  assign dataGroup_lo_lo_1981 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1982;
  assign dataGroup_lo_lo_1982 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1983;
  assign dataGroup_lo_lo_1983 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1984;
  assign dataGroup_lo_lo_1984 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1985;
  assign dataGroup_lo_lo_1985 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1986;
  assign dataGroup_lo_lo_1986 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1987;
  assign dataGroup_lo_lo_1987 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1988;
  assign dataGroup_lo_lo_1988 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1989;
  assign dataGroup_lo_lo_1989 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1990;
  assign dataGroup_lo_lo_1990 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1991;
  assign dataGroup_lo_lo_1991 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1992;
  assign dataGroup_lo_lo_1992 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1993;
  assign dataGroup_lo_lo_1993 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1994;
  assign dataGroup_lo_lo_1994 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1995;
  assign dataGroup_lo_lo_1995 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1996;
  assign dataGroup_lo_lo_1996 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1997;
  assign dataGroup_lo_lo_1997 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1998;
  assign dataGroup_lo_lo_1998 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_1999;
  assign dataGroup_lo_lo_1999 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2000;
  assign dataGroup_lo_lo_2000 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2001;
  assign dataGroup_lo_lo_2001 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2002;
  assign dataGroup_lo_lo_2002 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2003;
  assign dataGroup_lo_lo_2003 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2004;
  assign dataGroup_lo_lo_2004 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2005;
  assign dataGroup_lo_lo_2005 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2006;
  assign dataGroup_lo_lo_2006 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2007;
  assign dataGroup_lo_lo_2007 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2008;
  assign dataGroup_lo_lo_2008 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2009;
  assign dataGroup_lo_lo_2009 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2010;
  assign dataGroup_lo_lo_2010 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2011;
  assign dataGroup_lo_lo_2011 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2012;
  assign dataGroup_lo_lo_2012 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2013;
  assign dataGroup_lo_lo_2013 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2014;
  assign dataGroup_lo_lo_2014 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2015;
  assign dataGroup_lo_lo_2015 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2016;
  assign dataGroup_lo_lo_2016 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2017;
  assign dataGroup_lo_lo_2017 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2018;
  assign dataGroup_lo_lo_2018 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2019;
  assign dataGroup_lo_lo_2019 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2020;
  assign dataGroup_lo_lo_2020 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2021;
  assign dataGroup_lo_lo_2021 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2022;
  assign dataGroup_lo_lo_2022 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2023;
  assign dataGroup_lo_lo_2023 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2024;
  assign dataGroup_lo_lo_2024 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2025;
  assign dataGroup_lo_lo_2025 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2026;
  assign dataGroup_lo_lo_2026 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2027;
  assign dataGroup_lo_lo_2027 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2028;
  assign dataGroup_lo_lo_2028 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2029;
  assign dataGroup_lo_lo_2029 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2030;
  assign dataGroup_lo_lo_2030 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2031;
  assign dataGroup_lo_lo_2031 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2032;
  assign dataGroup_lo_lo_2032 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2033;
  assign dataGroup_lo_lo_2033 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2034;
  assign dataGroup_lo_lo_2034 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2035;
  assign dataGroup_lo_lo_2035 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2036;
  assign dataGroup_lo_lo_2036 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2037;
  assign dataGroup_lo_lo_2037 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2038;
  assign dataGroup_lo_lo_2038 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2039;
  assign dataGroup_lo_lo_2039 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2040;
  assign dataGroup_lo_lo_2040 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2041;
  assign dataGroup_lo_lo_2041 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2042;
  assign dataGroup_lo_lo_2042 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2043;
  assign dataGroup_lo_lo_2043 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2044;
  assign dataGroup_lo_lo_2044 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2045;
  assign dataGroup_lo_lo_2045 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2046;
  assign dataGroup_lo_lo_2046 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2047;
  assign dataGroup_lo_lo_2047 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2048;
  assign dataGroup_lo_lo_2048 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2049;
  assign dataGroup_lo_lo_2049 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2050;
  assign dataGroup_lo_lo_2050 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2051;
  assign dataGroup_lo_lo_2051 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2052;
  assign dataGroup_lo_lo_2052 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2053;
  assign dataGroup_lo_lo_2053 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2054;
  assign dataGroup_lo_lo_2054 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2055;
  assign dataGroup_lo_lo_2055 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2056;
  assign dataGroup_lo_lo_2056 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2057;
  assign dataGroup_lo_lo_2057 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2058;
  assign dataGroup_lo_lo_2058 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2059;
  assign dataGroup_lo_lo_2059 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2060;
  assign dataGroup_lo_lo_2060 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2061;
  assign dataGroup_lo_lo_2061 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2062;
  assign dataGroup_lo_lo_2062 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2063;
  assign dataGroup_lo_lo_2063 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2064;
  assign dataGroup_lo_lo_2064 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2065;
  assign dataGroup_lo_lo_2065 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2066;
  assign dataGroup_lo_lo_2066 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2067;
  assign dataGroup_lo_lo_2067 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2068;
  assign dataGroup_lo_lo_2068 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2069;
  assign dataGroup_lo_lo_2069 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2070;
  assign dataGroup_lo_lo_2070 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2071;
  assign dataGroup_lo_lo_2071 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2072;
  assign dataGroup_lo_lo_2072 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2073;
  assign dataGroup_lo_lo_2073 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2074;
  assign dataGroup_lo_lo_2074 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2075;
  assign dataGroup_lo_lo_2075 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2076;
  assign dataGroup_lo_lo_2076 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2077;
  assign dataGroup_lo_lo_2077 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2078;
  assign dataGroup_lo_lo_2078 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2079;
  assign dataGroup_lo_lo_2079 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2080;
  assign dataGroup_lo_lo_2080 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2081;
  assign dataGroup_lo_lo_2081 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2082;
  assign dataGroup_lo_lo_2082 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2083;
  assign dataGroup_lo_lo_2083 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2084;
  assign dataGroup_lo_lo_2084 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2085;
  assign dataGroup_lo_lo_2085 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2086;
  assign dataGroup_lo_lo_2086 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2087;
  assign dataGroup_lo_lo_2087 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2088;
  assign dataGroup_lo_lo_2088 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2089;
  assign dataGroup_lo_lo_2089 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2090;
  assign dataGroup_lo_lo_2090 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2091;
  assign dataGroup_lo_lo_2091 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2092;
  assign dataGroup_lo_lo_2092 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2093;
  assign dataGroup_lo_lo_2093 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2094;
  assign dataGroup_lo_lo_2094 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2095;
  assign dataGroup_lo_lo_2095 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2096;
  assign dataGroup_lo_lo_2096 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2097;
  assign dataGroup_lo_lo_2097 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2098;
  assign dataGroup_lo_lo_2098 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2099;
  assign dataGroup_lo_lo_2099 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2100;
  assign dataGroup_lo_lo_2100 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2101;
  assign dataGroup_lo_lo_2101 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2102;
  assign dataGroup_lo_lo_2102 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2103;
  assign dataGroup_lo_lo_2103 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2104;
  assign dataGroup_lo_lo_2104 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2105;
  assign dataGroup_lo_lo_2105 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2106;
  assign dataGroup_lo_lo_2106 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2107;
  assign dataGroup_lo_lo_2107 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2108;
  assign dataGroup_lo_lo_2108 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2109;
  assign dataGroup_lo_lo_2109 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2110;
  assign dataGroup_lo_lo_2110 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2111;
  assign dataGroup_lo_lo_2111 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2112;
  assign dataGroup_lo_lo_2112 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2113;
  assign dataGroup_lo_lo_2113 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2114;
  assign dataGroup_lo_lo_2114 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2115;
  assign dataGroup_lo_lo_2115 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2116;
  assign dataGroup_lo_lo_2116 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2117;
  assign dataGroup_lo_lo_2117 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2118;
  assign dataGroup_lo_lo_2118 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2119;
  assign dataGroup_lo_lo_2119 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2120;
  assign dataGroup_lo_lo_2120 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2121;
  assign dataGroup_lo_lo_2121 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2122;
  assign dataGroup_lo_lo_2122 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2123;
  assign dataGroup_lo_lo_2123 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2124;
  assign dataGroup_lo_lo_2124 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2125;
  assign dataGroup_lo_lo_2125 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2126;
  assign dataGroup_lo_lo_2126 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2127;
  assign dataGroup_lo_lo_2127 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2128;
  assign dataGroup_lo_lo_2128 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2129;
  assign dataGroup_lo_lo_2129 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2130;
  assign dataGroup_lo_lo_2130 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2131;
  assign dataGroup_lo_lo_2131 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2132;
  assign dataGroup_lo_lo_2132 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2133;
  assign dataGroup_lo_lo_2133 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2134;
  assign dataGroup_lo_lo_2134 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2135;
  assign dataGroup_lo_lo_2135 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2136;
  assign dataGroup_lo_lo_2136 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2137;
  assign dataGroup_lo_lo_2137 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2138;
  assign dataGroup_lo_lo_2138 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2139;
  assign dataGroup_lo_lo_2139 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2140;
  assign dataGroup_lo_lo_2140 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2141;
  assign dataGroup_lo_lo_2141 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2142;
  assign dataGroup_lo_lo_2142 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2143;
  assign dataGroup_lo_lo_2143 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2144;
  assign dataGroup_lo_lo_2144 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2145;
  assign dataGroup_lo_lo_2145 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2146;
  assign dataGroup_lo_lo_2146 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2147;
  assign dataGroup_lo_lo_2147 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2148;
  assign dataGroup_lo_lo_2148 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2149;
  assign dataGroup_lo_lo_2149 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2150;
  assign dataGroup_lo_lo_2150 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2151;
  assign dataGroup_lo_lo_2151 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2152;
  assign dataGroup_lo_lo_2152 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2153;
  assign dataGroup_lo_lo_2153 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2154;
  assign dataGroup_lo_lo_2154 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2155;
  assign dataGroup_lo_lo_2155 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2156;
  assign dataGroup_lo_lo_2156 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2157;
  assign dataGroup_lo_lo_2157 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2158;
  assign dataGroup_lo_lo_2158 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2159;
  assign dataGroup_lo_lo_2159 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2160;
  assign dataGroup_lo_lo_2160 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2161;
  assign dataGroup_lo_lo_2161 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2162;
  assign dataGroup_lo_lo_2162 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2163;
  assign dataGroup_lo_lo_2163 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2164;
  assign dataGroup_lo_lo_2164 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2165;
  assign dataGroup_lo_lo_2165 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2166;
  assign dataGroup_lo_lo_2166 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2167;
  assign dataGroup_lo_lo_2167 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2168;
  assign dataGroup_lo_lo_2168 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2169;
  assign dataGroup_lo_lo_2169 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2170;
  assign dataGroup_lo_lo_2170 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2171;
  assign dataGroup_lo_lo_2171 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2172;
  assign dataGroup_lo_lo_2172 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2173;
  assign dataGroup_lo_lo_2173 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2174;
  assign dataGroup_lo_lo_2174 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2175;
  assign dataGroup_lo_lo_2175 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2176;
  assign dataGroup_lo_lo_2176 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2177;
  assign dataGroup_lo_lo_2177 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2178;
  assign dataGroup_lo_lo_2178 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2179;
  assign dataGroup_lo_lo_2179 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2180;
  assign dataGroup_lo_lo_2180 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2181;
  assign dataGroup_lo_lo_2181 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2182;
  assign dataGroup_lo_lo_2182 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2183;
  assign dataGroup_lo_lo_2183 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2184;
  assign dataGroup_lo_lo_2184 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2185;
  assign dataGroup_lo_lo_2185 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2186;
  assign dataGroup_lo_lo_2186 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2187;
  assign dataGroup_lo_lo_2187 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2188;
  assign dataGroup_lo_lo_2188 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2189;
  assign dataGroup_lo_lo_2189 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2190;
  assign dataGroup_lo_lo_2190 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2191;
  assign dataGroup_lo_lo_2191 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2192;
  assign dataGroup_lo_lo_2192 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2193;
  assign dataGroup_lo_lo_2193 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2194;
  assign dataGroup_lo_lo_2194 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2195;
  assign dataGroup_lo_lo_2195 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2196;
  assign dataGroup_lo_lo_2196 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2197;
  assign dataGroup_lo_lo_2197 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2198;
  assign dataGroup_lo_lo_2198 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2199;
  assign dataGroup_lo_lo_2199 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2200;
  assign dataGroup_lo_lo_2200 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2201;
  assign dataGroup_lo_lo_2201 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2202;
  assign dataGroup_lo_lo_2202 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2203;
  assign dataGroup_lo_lo_2203 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2204;
  assign dataGroup_lo_lo_2204 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2205;
  assign dataGroup_lo_lo_2205 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2206;
  assign dataGroup_lo_lo_2206 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2207;
  assign dataGroup_lo_lo_2207 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2208;
  assign dataGroup_lo_lo_2208 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2209;
  assign dataGroup_lo_lo_2209 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2210;
  assign dataGroup_lo_lo_2210 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2211;
  assign dataGroup_lo_lo_2211 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2212;
  assign dataGroup_lo_lo_2212 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2213;
  assign dataGroup_lo_lo_2213 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2214;
  assign dataGroup_lo_lo_2214 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2215;
  assign dataGroup_lo_lo_2215 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2216;
  assign dataGroup_lo_lo_2216 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2217;
  assign dataGroup_lo_lo_2217 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2218;
  assign dataGroup_lo_lo_2218 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2219;
  assign dataGroup_lo_lo_2219 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2220;
  assign dataGroup_lo_lo_2220 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2221;
  assign dataGroup_lo_lo_2221 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2222;
  assign dataGroup_lo_lo_2222 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2223;
  assign dataGroup_lo_lo_2223 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2224;
  assign dataGroup_lo_lo_2224 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2225;
  assign dataGroup_lo_lo_2225 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2226;
  assign dataGroup_lo_lo_2226 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2227;
  assign dataGroup_lo_lo_2227 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2228;
  assign dataGroup_lo_lo_2228 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2229;
  assign dataGroup_lo_lo_2229 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2230;
  assign dataGroup_lo_lo_2230 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2231;
  assign dataGroup_lo_lo_2231 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2232;
  assign dataGroup_lo_lo_2232 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2233;
  assign dataGroup_lo_lo_2233 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2234;
  assign dataGroup_lo_lo_2234 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2235;
  assign dataGroup_lo_lo_2235 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2236;
  assign dataGroup_lo_lo_2236 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2237;
  assign dataGroup_lo_lo_2237 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2238;
  assign dataGroup_lo_lo_2238 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2239;
  assign dataGroup_lo_lo_2239 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2240;
  assign dataGroup_lo_lo_2240 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2241;
  assign dataGroup_lo_lo_2241 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2242;
  assign dataGroup_lo_lo_2242 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2243;
  assign dataGroup_lo_lo_2243 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2244;
  assign dataGroup_lo_lo_2244 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2245;
  assign dataGroup_lo_lo_2245 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2246;
  assign dataGroup_lo_lo_2246 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2247;
  assign dataGroup_lo_lo_2247 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2248;
  assign dataGroup_lo_lo_2248 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2249;
  assign dataGroup_lo_lo_2249 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2250;
  assign dataGroup_lo_lo_2250 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2251;
  assign dataGroup_lo_lo_2251 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2252;
  assign dataGroup_lo_lo_2252 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2253;
  assign dataGroup_lo_lo_2253 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2254;
  assign dataGroup_lo_lo_2254 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2255;
  assign dataGroup_lo_lo_2255 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2256;
  assign dataGroup_lo_lo_2256 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2257;
  assign dataGroup_lo_lo_2257 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2258;
  assign dataGroup_lo_lo_2258 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2259;
  assign dataGroup_lo_lo_2259 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2260;
  assign dataGroup_lo_lo_2260 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2261;
  assign dataGroup_lo_lo_2261 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2262;
  assign dataGroup_lo_lo_2262 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2263;
  assign dataGroup_lo_lo_2263 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2264;
  assign dataGroup_lo_lo_2264 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2265;
  assign dataGroup_lo_lo_2265 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2266;
  assign dataGroup_lo_lo_2266 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2267;
  assign dataGroup_lo_lo_2267 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2268;
  assign dataGroup_lo_lo_2268 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2269;
  assign dataGroup_lo_lo_2269 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2270;
  assign dataGroup_lo_lo_2270 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2271;
  assign dataGroup_lo_lo_2271 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2272;
  assign dataGroup_lo_lo_2272 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2273;
  assign dataGroup_lo_lo_2273 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2274;
  assign dataGroup_lo_lo_2274 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2275;
  assign dataGroup_lo_lo_2275 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2276;
  assign dataGroup_lo_lo_2276 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2277;
  assign dataGroup_lo_lo_2277 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2278;
  assign dataGroup_lo_lo_2278 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2279;
  assign dataGroup_lo_lo_2279 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2280;
  assign dataGroup_lo_lo_2280 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2281;
  assign dataGroup_lo_lo_2281 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2282;
  assign dataGroup_lo_lo_2282 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2283;
  assign dataGroup_lo_lo_2283 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2284;
  assign dataGroup_lo_lo_2284 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2285;
  assign dataGroup_lo_lo_2285 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2286;
  assign dataGroup_lo_lo_2286 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2287;
  assign dataGroup_lo_lo_2287 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2288;
  assign dataGroup_lo_lo_2288 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2289;
  assign dataGroup_lo_lo_2289 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2290;
  assign dataGroup_lo_lo_2290 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2291;
  assign dataGroup_lo_lo_2291 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2292;
  assign dataGroup_lo_lo_2292 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2293;
  assign dataGroup_lo_lo_2293 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2294;
  assign dataGroup_lo_lo_2294 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2295;
  assign dataGroup_lo_lo_2295 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2296;
  assign dataGroup_lo_lo_2296 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2297;
  assign dataGroup_lo_lo_2297 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2298;
  assign dataGroup_lo_lo_2298 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2299;
  assign dataGroup_lo_lo_2299 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2300;
  assign dataGroup_lo_lo_2300 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2301;
  assign dataGroup_lo_lo_2301 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2302;
  assign dataGroup_lo_lo_2302 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2303;
  assign dataGroup_lo_lo_2303 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2304;
  assign dataGroup_lo_lo_2304 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2305;
  assign dataGroup_lo_lo_2305 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2306;
  assign dataGroup_lo_lo_2306 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2307;
  assign dataGroup_lo_lo_2307 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2308;
  assign dataGroup_lo_lo_2308 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2309;
  assign dataGroup_lo_lo_2309 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2310;
  assign dataGroup_lo_lo_2310 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2311;
  assign dataGroup_lo_lo_2311 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2312;
  assign dataGroup_lo_lo_2312 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2313;
  assign dataGroup_lo_lo_2313 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2314;
  assign dataGroup_lo_lo_2314 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2315;
  assign dataGroup_lo_lo_2315 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2316;
  assign dataGroup_lo_lo_2316 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2317;
  assign dataGroup_lo_lo_2317 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2318;
  assign dataGroup_lo_lo_2318 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2319;
  assign dataGroup_lo_lo_2319 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2320;
  assign dataGroup_lo_lo_2320 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2321;
  assign dataGroup_lo_lo_2321 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2322;
  assign dataGroup_lo_lo_2322 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2323;
  assign dataGroup_lo_lo_2323 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2324;
  assign dataGroup_lo_lo_2324 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2325;
  assign dataGroup_lo_lo_2325 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2326;
  assign dataGroup_lo_lo_2326 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2327;
  assign dataGroup_lo_lo_2327 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2328;
  assign dataGroup_lo_lo_2328 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2329;
  assign dataGroup_lo_lo_2329 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2330;
  assign dataGroup_lo_lo_2330 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2331;
  assign dataGroup_lo_lo_2331 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2332;
  assign dataGroup_lo_lo_2332 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2333;
  assign dataGroup_lo_lo_2333 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2334;
  assign dataGroup_lo_lo_2334 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2335;
  assign dataGroup_lo_lo_2335 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2336;
  assign dataGroup_lo_lo_2336 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2337;
  assign dataGroup_lo_lo_2337 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2338;
  assign dataGroup_lo_lo_2338 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2339;
  assign dataGroup_lo_lo_2339 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2340;
  assign dataGroup_lo_lo_2340 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2341;
  assign dataGroup_lo_lo_2341 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2342;
  assign dataGroup_lo_lo_2342 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2343;
  assign dataGroup_lo_lo_2343 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2344;
  assign dataGroup_lo_lo_2344 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2345;
  assign dataGroup_lo_lo_2345 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2346;
  assign dataGroup_lo_lo_2346 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2347;
  assign dataGroup_lo_lo_2347 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2348;
  assign dataGroup_lo_lo_2348 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2349;
  assign dataGroup_lo_lo_2349 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2350;
  assign dataGroup_lo_lo_2350 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2351;
  assign dataGroup_lo_lo_2351 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2352;
  assign dataGroup_lo_lo_2352 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2353;
  assign dataGroup_lo_lo_2353 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2354;
  assign dataGroup_lo_lo_2354 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2355;
  assign dataGroup_lo_lo_2355 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2356;
  assign dataGroup_lo_lo_2356 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2357;
  assign dataGroup_lo_lo_2357 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2358;
  assign dataGroup_lo_lo_2358 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2359;
  assign dataGroup_lo_lo_2359 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2360;
  assign dataGroup_lo_lo_2360 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2361;
  assign dataGroup_lo_lo_2361 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2362;
  assign dataGroup_lo_lo_2362 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2363;
  assign dataGroup_lo_lo_2363 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2364;
  assign dataGroup_lo_lo_2364 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2365;
  assign dataGroup_lo_lo_2365 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2366;
  assign dataGroup_lo_lo_2366 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2367;
  assign dataGroup_lo_lo_2367 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2368;
  assign dataGroup_lo_lo_2368 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2369;
  assign dataGroup_lo_lo_2369 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2370;
  assign dataGroup_lo_lo_2370 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2371;
  assign dataGroup_lo_lo_2371 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2372;
  assign dataGroup_lo_lo_2372 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2373;
  assign dataGroup_lo_lo_2373 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2374;
  assign dataGroup_lo_lo_2374 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2375;
  assign dataGroup_lo_lo_2375 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2376;
  assign dataGroup_lo_lo_2376 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2377;
  assign dataGroup_lo_lo_2377 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2378;
  assign dataGroup_lo_lo_2378 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2379;
  assign dataGroup_lo_lo_2379 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2380;
  assign dataGroup_lo_lo_2380 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2381;
  assign dataGroup_lo_lo_2381 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2382;
  assign dataGroup_lo_lo_2382 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2383;
  assign dataGroup_lo_lo_2383 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2384;
  assign dataGroup_lo_lo_2384 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2385;
  assign dataGroup_lo_lo_2385 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2386;
  assign dataGroup_lo_lo_2386 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2387;
  assign dataGroup_lo_lo_2387 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2388;
  assign dataGroup_lo_lo_2388 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2389;
  assign dataGroup_lo_lo_2389 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2390;
  assign dataGroup_lo_lo_2390 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2391;
  assign dataGroup_lo_lo_2391 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2392;
  assign dataGroup_lo_lo_2392 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2393;
  assign dataGroup_lo_lo_2393 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2394;
  assign dataGroup_lo_lo_2394 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2395;
  assign dataGroup_lo_lo_2395 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2396;
  assign dataGroup_lo_lo_2396 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2397;
  assign dataGroup_lo_lo_2397 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2398;
  assign dataGroup_lo_lo_2398 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2399;
  assign dataGroup_lo_lo_2399 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2400;
  assign dataGroup_lo_lo_2400 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2401;
  assign dataGroup_lo_lo_2401 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2402;
  assign dataGroup_lo_lo_2402 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2403;
  assign dataGroup_lo_lo_2403 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2404;
  assign dataGroup_lo_lo_2404 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2405;
  assign dataGroup_lo_lo_2405 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2406;
  assign dataGroup_lo_lo_2406 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2407;
  assign dataGroup_lo_lo_2407 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2408;
  assign dataGroup_lo_lo_2408 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2409;
  assign dataGroup_lo_lo_2409 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2410;
  assign dataGroup_lo_lo_2410 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2411;
  assign dataGroup_lo_lo_2411 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2412;
  assign dataGroup_lo_lo_2412 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2413;
  assign dataGroup_lo_lo_2413 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2414;
  assign dataGroup_lo_lo_2414 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2415;
  assign dataGroup_lo_lo_2415 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2416;
  assign dataGroup_lo_lo_2416 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2417;
  assign dataGroup_lo_lo_2417 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2418;
  assign dataGroup_lo_lo_2418 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2419;
  assign dataGroup_lo_lo_2419 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2420;
  assign dataGroup_lo_lo_2420 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2421;
  assign dataGroup_lo_lo_2421 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2422;
  assign dataGroup_lo_lo_2422 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2423;
  assign dataGroup_lo_lo_2423 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2424;
  assign dataGroup_lo_lo_2424 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2425;
  assign dataGroup_lo_lo_2425 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2426;
  assign dataGroup_lo_lo_2426 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2427;
  assign dataGroup_lo_lo_2427 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2428;
  assign dataGroup_lo_lo_2428 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2429;
  assign dataGroup_lo_lo_2429 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2430;
  assign dataGroup_lo_lo_2430 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2431;
  assign dataGroup_lo_lo_2431 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2432;
  assign dataGroup_lo_lo_2432 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2433;
  assign dataGroup_lo_lo_2433 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2434;
  assign dataGroup_lo_lo_2434 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2435;
  assign dataGroup_lo_lo_2435 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2436;
  assign dataGroup_lo_lo_2436 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2437;
  assign dataGroup_lo_lo_2437 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2438;
  assign dataGroup_lo_lo_2438 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2439;
  assign dataGroup_lo_lo_2439 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2440;
  assign dataGroup_lo_lo_2440 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2441;
  assign dataGroup_lo_lo_2441 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2442;
  assign dataGroup_lo_lo_2442 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2443;
  assign dataGroup_lo_lo_2443 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2444;
  assign dataGroup_lo_lo_2444 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2445;
  assign dataGroup_lo_lo_2445 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2446;
  assign dataGroup_lo_lo_2446 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2447;
  assign dataGroup_lo_lo_2447 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2448;
  assign dataGroup_lo_lo_2448 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2449;
  assign dataGroup_lo_lo_2449 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2450;
  assign dataGroup_lo_lo_2450 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2451;
  assign dataGroup_lo_lo_2451 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2452;
  assign dataGroup_lo_lo_2452 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2453;
  assign dataGroup_lo_lo_2453 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2454;
  assign dataGroup_lo_lo_2454 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2455;
  assign dataGroup_lo_lo_2455 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2456;
  assign dataGroup_lo_lo_2456 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2457;
  assign dataGroup_lo_lo_2457 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2458;
  assign dataGroup_lo_lo_2458 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2459;
  assign dataGroup_lo_lo_2459 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2460;
  assign dataGroup_lo_lo_2460 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2461;
  assign dataGroup_lo_lo_2461 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2462;
  assign dataGroup_lo_lo_2462 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2463;
  assign dataGroup_lo_lo_2463 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2464;
  assign dataGroup_lo_lo_2464 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2465;
  assign dataGroup_lo_lo_2465 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2466;
  assign dataGroup_lo_lo_2466 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2467;
  assign dataGroup_lo_lo_2467 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2468;
  assign dataGroup_lo_lo_2468 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2469;
  assign dataGroup_lo_lo_2469 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2470;
  assign dataGroup_lo_lo_2470 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2471;
  assign dataGroup_lo_lo_2471 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2472;
  assign dataGroup_lo_lo_2472 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2473;
  assign dataGroup_lo_lo_2473 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2474;
  assign dataGroup_lo_lo_2474 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2475;
  assign dataGroup_lo_lo_2475 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2476;
  assign dataGroup_lo_lo_2476 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2477;
  assign dataGroup_lo_lo_2477 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2478;
  assign dataGroup_lo_lo_2478 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2479;
  assign dataGroup_lo_lo_2479 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2480;
  assign dataGroup_lo_lo_2480 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2481;
  assign dataGroup_lo_lo_2481 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2482;
  assign dataGroup_lo_lo_2482 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2483;
  assign dataGroup_lo_lo_2483 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2484;
  assign dataGroup_lo_lo_2484 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2485;
  assign dataGroup_lo_lo_2485 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2486;
  assign dataGroup_lo_lo_2486 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2487;
  assign dataGroup_lo_lo_2487 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2488;
  assign dataGroup_lo_lo_2488 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2489;
  assign dataGroup_lo_lo_2489 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2490;
  assign dataGroup_lo_lo_2490 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2491;
  assign dataGroup_lo_lo_2491 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2492;
  assign dataGroup_lo_lo_2492 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2493;
  assign dataGroup_lo_lo_2493 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2494;
  assign dataGroup_lo_lo_2494 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2495;
  assign dataGroup_lo_lo_2495 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2496;
  assign dataGroup_lo_lo_2496 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2497;
  assign dataGroup_lo_lo_2497 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2498;
  assign dataGroup_lo_lo_2498 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2499;
  assign dataGroup_lo_lo_2499 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2500;
  assign dataGroup_lo_lo_2500 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2501;
  assign dataGroup_lo_lo_2501 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2502;
  assign dataGroup_lo_lo_2502 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2503;
  assign dataGroup_lo_lo_2503 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2504;
  assign dataGroup_lo_lo_2504 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2505;
  assign dataGroup_lo_lo_2505 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2506;
  assign dataGroup_lo_lo_2506 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2507;
  assign dataGroup_lo_lo_2507 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2508;
  assign dataGroup_lo_lo_2508 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2509;
  assign dataGroup_lo_lo_2509 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2510;
  assign dataGroup_lo_lo_2510 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2511;
  assign dataGroup_lo_lo_2511 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2512;
  assign dataGroup_lo_lo_2512 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2513;
  assign dataGroup_lo_lo_2513 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2514;
  assign dataGroup_lo_lo_2514 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2515;
  assign dataGroup_lo_lo_2515 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2516;
  assign dataGroup_lo_lo_2516 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2517;
  assign dataGroup_lo_lo_2517 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2518;
  assign dataGroup_lo_lo_2518 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2519;
  assign dataGroup_lo_lo_2519 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2520;
  assign dataGroup_lo_lo_2520 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2521;
  assign dataGroup_lo_lo_2521 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2522;
  assign dataGroup_lo_lo_2522 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2523;
  assign dataGroup_lo_lo_2523 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2524;
  assign dataGroup_lo_lo_2524 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2525;
  assign dataGroup_lo_lo_2525 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2526;
  assign dataGroup_lo_lo_2526 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2527;
  assign dataGroup_lo_lo_2527 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2528;
  assign dataGroup_lo_lo_2528 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2529;
  assign dataGroup_lo_lo_2529 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2530;
  assign dataGroup_lo_lo_2530 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2531;
  assign dataGroup_lo_lo_2531 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2532;
  assign dataGroup_lo_lo_2532 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2533;
  assign dataGroup_lo_lo_2533 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2534;
  assign dataGroup_lo_lo_2534 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2535;
  assign dataGroup_lo_lo_2535 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2536;
  assign dataGroup_lo_lo_2536 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2537;
  assign dataGroup_lo_lo_2537 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2538;
  assign dataGroup_lo_lo_2538 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2539;
  assign dataGroup_lo_lo_2539 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2540;
  assign dataGroup_lo_lo_2540 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2541;
  assign dataGroup_lo_lo_2541 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2542;
  assign dataGroup_lo_lo_2542 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2543;
  assign dataGroup_lo_lo_2543 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2544;
  assign dataGroup_lo_lo_2544 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2545;
  assign dataGroup_lo_lo_2545 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2546;
  assign dataGroup_lo_lo_2546 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2547;
  assign dataGroup_lo_lo_2547 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2548;
  assign dataGroup_lo_lo_2548 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2549;
  assign dataGroup_lo_lo_2549 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2550;
  assign dataGroup_lo_lo_2550 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2551;
  assign dataGroup_lo_lo_2551 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2552;
  assign dataGroup_lo_lo_2552 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2553;
  assign dataGroup_lo_lo_2553 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2554;
  assign dataGroup_lo_lo_2554 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2555;
  assign dataGroup_lo_lo_2555 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2556;
  assign dataGroup_lo_lo_2556 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2557;
  assign dataGroup_lo_lo_2557 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2558;
  assign dataGroup_lo_lo_2558 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2559;
  assign dataGroup_lo_lo_2559 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2560;
  assign dataGroup_lo_lo_2560 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2561;
  assign dataGroup_lo_lo_2561 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2562;
  assign dataGroup_lo_lo_2562 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2563;
  assign dataGroup_lo_lo_2563 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2564;
  assign dataGroup_lo_lo_2564 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2565;
  assign dataGroup_lo_lo_2565 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2566;
  assign dataGroup_lo_lo_2566 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2567;
  assign dataGroup_lo_lo_2567 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2568;
  assign dataGroup_lo_lo_2568 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2569;
  assign dataGroup_lo_lo_2569 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2570;
  assign dataGroup_lo_lo_2570 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2571;
  assign dataGroup_lo_lo_2571 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2572;
  assign dataGroup_lo_lo_2572 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2573;
  assign dataGroup_lo_lo_2573 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2574;
  assign dataGroup_lo_lo_2574 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2575;
  assign dataGroup_lo_lo_2575 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2576;
  assign dataGroup_lo_lo_2576 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2577;
  assign dataGroup_lo_lo_2577 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2578;
  assign dataGroup_lo_lo_2578 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2579;
  assign dataGroup_lo_lo_2579 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2580;
  assign dataGroup_lo_lo_2580 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2581;
  assign dataGroup_lo_lo_2581 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2582;
  assign dataGroup_lo_lo_2582 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2583;
  assign dataGroup_lo_lo_2583 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2584;
  assign dataGroup_lo_lo_2584 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2585;
  assign dataGroup_lo_lo_2585 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2586;
  assign dataGroup_lo_lo_2586 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2587;
  assign dataGroup_lo_lo_2587 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2588;
  assign dataGroup_lo_lo_2588 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2589;
  assign dataGroup_lo_lo_2589 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2590;
  assign dataGroup_lo_lo_2590 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2591;
  assign dataGroup_lo_lo_2591 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2592;
  assign dataGroup_lo_lo_2592 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2593;
  assign dataGroup_lo_lo_2593 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2594;
  assign dataGroup_lo_lo_2594 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2595;
  assign dataGroup_lo_lo_2595 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2596;
  assign dataGroup_lo_lo_2596 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2597;
  assign dataGroup_lo_lo_2597 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2598;
  assign dataGroup_lo_lo_2598 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2599;
  assign dataGroup_lo_lo_2599 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2600;
  assign dataGroup_lo_lo_2600 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2601;
  assign dataGroup_lo_lo_2601 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2602;
  assign dataGroup_lo_lo_2602 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2603;
  assign dataGroup_lo_lo_2603 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2604;
  assign dataGroup_lo_lo_2604 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2605;
  assign dataGroup_lo_lo_2605 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2606;
  assign dataGroup_lo_lo_2606 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2607;
  assign dataGroup_lo_lo_2607 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2608;
  assign dataGroup_lo_lo_2608 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2609;
  assign dataGroup_lo_lo_2609 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2610;
  assign dataGroup_lo_lo_2610 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2611;
  assign dataGroup_lo_lo_2611 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2612;
  assign dataGroup_lo_lo_2612 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2613;
  assign dataGroup_lo_lo_2613 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2614;
  assign dataGroup_lo_lo_2614 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2615;
  assign dataGroup_lo_lo_2615 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2616;
  assign dataGroup_lo_lo_2616 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2617;
  assign dataGroup_lo_lo_2617 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2618;
  assign dataGroup_lo_lo_2618 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2619;
  assign dataGroup_lo_lo_2619 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2620;
  assign dataGroup_lo_lo_2620 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2621;
  assign dataGroup_lo_lo_2621 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2622;
  assign dataGroup_lo_lo_2622 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2623;
  assign dataGroup_lo_lo_2623 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2624;
  assign dataGroup_lo_lo_2624 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2625;
  assign dataGroup_lo_lo_2625 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2626;
  assign dataGroup_lo_lo_2626 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2627;
  assign dataGroup_lo_lo_2627 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2628;
  assign dataGroup_lo_lo_2628 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2629;
  assign dataGroup_lo_lo_2629 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2630;
  assign dataGroup_lo_lo_2630 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2631;
  assign dataGroup_lo_lo_2631 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2632;
  assign dataGroup_lo_lo_2632 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2633;
  assign dataGroup_lo_lo_2633 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2634;
  assign dataGroup_lo_lo_2634 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2635;
  assign dataGroup_lo_lo_2635 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2636;
  assign dataGroup_lo_lo_2636 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2637;
  assign dataGroup_lo_lo_2637 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2638;
  assign dataGroup_lo_lo_2638 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2639;
  assign dataGroup_lo_lo_2639 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2640;
  assign dataGroup_lo_lo_2640 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2641;
  assign dataGroup_lo_lo_2641 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2642;
  assign dataGroup_lo_lo_2642 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2643;
  assign dataGroup_lo_lo_2643 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2644;
  assign dataGroup_lo_lo_2644 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2645;
  assign dataGroup_lo_lo_2645 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2646;
  assign dataGroup_lo_lo_2646 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2647;
  assign dataGroup_lo_lo_2647 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2648;
  assign dataGroup_lo_lo_2648 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2649;
  assign dataGroup_lo_lo_2649 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2650;
  assign dataGroup_lo_lo_2650 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2651;
  assign dataGroup_lo_lo_2651 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2652;
  assign dataGroup_lo_lo_2652 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2653;
  assign dataGroup_lo_lo_2653 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2654;
  assign dataGroup_lo_lo_2654 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2655;
  assign dataGroup_lo_lo_2655 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2656;
  assign dataGroup_lo_lo_2656 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2657;
  assign dataGroup_lo_lo_2657 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2658;
  assign dataGroup_lo_lo_2658 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2659;
  assign dataGroup_lo_lo_2659 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2660;
  assign dataGroup_lo_lo_2660 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2661;
  assign dataGroup_lo_lo_2661 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2662;
  assign dataGroup_lo_lo_2662 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2663;
  assign dataGroup_lo_lo_2663 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2664;
  assign dataGroup_lo_lo_2664 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2665;
  assign dataGroup_lo_lo_2665 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2666;
  assign dataGroup_lo_lo_2666 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2667;
  assign dataGroup_lo_lo_2667 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2668;
  assign dataGroup_lo_lo_2668 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2669;
  assign dataGroup_lo_lo_2669 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2670;
  assign dataGroup_lo_lo_2670 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2671;
  assign dataGroup_lo_lo_2671 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2672;
  assign dataGroup_lo_lo_2672 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2673;
  assign dataGroup_lo_lo_2673 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2674;
  assign dataGroup_lo_lo_2674 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2675;
  assign dataGroup_lo_lo_2675 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2676;
  assign dataGroup_lo_lo_2676 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2677;
  assign dataGroup_lo_lo_2677 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2678;
  assign dataGroup_lo_lo_2678 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2679;
  assign dataGroup_lo_lo_2679 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2680;
  assign dataGroup_lo_lo_2680 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2681;
  assign dataGroup_lo_lo_2681 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2682;
  assign dataGroup_lo_lo_2682 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2683;
  assign dataGroup_lo_lo_2683 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2684;
  assign dataGroup_lo_lo_2684 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2685;
  assign dataGroup_lo_lo_2685 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2686;
  assign dataGroup_lo_lo_2686 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2687;
  assign dataGroup_lo_lo_2687 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2688;
  assign dataGroup_lo_lo_2688 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2689;
  assign dataGroup_lo_lo_2689 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2690;
  assign dataGroup_lo_lo_2690 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2691;
  assign dataGroup_lo_lo_2691 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2692;
  assign dataGroup_lo_lo_2692 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2693;
  assign dataGroup_lo_lo_2693 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2694;
  assign dataGroup_lo_lo_2694 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2695;
  assign dataGroup_lo_lo_2695 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2696;
  assign dataGroup_lo_lo_2696 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2697;
  assign dataGroup_lo_lo_2697 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2698;
  assign dataGroup_lo_lo_2698 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2699;
  assign dataGroup_lo_lo_2699 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2700;
  assign dataGroup_lo_lo_2700 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2701;
  assign dataGroup_lo_lo_2701 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2702;
  assign dataGroup_lo_lo_2702 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2703;
  assign dataGroup_lo_lo_2703 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2704;
  assign dataGroup_lo_lo_2704 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2705;
  assign dataGroup_lo_lo_2705 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2706;
  assign dataGroup_lo_lo_2706 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2707;
  assign dataGroup_lo_lo_2707 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2708;
  assign dataGroup_lo_lo_2708 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2709;
  assign dataGroup_lo_lo_2709 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2710;
  assign dataGroup_lo_lo_2710 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2711;
  assign dataGroup_lo_lo_2711 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2712;
  assign dataGroup_lo_lo_2712 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2713;
  assign dataGroup_lo_lo_2713 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2714;
  assign dataGroup_lo_lo_2714 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2715;
  assign dataGroup_lo_lo_2715 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2716;
  assign dataGroup_lo_lo_2716 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2717;
  assign dataGroup_lo_lo_2717 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2718;
  assign dataGroup_lo_lo_2718 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2719;
  assign dataGroup_lo_lo_2719 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2720;
  assign dataGroup_lo_lo_2720 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2721;
  assign dataGroup_lo_lo_2721 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2722;
  assign dataGroup_lo_lo_2722 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2723;
  assign dataGroup_lo_lo_2723 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2724;
  assign dataGroup_lo_lo_2724 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2725;
  assign dataGroup_lo_lo_2725 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2726;
  assign dataGroup_lo_lo_2726 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2727;
  assign dataGroup_lo_lo_2727 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2728;
  assign dataGroup_lo_lo_2728 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2729;
  assign dataGroup_lo_lo_2729 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2730;
  assign dataGroup_lo_lo_2730 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2731;
  assign dataGroup_lo_lo_2731 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2732;
  assign dataGroup_lo_lo_2732 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2733;
  assign dataGroup_lo_lo_2733 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2734;
  assign dataGroup_lo_lo_2734 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2735;
  assign dataGroup_lo_lo_2735 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2736;
  assign dataGroup_lo_lo_2736 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2737;
  assign dataGroup_lo_lo_2737 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2738;
  assign dataGroup_lo_lo_2738 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2739;
  assign dataGroup_lo_lo_2739 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2740;
  assign dataGroup_lo_lo_2740 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2741;
  assign dataGroup_lo_lo_2741 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2742;
  assign dataGroup_lo_lo_2742 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2743;
  assign dataGroup_lo_lo_2743 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2744;
  assign dataGroup_lo_lo_2744 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2745;
  assign dataGroup_lo_lo_2745 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2746;
  assign dataGroup_lo_lo_2746 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2747;
  assign dataGroup_lo_lo_2747 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2748;
  assign dataGroup_lo_lo_2748 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2749;
  assign dataGroup_lo_lo_2749 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2750;
  assign dataGroup_lo_lo_2750 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2751;
  assign dataGroup_lo_lo_2751 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2752;
  assign dataGroup_lo_lo_2752 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2753;
  assign dataGroup_lo_lo_2753 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2754;
  assign dataGroup_lo_lo_2754 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2755;
  assign dataGroup_lo_lo_2755 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2756;
  assign dataGroup_lo_lo_2756 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2757;
  assign dataGroup_lo_lo_2757 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2758;
  assign dataGroup_lo_lo_2758 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2759;
  assign dataGroup_lo_lo_2759 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2760;
  assign dataGroup_lo_lo_2760 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2761;
  assign dataGroup_lo_lo_2761 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2762;
  assign dataGroup_lo_lo_2762 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2763;
  assign dataGroup_lo_lo_2763 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2764;
  assign dataGroup_lo_lo_2764 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2765;
  assign dataGroup_lo_lo_2765 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2766;
  assign dataGroup_lo_lo_2766 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2767;
  assign dataGroup_lo_lo_2767 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2768;
  assign dataGroup_lo_lo_2768 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2769;
  assign dataGroup_lo_lo_2769 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2770;
  assign dataGroup_lo_lo_2770 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2771;
  assign dataGroup_lo_lo_2771 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2772;
  assign dataGroup_lo_lo_2772 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2773;
  assign dataGroup_lo_lo_2773 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2774;
  assign dataGroup_lo_lo_2774 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2775;
  assign dataGroup_lo_lo_2775 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2776;
  assign dataGroup_lo_lo_2776 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2777;
  assign dataGroup_lo_lo_2777 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2778;
  assign dataGroup_lo_lo_2778 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2779;
  assign dataGroup_lo_lo_2779 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2780;
  assign dataGroup_lo_lo_2780 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2781;
  assign dataGroup_lo_lo_2781 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2782;
  assign dataGroup_lo_lo_2782 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2783;
  assign dataGroup_lo_lo_2783 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2784;
  assign dataGroup_lo_lo_2784 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2785;
  assign dataGroup_lo_lo_2785 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2786;
  assign dataGroup_lo_lo_2786 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2787;
  assign dataGroup_lo_lo_2787 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2788;
  assign dataGroup_lo_lo_2788 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2789;
  assign dataGroup_lo_lo_2789 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2790;
  assign dataGroup_lo_lo_2790 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2791;
  assign dataGroup_lo_lo_2791 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2792;
  assign dataGroup_lo_lo_2792 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2793;
  assign dataGroup_lo_lo_2793 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2794;
  assign dataGroup_lo_lo_2794 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2795;
  assign dataGroup_lo_lo_2795 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2796;
  assign dataGroup_lo_lo_2796 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2797;
  assign dataGroup_lo_lo_2797 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2798;
  assign dataGroup_lo_lo_2798 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2799;
  assign dataGroup_lo_lo_2799 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2800;
  assign dataGroup_lo_lo_2800 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2801;
  assign dataGroup_lo_lo_2801 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2802;
  assign dataGroup_lo_lo_2802 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2803;
  assign dataGroup_lo_lo_2803 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2804;
  assign dataGroup_lo_lo_2804 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2805;
  assign dataGroup_lo_lo_2805 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2806;
  assign dataGroup_lo_lo_2806 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2807;
  assign dataGroup_lo_lo_2807 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2808;
  assign dataGroup_lo_lo_2808 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2809;
  assign dataGroup_lo_lo_2809 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2810;
  assign dataGroup_lo_lo_2810 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2811;
  assign dataGroup_lo_lo_2811 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2812;
  assign dataGroup_lo_lo_2812 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2813;
  assign dataGroup_lo_lo_2813 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2814;
  assign dataGroup_lo_lo_2814 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2815;
  assign dataGroup_lo_lo_2815 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2816;
  assign dataGroup_lo_lo_2816 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2817;
  assign dataGroup_lo_lo_2817 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2818;
  assign dataGroup_lo_lo_2818 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2819;
  assign dataGroup_lo_lo_2819 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2820;
  assign dataGroup_lo_lo_2820 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2821;
  assign dataGroup_lo_lo_2821 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2822;
  assign dataGroup_lo_lo_2822 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2823;
  assign dataGroup_lo_lo_2823 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2824;
  assign dataGroup_lo_lo_2824 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2825;
  assign dataGroup_lo_lo_2825 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2826;
  assign dataGroup_lo_lo_2826 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2827;
  assign dataGroup_lo_lo_2827 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2828;
  assign dataGroup_lo_lo_2828 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2829;
  assign dataGroup_lo_lo_2829 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2830;
  assign dataGroup_lo_lo_2830 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2831;
  assign dataGroup_lo_lo_2831 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2832;
  assign dataGroup_lo_lo_2832 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2833;
  assign dataGroup_lo_lo_2833 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2834;
  assign dataGroup_lo_lo_2834 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2835;
  assign dataGroup_lo_lo_2835 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2836;
  assign dataGroup_lo_lo_2836 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2837;
  assign dataGroup_lo_lo_2837 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2838;
  assign dataGroup_lo_lo_2838 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2839;
  assign dataGroup_lo_lo_2839 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2840;
  assign dataGroup_lo_lo_2840 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2841;
  assign dataGroup_lo_lo_2841 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2842;
  assign dataGroup_lo_lo_2842 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2843;
  assign dataGroup_lo_lo_2843 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2844;
  assign dataGroup_lo_lo_2844 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2845;
  assign dataGroup_lo_lo_2845 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2846;
  assign dataGroup_lo_lo_2846 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2847;
  assign dataGroup_lo_lo_2847 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2848;
  assign dataGroup_lo_lo_2848 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2849;
  assign dataGroup_lo_lo_2849 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2850;
  assign dataGroup_lo_lo_2850 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2851;
  assign dataGroup_lo_lo_2851 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2852;
  assign dataGroup_lo_lo_2852 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2853;
  assign dataGroup_lo_lo_2853 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2854;
  assign dataGroup_lo_lo_2854 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2855;
  assign dataGroup_lo_lo_2855 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2856;
  assign dataGroup_lo_lo_2856 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2857;
  assign dataGroup_lo_lo_2857 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2858;
  assign dataGroup_lo_lo_2858 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2859;
  assign dataGroup_lo_lo_2859 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2860;
  assign dataGroup_lo_lo_2860 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2861;
  assign dataGroup_lo_lo_2861 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2862;
  assign dataGroup_lo_lo_2862 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2863;
  assign dataGroup_lo_lo_2863 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2864;
  assign dataGroup_lo_lo_2864 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2865;
  assign dataGroup_lo_lo_2865 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2866;
  assign dataGroup_lo_lo_2866 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2867;
  assign dataGroup_lo_lo_2867 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2868;
  assign dataGroup_lo_lo_2868 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2869;
  assign dataGroup_lo_lo_2869 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2870;
  assign dataGroup_lo_lo_2870 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2871;
  assign dataGroup_lo_lo_2871 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2872;
  assign dataGroup_lo_lo_2872 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2873;
  assign dataGroup_lo_lo_2873 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2874;
  assign dataGroup_lo_lo_2874 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2875;
  assign dataGroup_lo_lo_2875 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2876;
  assign dataGroup_lo_lo_2876 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2877;
  assign dataGroup_lo_lo_2877 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2878;
  assign dataGroup_lo_lo_2878 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2879;
  assign dataGroup_lo_lo_2879 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2880;
  assign dataGroup_lo_lo_2880 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2881;
  assign dataGroup_lo_lo_2881 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2882;
  assign dataGroup_lo_lo_2882 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2883;
  assign dataGroup_lo_lo_2883 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2884;
  assign dataGroup_lo_lo_2884 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2885;
  assign dataGroup_lo_lo_2885 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2886;
  assign dataGroup_lo_lo_2886 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2887;
  assign dataGroup_lo_lo_2887 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2888;
  assign dataGroup_lo_lo_2888 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2889;
  assign dataGroup_lo_lo_2889 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2890;
  assign dataGroup_lo_lo_2890 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2891;
  assign dataGroup_lo_lo_2891 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2892;
  assign dataGroup_lo_lo_2892 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2893;
  assign dataGroup_lo_lo_2893 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2894;
  assign dataGroup_lo_lo_2894 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2895;
  assign dataGroup_lo_lo_2895 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2896;
  assign dataGroup_lo_lo_2896 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2897;
  assign dataGroup_lo_lo_2897 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2898;
  assign dataGroup_lo_lo_2898 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2899;
  assign dataGroup_lo_lo_2899 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2900;
  assign dataGroup_lo_lo_2900 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2901;
  assign dataGroup_lo_lo_2901 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2902;
  assign dataGroup_lo_lo_2902 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2903;
  assign dataGroup_lo_lo_2903 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2904;
  assign dataGroup_lo_lo_2904 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2905;
  assign dataGroup_lo_lo_2905 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2906;
  assign dataGroup_lo_lo_2906 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2907;
  assign dataGroup_lo_lo_2907 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2908;
  assign dataGroup_lo_lo_2908 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2909;
  assign dataGroup_lo_lo_2909 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2910;
  assign dataGroup_lo_lo_2910 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2911;
  assign dataGroup_lo_lo_2911 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2912;
  assign dataGroup_lo_lo_2912 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2913;
  assign dataGroup_lo_lo_2913 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2914;
  assign dataGroup_lo_lo_2914 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2915;
  assign dataGroup_lo_lo_2915 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2916;
  assign dataGroup_lo_lo_2916 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2917;
  assign dataGroup_lo_lo_2917 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2918;
  assign dataGroup_lo_lo_2918 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2919;
  assign dataGroup_lo_lo_2919 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2920;
  assign dataGroup_lo_lo_2920 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2921;
  assign dataGroup_lo_lo_2921 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2922;
  assign dataGroup_lo_lo_2922 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2923;
  assign dataGroup_lo_lo_2923 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2924;
  assign dataGroup_lo_lo_2924 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2925;
  assign dataGroup_lo_lo_2925 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2926;
  assign dataGroup_lo_lo_2926 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2927;
  assign dataGroup_lo_lo_2927 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2928;
  assign dataGroup_lo_lo_2928 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2929;
  assign dataGroup_lo_lo_2929 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2930;
  assign dataGroup_lo_lo_2930 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2931;
  assign dataGroup_lo_lo_2931 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2932;
  assign dataGroup_lo_lo_2932 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2933;
  assign dataGroup_lo_lo_2933 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2934;
  assign dataGroup_lo_lo_2934 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2935;
  assign dataGroup_lo_lo_2935 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2936;
  assign dataGroup_lo_lo_2936 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2937;
  assign dataGroup_lo_lo_2937 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2938;
  assign dataGroup_lo_lo_2938 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2939;
  assign dataGroup_lo_lo_2939 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2940;
  assign dataGroup_lo_lo_2940 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2941;
  assign dataGroup_lo_lo_2941 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2942;
  assign dataGroup_lo_lo_2942 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2943;
  assign dataGroup_lo_lo_2943 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2944;
  assign dataGroup_lo_lo_2944 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2945;
  assign dataGroup_lo_lo_2945 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2946;
  assign dataGroup_lo_lo_2946 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2947;
  assign dataGroup_lo_lo_2947 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2948;
  assign dataGroup_lo_lo_2948 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2949;
  assign dataGroup_lo_lo_2949 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2950;
  assign dataGroup_lo_lo_2950 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2951;
  assign dataGroup_lo_lo_2951 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2952;
  assign dataGroup_lo_lo_2952 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2953;
  assign dataGroup_lo_lo_2953 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2954;
  assign dataGroup_lo_lo_2954 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2955;
  assign dataGroup_lo_lo_2955 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2956;
  assign dataGroup_lo_lo_2956 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2957;
  assign dataGroup_lo_lo_2957 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2958;
  assign dataGroup_lo_lo_2958 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2959;
  assign dataGroup_lo_lo_2959 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2960;
  assign dataGroup_lo_lo_2960 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2961;
  assign dataGroup_lo_lo_2961 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2962;
  assign dataGroup_lo_lo_2962 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2963;
  assign dataGroup_lo_lo_2963 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2964;
  assign dataGroup_lo_lo_2964 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2965;
  assign dataGroup_lo_lo_2965 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2966;
  assign dataGroup_lo_lo_2966 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2967;
  assign dataGroup_lo_lo_2967 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2968;
  assign dataGroup_lo_lo_2968 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2969;
  assign dataGroup_lo_lo_2969 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2970;
  assign dataGroup_lo_lo_2970 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2971;
  assign dataGroup_lo_lo_2971 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2972;
  assign dataGroup_lo_lo_2972 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2973;
  assign dataGroup_lo_lo_2973 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2974;
  assign dataGroup_lo_lo_2974 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2975;
  assign dataGroup_lo_lo_2975 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2976;
  assign dataGroup_lo_lo_2976 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2977;
  assign dataGroup_lo_lo_2977 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2978;
  assign dataGroup_lo_lo_2978 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2979;
  assign dataGroup_lo_lo_2979 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2980;
  assign dataGroup_lo_lo_2980 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2981;
  assign dataGroup_lo_lo_2981 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2982;
  assign dataGroup_lo_lo_2982 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2983;
  assign dataGroup_lo_lo_2983 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2984;
  assign dataGroup_lo_lo_2984 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2985;
  assign dataGroup_lo_lo_2985 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2986;
  assign dataGroup_lo_lo_2986 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2987;
  assign dataGroup_lo_lo_2987 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2988;
  assign dataGroup_lo_lo_2988 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2989;
  assign dataGroup_lo_lo_2989 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2990;
  assign dataGroup_lo_lo_2990 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2991;
  assign dataGroup_lo_lo_2991 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2992;
  assign dataGroup_lo_lo_2992 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2993;
  assign dataGroup_lo_lo_2993 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2994;
  assign dataGroup_lo_lo_2994 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2995;
  assign dataGroup_lo_lo_2995 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2996;
  assign dataGroup_lo_lo_2996 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2997;
  assign dataGroup_lo_lo_2997 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2998;
  assign dataGroup_lo_lo_2998 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_2999;
  assign dataGroup_lo_lo_2999 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3000;
  assign dataGroup_lo_lo_3000 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3001;
  assign dataGroup_lo_lo_3001 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3002;
  assign dataGroup_lo_lo_3002 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3003;
  assign dataGroup_lo_lo_3003 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3004;
  assign dataGroup_lo_lo_3004 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3005;
  assign dataGroup_lo_lo_3005 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3006;
  assign dataGroup_lo_lo_3006 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3007;
  assign dataGroup_lo_lo_3007 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3008;
  assign dataGroup_lo_lo_3008 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3009;
  assign dataGroup_lo_lo_3009 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3010;
  assign dataGroup_lo_lo_3010 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3011;
  assign dataGroup_lo_lo_3011 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3012;
  assign dataGroup_lo_lo_3012 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3013;
  assign dataGroup_lo_lo_3013 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3014;
  assign dataGroup_lo_lo_3014 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3015;
  assign dataGroup_lo_lo_3015 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3016;
  assign dataGroup_lo_lo_3016 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3017;
  assign dataGroup_lo_lo_3017 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3018;
  assign dataGroup_lo_lo_3018 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3019;
  assign dataGroup_lo_lo_3019 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3020;
  assign dataGroup_lo_lo_3020 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3021;
  assign dataGroup_lo_lo_3021 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3022;
  assign dataGroup_lo_lo_3022 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3023;
  assign dataGroup_lo_lo_3023 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3024;
  assign dataGroup_lo_lo_3024 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3025;
  assign dataGroup_lo_lo_3025 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3026;
  assign dataGroup_lo_lo_3026 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3027;
  assign dataGroup_lo_lo_3027 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3028;
  assign dataGroup_lo_lo_3028 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3029;
  assign dataGroup_lo_lo_3029 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3030;
  assign dataGroup_lo_lo_3030 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3031;
  assign dataGroup_lo_lo_3031 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3032;
  assign dataGroup_lo_lo_3032 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3033;
  assign dataGroup_lo_lo_3033 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3034;
  assign dataGroup_lo_lo_3034 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3035;
  assign dataGroup_lo_lo_3035 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3036;
  assign dataGroup_lo_lo_3036 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3037;
  assign dataGroup_lo_lo_3037 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3038;
  assign dataGroup_lo_lo_3038 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3039;
  assign dataGroup_lo_lo_3039 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3040;
  assign dataGroup_lo_lo_3040 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3041;
  assign dataGroup_lo_lo_3041 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3042;
  assign dataGroup_lo_lo_3042 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3043;
  assign dataGroup_lo_lo_3043 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3044;
  assign dataGroup_lo_lo_3044 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3045;
  assign dataGroup_lo_lo_3045 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3046;
  assign dataGroup_lo_lo_3046 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3047;
  assign dataGroup_lo_lo_3047 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3048;
  assign dataGroup_lo_lo_3048 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3049;
  assign dataGroup_lo_lo_3049 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3050;
  assign dataGroup_lo_lo_3050 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3051;
  assign dataGroup_lo_lo_3051 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3052;
  assign dataGroup_lo_lo_3052 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3053;
  assign dataGroup_lo_lo_3053 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3054;
  assign dataGroup_lo_lo_3054 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3055;
  assign dataGroup_lo_lo_3055 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3056;
  assign dataGroup_lo_lo_3056 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3057;
  assign dataGroup_lo_lo_3057 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3058;
  assign dataGroup_lo_lo_3058 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3059;
  assign dataGroup_lo_lo_3059 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3060;
  assign dataGroup_lo_lo_3060 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3061;
  assign dataGroup_lo_lo_3061 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3062;
  assign dataGroup_lo_lo_3062 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3063;
  assign dataGroup_lo_lo_3063 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3064;
  assign dataGroup_lo_lo_3064 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3065;
  assign dataGroup_lo_lo_3065 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3066;
  assign dataGroup_lo_lo_3066 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3067;
  assign dataGroup_lo_lo_3067 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3068;
  assign dataGroup_lo_lo_3068 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3069;
  assign dataGroup_lo_lo_3069 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3070;
  assign dataGroup_lo_lo_3070 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3071;
  assign dataGroup_lo_lo_3071 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3072;
  assign dataGroup_lo_lo_3072 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3073;
  assign dataGroup_lo_lo_3073 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3074;
  assign dataGroup_lo_lo_3074 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3075;
  assign dataGroup_lo_lo_3075 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3076;
  assign dataGroup_lo_lo_3076 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3077;
  assign dataGroup_lo_lo_3077 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3078;
  assign dataGroup_lo_lo_3078 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3079;
  assign dataGroup_lo_lo_3079 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3080;
  assign dataGroup_lo_lo_3080 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3081;
  assign dataGroup_lo_lo_3081 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3082;
  assign dataGroup_lo_lo_3082 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3083;
  assign dataGroup_lo_lo_3083 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3084;
  assign dataGroup_lo_lo_3084 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3085;
  assign dataGroup_lo_lo_3085 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3086;
  assign dataGroup_lo_lo_3086 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3087;
  assign dataGroup_lo_lo_3087 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3088;
  assign dataGroup_lo_lo_3088 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3089;
  assign dataGroup_lo_lo_3089 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3090;
  assign dataGroup_lo_lo_3090 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3091;
  assign dataGroup_lo_lo_3091 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3092;
  assign dataGroup_lo_lo_3092 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3093;
  assign dataGroup_lo_lo_3093 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3094;
  assign dataGroup_lo_lo_3094 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3095;
  assign dataGroup_lo_lo_3095 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3096;
  assign dataGroup_lo_lo_3096 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3097;
  assign dataGroup_lo_lo_3097 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3098;
  assign dataGroup_lo_lo_3098 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3099;
  assign dataGroup_lo_lo_3099 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3100;
  assign dataGroup_lo_lo_3100 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3101;
  assign dataGroup_lo_lo_3101 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3102;
  assign dataGroup_lo_lo_3102 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3103;
  assign dataGroup_lo_lo_3103 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3104;
  assign dataGroup_lo_lo_3104 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3105;
  assign dataGroup_lo_lo_3105 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3106;
  assign dataGroup_lo_lo_3106 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3107;
  assign dataGroup_lo_lo_3107 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3108;
  assign dataGroup_lo_lo_3108 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3109;
  assign dataGroup_lo_lo_3109 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3110;
  assign dataGroup_lo_lo_3110 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3111;
  assign dataGroup_lo_lo_3111 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3112;
  assign dataGroup_lo_lo_3112 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3113;
  assign dataGroup_lo_lo_3113 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3114;
  assign dataGroup_lo_lo_3114 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3115;
  assign dataGroup_lo_lo_3115 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3116;
  assign dataGroup_lo_lo_3116 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3117;
  assign dataGroup_lo_lo_3117 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3118;
  assign dataGroup_lo_lo_3118 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3119;
  assign dataGroup_lo_lo_3119 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3120;
  assign dataGroup_lo_lo_3120 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3121;
  assign dataGroup_lo_lo_3121 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3122;
  assign dataGroup_lo_lo_3122 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3123;
  assign dataGroup_lo_lo_3123 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3124;
  assign dataGroup_lo_lo_3124 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3125;
  assign dataGroup_lo_lo_3125 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3126;
  assign dataGroup_lo_lo_3126 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3127;
  assign dataGroup_lo_lo_3127 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3128;
  assign dataGroup_lo_lo_3128 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3129;
  assign dataGroup_lo_lo_3129 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3130;
  assign dataGroup_lo_lo_3130 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3131;
  assign dataGroup_lo_lo_3131 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3132;
  assign dataGroup_lo_lo_3132 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3133;
  assign dataGroup_lo_lo_3133 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3134;
  assign dataGroup_lo_lo_3134 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3135;
  assign dataGroup_lo_lo_3135 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3136;
  assign dataGroup_lo_lo_3136 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3137;
  assign dataGroup_lo_lo_3137 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3138;
  assign dataGroup_lo_lo_3138 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3139;
  assign dataGroup_lo_lo_3139 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3140;
  assign dataGroup_lo_lo_3140 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3141;
  assign dataGroup_lo_lo_3141 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3142;
  assign dataGroup_lo_lo_3142 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3143;
  assign dataGroup_lo_lo_3143 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3144;
  assign dataGroup_lo_lo_3144 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3145;
  assign dataGroup_lo_lo_3145 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3146;
  assign dataGroup_lo_lo_3146 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3147;
  assign dataGroup_lo_lo_3147 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3148;
  assign dataGroup_lo_lo_3148 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3149;
  assign dataGroup_lo_lo_3149 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3150;
  assign dataGroup_lo_lo_3150 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3151;
  assign dataGroup_lo_lo_3151 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3152;
  assign dataGroup_lo_lo_3152 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3153;
  assign dataGroup_lo_lo_3153 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3154;
  assign dataGroup_lo_lo_3154 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3155;
  assign dataGroup_lo_lo_3155 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3156;
  assign dataGroup_lo_lo_3156 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3157;
  assign dataGroup_lo_lo_3157 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3158;
  assign dataGroup_lo_lo_3158 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3159;
  assign dataGroup_lo_lo_3159 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3160;
  assign dataGroup_lo_lo_3160 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3161;
  assign dataGroup_lo_lo_3161 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3162;
  assign dataGroup_lo_lo_3162 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3163;
  assign dataGroup_lo_lo_3163 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3164;
  assign dataGroup_lo_lo_3164 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3165;
  assign dataGroup_lo_lo_3165 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3166;
  assign dataGroup_lo_lo_3166 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3167;
  assign dataGroup_lo_lo_3167 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3168;
  assign dataGroup_lo_lo_3168 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3169;
  assign dataGroup_lo_lo_3169 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3170;
  assign dataGroup_lo_lo_3170 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3171;
  assign dataGroup_lo_lo_3171 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3172;
  assign dataGroup_lo_lo_3172 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3173;
  assign dataGroup_lo_lo_3173 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3174;
  assign dataGroup_lo_lo_3174 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3175;
  assign dataGroup_lo_lo_3175 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3176;
  assign dataGroup_lo_lo_3176 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3177;
  assign dataGroup_lo_lo_3177 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3178;
  assign dataGroup_lo_lo_3178 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3179;
  assign dataGroup_lo_lo_3179 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3180;
  assign dataGroup_lo_lo_3180 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3181;
  assign dataGroup_lo_lo_3181 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3182;
  assign dataGroup_lo_lo_3182 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3183;
  assign dataGroup_lo_lo_3183 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3184;
  assign dataGroup_lo_lo_3184 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3185;
  assign dataGroup_lo_lo_3185 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3186;
  assign dataGroup_lo_lo_3186 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3187;
  assign dataGroup_lo_lo_3187 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3188;
  assign dataGroup_lo_lo_3188 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3189;
  assign dataGroup_lo_lo_3189 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3190;
  assign dataGroup_lo_lo_3190 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3191;
  assign dataGroup_lo_lo_3191 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3192;
  assign dataGroup_lo_lo_3192 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3193;
  assign dataGroup_lo_lo_3193 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3194;
  assign dataGroup_lo_lo_3194 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3195;
  assign dataGroup_lo_lo_3195 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3196;
  assign dataGroup_lo_lo_3196 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3197;
  assign dataGroup_lo_lo_3197 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3198;
  assign dataGroup_lo_lo_3198 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3199;
  assign dataGroup_lo_lo_3199 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3200;
  assign dataGroup_lo_lo_3200 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3201;
  assign dataGroup_lo_lo_3201 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3202;
  assign dataGroup_lo_lo_3202 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3203;
  assign dataGroup_lo_lo_3203 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3204;
  assign dataGroup_lo_lo_3204 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3205;
  assign dataGroup_lo_lo_3205 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3206;
  assign dataGroup_lo_lo_3206 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3207;
  assign dataGroup_lo_lo_3207 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3208;
  assign dataGroup_lo_lo_3208 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3209;
  assign dataGroup_lo_lo_3209 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3210;
  assign dataGroup_lo_lo_3210 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3211;
  assign dataGroup_lo_lo_3211 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3212;
  assign dataGroup_lo_lo_3212 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3213;
  assign dataGroup_lo_lo_3213 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3214;
  assign dataGroup_lo_lo_3214 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3215;
  assign dataGroup_lo_lo_3215 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3216;
  assign dataGroup_lo_lo_3216 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3217;
  assign dataGroup_lo_lo_3217 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3218;
  assign dataGroup_lo_lo_3218 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3219;
  assign dataGroup_lo_lo_3219 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3220;
  assign dataGroup_lo_lo_3220 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3221;
  assign dataGroup_lo_lo_3221 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3222;
  assign dataGroup_lo_lo_3222 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3223;
  assign dataGroup_lo_lo_3223 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3224;
  assign dataGroup_lo_lo_3224 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3225;
  assign dataGroup_lo_lo_3225 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3226;
  assign dataGroup_lo_lo_3226 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3227;
  assign dataGroup_lo_lo_3227 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3228;
  assign dataGroup_lo_lo_3228 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3229;
  assign dataGroup_lo_lo_3229 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3230;
  assign dataGroup_lo_lo_3230 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3231;
  assign dataGroup_lo_lo_3231 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3232;
  assign dataGroup_lo_lo_3232 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3233;
  assign dataGroup_lo_lo_3233 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3234;
  assign dataGroup_lo_lo_3234 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3235;
  assign dataGroup_lo_lo_3235 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3236;
  assign dataGroup_lo_lo_3236 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3237;
  assign dataGroup_lo_lo_3237 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3238;
  assign dataGroup_lo_lo_3238 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3239;
  assign dataGroup_lo_lo_3239 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3240;
  assign dataGroup_lo_lo_3240 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3241;
  assign dataGroup_lo_lo_3241 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3242;
  assign dataGroup_lo_lo_3242 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3243;
  assign dataGroup_lo_lo_3243 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3244;
  assign dataGroup_lo_lo_3244 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3245;
  assign dataGroup_lo_lo_3245 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3246;
  assign dataGroup_lo_lo_3246 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3247;
  assign dataGroup_lo_lo_3247 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3248;
  assign dataGroup_lo_lo_3248 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3249;
  assign dataGroup_lo_lo_3249 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3250;
  assign dataGroup_lo_lo_3250 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3251;
  assign dataGroup_lo_lo_3251 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3252;
  assign dataGroup_lo_lo_3252 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3253;
  assign dataGroup_lo_lo_3253 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3254;
  assign dataGroup_lo_lo_3254 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3255;
  assign dataGroup_lo_lo_3255 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3256;
  assign dataGroup_lo_lo_3256 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3257;
  assign dataGroup_lo_lo_3257 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3258;
  assign dataGroup_lo_lo_3258 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3259;
  assign dataGroup_lo_lo_3259 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3260;
  assign dataGroup_lo_lo_3260 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3261;
  assign dataGroup_lo_lo_3261 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3262;
  assign dataGroup_lo_lo_3262 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3263;
  assign dataGroup_lo_lo_3263 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3264;
  assign dataGroup_lo_lo_3264 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3265;
  assign dataGroup_lo_lo_3265 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3266;
  assign dataGroup_lo_lo_3266 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3267;
  assign dataGroup_lo_lo_3267 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3268;
  assign dataGroup_lo_lo_3268 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3269;
  assign dataGroup_lo_lo_3269 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3270;
  assign dataGroup_lo_lo_3270 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3271;
  assign dataGroup_lo_lo_3271 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3272;
  assign dataGroup_lo_lo_3272 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3273;
  assign dataGroup_lo_lo_3273 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3274;
  assign dataGroup_lo_lo_3274 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3275;
  assign dataGroup_lo_lo_3275 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3276;
  assign dataGroup_lo_lo_3276 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3277;
  assign dataGroup_lo_lo_3277 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3278;
  assign dataGroup_lo_lo_3278 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3279;
  assign dataGroup_lo_lo_3279 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3280;
  assign dataGroup_lo_lo_3280 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3281;
  assign dataGroup_lo_lo_3281 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3282;
  assign dataGroup_lo_lo_3282 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3283;
  assign dataGroup_lo_lo_3283 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3284;
  assign dataGroup_lo_lo_3284 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3285;
  assign dataGroup_lo_lo_3285 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3286;
  assign dataGroup_lo_lo_3286 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3287;
  assign dataGroup_lo_lo_3287 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3288;
  assign dataGroup_lo_lo_3288 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3289;
  assign dataGroup_lo_lo_3289 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3290;
  assign dataGroup_lo_lo_3290 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3291;
  assign dataGroup_lo_lo_3291 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3292;
  assign dataGroup_lo_lo_3292 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3293;
  assign dataGroup_lo_lo_3293 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3294;
  assign dataGroup_lo_lo_3294 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3295;
  assign dataGroup_lo_lo_3295 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3296;
  assign dataGroup_lo_lo_3296 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3297;
  assign dataGroup_lo_lo_3297 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3298;
  assign dataGroup_lo_lo_3298 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3299;
  assign dataGroup_lo_lo_3299 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3300;
  assign dataGroup_lo_lo_3300 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3301;
  assign dataGroup_lo_lo_3301 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3302;
  assign dataGroup_lo_lo_3302 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3303;
  assign dataGroup_lo_lo_3303 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3304;
  assign dataGroup_lo_lo_3304 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3305;
  assign dataGroup_lo_lo_3305 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3306;
  assign dataGroup_lo_lo_3306 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3307;
  assign dataGroup_lo_lo_3307 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3308;
  assign dataGroup_lo_lo_3308 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3309;
  assign dataGroup_lo_lo_3309 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3310;
  assign dataGroup_lo_lo_3310 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3311;
  assign dataGroup_lo_lo_3311 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3312;
  assign dataGroup_lo_lo_3312 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3313;
  assign dataGroup_lo_lo_3313 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3314;
  assign dataGroup_lo_lo_3314 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3315;
  assign dataGroup_lo_lo_3315 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3316;
  assign dataGroup_lo_lo_3316 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3317;
  assign dataGroup_lo_lo_3317 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3318;
  assign dataGroup_lo_lo_3318 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3319;
  assign dataGroup_lo_lo_3319 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3320;
  assign dataGroup_lo_lo_3320 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3321;
  assign dataGroup_lo_lo_3321 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3322;
  assign dataGroup_lo_lo_3322 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3323;
  assign dataGroup_lo_lo_3323 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3324;
  assign dataGroup_lo_lo_3324 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3325;
  assign dataGroup_lo_lo_3325 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3326;
  assign dataGroup_lo_lo_3326 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3327;
  assign dataGroup_lo_lo_3327 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3328;
  assign dataGroup_lo_lo_3328 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3329;
  assign dataGroup_lo_lo_3329 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3330;
  assign dataGroup_lo_lo_3330 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3331;
  assign dataGroup_lo_lo_3331 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3332;
  assign dataGroup_lo_lo_3332 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3333;
  assign dataGroup_lo_lo_3333 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3334;
  assign dataGroup_lo_lo_3334 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3335;
  assign dataGroup_lo_lo_3335 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3336;
  assign dataGroup_lo_lo_3336 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3337;
  assign dataGroup_lo_lo_3337 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3338;
  assign dataGroup_lo_lo_3338 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3339;
  assign dataGroup_lo_lo_3339 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3340;
  assign dataGroup_lo_lo_3340 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3341;
  assign dataGroup_lo_lo_3341 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3342;
  assign dataGroup_lo_lo_3342 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3343;
  assign dataGroup_lo_lo_3343 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3344;
  assign dataGroup_lo_lo_3344 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3345;
  assign dataGroup_lo_lo_3345 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3346;
  assign dataGroup_lo_lo_3346 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3347;
  assign dataGroup_lo_lo_3347 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3348;
  assign dataGroup_lo_lo_3348 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3349;
  assign dataGroup_lo_lo_3349 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3350;
  assign dataGroup_lo_lo_3350 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3351;
  assign dataGroup_lo_lo_3351 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3352;
  assign dataGroup_lo_lo_3352 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3353;
  assign dataGroup_lo_lo_3353 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3354;
  assign dataGroup_lo_lo_3354 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3355;
  assign dataGroup_lo_lo_3355 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3356;
  assign dataGroup_lo_lo_3356 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3357;
  assign dataGroup_lo_lo_3357 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3358;
  assign dataGroup_lo_lo_3358 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3359;
  assign dataGroup_lo_lo_3359 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3360;
  assign dataGroup_lo_lo_3360 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3361;
  assign dataGroup_lo_lo_3361 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3362;
  assign dataGroup_lo_lo_3362 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3363;
  assign dataGroup_lo_lo_3363 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3364;
  assign dataGroup_lo_lo_3364 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3365;
  assign dataGroup_lo_lo_3365 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3366;
  assign dataGroup_lo_lo_3366 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3367;
  assign dataGroup_lo_lo_3367 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3368;
  assign dataGroup_lo_lo_3368 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3369;
  assign dataGroup_lo_lo_3369 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3370;
  assign dataGroup_lo_lo_3370 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3371;
  assign dataGroup_lo_lo_3371 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3372;
  assign dataGroup_lo_lo_3372 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3373;
  assign dataGroup_lo_lo_3373 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3374;
  assign dataGroup_lo_lo_3374 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3375;
  assign dataGroup_lo_lo_3375 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3376;
  assign dataGroup_lo_lo_3376 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3377;
  assign dataGroup_lo_lo_3377 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3378;
  assign dataGroup_lo_lo_3378 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3379;
  assign dataGroup_lo_lo_3379 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3380;
  assign dataGroup_lo_lo_3380 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3381;
  assign dataGroup_lo_lo_3381 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3382;
  assign dataGroup_lo_lo_3382 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3383;
  assign dataGroup_lo_lo_3383 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3384;
  assign dataGroup_lo_lo_3384 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3385;
  assign dataGroup_lo_lo_3385 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3386;
  assign dataGroup_lo_lo_3386 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3387;
  assign dataGroup_lo_lo_3387 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3388;
  assign dataGroup_lo_lo_3388 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3389;
  assign dataGroup_lo_lo_3389 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3390;
  assign dataGroup_lo_lo_3390 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3391;
  assign dataGroup_lo_lo_3391 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3392;
  assign dataGroup_lo_lo_3392 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3393;
  assign dataGroup_lo_lo_3393 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3394;
  assign dataGroup_lo_lo_3394 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3395;
  assign dataGroup_lo_lo_3395 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3396;
  assign dataGroup_lo_lo_3396 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3397;
  assign dataGroup_lo_lo_3397 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3398;
  assign dataGroup_lo_lo_3398 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3399;
  assign dataGroup_lo_lo_3399 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3400;
  assign dataGroup_lo_lo_3400 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3401;
  assign dataGroup_lo_lo_3401 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3402;
  assign dataGroup_lo_lo_3402 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3403;
  assign dataGroup_lo_lo_3403 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3404;
  assign dataGroup_lo_lo_3404 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3405;
  assign dataGroup_lo_lo_3405 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3406;
  assign dataGroup_lo_lo_3406 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3407;
  assign dataGroup_lo_lo_3407 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3408;
  assign dataGroup_lo_lo_3408 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3409;
  assign dataGroup_lo_lo_3409 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3410;
  assign dataGroup_lo_lo_3410 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3411;
  assign dataGroup_lo_lo_3411 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3412;
  assign dataGroup_lo_lo_3412 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3413;
  assign dataGroup_lo_lo_3413 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3414;
  assign dataGroup_lo_lo_3414 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3415;
  assign dataGroup_lo_lo_3415 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3416;
  assign dataGroup_lo_lo_3416 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3417;
  assign dataGroup_lo_lo_3417 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3418;
  assign dataGroup_lo_lo_3418 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3419;
  assign dataGroup_lo_lo_3419 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3420;
  assign dataGroup_lo_lo_3420 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3421;
  assign dataGroup_lo_lo_3421 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3422;
  assign dataGroup_lo_lo_3422 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3423;
  assign dataGroup_lo_lo_3423 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3424;
  assign dataGroup_lo_lo_3424 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3425;
  assign dataGroup_lo_lo_3425 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3426;
  assign dataGroup_lo_lo_3426 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3427;
  assign dataGroup_lo_lo_3427 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3428;
  assign dataGroup_lo_lo_3428 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3429;
  assign dataGroup_lo_lo_3429 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3430;
  assign dataGroup_lo_lo_3430 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3431;
  assign dataGroup_lo_lo_3431 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3432;
  assign dataGroup_lo_lo_3432 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3433;
  assign dataGroup_lo_lo_3433 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3434;
  assign dataGroup_lo_lo_3434 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3435;
  assign dataGroup_lo_lo_3435 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3436;
  assign dataGroup_lo_lo_3436 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3437;
  assign dataGroup_lo_lo_3437 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3438;
  assign dataGroup_lo_lo_3438 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3439;
  assign dataGroup_lo_lo_3439 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3440;
  assign dataGroup_lo_lo_3440 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3441;
  assign dataGroup_lo_lo_3441 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3442;
  assign dataGroup_lo_lo_3442 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3443;
  assign dataGroup_lo_lo_3443 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3444;
  assign dataGroup_lo_lo_3444 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3445;
  assign dataGroup_lo_lo_3445 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3446;
  assign dataGroup_lo_lo_3446 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3447;
  assign dataGroup_lo_lo_3447 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3448;
  assign dataGroup_lo_lo_3448 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3449;
  assign dataGroup_lo_lo_3449 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3450;
  assign dataGroup_lo_lo_3450 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3451;
  assign dataGroup_lo_lo_3451 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3452;
  assign dataGroup_lo_lo_3452 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3453;
  assign dataGroup_lo_lo_3453 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3454;
  assign dataGroup_lo_lo_3454 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3455;
  assign dataGroup_lo_lo_3455 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3456;
  assign dataGroup_lo_lo_3456 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3457;
  assign dataGroup_lo_lo_3457 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3458;
  assign dataGroup_lo_lo_3458 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3459;
  assign dataGroup_lo_lo_3459 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3460;
  assign dataGroup_lo_lo_3460 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3461;
  assign dataGroup_lo_lo_3461 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3462;
  assign dataGroup_lo_lo_3462 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3463;
  assign dataGroup_lo_lo_3463 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3464;
  assign dataGroup_lo_lo_3464 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3465;
  assign dataGroup_lo_lo_3465 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3466;
  assign dataGroup_lo_lo_3466 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3467;
  assign dataGroup_lo_lo_3467 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3468;
  assign dataGroup_lo_lo_3468 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3469;
  assign dataGroup_lo_lo_3469 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3470;
  assign dataGroup_lo_lo_3470 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3471;
  assign dataGroup_lo_lo_3471 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3472;
  assign dataGroup_lo_lo_3472 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3473;
  assign dataGroup_lo_lo_3473 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3474;
  assign dataGroup_lo_lo_3474 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3475;
  assign dataGroup_lo_lo_3475 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3476;
  assign dataGroup_lo_lo_3476 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3477;
  assign dataGroup_lo_lo_3477 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3478;
  assign dataGroup_lo_lo_3478 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3479;
  assign dataGroup_lo_lo_3479 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3480;
  assign dataGroup_lo_lo_3480 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3481;
  assign dataGroup_lo_lo_3481 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3482;
  assign dataGroup_lo_lo_3482 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3483;
  assign dataGroup_lo_lo_3483 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3484;
  assign dataGroup_lo_lo_3484 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3485;
  assign dataGroup_lo_lo_3485 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3486;
  assign dataGroup_lo_lo_3486 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3487;
  assign dataGroup_lo_lo_3487 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3488;
  assign dataGroup_lo_lo_3488 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3489;
  assign dataGroup_lo_lo_3489 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3490;
  assign dataGroup_lo_lo_3490 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3491;
  assign dataGroup_lo_lo_3491 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3492;
  assign dataGroup_lo_lo_3492 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3493;
  assign dataGroup_lo_lo_3493 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3494;
  assign dataGroup_lo_lo_3494 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3495;
  assign dataGroup_lo_lo_3495 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3496;
  assign dataGroup_lo_lo_3496 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3497;
  assign dataGroup_lo_lo_3497 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3498;
  assign dataGroup_lo_lo_3498 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3499;
  assign dataGroup_lo_lo_3499 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3500;
  assign dataGroup_lo_lo_3500 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3501;
  assign dataGroup_lo_lo_3501 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3502;
  assign dataGroup_lo_lo_3502 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3503;
  assign dataGroup_lo_lo_3503 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3504;
  assign dataGroup_lo_lo_3504 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3505;
  assign dataGroup_lo_lo_3505 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3506;
  assign dataGroup_lo_lo_3506 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3507;
  assign dataGroup_lo_lo_3507 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3508;
  assign dataGroup_lo_lo_3508 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3509;
  assign dataGroup_lo_lo_3509 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3510;
  assign dataGroup_lo_lo_3510 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3511;
  assign dataGroup_lo_lo_3511 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3512;
  assign dataGroup_lo_lo_3512 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3513;
  assign dataGroup_lo_lo_3513 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3514;
  assign dataGroup_lo_lo_3514 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3515;
  assign dataGroup_lo_lo_3515 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3516;
  assign dataGroup_lo_lo_3516 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3517;
  assign dataGroup_lo_lo_3517 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3518;
  assign dataGroup_lo_lo_3518 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3519;
  assign dataGroup_lo_lo_3519 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3520;
  assign dataGroup_lo_lo_3520 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3521;
  assign dataGroup_lo_lo_3521 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3522;
  assign dataGroup_lo_lo_3522 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3523;
  assign dataGroup_lo_lo_3523 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3524;
  assign dataGroup_lo_lo_3524 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3525;
  assign dataGroup_lo_lo_3525 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3526;
  assign dataGroup_lo_lo_3526 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3527;
  assign dataGroup_lo_lo_3527 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3528;
  assign dataGroup_lo_lo_3528 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3529;
  assign dataGroup_lo_lo_3529 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3530;
  assign dataGroup_lo_lo_3530 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3531;
  assign dataGroup_lo_lo_3531 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3532;
  assign dataGroup_lo_lo_3532 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3533;
  assign dataGroup_lo_lo_3533 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3534;
  assign dataGroup_lo_lo_3534 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3535;
  assign dataGroup_lo_lo_3535 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3536;
  assign dataGroup_lo_lo_3536 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3537;
  assign dataGroup_lo_lo_3537 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3538;
  assign dataGroup_lo_lo_3538 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3539;
  assign dataGroup_lo_lo_3539 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3540;
  assign dataGroup_lo_lo_3540 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3541;
  assign dataGroup_lo_lo_3541 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3542;
  assign dataGroup_lo_lo_3542 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3543;
  assign dataGroup_lo_lo_3543 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3544;
  assign dataGroup_lo_lo_3544 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3545;
  assign dataGroup_lo_lo_3545 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3546;
  assign dataGroup_lo_lo_3546 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3547;
  assign dataGroup_lo_lo_3547 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3548;
  assign dataGroup_lo_lo_3548 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3549;
  assign dataGroup_lo_lo_3549 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3550;
  assign dataGroup_lo_lo_3550 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3551;
  assign dataGroup_lo_lo_3551 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3552;
  assign dataGroup_lo_lo_3552 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3553;
  assign dataGroup_lo_lo_3553 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3554;
  assign dataGroup_lo_lo_3554 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3555;
  assign dataGroup_lo_lo_3555 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3556;
  assign dataGroup_lo_lo_3556 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3557;
  assign dataGroup_lo_lo_3557 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3558;
  assign dataGroup_lo_lo_3558 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3559;
  assign dataGroup_lo_lo_3559 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3560;
  assign dataGroup_lo_lo_3560 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3561;
  assign dataGroup_lo_lo_3561 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3562;
  assign dataGroup_lo_lo_3562 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3563;
  assign dataGroup_lo_lo_3563 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3564;
  assign dataGroup_lo_lo_3564 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3565;
  assign dataGroup_lo_lo_3565 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3566;
  assign dataGroup_lo_lo_3566 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3567;
  assign dataGroup_lo_lo_3567 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3568;
  assign dataGroup_lo_lo_3568 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3569;
  assign dataGroup_lo_lo_3569 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3570;
  assign dataGroup_lo_lo_3570 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3571;
  assign dataGroup_lo_lo_3571 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3572;
  assign dataGroup_lo_lo_3572 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3573;
  assign dataGroup_lo_lo_3573 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3574;
  assign dataGroup_lo_lo_3574 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3575;
  assign dataGroup_lo_lo_3575 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3576;
  assign dataGroup_lo_lo_3576 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3577;
  assign dataGroup_lo_lo_3577 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3578;
  assign dataGroup_lo_lo_3578 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3579;
  assign dataGroup_lo_lo_3579 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3580;
  assign dataGroup_lo_lo_3580 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3581;
  assign dataGroup_lo_lo_3581 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3582;
  assign dataGroup_lo_lo_3582 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3583;
  assign dataGroup_lo_lo_3583 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3584;
  assign dataGroup_lo_lo_3584 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3585;
  assign dataGroup_lo_lo_3585 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3586;
  assign dataGroup_lo_lo_3586 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3587;
  assign dataGroup_lo_lo_3587 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3588;
  assign dataGroup_lo_lo_3588 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3589;
  assign dataGroup_lo_lo_3589 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3590;
  assign dataGroup_lo_lo_3590 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3591;
  assign dataGroup_lo_lo_3591 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3592;
  assign dataGroup_lo_lo_3592 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3593;
  assign dataGroup_lo_lo_3593 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3594;
  assign dataGroup_lo_lo_3594 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3595;
  assign dataGroup_lo_lo_3595 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3596;
  assign dataGroup_lo_lo_3596 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3597;
  assign dataGroup_lo_lo_3597 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3598;
  assign dataGroup_lo_lo_3598 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3599;
  assign dataGroup_lo_lo_3599 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3600;
  assign dataGroup_lo_lo_3600 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3601;
  assign dataGroup_lo_lo_3601 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3602;
  assign dataGroup_lo_lo_3602 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3603;
  assign dataGroup_lo_lo_3603 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3604;
  assign dataGroup_lo_lo_3604 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3605;
  assign dataGroup_lo_lo_3605 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3606;
  assign dataGroup_lo_lo_3606 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3607;
  assign dataGroup_lo_lo_3607 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3608;
  assign dataGroup_lo_lo_3608 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3609;
  assign dataGroup_lo_lo_3609 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3610;
  assign dataGroup_lo_lo_3610 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3611;
  assign dataGroup_lo_lo_3611 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3612;
  assign dataGroup_lo_lo_3612 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3613;
  assign dataGroup_lo_lo_3613 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3614;
  assign dataGroup_lo_lo_3614 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3615;
  assign dataGroup_lo_lo_3615 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3616;
  assign dataGroup_lo_lo_3616 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3617;
  assign dataGroup_lo_lo_3617 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3618;
  assign dataGroup_lo_lo_3618 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3619;
  assign dataGroup_lo_lo_3619 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3620;
  assign dataGroup_lo_lo_3620 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3621;
  assign dataGroup_lo_lo_3621 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3622;
  assign dataGroup_lo_lo_3622 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3623;
  assign dataGroup_lo_lo_3623 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3624;
  assign dataGroup_lo_lo_3624 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3625;
  assign dataGroup_lo_lo_3625 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3626;
  assign dataGroup_lo_lo_3626 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3627;
  assign dataGroup_lo_lo_3627 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3628;
  assign dataGroup_lo_lo_3628 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3629;
  assign dataGroup_lo_lo_3629 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3630;
  assign dataGroup_lo_lo_3630 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3631;
  assign dataGroup_lo_lo_3631 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3632;
  assign dataGroup_lo_lo_3632 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3633;
  assign dataGroup_lo_lo_3633 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3634;
  assign dataGroup_lo_lo_3634 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3635;
  assign dataGroup_lo_lo_3635 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3636;
  assign dataGroup_lo_lo_3636 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3637;
  assign dataGroup_lo_lo_3637 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3638;
  assign dataGroup_lo_lo_3638 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3639;
  assign dataGroup_lo_lo_3639 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3640;
  assign dataGroup_lo_lo_3640 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3641;
  assign dataGroup_lo_lo_3641 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3642;
  assign dataGroup_lo_lo_3642 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3643;
  assign dataGroup_lo_lo_3643 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3644;
  assign dataGroup_lo_lo_3644 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3645;
  assign dataGroup_lo_lo_3645 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3646;
  assign dataGroup_lo_lo_3646 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3647;
  assign dataGroup_lo_lo_3647 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3648;
  assign dataGroup_lo_lo_3648 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3649;
  assign dataGroup_lo_lo_3649 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3650;
  assign dataGroup_lo_lo_3650 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3651;
  assign dataGroup_lo_lo_3651 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3652;
  assign dataGroup_lo_lo_3652 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3653;
  assign dataGroup_lo_lo_3653 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3654;
  assign dataGroup_lo_lo_3654 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3655;
  assign dataGroup_lo_lo_3655 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3656;
  assign dataGroup_lo_lo_3656 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3657;
  assign dataGroup_lo_lo_3657 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3658;
  assign dataGroup_lo_lo_3658 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3659;
  assign dataGroup_lo_lo_3659 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3660;
  assign dataGroup_lo_lo_3660 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3661;
  assign dataGroup_lo_lo_3661 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3662;
  assign dataGroup_lo_lo_3662 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3663;
  assign dataGroup_lo_lo_3663 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3664;
  assign dataGroup_lo_lo_3664 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3665;
  assign dataGroup_lo_lo_3665 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3666;
  assign dataGroup_lo_lo_3666 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3667;
  assign dataGroup_lo_lo_3667 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3668;
  assign dataGroup_lo_lo_3668 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3669;
  assign dataGroup_lo_lo_3669 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3670;
  assign dataGroup_lo_lo_3670 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3671;
  assign dataGroup_lo_lo_3671 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3672;
  assign dataGroup_lo_lo_3672 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3673;
  assign dataGroup_lo_lo_3673 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3674;
  assign dataGroup_lo_lo_3674 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3675;
  assign dataGroup_lo_lo_3675 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3676;
  assign dataGroup_lo_lo_3676 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3677;
  assign dataGroup_lo_lo_3677 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3678;
  assign dataGroup_lo_lo_3678 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3679;
  assign dataGroup_lo_lo_3679 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3680;
  assign dataGroup_lo_lo_3680 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3681;
  assign dataGroup_lo_lo_3681 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3682;
  assign dataGroup_lo_lo_3682 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3683;
  assign dataGroup_lo_lo_3683 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3684;
  assign dataGroup_lo_lo_3684 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3685;
  assign dataGroup_lo_lo_3685 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3686;
  assign dataGroup_lo_lo_3686 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3687;
  assign dataGroup_lo_lo_3687 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3688;
  assign dataGroup_lo_lo_3688 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3689;
  assign dataGroup_lo_lo_3689 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3690;
  assign dataGroup_lo_lo_3690 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3691;
  assign dataGroup_lo_lo_3691 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3692;
  assign dataGroup_lo_lo_3692 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3693;
  assign dataGroup_lo_lo_3693 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3694;
  assign dataGroup_lo_lo_3694 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3695;
  assign dataGroup_lo_lo_3695 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3696;
  assign dataGroup_lo_lo_3696 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3697;
  assign dataGroup_lo_lo_3697 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3698;
  assign dataGroup_lo_lo_3698 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3699;
  assign dataGroup_lo_lo_3699 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3700;
  assign dataGroup_lo_lo_3700 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3701;
  assign dataGroup_lo_lo_3701 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3702;
  assign dataGroup_lo_lo_3702 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3703;
  assign dataGroup_lo_lo_3703 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3704;
  assign dataGroup_lo_lo_3704 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3705;
  assign dataGroup_lo_lo_3705 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3706;
  assign dataGroup_lo_lo_3706 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3707;
  assign dataGroup_lo_lo_3707 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3708;
  assign dataGroup_lo_lo_3708 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3709;
  assign dataGroup_lo_lo_3709 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3710;
  assign dataGroup_lo_lo_3710 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3711;
  assign dataGroup_lo_lo_3711 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3712;
  assign dataGroup_lo_lo_3712 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3713;
  assign dataGroup_lo_lo_3713 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3714;
  assign dataGroup_lo_lo_3714 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3715;
  assign dataGroup_lo_lo_3715 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3716;
  assign dataGroup_lo_lo_3716 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3717;
  assign dataGroup_lo_lo_3717 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3718;
  assign dataGroup_lo_lo_3718 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3719;
  assign dataGroup_lo_lo_3719 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3720;
  assign dataGroup_lo_lo_3720 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3721;
  assign dataGroup_lo_lo_3721 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3722;
  assign dataGroup_lo_lo_3722 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3723;
  assign dataGroup_lo_lo_3723 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3724;
  assign dataGroup_lo_lo_3724 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3725;
  assign dataGroup_lo_lo_3725 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3726;
  assign dataGroup_lo_lo_3726 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3727;
  assign dataGroup_lo_lo_3727 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3728;
  assign dataGroup_lo_lo_3728 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3729;
  assign dataGroup_lo_lo_3729 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3730;
  assign dataGroup_lo_lo_3730 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3731;
  assign dataGroup_lo_lo_3731 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3732;
  assign dataGroup_lo_lo_3732 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3733;
  assign dataGroup_lo_lo_3733 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3734;
  assign dataGroup_lo_lo_3734 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3735;
  assign dataGroup_lo_lo_3735 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3736;
  assign dataGroup_lo_lo_3736 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3737;
  assign dataGroup_lo_lo_3737 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3738;
  assign dataGroup_lo_lo_3738 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3739;
  assign dataGroup_lo_lo_3739 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3740;
  assign dataGroup_lo_lo_3740 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3741;
  assign dataGroup_lo_lo_3741 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3742;
  assign dataGroup_lo_lo_3742 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3743;
  assign dataGroup_lo_lo_3743 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3744;
  assign dataGroup_lo_lo_3744 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3745;
  assign dataGroup_lo_lo_3745 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3746;
  assign dataGroup_lo_lo_3746 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3747;
  assign dataGroup_lo_lo_3747 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3748;
  assign dataGroup_lo_lo_3748 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3749;
  assign dataGroup_lo_lo_3749 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3750;
  assign dataGroup_lo_lo_3750 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3751;
  assign dataGroup_lo_lo_3751 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3752;
  assign dataGroup_lo_lo_3752 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3753;
  assign dataGroup_lo_lo_3753 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3754;
  assign dataGroup_lo_lo_3754 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3755;
  assign dataGroup_lo_lo_3755 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3756;
  assign dataGroup_lo_lo_3756 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3757;
  assign dataGroup_lo_lo_3757 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3758;
  assign dataGroup_lo_lo_3758 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3759;
  assign dataGroup_lo_lo_3759 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3760;
  assign dataGroup_lo_lo_3760 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3761;
  assign dataGroup_lo_lo_3761 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3762;
  assign dataGroup_lo_lo_3762 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3763;
  assign dataGroup_lo_lo_3763 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3764;
  assign dataGroup_lo_lo_3764 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3765;
  assign dataGroup_lo_lo_3765 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3766;
  assign dataGroup_lo_lo_3766 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3767;
  assign dataGroup_lo_lo_3767 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3768;
  assign dataGroup_lo_lo_3768 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3769;
  assign dataGroup_lo_lo_3769 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3770;
  assign dataGroup_lo_lo_3770 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3771;
  assign dataGroup_lo_lo_3771 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3772;
  assign dataGroup_lo_lo_3772 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3773;
  assign dataGroup_lo_lo_3773 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3774;
  assign dataGroup_lo_lo_3774 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3775;
  assign dataGroup_lo_lo_3775 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3776;
  assign dataGroup_lo_lo_3776 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3777;
  assign dataGroup_lo_lo_3777 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3778;
  assign dataGroup_lo_lo_3778 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3779;
  assign dataGroup_lo_lo_3779 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3780;
  assign dataGroup_lo_lo_3780 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3781;
  assign dataGroup_lo_lo_3781 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3782;
  assign dataGroup_lo_lo_3782 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3783;
  assign dataGroup_lo_lo_3783 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3784;
  assign dataGroup_lo_lo_3784 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3785;
  assign dataGroup_lo_lo_3785 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3786;
  assign dataGroup_lo_lo_3786 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3787;
  assign dataGroup_lo_lo_3787 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3788;
  assign dataGroup_lo_lo_3788 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3789;
  assign dataGroup_lo_lo_3789 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3790;
  assign dataGroup_lo_lo_3790 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3791;
  assign dataGroup_lo_lo_3791 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3792;
  assign dataGroup_lo_lo_3792 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3793;
  assign dataGroup_lo_lo_3793 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3794;
  assign dataGroup_lo_lo_3794 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3795;
  assign dataGroup_lo_lo_3795 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3796;
  assign dataGroup_lo_lo_3796 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3797;
  assign dataGroup_lo_lo_3797 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3798;
  assign dataGroup_lo_lo_3798 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3799;
  assign dataGroup_lo_lo_3799 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3800;
  assign dataGroup_lo_lo_3800 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3801;
  assign dataGroup_lo_lo_3801 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3802;
  assign dataGroup_lo_lo_3802 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3803;
  assign dataGroup_lo_lo_3803 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3804;
  assign dataGroup_lo_lo_3804 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3805;
  assign dataGroup_lo_lo_3805 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3806;
  assign dataGroup_lo_lo_3806 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3807;
  assign dataGroup_lo_lo_3807 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3808;
  assign dataGroup_lo_lo_3808 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3809;
  assign dataGroup_lo_lo_3809 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3810;
  assign dataGroup_lo_lo_3810 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3811;
  assign dataGroup_lo_lo_3811 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3812;
  assign dataGroup_lo_lo_3812 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3813;
  assign dataGroup_lo_lo_3813 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3814;
  assign dataGroup_lo_lo_3814 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3815;
  assign dataGroup_lo_lo_3815 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3816;
  assign dataGroup_lo_lo_3816 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3817;
  assign dataGroup_lo_lo_3817 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3818;
  assign dataGroup_lo_lo_3818 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3819;
  assign dataGroup_lo_lo_3819 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3820;
  assign dataGroup_lo_lo_3820 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3821;
  assign dataGroup_lo_lo_3821 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3822;
  assign dataGroup_lo_lo_3822 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3823;
  assign dataGroup_lo_lo_3823 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3824;
  assign dataGroup_lo_lo_3824 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3825;
  assign dataGroup_lo_lo_3825 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3826;
  assign dataGroup_lo_lo_3826 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3827;
  assign dataGroup_lo_lo_3827 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3828;
  assign dataGroup_lo_lo_3828 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3829;
  assign dataGroup_lo_lo_3829 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3830;
  assign dataGroup_lo_lo_3830 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3831;
  assign dataGroup_lo_lo_3831 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3832;
  assign dataGroup_lo_lo_3832 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3833;
  assign dataGroup_lo_lo_3833 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3834;
  assign dataGroup_lo_lo_3834 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3835;
  assign dataGroup_lo_lo_3835 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3836;
  assign dataGroup_lo_lo_3836 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3837;
  assign dataGroup_lo_lo_3837 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3838;
  assign dataGroup_lo_lo_3838 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3839;
  assign dataGroup_lo_lo_3839 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3840;
  assign dataGroup_lo_lo_3840 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3841;
  assign dataGroup_lo_lo_3841 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3842;
  assign dataGroup_lo_lo_3842 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3843;
  assign dataGroup_lo_lo_3843 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3844;
  assign dataGroup_lo_lo_3844 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3845;
  assign dataGroup_lo_lo_3845 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3846;
  assign dataGroup_lo_lo_3846 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3847;
  assign dataGroup_lo_lo_3847 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3848;
  assign dataGroup_lo_lo_3848 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3849;
  assign dataGroup_lo_lo_3849 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3850;
  assign dataGroup_lo_lo_3850 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3851;
  assign dataGroup_lo_lo_3851 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3852;
  assign dataGroup_lo_lo_3852 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3853;
  assign dataGroup_lo_lo_3853 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3854;
  assign dataGroup_lo_lo_3854 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3855;
  assign dataGroup_lo_lo_3855 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3856;
  assign dataGroup_lo_lo_3856 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3857;
  assign dataGroup_lo_lo_3857 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3858;
  assign dataGroup_lo_lo_3858 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3859;
  assign dataGroup_lo_lo_3859 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3860;
  assign dataGroup_lo_lo_3860 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3861;
  assign dataGroup_lo_lo_3861 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3862;
  assign dataGroup_lo_lo_3862 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3863;
  assign dataGroup_lo_lo_3863 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3864;
  assign dataGroup_lo_lo_3864 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3865;
  assign dataGroup_lo_lo_3865 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3866;
  assign dataGroup_lo_lo_3866 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3867;
  assign dataGroup_lo_lo_3867 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3868;
  assign dataGroup_lo_lo_3868 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3869;
  assign dataGroup_lo_lo_3869 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3870;
  assign dataGroup_lo_lo_3870 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3871;
  assign dataGroup_lo_lo_3871 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3872;
  assign dataGroup_lo_lo_3872 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3873;
  assign dataGroup_lo_lo_3873 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3874;
  assign dataGroup_lo_lo_3874 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3875;
  assign dataGroup_lo_lo_3875 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3876;
  assign dataGroup_lo_lo_3876 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3877;
  assign dataGroup_lo_lo_3877 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3878;
  assign dataGroup_lo_lo_3878 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3879;
  assign dataGroup_lo_lo_3879 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3880;
  assign dataGroup_lo_lo_3880 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3881;
  assign dataGroup_lo_lo_3881 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3882;
  assign dataGroup_lo_lo_3882 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3883;
  assign dataGroup_lo_lo_3883 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3884;
  assign dataGroup_lo_lo_3884 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3885;
  assign dataGroup_lo_lo_3885 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3886;
  assign dataGroup_lo_lo_3886 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3887;
  assign dataGroup_lo_lo_3887 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3888;
  assign dataGroup_lo_lo_3888 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3889;
  assign dataGroup_lo_lo_3889 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3890;
  assign dataGroup_lo_lo_3890 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3891;
  assign dataGroup_lo_lo_3891 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3892;
  assign dataGroup_lo_lo_3892 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3893;
  assign dataGroup_lo_lo_3893 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3894;
  assign dataGroup_lo_lo_3894 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3895;
  assign dataGroup_lo_lo_3895 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3896;
  assign dataGroup_lo_lo_3896 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3897;
  assign dataGroup_lo_lo_3897 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3898;
  assign dataGroup_lo_lo_3898 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3899;
  assign dataGroup_lo_lo_3899 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3900;
  assign dataGroup_lo_lo_3900 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3901;
  assign dataGroup_lo_lo_3901 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3902;
  assign dataGroup_lo_lo_3902 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3903;
  assign dataGroup_lo_lo_3903 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3904;
  assign dataGroup_lo_lo_3904 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3905;
  assign dataGroup_lo_lo_3905 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3906;
  assign dataGroup_lo_lo_3906 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3907;
  assign dataGroup_lo_lo_3907 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3908;
  assign dataGroup_lo_lo_3908 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3909;
  assign dataGroup_lo_lo_3909 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3910;
  assign dataGroup_lo_lo_3910 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3911;
  assign dataGroup_lo_lo_3911 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3912;
  assign dataGroup_lo_lo_3912 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3913;
  assign dataGroup_lo_lo_3913 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3914;
  assign dataGroup_lo_lo_3914 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3915;
  assign dataGroup_lo_lo_3915 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3916;
  assign dataGroup_lo_lo_3916 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3917;
  assign dataGroup_lo_lo_3917 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3918;
  assign dataGroup_lo_lo_3918 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3919;
  assign dataGroup_lo_lo_3919 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3920;
  assign dataGroup_lo_lo_3920 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3921;
  assign dataGroup_lo_lo_3921 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3922;
  assign dataGroup_lo_lo_3922 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3923;
  assign dataGroup_lo_lo_3923 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3924;
  assign dataGroup_lo_lo_3924 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3925;
  assign dataGroup_lo_lo_3925 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3926;
  assign dataGroup_lo_lo_3926 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3927;
  assign dataGroup_lo_lo_3927 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3928;
  assign dataGroup_lo_lo_3928 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3929;
  assign dataGroup_lo_lo_3929 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3930;
  assign dataGroup_lo_lo_3930 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3931;
  assign dataGroup_lo_lo_3931 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3932;
  assign dataGroup_lo_lo_3932 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3933;
  assign dataGroup_lo_lo_3933 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3934;
  assign dataGroup_lo_lo_3934 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3935;
  assign dataGroup_lo_lo_3935 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3936;
  assign dataGroup_lo_lo_3936 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3937;
  assign dataGroup_lo_lo_3937 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3938;
  assign dataGroup_lo_lo_3938 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3939;
  assign dataGroup_lo_lo_3939 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3940;
  assign dataGroup_lo_lo_3940 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3941;
  assign dataGroup_lo_lo_3941 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3942;
  assign dataGroup_lo_lo_3942 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3943;
  assign dataGroup_lo_lo_3943 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3944;
  assign dataGroup_lo_lo_3944 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3945;
  assign dataGroup_lo_lo_3945 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3946;
  assign dataGroup_lo_lo_3946 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3947;
  assign dataGroup_lo_lo_3947 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3948;
  assign dataGroup_lo_lo_3948 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3949;
  assign dataGroup_lo_lo_3949 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3950;
  assign dataGroup_lo_lo_3950 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3951;
  assign dataGroup_lo_lo_3951 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3952;
  assign dataGroup_lo_lo_3952 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3953;
  assign dataGroup_lo_lo_3953 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3954;
  assign dataGroup_lo_lo_3954 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3955;
  assign dataGroup_lo_lo_3955 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3956;
  assign dataGroup_lo_lo_3956 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3957;
  assign dataGroup_lo_lo_3957 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3958;
  assign dataGroup_lo_lo_3958 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3959;
  assign dataGroup_lo_lo_3959 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3960;
  assign dataGroup_lo_lo_3960 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3961;
  assign dataGroup_lo_lo_3961 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3962;
  assign dataGroup_lo_lo_3962 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3963;
  assign dataGroup_lo_lo_3963 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3964;
  assign dataGroup_lo_lo_3964 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3965;
  assign dataGroup_lo_lo_3965 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3966;
  assign dataGroup_lo_lo_3966 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3967;
  assign dataGroup_lo_lo_3967 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3968;
  assign dataGroup_lo_lo_3968 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3969;
  assign dataGroup_lo_lo_3969 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3970;
  assign dataGroup_lo_lo_3970 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3971;
  assign dataGroup_lo_lo_3971 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3972;
  assign dataGroup_lo_lo_3972 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3973;
  assign dataGroup_lo_lo_3973 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3974;
  assign dataGroup_lo_lo_3974 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3975;
  assign dataGroup_lo_lo_3975 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3976;
  assign dataGroup_lo_lo_3976 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3977;
  assign dataGroup_lo_lo_3977 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3978;
  assign dataGroup_lo_lo_3978 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3979;
  assign dataGroup_lo_lo_3979 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3980;
  assign dataGroup_lo_lo_3980 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3981;
  assign dataGroup_lo_lo_3981 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3982;
  assign dataGroup_lo_lo_3982 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3983;
  assign dataGroup_lo_lo_3983 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3984;
  assign dataGroup_lo_lo_3984 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3985;
  assign dataGroup_lo_lo_3985 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3986;
  assign dataGroup_lo_lo_3986 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3987;
  assign dataGroup_lo_lo_3987 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3988;
  assign dataGroup_lo_lo_3988 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3989;
  assign dataGroup_lo_lo_3989 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3990;
  assign dataGroup_lo_lo_3990 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3991;
  assign dataGroup_lo_lo_3991 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3992;
  assign dataGroup_lo_lo_3992 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3993;
  assign dataGroup_lo_lo_3993 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3994;
  assign dataGroup_lo_lo_3994 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3995;
  assign dataGroup_lo_lo_3995 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3996;
  assign dataGroup_lo_lo_3996 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3997;
  assign dataGroup_lo_lo_3997 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3998;
  assign dataGroup_lo_lo_3998 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_3999;
  assign dataGroup_lo_lo_3999 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4000;
  assign dataGroup_lo_lo_4000 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4001;
  assign dataGroup_lo_lo_4001 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4002;
  assign dataGroup_lo_lo_4002 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4003;
  assign dataGroup_lo_lo_4003 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4004;
  assign dataGroup_lo_lo_4004 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4005;
  assign dataGroup_lo_lo_4005 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4006;
  assign dataGroup_lo_lo_4006 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4007;
  assign dataGroup_lo_lo_4007 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4008;
  assign dataGroup_lo_lo_4008 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4009;
  assign dataGroup_lo_lo_4009 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4010;
  assign dataGroup_lo_lo_4010 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4011;
  assign dataGroup_lo_lo_4011 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4012;
  assign dataGroup_lo_lo_4012 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4013;
  assign dataGroup_lo_lo_4013 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4014;
  assign dataGroup_lo_lo_4014 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4015;
  assign dataGroup_lo_lo_4015 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4016;
  assign dataGroup_lo_lo_4016 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4017;
  assign dataGroup_lo_lo_4017 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4018;
  assign dataGroup_lo_lo_4018 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4019;
  assign dataGroup_lo_lo_4019 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4020;
  assign dataGroup_lo_lo_4020 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4021;
  assign dataGroup_lo_lo_4021 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4022;
  assign dataGroup_lo_lo_4022 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4023;
  assign dataGroup_lo_lo_4023 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4024;
  assign dataGroup_lo_lo_4024 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4025;
  assign dataGroup_lo_lo_4025 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4026;
  assign dataGroup_lo_lo_4026 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4027;
  assign dataGroup_lo_lo_4027 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4028;
  assign dataGroup_lo_lo_4028 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4029;
  assign dataGroup_lo_lo_4029 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4030;
  assign dataGroup_lo_lo_4030 = _GEN_5;
  wire [1023:0] dataGroup_lo_lo_4031;
  assign dataGroup_lo_lo_4031 = _GEN_5;
  wire [1023:0] _GEN_6 = {dataSelect_3, dataSelect_2};
  wire [1023:0] dataGroup_lo_hi;
  assign dataGroup_lo_hi = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1;
  assign dataGroup_lo_hi_1 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2;
  assign dataGroup_lo_hi_2 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3;
  assign dataGroup_lo_hi_3 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4;
  assign dataGroup_lo_hi_4 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_5;
  assign dataGroup_lo_hi_5 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_6;
  assign dataGroup_lo_hi_6 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_7;
  assign dataGroup_lo_hi_7 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_8;
  assign dataGroup_lo_hi_8 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_9;
  assign dataGroup_lo_hi_9 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_10;
  assign dataGroup_lo_hi_10 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_11;
  assign dataGroup_lo_hi_11 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_12;
  assign dataGroup_lo_hi_12 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_13;
  assign dataGroup_lo_hi_13 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_14;
  assign dataGroup_lo_hi_14 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_15;
  assign dataGroup_lo_hi_15 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_16;
  assign dataGroup_lo_hi_16 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_17;
  assign dataGroup_lo_hi_17 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_18;
  assign dataGroup_lo_hi_18 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_19;
  assign dataGroup_lo_hi_19 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_20;
  assign dataGroup_lo_hi_20 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_21;
  assign dataGroup_lo_hi_21 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_22;
  assign dataGroup_lo_hi_22 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_23;
  assign dataGroup_lo_hi_23 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_24;
  assign dataGroup_lo_hi_24 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_25;
  assign dataGroup_lo_hi_25 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_26;
  assign dataGroup_lo_hi_26 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_27;
  assign dataGroup_lo_hi_27 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_28;
  assign dataGroup_lo_hi_28 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_29;
  assign dataGroup_lo_hi_29 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_30;
  assign dataGroup_lo_hi_30 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_31;
  assign dataGroup_lo_hi_31 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_32;
  assign dataGroup_lo_hi_32 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_33;
  assign dataGroup_lo_hi_33 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_34;
  assign dataGroup_lo_hi_34 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_35;
  assign dataGroup_lo_hi_35 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_36;
  assign dataGroup_lo_hi_36 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_37;
  assign dataGroup_lo_hi_37 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_38;
  assign dataGroup_lo_hi_38 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_39;
  assign dataGroup_lo_hi_39 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_40;
  assign dataGroup_lo_hi_40 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_41;
  assign dataGroup_lo_hi_41 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_42;
  assign dataGroup_lo_hi_42 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_43;
  assign dataGroup_lo_hi_43 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_44;
  assign dataGroup_lo_hi_44 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_45;
  assign dataGroup_lo_hi_45 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_46;
  assign dataGroup_lo_hi_46 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_47;
  assign dataGroup_lo_hi_47 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_48;
  assign dataGroup_lo_hi_48 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_49;
  assign dataGroup_lo_hi_49 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_50;
  assign dataGroup_lo_hi_50 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_51;
  assign dataGroup_lo_hi_51 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_52;
  assign dataGroup_lo_hi_52 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_53;
  assign dataGroup_lo_hi_53 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_54;
  assign dataGroup_lo_hi_54 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_55;
  assign dataGroup_lo_hi_55 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_56;
  assign dataGroup_lo_hi_56 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_57;
  assign dataGroup_lo_hi_57 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_58;
  assign dataGroup_lo_hi_58 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_59;
  assign dataGroup_lo_hi_59 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_60;
  assign dataGroup_lo_hi_60 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_61;
  assign dataGroup_lo_hi_61 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_62;
  assign dataGroup_lo_hi_62 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_63;
  assign dataGroup_lo_hi_63 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_64;
  assign dataGroup_lo_hi_64 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_65;
  assign dataGroup_lo_hi_65 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_66;
  assign dataGroup_lo_hi_66 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_67;
  assign dataGroup_lo_hi_67 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_68;
  assign dataGroup_lo_hi_68 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_69;
  assign dataGroup_lo_hi_69 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_70;
  assign dataGroup_lo_hi_70 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_71;
  assign dataGroup_lo_hi_71 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_72;
  assign dataGroup_lo_hi_72 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_73;
  assign dataGroup_lo_hi_73 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_74;
  assign dataGroup_lo_hi_74 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_75;
  assign dataGroup_lo_hi_75 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_76;
  assign dataGroup_lo_hi_76 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_77;
  assign dataGroup_lo_hi_77 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_78;
  assign dataGroup_lo_hi_78 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_79;
  assign dataGroup_lo_hi_79 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_80;
  assign dataGroup_lo_hi_80 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_81;
  assign dataGroup_lo_hi_81 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_82;
  assign dataGroup_lo_hi_82 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_83;
  assign dataGroup_lo_hi_83 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_84;
  assign dataGroup_lo_hi_84 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_85;
  assign dataGroup_lo_hi_85 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_86;
  assign dataGroup_lo_hi_86 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_87;
  assign dataGroup_lo_hi_87 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_88;
  assign dataGroup_lo_hi_88 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_89;
  assign dataGroup_lo_hi_89 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_90;
  assign dataGroup_lo_hi_90 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_91;
  assign dataGroup_lo_hi_91 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_92;
  assign dataGroup_lo_hi_92 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_93;
  assign dataGroup_lo_hi_93 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_94;
  assign dataGroup_lo_hi_94 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_95;
  assign dataGroup_lo_hi_95 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_96;
  assign dataGroup_lo_hi_96 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_97;
  assign dataGroup_lo_hi_97 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_98;
  assign dataGroup_lo_hi_98 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_99;
  assign dataGroup_lo_hi_99 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_100;
  assign dataGroup_lo_hi_100 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_101;
  assign dataGroup_lo_hi_101 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_102;
  assign dataGroup_lo_hi_102 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_103;
  assign dataGroup_lo_hi_103 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_104;
  assign dataGroup_lo_hi_104 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_105;
  assign dataGroup_lo_hi_105 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_106;
  assign dataGroup_lo_hi_106 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_107;
  assign dataGroup_lo_hi_107 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_108;
  assign dataGroup_lo_hi_108 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_109;
  assign dataGroup_lo_hi_109 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_110;
  assign dataGroup_lo_hi_110 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_111;
  assign dataGroup_lo_hi_111 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_112;
  assign dataGroup_lo_hi_112 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_113;
  assign dataGroup_lo_hi_113 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_114;
  assign dataGroup_lo_hi_114 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_115;
  assign dataGroup_lo_hi_115 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_116;
  assign dataGroup_lo_hi_116 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_117;
  assign dataGroup_lo_hi_117 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_118;
  assign dataGroup_lo_hi_118 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_119;
  assign dataGroup_lo_hi_119 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_120;
  assign dataGroup_lo_hi_120 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_121;
  assign dataGroup_lo_hi_121 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_122;
  assign dataGroup_lo_hi_122 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_123;
  assign dataGroup_lo_hi_123 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_124;
  assign dataGroup_lo_hi_124 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_125;
  assign dataGroup_lo_hi_125 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_126;
  assign dataGroup_lo_hi_126 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_127;
  assign dataGroup_lo_hi_127 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_128;
  assign dataGroup_lo_hi_128 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_129;
  assign dataGroup_lo_hi_129 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_130;
  assign dataGroup_lo_hi_130 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_131;
  assign dataGroup_lo_hi_131 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_132;
  assign dataGroup_lo_hi_132 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_133;
  assign dataGroup_lo_hi_133 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_134;
  assign dataGroup_lo_hi_134 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_135;
  assign dataGroup_lo_hi_135 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_136;
  assign dataGroup_lo_hi_136 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_137;
  assign dataGroup_lo_hi_137 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_138;
  assign dataGroup_lo_hi_138 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_139;
  assign dataGroup_lo_hi_139 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_140;
  assign dataGroup_lo_hi_140 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_141;
  assign dataGroup_lo_hi_141 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_142;
  assign dataGroup_lo_hi_142 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_143;
  assign dataGroup_lo_hi_143 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_144;
  assign dataGroup_lo_hi_144 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_145;
  assign dataGroup_lo_hi_145 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_146;
  assign dataGroup_lo_hi_146 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_147;
  assign dataGroup_lo_hi_147 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_148;
  assign dataGroup_lo_hi_148 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_149;
  assign dataGroup_lo_hi_149 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_150;
  assign dataGroup_lo_hi_150 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_151;
  assign dataGroup_lo_hi_151 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_152;
  assign dataGroup_lo_hi_152 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_153;
  assign dataGroup_lo_hi_153 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_154;
  assign dataGroup_lo_hi_154 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_155;
  assign dataGroup_lo_hi_155 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_156;
  assign dataGroup_lo_hi_156 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_157;
  assign dataGroup_lo_hi_157 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_158;
  assign dataGroup_lo_hi_158 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_159;
  assign dataGroup_lo_hi_159 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_160;
  assign dataGroup_lo_hi_160 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_161;
  assign dataGroup_lo_hi_161 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_162;
  assign dataGroup_lo_hi_162 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_163;
  assign dataGroup_lo_hi_163 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_164;
  assign dataGroup_lo_hi_164 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_165;
  assign dataGroup_lo_hi_165 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_166;
  assign dataGroup_lo_hi_166 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_167;
  assign dataGroup_lo_hi_167 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_168;
  assign dataGroup_lo_hi_168 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_169;
  assign dataGroup_lo_hi_169 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_170;
  assign dataGroup_lo_hi_170 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_171;
  assign dataGroup_lo_hi_171 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_172;
  assign dataGroup_lo_hi_172 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_173;
  assign dataGroup_lo_hi_173 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_174;
  assign dataGroup_lo_hi_174 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_175;
  assign dataGroup_lo_hi_175 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_176;
  assign dataGroup_lo_hi_176 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_177;
  assign dataGroup_lo_hi_177 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_178;
  assign dataGroup_lo_hi_178 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_179;
  assign dataGroup_lo_hi_179 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_180;
  assign dataGroup_lo_hi_180 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_181;
  assign dataGroup_lo_hi_181 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_182;
  assign dataGroup_lo_hi_182 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_183;
  assign dataGroup_lo_hi_183 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_184;
  assign dataGroup_lo_hi_184 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_185;
  assign dataGroup_lo_hi_185 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_186;
  assign dataGroup_lo_hi_186 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_187;
  assign dataGroup_lo_hi_187 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_188;
  assign dataGroup_lo_hi_188 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_189;
  assign dataGroup_lo_hi_189 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_190;
  assign dataGroup_lo_hi_190 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_191;
  assign dataGroup_lo_hi_191 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_192;
  assign dataGroup_lo_hi_192 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_193;
  assign dataGroup_lo_hi_193 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_194;
  assign dataGroup_lo_hi_194 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_195;
  assign dataGroup_lo_hi_195 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_196;
  assign dataGroup_lo_hi_196 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_197;
  assign dataGroup_lo_hi_197 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_198;
  assign dataGroup_lo_hi_198 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_199;
  assign dataGroup_lo_hi_199 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_200;
  assign dataGroup_lo_hi_200 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_201;
  assign dataGroup_lo_hi_201 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_202;
  assign dataGroup_lo_hi_202 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_203;
  assign dataGroup_lo_hi_203 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_204;
  assign dataGroup_lo_hi_204 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_205;
  assign dataGroup_lo_hi_205 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_206;
  assign dataGroup_lo_hi_206 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_207;
  assign dataGroup_lo_hi_207 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_208;
  assign dataGroup_lo_hi_208 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_209;
  assign dataGroup_lo_hi_209 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_210;
  assign dataGroup_lo_hi_210 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_211;
  assign dataGroup_lo_hi_211 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_212;
  assign dataGroup_lo_hi_212 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_213;
  assign dataGroup_lo_hi_213 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_214;
  assign dataGroup_lo_hi_214 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_215;
  assign dataGroup_lo_hi_215 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_216;
  assign dataGroup_lo_hi_216 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_217;
  assign dataGroup_lo_hi_217 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_218;
  assign dataGroup_lo_hi_218 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_219;
  assign dataGroup_lo_hi_219 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_220;
  assign dataGroup_lo_hi_220 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_221;
  assign dataGroup_lo_hi_221 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_222;
  assign dataGroup_lo_hi_222 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_223;
  assign dataGroup_lo_hi_223 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_224;
  assign dataGroup_lo_hi_224 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_225;
  assign dataGroup_lo_hi_225 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_226;
  assign dataGroup_lo_hi_226 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_227;
  assign dataGroup_lo_hi_227 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_228;
  assign dataGroup_lo_hi_228 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_229;
  assign dataGroup_lo_hi_229 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_230;
  assign dataGroup_lo_hi_230 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_231;
  assign dataGroup_lo_hi_231 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_232;
  assign dataGroup_lo_hi_232 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_233;
  assign dataGroup_lo_hi_233 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_234;
  assign dataGroup_lo_hi_234 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_235;
  assign dataGroup_lo_hi_235 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_236;
  assign dataGroup_lo_hi_236 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_237;
  assign dataGroup_lo_hi_237 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_238;
  assign dataGroup_lo_hi_238 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_239;
  assign dataGroup_lo_hi_239 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_240;
  assign dataGroup_lo_hi_240 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_241;
  assign dataGroup_lo_hi_241 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_242;
  assign dataGroup_lo_hi_242 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_243;
  assign dataGroup_lo_hi_243 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_244;
  assign dataGroup_lo_hi_244 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_245;
  assign dataGroup_lo_hi_245 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_246;
  assign dataGroup_lo_hi_246 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_247;
  assign dataGroup_lo_hi_247 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_248;
  assign dataGroup_lo_hi_248 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_249;
  assign dataGroup_lo_hi_249 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_250;
  assign dataGroup_lo_hi_250 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_251;
  assign dataGroup_lo_hi_251 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_252;
  assign dataGroup_lo_hi_252 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_253;
  assign dataGroup_lo_hi_253 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_254;
  assign dataGroup_lo_hi_254 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_255;
  assign dataGroup_lo_hi_255 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_256;
  assign dataGroup_lo_hi_256 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_257;
  assign dataGroup_lo_hi_257 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_258;
  assign dataGroup_lo_hi_258 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_259;
  assign dataGroup_lo_hi_259 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_260;
  assign dataGroup_lo_hi_260 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_261;
  assign dataGroup_lo_hi_261 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_262;
  assign dataGroup_lo_hi_262 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_263;
  assign dataGroup_lo_hi_263 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_264;
  assign dataGroup_lo_hi_264 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_265;
  assign dataGroup_lo_hi_265 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_266;
  assign dataGroup_lo_hi_266 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_267;
  assign dataGroup_lo_hi_267 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_268;
  assign dataGroup_lo_hi_268 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_269;
  assign dataGroup_lo_hi_269 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_270;
  assign dataGroup_lo_hi_270 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_271;
  assign dataGroup_lo_hi_271 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_272;
  assign dataGroup_lo_hi_272 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_273;
  assign dataGroup_lo_hi_273 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_274;
  assign dataGroup_lo_hi_274 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_275;
  assign dataGroup_lo_hi_275 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_276;
  assign dataGroup_lo_hi_276 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_277;
  assign dataGroup_lo_hi_277 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_278;
  assign dataGroup_lo_hi_278 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_279;
  assign dataGroup_lo_hi_279 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_280;
  assign dataGroup_lo_hi_280 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_281;
  assign dataGroup_lo_hi_281 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_282;
  assign dataGroup_lo_hi_282 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_283;
  assign dataGroup_lo_hi_283 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_284;
  assign dataGroup_lo_hi_284 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_285;
  assign dataGroup_lo_hi_285 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_286;
  assign dataGroup_lo_hi_286 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_287;
  assign dataGroup_lo_hi_287 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_288;
  assign dataGroup_lo_hi_288 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_289;
  assign dataGroup_lo_hi_289 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_290;
  assign dataGroup_lo_hi_290 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_291;
  assign dataGroup_lo_hi_291 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_292;
  assign dataGroup_lo_hi_292 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_293;
  assign dataGroup_lo_hi_293 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_294;
  assign dataGroup_lo_hi_294 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_295;
  assign dataGroup_lo_hi_295 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_296;
  assign dataGroup_lo_hi_296 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_297;
  assign dataGroup_lo_hi_297 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_298;
  assign dataGroup_lo_hi_298 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_299;
  assign dataGroup_lo_hi_299 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_300;
  assign dataGroup_lo_hi_300 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_301;
  assign dataGroup_lo_hi_301 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_302;
  assign dataGroup_lo_hi_302 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_303;
  assign dataGroup_lo_hi_303 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_304;
  assign dataGroup_lo_hi_304 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_305;
  assign dataGroup_lo_hi_305 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_306;
  assign dataGroup_lo_hi_306 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_307;
  assign dataGroup_lo_hi_307 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_308;
  assign dataGroup_lo_hi_308 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_309;
  assign dataGroup_lo_hi_309 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_310;
  assign dataGroup_lo_hi_310 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_311;
  assign dataGroup_lo_hi_311 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_312;
  assign dataGroup_lo_hi_312 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_313;
  assign dataGroup_lo_hi_313 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_314;
  assign dataGroup_lo_hi_314 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_315;
  assign dataGroup_lo_hi_315 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_316;
  assign dataGroup_lo_hi_316 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_317;
  assign dataGroup_lo_hi_317 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_318;
  assign dataGroup_lo_hi_318 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_319;
  assign dataGroup_lo_hi_319 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_320;
  assign dataGroup_lo_hi_320 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_321;
  assign dataGroup_lo_hi_321 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_322;
  assign dataGroup_lo_hi_322 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_323;
  assign dataGroup_lo_hi_323 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_324;
  assign dataGroup_lo_hi_324 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_325;
  assign dataGroup_lo_hi_325 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_326;
  assign dataGroup_lo_hi_326 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_327;
  assign dataGroup_lo_hi_327 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_328;
  assign dataGroup_lo_hi_328 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_329;
  assign dataGroup_lo_hi_329 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_330;
  assign dataGroup_lo_hi_330 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_331;
  assign dataGroup_lo_hi_331 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_332;
  assign dataGroup_lo_hi_332 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_333;
  assign dataGroup_lo_hi_333 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_334;
  assign dataGroup_lo_hi_334 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_335;
  assign dataGroup_lo_hi_335 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_336;
  assign dataGroup_lo_hi_336 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_337;
  assign dataGroup_lo_hi_337 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_338;
  assign dataGroup_lo_hi_338 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_339;
  assign dataGroup_lo_hi_339 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_340;
  assign dataGroup_lo_hi_340 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_341;
  assign dataGroup_lo_hi_341 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_342;
  assign dataGroup_lo_hi_342 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_343;
  assign dataGroup_lo_hi_343 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_344;
  assign dataGroup_lo_hi_344 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_345;
  assign dataGroup_lo_hi_345 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_346;
  assign dataGroup_lo_hi_346 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_347;
  assign dataGroup_lo_hi_347 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_348;
  assign dataGroup_lo_hi_348 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_349;
  assign dataGroup_lo_hi_349 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_350;
  assign dataGroup_lo_hi_350 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_351;
  assign dataGroup_lo_hi_351 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_352;
  assign dataGroup_lo_hi_352 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_353;
  assign dataGroup_lo_hi_353 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_354;
  assign dataGroup_lo_hi_354 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_355;
  assign dataGroup_lo_hi_355 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_356;
  assign dataGroup_lo_hi_356 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_357;
  assign dataGroup_lo_hi_357 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_358;
  assign dataGroup_lo_hi_358 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_359;
  assign dataGroup_lo_hi_359 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_360;
  assign dataGroup_lo_hi_360 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_361;
  assign dataGroup_lo_hi_361 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_362;
  assign dataGroup_lo_hi_362 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_363;
  assign dataGroup_lo_hi_363 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_364;
  assign dataGroup_lo_hi_364 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_365;
  assign dataGroup_lo_hi_365 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_366;
  assign dataGroup_lo_hi_366 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_367;
  assign dataGroup_lo_hi_367 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_368;
  assign dataGroup_lo_hi_368 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_369;
  assign dataGroup_lo_hi_369 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_370;
  assign dataGroup_lo_hi_370 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_371;
  assign dataGroup_lo_hi_371 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_372;
  assign dataGroup_lo_hi_372 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_373;
  assign dataGroup_lo_hi_373 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_374;
  assign dataGroup_lo_hi_374 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_375;
  assign dataGroup_lo_hi_375 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_376;
  assign dataGroup_lo_hi_376 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_377;
  assign dataGroup_lo_hi_377 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_378;
  assign dataGroup_lo_hi_378 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_379;
  assign dataGroup_lo_hi_379 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_380;
  assign dataGroup_lo_hi_380 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_381;
  assign dataGroup_lo_hi_381 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_382;
  assign dataGroup_lo_hi_382 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_383;
  assign dataGroup_lo_hi_383 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_384;
  assign dataGroup_lo_hi_384 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_385;
  assign dataGroup_lo_hi_385 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_386;
  assign dataGroup_lo_hi_386 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_387;
  assign dataGroup_lo_hi_387 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_388;
  assign dataGroup_lo_hi_388 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_389;
  assign dataGroup_lo_hi_389 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_390;
  assign dataGroup_lo_hi_390 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_391;
  assign dataGroup_lo_hi_391 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_392;
  assign dataGroup_lo_hi_392 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_393;
  assign dataGroup_lo_hi_393 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_394;
  assign dataGroup_lo_hi_394 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_395;
  assign dataGroup_lo_hi_395 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_396;
  assign dataGroup_lo_hi_396 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_397;
  assign dataGroup_lo_hi_397 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_398;
  assign dataGroup_lo_hi_398 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_399;
  assign dataGroup_lo_hi_399 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_400;
  assign dataGroup_lo_hi_400 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_401;
  assign dataGroup_lo_hi_401 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_402;
  assign dataGroup_lo_hi_402 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_403;
  assign dataGroup_lo_hi_403 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_404;
  assign dataGroup_lo_hi_404 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_405;
  assign dataGroup_lo_hi_405 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_406;
  assign dataGroup_lo_hi_406 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_407;
  assign dataGroup_lo_hi_407 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_408;
  assign dataGroup_lo_hi_408 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_409;
  assign dataGroup_lo_hi_409 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_410;
  assign dataGroup_lo_hi_410 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_411;
  assign dataGroup_lo_hi_411 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_412;
  assign dataGroup_lo_hi_412 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_413;
  assign dataGroup_lo_hi_413 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_414;
  assign dataGroup_lo_hi_414 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_415;
  assign dataGroup_lo_hi_415 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_416;
  assign dataGroup_lo_hi_416 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_417;
  assign dataGroup_lo_hi_417 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_418;
  assign dataGroup_lo_hi_418 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_419;
  assign dataGroup_lo_hi_419 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_420;
  assign dataGroup_lo_hi_420 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_421;
  assign dataGroup_lo_hi_421 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_422;
  assign dataGroup_lo_hi_422 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_423;
  assign dataGroup_lo_hi_423 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_424;
  assign dataGroup_lo_hi_424 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_425;
  assign dataGroup_lo_hi_425 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_426;
  assign dataGroup_lo_hi_426 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_427;
  assign dataGroup_lo_hi_427 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_428;
  assign dataGroup_lo_hi_428 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_429;
  assign dataGroup_lo_hi_429 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_430;
  assign dataGroup_lo_hi_430 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_431;
  assign dataGroup_lo_hi_431 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_432;
  assign dataGroup_lo_hi_432 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_433;
  assign dataGroup_lo_hi_433 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_434;
  assign dataGroup_lo_hi_434 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_435;
  assign dataGroup_lo_hi_435 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_436;
  assign dataGroup_lo_hi_436 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_437;
  assign dataGroup_lo_hi_437 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_438;
  assign dataGroup_lo_hi_438 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_439;
  assign dataGroup_lo_hi_439 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_440;
  assign dataGroup_lo_hi_440 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_441;
  assign dataGroup_lo_hi_441 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_442;
  assign dataGroup_lo_hi_442 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_443;
  assign dataGroup_lo_hi_443 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_444;
  assign dataGroup_lo_hi_444 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_445;
  assign dataGroup_lo_hi_445 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_446;
  assign dataGroup_lo_hi_446 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_447;
  assign dataGroup_lo_hi_447 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_448;
  assign dataGroup_lo_hi_448 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_449;
  assign dataGroup_lo_hi_449 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_450;
  assign dataGroup_lo_hi_450 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_451;
  assign dataGroup_lo_hi_451 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_452;
  assign dataGroup_lo_hi_452 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_453;
  assign dataGroup_lo_hi_453 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_454;
  assign dataGroup_lo_hi_454 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_455;
  assign dataGroup_lo_hi_455 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_456;
  assign dataGroup_lo_hi_456 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_457;
  assign dataGroup_lo_hi_457 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_458;
  assign dataGroup_lo_hi_458 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_459;
  assign dataGroup_lo_hi_459 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_460;
  assign dataGroup_lo_hi_460 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_461;
  assign dataGroup_lo_hi_461 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_462;
  assign dataGroup_lo_hi_462 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_463;
  assign dataGroup_lo_hi_463 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_464;
  assign dataGroup_lo_hi_464 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_465;
  assign dataGroup_lo_hi_465 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_466;
  assign dataGroup_lo_hi_466 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_467;
  assign dataGroup_lo_hi_467 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_468;
  assign dataGroup_lo_hi_468 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_469;
  assign dataGroup_lo_hi_469 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_470;
  assign dataGroup_lo_hi_470 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_471;
  assign dataGroup_lo_hi_471 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_472;
  assign dataGroup_lo_hi_472 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_473;
  assign dataGroup_lo_hi_473 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_474;
  assign dataGroup_lo_hi_474 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_475;
  assign dataGroup_lo_hi_475 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_476;
  assign dataGroup_lo_hi_476 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_477;
  assign dataGroup_lo_hi_477 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_478;
  assign dataGroup_lo_hi_478 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_479;
  assign dataGroup_lo_hi_479 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_480;
  assign dataGroup_lo_hi_480 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_481;
  assign dataGroup_lo_hi_481 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_482;
  assign dataGroup_lo_hi_482 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_483;
  assign dataGroup_lo_hi_483 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_484;
  assign dataGroup_lo_hi_484 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_485;
  assign dataGroup_lo_hi_485 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_486;
  assign dataGroup_lo_hi_486 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_487;
  assign dataGroup_lo_hi_487 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_488;
  assign dataGroup_lo_hi_488 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_489;
  assign dataGroup_lo_hi_489 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_490;
  assign dataGroup_lo_hi_490 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_491;
  assign dataGroup_lo_hi_491 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_492;
  assign dataGroup_lo_hi_492 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_493;
  assign dataGroup_lo_hi_493 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_494;
  assign dataGroup_lo_hi_494 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_495;
  assign dataGroup_lo_hi_495 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_496;
  assign dataGroup_lo_hi_496 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_497;
  assign dataGroup_lo_hi_497 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_498;
  assign dataGroup_lo_hi_498 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_499;
  assign dataGroup_lo_hi_499 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_500;
  assign dataGroup_lo_hi_500 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_501;
  assign dataGroup_lo_hi_501 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_502;
  assign dataGroup_lo_hi_502 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_503;
  assign dataGroup_lo_hi_503 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_504;
  assign dataGroup_lo_hi_504 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_505;
  assign dataGroup_lo_hi_505 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_506;
  assign dataGroup_lo_hi_506 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_507;
  assign dataGroup_lo_hi_507 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_508;
  assign dataGroup_lo_hi_508 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_509;
  assign dataGroup_lo_hi_509 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_510;
  assign dataGroup_lo_hi_510 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_511;
  assign dataGroup_lo_hi_511 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_512;
  assign dataGroup_lo_hi_512 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_513;
  assign dataGroup_lo_hi_513 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_514;
  assign dataGroup_lo_hi_514 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_515;
  assign dataGroup_lo_hi_515 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_516;
  assign dataGroup_lo_hi_516 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_517;
  assign dataGroup_lo_hi_517 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_518;
  assign dataGroup_lo_hi_518 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_519;
  assign dataGroup_lo_hi_519 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_520;
  assign dataGroup_lo_hi_520 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_521;
  assign dataGroup_lo_hi_521 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_522;
  assign dataGroup_lo_hi_522 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_523;
  assign dataGroup_lo_hi_523 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_524;
  assign dataGroup_lo_hi_524 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_525;
  assign dataGroup_lo_hi_525 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_526;
  assign dataGroup_lo_hi_526 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_527;
  assign dataGroup_lo_hi_527 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_528;
  assign dataGroup_lo_hi_528 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_529;
  assign dataGroup_lo_hi_529 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_530;
  assign dataGroup_lo_hi_530 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_531;
  assign dataGroup_lo_hi_531 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_532;
  assign dataGroup_lo_hi_532 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_533;
  assign dataGroup_lo_hi_533 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_534;
  assign dataGroup_lo_hi_534 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_535;
  assign dataGroup_lo_hi_535 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_536;
  assign dataGroup_lo_hi_536 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_537;
  assign dataGroup_lo_hi_537 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_538;
  assign dataGroup_lo_hi_538 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_539;
  assign dataGroup_lo_hi_539 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_540;
  assign dataGroup_lo_hi_540 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_541;
  assign dataGroup_lo_hi_541 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_542;
  assign dataGroup_lo_hi_542 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_543;
  assign dataGroup_lo_hi_543 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_544;
  assign dataGroup_lo_hi_544 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_545;
  assign dataGroup_lo_hi_545 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_546;
  assign dataGroup_lo_hi_546 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_547;
  assign dataGroup_lo_hi_547 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_548;
  assign dataGroup_lo_hi_548 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_549;
  assign dataGroup_lo_hi_549 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_550;
  assign dataGroup_lo_hi_550 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_551;
  assign dataGroup_lo_hi_551 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_552;
  assign dataGroup_lo_hi_552 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_553;
  assign dataGroup_lo_hi_553 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_554;
  assign dataGroup_lo_hi_554 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_555;
  assign dataGroup_lo_hi_555 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_556;
  assign dataGroup_lo_hi_556 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_557;
  assign dataGroup_lo_hi_557 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_558;
  assign dataGroup_lo_hi_558 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_559;
  assign dataGroup_lo_hi_559 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_560;
  assign dataGroup_lo_hi_560 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_561;
  assign dataGroup_lo_hi_561 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_562;
  assign dataGroup_lo_hi_562 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_563;
  assign dataGroup_lo_hi_563 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_564;
  assign dataGroup_lo_hi_564 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_565;
  assign dataGroup_lo_hi_565 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_566;
  assign dataGroup_lo_hi_566 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_567;
  assign dataGroup_lo_hi_567 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_568;
  assign dataGroup_lo_hi_568 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_569;
  assign dataGroup_lo_hi_569 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_570;
  assign dataGroup_lo_hi_570 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_571;
  assign dataGroup_lo_hi_571 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_572;
  assign dataGroup_lo_hi_572 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_573;
  assign dataGroup_lo_hi_573 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_574;
  assign dataGroup_lo_hi_574 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_575;
  assign dataGroup_lo_hi_575 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_576;
  assign dataGroup_lo_hi_576 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_577;
  assign dataGroup_lo_hi_577 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_578;
  assign dataGroup_lo_hi_578 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_579;
  assign dataGroup_lo_hi_579 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_580;
  assign dataGroup_lo_hi_580 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_581;
  assign dataGroup_lo_hi_581 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_582;
  assign dataGroup_lo_hi_582 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_583;
  assign dataGroup_lo_hi_583 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_584;
  assign dataGroup_lo_hi_584 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_585;
  assign dataGroup_lo_hi_585 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_586;
  assign dataGroup_lo_hi_586 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_587;
  assign dataGroup_lo_hi_587 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_588;
  assign dataGroup_lo_hi_588 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_589;
  assign dataGroup_lo_hi_589 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_590;
  assign dataGroup_lo_hi_590 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_591;
  assign dataGroup_lo_hi_591 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_592;
  assign dataGroup_lo_hi_592 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_593;
  assign dataGroup_lo_hi_593 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_594;
  assign dataGroup_lo_hi_594 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_595;
  assign dataGroup_lo_hi_595 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_596;
  assign dataGroup_lo_hi_596 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_597;
  assign dataGroup_lo_hi_597 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_598;
  assign dataGroup_lo_hi_598 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_599;
  assign dataGroup_lo_hi_599 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_600;
  assign dataGroup_lo_hi_600 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_601;
  assign dataGroup_lo_hi_601 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_602;
  assign dataGroup_lo_hi_602 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_603;
  assign dataGroup_lo_hi_603 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_604;
  assign dataGroup_lo_hi_604 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_605;
  assign dataGroup_lo_hi_605 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_606;
  assign dataGroup_lo_hi_606 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_607;
  assign dataGroup_lo_hi_607 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_608;
  assign dataGroup_lo_hi_608 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_609;
  assign dataGroup_lo_hi_609 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_610;
  assign dataGroup_lo_hi_610 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_611;
  assign dataGroup_lo_hi_611 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_612;
  assign dataGroup_lo_hi_612 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_613;
  assign dataGroup_lo_hi_613 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_614;
  assign dataGroup_lo_hi_614 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_615;
  assign dataGroup_lo_hi_615 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_616;
  assign dataGroup_lo_hi_616 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_617;
  assign dataGroup_lo_hi_617 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_618;
  assign dataGroup_lo_hi_618 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_619;
  assign dataGroup_lo_hi_619 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_620;
  assign dataGroup_lo_hi_620 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_621;
  assign dataGroup_lo_hi_621 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_622;
  assign dataGroup_lo_hi_622 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_623;
  assign dataGroup_lo_hi_623 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_624;
  assign dataGroup_lo_hi_624 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_625;
  assign dataGroup_lo_hi_625 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_626;
  assign dataGroup_lo_hi_626 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_627;
  assign dataGroup_lo_hi_627 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_628;
  assign dataGroup_lo_hi_628 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_629;
  assign dataGroup_lo_hi_629 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_630;
  assign dataGroup_lo_hi_630 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_631;
  assign dataGroup_lo_hi_631 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_632;
  assign dataGroup_lo_hi_632 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_633;
  assign dataGroup_lo_hi_633 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_634;
  assign dataGroup_lo_hi_634 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_635;
  assign dataGroup_lo_hi_635 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_636;
  assign dataGroup_lo_hi_636 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_637;
  assign dataGroup_lo_hi_637 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_638;
  assign dataGroup_lo_hi_638 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_639;
  assign dataGroup_lo_hi_639 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_640;
  assign dataGroup_lo_hi_640 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_641;
  assign dataGroup_lo_hi_641 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_642;
  assign dataGroup_lo_hi_642 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_643;
  assign dataGroup_lo_hi_643 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_644;
  assign dataGroup_lo_hi_644 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_645;
  assign dataGroup_lo_hi_645 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_646;
  assign dataGroup_lo_hi_646 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_647;
  assign dataGroup_lo_hi_647 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_648;
  assign dataGroup_lo_hi_648 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_649;
  assign dataGroup_lo_hi_649 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_650;
  assign dataGroup_lo_hi_650 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_651;
  assign dataGroup_lo_hi_651 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_652;
  assign dataGroup_lo_hi_652 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_653;
  assign dataGroup_lo_hi_653 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_654;
  assign dataGroup_lo_hi_654 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_655;
  assign dataGroup_lo_hi_655 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_656;
  assign dataGroup_lo_hi_656 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_657;
  assign dataGroup_lo_hi_657 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_658;
  assign dataGroup_lo_hi_658 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_659;
  assign dataGroup_lo_hi_659 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_660;
  assign dataGroup_lo_hi_660 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_661;
  assign dataGroup_lo_hi_661 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_662;
  assign dataGroup_lo_hi_662 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_663;
  assign dataGroup_lo_hi_663 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_664;
  assign dataGroup_lo_hi_664 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_665;
  assign dataGroup_lo_hi_665 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_666;
  assign dataGroup_lo_hi_666 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_667;
  assign dataGroup_lo_hi_667 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_668;
  assign dataGroup_lo_hi_668 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_669;
  assign dataGroup_lo_hi_669 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_670;
  assign dataGroup_lo_hi_670 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_671;
  assign dataGroup_lo_hi_671 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_672;
  assign dataGroup_lo_hi_672 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_673;
  assign dataGroup_lo_hi_673 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_674;
  assign dataGroup_lo_hi_674 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_675;
  assign dataGroup_lo_hi_675 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_676;
  assign dataGroup_lo_hi_676 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_677;
  assign dataGroup_lo_hi_677 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_678;
  assign dataGroup_lo_hi_678 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_679;
  assign dataGroup_lo_hi_679 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_680;
  assign dataGroup_lo_hi_680 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_681;
  assign dataGroup_lo_hi_681 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_682;
  assign dataGroup_lo_hi_682 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_683;
  assign dataGroup_lo_hi_683 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_684;
  assign dataGroup_lo_hi_684 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_685;
  assign dataGroup_lo_hi_685 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_686;
  assign dataGroup_lo_hi_686 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_687;
  assign dataGroup_lo_hi_687 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_688;
  assign dataGroup_lo_hi_688 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_689;
  assign dataGroup_lo_hi_689 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_690;
  assign dataGroup_lo_hi_690 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_691;
  assign dataGroup_lo_hi_691 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_692;
  assign dataGroup_lo_hi_692 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_693;
  assign dataGroup_lo_hi_693 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_694;
  assign dataGroup_lo_hi_694 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_695;
  assign dataGroup_lo_hi_695 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_696;
  assign dataGroup_lo_hi_696 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_697;
  assign dataGroup_lo_hi_697 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_698;
  assign dataGroup_lo_hi_698 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_699;
  assign dataGroup_lo_hi_699 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_700;
  assign dataGroup_lo_hi_700 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_701;
  assign dataGroup_lo_hi_701 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_702;
  assign dataGroup_lo_hi_702 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_703;
  assign dataGroup_lo_hi_703 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_704;
  assign dataGroup_lo_hi_704 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_705;
  assign dataGroup_lo_hi_705 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_706;
  assign dataGroup_lo_hi_706 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_707;
  assign dataGroup_lo_hi_707 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_708;
  assign dataGroup_lo_hi_708 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_709;
  assign dataGroup_lo_hi_709 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_710;
  assign dataGroup_lo_hi_710 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_711;
  assign dataGroup_lo_hi_711 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_712;
  assign dataGroup_lo_hi_712 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_713;
  assign dataGroup_lo_hi_713 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_714;
  assign dataGroup_lo_hi_714 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_715;
  assign dataGroup_lo_hi_715 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_716;
  assign dataGroup_lo_hi_716 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_717;
  assign dataGroup_lo_hi_717 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_718;
  assign dataGroup_lo_hi_718 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_719;
  assign dataGroup_lo_hi_719 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_720;
  assign dataGroup_lo_hi_720 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_721;
  assign dataGroup_lo_hi_721 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_722;
  assign dataGroup_lo_hi_722 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_723;
  assign dataGroup_lo_hi_723 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_724;
  assign dataGroup_lo_hi_724 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_725;
  assign dataGroup_lo_hi_725 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_726;
  assign dataGroup_lo_hi_726 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_727;
  assign dataGroup_lo_hi_727 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_728;
  assign dataGroup_lo_hi_728 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_729;
  assign dataGroup_lo_hi_729 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_730;
  assign dataGroup_lo_hi_730 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_731;
  assign dataGroup_lo_hi_731 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_732;
  assign dataGroup_lo_hi_732 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_733;
  assign dataGroup_lo_hi_733 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_734;
  assign dataGroup_lo_hi_734 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_735;
  assign dataGroup_lo_hi_735 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_736;
  assign dataGroup_lo_hi_736 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_737;
  assign dataGroup_lo_hi_737 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_738;
  assign dataGroup_lo_hi_738 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_739;
  assign dataGroup_lo_hi_739 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_740;
  assign dataGroup_lo_hi_740 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_741;
  assign dataGroup_lo_hi_741 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_742;
  assign dataGroup_lo_hi_742 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_743;
  assign dataGroup_lo_hi_743 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_744;
  assign dataGroup_lo_hi_744 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_745;
  assign dataGroup_lo_hi_745 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_746;
  assign dataGroup_lo_hi_746 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_747;
  assign dataGroup_lo_hi_747 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_748;
  assign dataGroup_lo_hi_748 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_749;
  assign dataGroup_lo_hi_749 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_750;
  assign dataGroup_lo_hi_750 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_751;
  assign dataGroup_lo_hi_751 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_752;
  assign dataGroup_lo_hi_752 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_753;
  assign dataGroup_lo_hi_753 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_754;
  assign dataGroup_lo_hi_754 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_755;
  assign dataGroup_lo_hi_755 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_756;
  assign dataGroup_lo_hi_756 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_757;
  assign dataGroup_lo_hi_757 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_758;
  assign dataGroup_lo_hi_758 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_759;
  assign dataGroup_lo_hi_759 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_760;
  assign dataGroup_lo_hi_760 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_761;
  assign dataGroup_lo_hi_761 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_762;
  assign dataGroup_lo_hi_762 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_763;
  assign dataGroup_lo_hi_763 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_764;
  assign dataGroup_lo_hi_764 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_765;
  assign dataGroup_lo_hi_765 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_766;
  assign dataGroup_lo_hi_766 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_767;
  assign dataGroup_lo_hi_767 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_768;
  assign dataGroup_lo_hi_768 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_769;
  assign dataGroup_lo_hi_769 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_770;
  assign dataGroup_lo_hi_770 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_771;
  assign dataGroup_lo_hi_771 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_772;
  assign dataGroup_lo_hi_772 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_773;
  assign dataGroup_lo_hi_773 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_774;
  assign dataGroup_lo_hi_774 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_775;
  assign dataGroup_lo_hi_775 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_776;
  assign dataGroup_lo_hi_776 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_777;
  assign dataGroup_lo_hi_777 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_778;
  assign dataGroup_lo_hi_778 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_779;
  assign dataGroup_lo_hi_779 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_780;
  assign dataGroup_lo_hi_780 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_781;
  assign dataGroup_lo_hi_781 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_782;
  assign dataGroup_lo_hi_782 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_783;
  assign dataGroup_lo_hi_783 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_784;
  assign dataGroup_lo_hi_784 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_785;
  assign dataGroup_lo_hi_785 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_786;
  assign dataGroup_lo_hi_786 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_787;
  assign dataGroup_lo_hi_787 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_788;
  assign dataGroup_lo_hi_788 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_789;
  assign dataGroup_lo_hi_789 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_790;
  assign dataGroup_lo_hi_790 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_791;
  assign dataGroup_lo_hi_791 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_792;
  assign dataGroup_lo_hi_792 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_793;
  assign dataGroup_lo_hi_793 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_794;
  assign dataGroup_lo_hi_794 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_795;
  assign dataGroup_lo_hi_795 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_796;
  assign dataGroup_lo_hi_796 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_797;
  assign dataGroup_lo_hi_797 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_798;
  assign dataGroup_lo_hi_798 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_799;
  assign dataGroup_lo_hi_799 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_800;
  assign dataGroup_lo_hi_800 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_801;
  assign dataGroup_lo_hi_801 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_802;
  assign dataGroup_lo_hi_802 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_803;
  assign dataGroup_lo_hi_803 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_804;
  assign dataGroup_lo_hi_804 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_805;
  assign dataGroup_lo_hi_805 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_806;
  assign dataGroup_lo_hi_806 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_807;
  assign dataGroup_lo_hi_807 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_808;
  assign dataGroup_lo_hi_808 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_809;
  assign dataGroup_lo_hi_809 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_810;
  assign dataGroup_lo_hi_810 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_811;
  assign dataGroup_lo_hi_811 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_812;
  assign dataGroup_lo_hi_812 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_813;
  assign dataGroup_lo_hi_813 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_814;
  assign dataGroup_lo_hi_814 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_815;
  assign dataGroup_lo_hi_815 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_816;
  assign dataGroup_lo_hi_816 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_817;
  assign dataGroup_lo_hi_817 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_818;
  assign dataGroup_lo_hi_818 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_819;
  assign dataGroup_lo_hi_819 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_820;
  assign dataGroup_lo_hi_820 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_821;
  assign dataGroup_lo_hi_821 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_822;
  assign dataGroup_lo_hi_822 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_823;
  assign dataGroup_lo_hi_823 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_824;
  assign dataGroup_lo_hi_824 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_825;
  assign dataGroup_lo_hi_825 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_826;
  assign dataGroup_lo_hi_826 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_827;
  assign dataGroup_lo_hi_827 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_828;
  assign dataGroup_lo_hi_828 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_829;
  assign dataGroup_lo_hi_829 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_830;
  assign dataGroup_lo_hi_830 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_831;
  assign dataGroup_lo_hi_831 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_832;
  assign dataGroup_lo_hi_832 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_833;
  assign dataGroup_lo_hi_833 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_834;
  assign dataGroup_lo_hi_834 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_835;
  assign dataGroup_lo_hi_835 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_836;
  assign dataGroup_lo_hi_836 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_837;
  assign dataGroup_lo_hi_837 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_838;
  assign dataGroup_lo_hi_838 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_839;
  assign dataGroup_lo_hi_839 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_840;
  assign dataGroup_lo_hi_840 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_841;
  assign dataGroup_lo_hi_841 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_842;
  assign dataGroup_lo_hi_842 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_843;
  assign dataGroup_lo_hi_843 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_844;
  assign dataGroup_lo_hi_844 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_845;
  assign dataGroup_lo_hi_845 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_846;
  assign dataGroup_lo_hi_846 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_847;
  assign dataGroup_lo_hi_847 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_848;
  assign dataGroup_lo_hi_848 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_849;
  assign dataGroup_lo_hi_849 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_850;
  assign dataGroup_lo_hi_850 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_851;
  assign dataGroup_lo_hi_851 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_852;
  assign dataGroup_lo_hi_852 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_853;
  assign dataGroup_lo_hi_853 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_854;
  assign dataGroup_lo_hi_854 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_855;
  assign dataGroup_lo_hi_855 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_856;
  assign dataGroup_lo_hi_856 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_857;
  assign dataGroup_lo_hi_857 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_858;
  assign dataGroup_lo_hi_858 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_859;
  assign dataGroup_lo_hi_859 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_860;
  assign dataGroup_lo_hi_860 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_861;
  assign dataGroup_lo_hi_861 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_862;
  assign dataGroup_lo_hi_862 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_863;
  assign dataGroup_lo_hi_863 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_864;
  assign dataGroup_lo_hi_864 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_865;
  assign dataGroup_lo_hi_865 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_866;
  assign dataGroup_lo_hi_866 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_867;
  assign dataGroup_lo_hi_867 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_868;
  assign dataGroup_lo_hi_868 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_869;
  assign dataGroup_lo_hi_869 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_870;
  assign dataGroup_lo_hi_870 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_871;
  assign dataGroup_lo_hi_871 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_872;
  assign dataGroup_lo_hi_872 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_873;
  assign dataGroup_lo_hi_873 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_874;
  assign dataGroup_lo_hi_874 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_875;
  assign dataGroup_lo_hi_875 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_876;
  assign dataGroup_lo_hi_876 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_877;
  assign dataGroup_lo_hi_877 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_878;
  assign dataGroup_lo_hi_878 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_879;
  assign dataGroup_lo_hi_879 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_880;
  assign dataGroup_lo_hi_880 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_881;
  assign dataGroup_lo_hi_881 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_882;
  assign dataGroup_lo_hi_882 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_883;
  assign dataGroup_lo_hi_883 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_884;
  assign dataGroup_lo_hi_884 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_885;
  assign dataGroup_lo_hi_885 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_886;
  assign dataGroup_lo_hi_886 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_887;
  assign dataGroup_lo_hi_887 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_888;
  assign dataGroup_lo_hi_888 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_889;
  assign dataGroup_lo_hi_889 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_890;
  assign dataGroup_lo_hi_890 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_891;
  assign dataGroup_lo_hi_891 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_892;
  assign dataGroup_lo_hi_892 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_893;
  assign dataGroup_lo_hi_893 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_894;
  assign dataGroup_lo_hi_894 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_895;
  assign dataGroup_lo_hi_895 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_896;
  assign dataGroup_lo_hi_896 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_897;
  assign dataGroup_lo_hi_897 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_898;
  assign dataGroup_lo_hi_898 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_899;
  assign dataGroup_lo_hi_899 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_900;
  assign dataGroup_lo_hi_900 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_901;
  assign dataGroup_lo_hi_901 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_902;
  assign dataGroup_lo_hi_902 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_903;
  assign dataGroup_lo_hi_903 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_904;
  assign dataGroup_lo_hi_904 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_905;
  assign dataGroup_lo_hi_905 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_906;
  assign dataGroup_lo_hi_906 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_907;
  assign dataGroup_lo_hi_907 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_908;
  assign dataGroup_lo_hi_908 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_909;
  assign dataGroup_lo_hi_909 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_910;
  assign dataGroup_lo_hi_910 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_911;
  assign dataGroup_lo_hi_911 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_912;
  assign dataGroup_lo_hi_912 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_913;
  assign dataGroup_lo_hi_913 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_914;
  assign dataGroup_lo_hi_914 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_915;
  assign dataGroup_lo_hi_915 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_916;
  assign dataGroup_lo_hi_916 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_917;
  assign dataGroup_lo_hi_917 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_918;
  assign dataGroup_lo_hi_918 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_919;
  assign dataGroup_lo_hi_919 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_920;
  assign dataGroup_lo_hi_920 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_921;
  assign dataGroup_lo_hi_921 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_922;
  assign dataGroup_lo_hi_922 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_923;
  assign dataGroup_lo_hi_923 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_924;
  assign dataGroup_lo_hi_924 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_925;
  assign dataGroup_lo_hi_925 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_926;
  assign dataGroup_lo_hi_926 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_927;
  assign dataGroup_lo_hi_927 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_928;
  assign dataGroup_lo_hi_928 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_929;
  assign dataGroup_lo_hi_929 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_930;
  assign dataGroup_lo_hi_930 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_931;
  assign dataGroup_lo_hi_931 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_932;
  assign dataGroup_lo_hi_932 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_933;
  assign dataGroup_lo_hi_933 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_934;
  assign dataGroup_lo_hi_934 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_935;
  assign dataGroup_lo_hi_935 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_936;
  assign dataGroup_lo_hi_936 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_937;
  assign dataGroup_lo_hi_937 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_938;
  assign dataGroup_lo_hi_938 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_939;
  assign dataGroup_lo_hi_939 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_940;
  assign dataGroup_lo_hi_940 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_941;
  assign dataGroup_lo_hi_941 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_942;
  assign dataGroup_lo_hi_942 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_943;
  assign dataGroup_lo_hi_943 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_944;
  assign dataGroup_lo_hi_944 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_945;
  assign dataGroup_lo_hi_945 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_946;
  assign dataGroup_lo_hi_946 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_947;
  assign dataGroup_lo_hi_947 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_948;
  assign dataGroup_lo_hi_948 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_949;
  assign dataGroup_lo_hi_949 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_950;
  assign dataGroup_lo_hi_950 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_951;
  assign dataGroup_lo_hi_951 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_952;
  assign dataGroup_lo_hi_952 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_953;
  assign dataGroup_lo_hi_953 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_954;
  assign dataGroup_lo_hi_954 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_955;
  assign dataGroup_lo_hi_955 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_956;
  assign dataGroup_lo_hi_956 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_957;
  assign dataGroup_lo_hi_957 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_958;
  assign dataGroup_lo_hi_958 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_959;
  assign dataGroup_lo_hi_959 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_960;
  assign dataGroup_lo_hi_960 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_961;
  assign dataGroup_lo_hi_961 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_962;
  assign dataGroup_lo_hi_962 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_963;
  assign dataGroup_lo_hi_963 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_964;
  assign dataGroup_lo_hi_964 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_965;
  assign dataGroup_lo_hi_965 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_966;
  assign dataGroup_lo_hi_966 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_967;
  assign dataGroup_lo_hi_967 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_968;
  assign dataGroup_lo_hi_968 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_969;
  assign dataGroup_lo_hi_969 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_970;
  assign dataGroup_lo_hi_970 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_971;
  assign dataGroup_lo_hi_971 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_972;
  assign dataGroup_lo_hi_972 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_973;
  assign dataGroup_lo_hi_973 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_974;
  assign dataGroup_lo_hi_974 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_975;
  assign dataGroup_lo_hi_975 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_976;
  assign dataGroup_lo_hi_976 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_977;
  assign dataGroup_lo_hi_977 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_978;
  assign dataGroup_lo_hi_978 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_979;
  assign dataGroup_lo_hi_979 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_980;
  assign dataGroup_lo_hi_980 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_981;
  assign dataGroup_lo_hi_981 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_982;
  assign dataGroup_lo_hi_982 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_983;
  assign dataGroup_lo_hi_983 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_984;
  assign dataGroup_lo_hi_984 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_985;
  assign dataGroup_lo_hi_985 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_986;
  assign dataGroup_lo_hi_986 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_987;
  assign dataGroup_lo_hi_987 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_988;
  assign dataGroup_lo_hi_988 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_989;
  assign dataGroup_lo_hi_989 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_990;
  assign dataGroup_lo_hi_990 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_991;
  assign dataGroup_lo_hi_991 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_992;
  assign dataGroup_lo_hi_992 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_993;
  assign dataGroup_lo_hi_993 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_994;
  assign dataGroup_lo_hi_994 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_995;
  assign dataGroup_lo_hi_995 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_996;
  assign dataGroup_lo_hi_996 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_997;
  assign dataGroup_lo_hi_997 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_998;
  assign dataGroup_lo_hi_998 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_999;
  assign dataGroup_lo_hi_999 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1000;
  assign dataGroup_lo_hi_1000 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1001;
  assign dataGroup_lo_hi_1001 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1002;
  assign dataGroup_lo_hi_1002 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1003;
  assign dataGroup_lo_hi_1003 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1004;
  assign dataGroup_lo_hi_1004 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1005;
  assign dataGroup_lo_hi_1005 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1006;
  assign dataGroup_lo_hi_1006 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1007;
  assign dataGroup_lo_hi_1007 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1008;
  assign dataGroup_lo_hi_1008 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1009;
  assign dataGroup_lo_hi_1009 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1010;
  assign dataGroup_lo_hi_1010 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1011;
  assign dataGroup_lo_hi_1011 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1012;
  assign dataGroup_lo_hi_1012 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1013;
  assign dataGroup_lo_hi_1013 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1014;
  assign dataGroup_lo_hi_1014 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1015;
  assign dataGroup_lo_hi_1015 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1016;
  assign dataGroup_lo_hi_1016 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1017;
  assign dataGroup_lo_hi_1017 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1018;
  assign dataGroup_lo_hi_1018 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1019;
  assign dataGroup_lo_hi_1019 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1020;
  assign dataGroup_lo_hi_1020 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1021;
  assign dataGroup_lo_hi_1021 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1022;
  assign dataGroup_lo_hi_1022 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1023;
  assign dataGroup_lo_hi_1023 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1024;
  assign dataGroup_lo_hi_1024 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1025;
  assign dataGroup_lo_hi_1025 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1026;
  assign dataGroup_lo_hi_1026 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1027;
  assign dataGroup_lo_hi_1027 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1028;
  assign dataGroup_lo_hi_1028 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1029;
  assign dataGroup_lo_hi_1029 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1030;
  assign dataGroup_lo_hi_1030 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1031;
  assign dataGroup_lo_hi_1031 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1032;
  assign dataGroup_lo_hi_1032 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1033;
  assign dataGroup_lo_hi_1033 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1034;
  assign dataGroup_lo_hi_1034 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1035;
  assign dataGroup_lo_hi_1035 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1036;
  assign dataGroup_lo_hi_1036 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1037;
  assign dataGroup_lo_hi_1037 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1038;
  assign dataGroup_lo_hi_1038 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1039;
  assign dataGroup_lo_hi_1039 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1040;
  assign dataGroup_lo_hi_1040 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1041;
  assign dataGroup_lo_hi_1041 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1042;
  assign dataGroup_lo_hi_1042 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1043;
  assign dataGroup_lo_hi_1043 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1044;
  assign dataGroup_lo_hi_1044 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1045;
  assign dataGroup_lo_hi_1045 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1046;
  assign dataGroup_lo_hi_1046 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1047;
  assign dataGroup_lo_hi_1047 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1048;
  assign dataGroup_lo_hi_1048 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1049;
  assign dataGroup_lo_hi_1049 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1050;
  assign dataGroup_lo_hi_1050 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1051;
  assign dataGroup_lo_hi_1051 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1052;
  assign dataGroup_lo_hi_1052 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1053;
  assign dataGroup_lo_hi_1053 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1054;
  assign dataGroup_lo_hi_1054 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1055;
  assign dataGroup_lo_hi_1055 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1056;
  assign dataGroup_lo_hi_1056 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1057;
  assign dataGroup_lo_hi_1057 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1058;
  assign dataGroup_lo_hi_1058 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1059;
  assign dataGroup_lo_hi_1059 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1060;
  assign dataGroup_lo_hi_1060 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1061;
  assign dataGroup_lo_hi_1061 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1062;
  assign dataGroup_lo_hi_1062 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1063;
  assign dataGroup_lo_hi_1063 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1064;
  assign dataGroup_lo_hi_1064 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1065;
  assign dataGroup_lo_hi_1065 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1066;
  assign dataGroup_lo_hi_1066 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1067;
  assign dataGroup_lo_hi_1067 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1068;
  assign dataGroup_lo_hi_1068 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1069;
  assign dataGroup_lo_hi_1069 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1070;
  assign dataGroup_lo_hi_1070 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1071;
  assign dataGroup_lo_hi_1071 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1072;
  assign dataGroup_lo_hi_1072 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1073;
  assign dataGroup_lo_hi_1073 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1074;
  assign dataGroup_lo_hi_1074 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1075;
  assign dataGroup_lo_hi_1075 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1076;
  assign dataGroup_lo_hi_1076 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1077;
  assign dataGroup_lo_hi_1077 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1078;
  assign dataGroup_lo_hi_1078 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1079;
  assign dataGroup_lo_hi_1079 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1080;
  assign dataGroup_lo_hi_1080 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1081;
  assign dataGroup_lo_hi_1081 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1082;
  assign dataGroup_lo_hi_1082 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1083;
  assign dataGroup_lo_hi_1083 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1084;
  assign dataGroup_lo_hi_1084 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1085;
  assign dataGroup_lo_hi_1085 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1086;
  assign dataGroup_lo_hi_1086 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1087;
  assign dataGroup_lo_hi_1087 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1088;
  assign dataGroup_lo_hi_1088 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1089;
  assign dataGroup_lo_hi_1089 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1090;
  assign dataGroup_lo_hi_1090 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1091;
  assign dataGroup_lo_hi_1091 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1092;
  assign dataGroup_lo_hi_1092 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1093;
  assign dataGroup_lo_hi_1093 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1094;
  assign dataGroup_lo_hi_1094 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1095;
  assign dataGroup_lo_hi_1095 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1096;
  assign dataGroup_lo_hi_1096 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1097;
  assign dataGroup_lo_hi_1097 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1098;
  assign dataGroup_lo_hi_1098 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1099;
  assign dataGroup_lo_hi_1099 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1100;
  assign dataGroup_lo_hi_1100 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1101;
  assign dataGroup_lo_hi_1101 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1102;
  assign dataGroup_lo_hi_1102 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1103;
  assign dataGroup_lo_hi_1103 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1104;
  assign dataGroup_lo_hi_1104 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1105;
  assign dataGroup_lo_hi_1105 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1106;
  assign dataGroup_lo_hi_1106 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1107;
  assign dataGroup_lo_hi_1107 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1108;
  assign dataGroup_lo_hi_1108 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1109;
  assign dataGroup_lo_hi_1109 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1110;
  assign dataGroup_lo_hi_1110 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1111;
  assign dataGroup_lo_hi_1111 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1112;
  assign dataGroup_lo_hi_1112 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1113;
  assign dataGroup_lo_hi_1113 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1114;
  assign dataGroup_lo_hi_1114 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1115;
  assign dataGroup_lo_hi_1115 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1116;
  assign dataGroup_lo_hi_1116 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1117;
  assign dataGroup_lo_hi_1117 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1118;
  assign dataGroup_lo_hi_1118 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1119;
  assign dataGroup_lo_hi_1119 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1120;
  assign dataGroup_lo_hi_1120 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1121;
  assign dataGroup_lo_hi_1121 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1122;
  assign dataGroup_lo_hi_1122 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1123;
  assign dataGroup_lo_hi_1123 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1124;
  assign dataGroup_lo_hi_1124 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1125;
  assign dataGroup_lo_hi_1125 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1126;
  assign dataGroup_lo_hi_1126 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1127;
  assign dataGroup_lo_hi_1127 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1128;
  assign dataGroup_lo_hi_1128 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1129;
  assign dataGroup_lo_hi_1129 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1130;
  assign dataGroup_lo_hi_1130 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1131;
  assign dataGroup_lo_hi_1131 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1132;
  assign dataGroup_lo_hi_1132 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1133;
  assign dataGroup_lo_hi_1133 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1134;
  assign dataGroup_lo_hi_1134 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1135;
  assign dataGroup_lo_hi_1135 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1136;
  assign dataGroup_lo_hi_1136 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1137;
  assign dataGroup_lo_hi_1137 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1138;
  assign dataGroup_lo_hi_1138 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1139;
  assign dataGroup_lo_hi_1139 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1140;
  assign dataGroup_lo_hi_1140 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1141;
  assign dataGroup_lo_hi_1141 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1142;
  assign dataGroup_lo_hi_1142 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1143;
  assign dataGroup_lo_hi_1143 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1144;
  assign dataGroup_lo_hi_1144 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1145;
  assign dataGroup_lo_hi_1145 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1146;
  assign dataGroup_lo_hi_1146 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1147;
  assign dataGroup_lo_hi_1147 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1148;
  assign dataGroup_lo_hi_1148 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1149;
  assign dataGroup_lo_hi_1149 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1150;
  assign dataGroup_lo_hi_1150 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1151;
  assign dataGroup_lo_hi_1151 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1152;
  assign dataGroup_lo_hi_1152 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1153;
  assign dataGroup_lo_hi_1153 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1154;
  assign dataGroup_lo_hi_1154 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1155;
  assign dataGroup_lo_hi_1155 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1156;
  assign dataGroup_lo_hi_1156 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1157;
  assign dataGroup_lo_hi_1157 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1158;
  assign dataGroup_lo_hi_1158 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1159;
  assign dataGroup_lo_hi_1159 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1160;
  assign dataGroup_lo_hi_1160 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1161;
  assign dataGroup_lo_hi_1161 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1162;
  assign dataGroup_lo_hi_1162 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1163;
  assign dataGroup_lo_hi_1163 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1164;
  assign dataGroup_lo_hi_1164 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1165;
  assign dataGroup_lo_hi_1165 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1166;
  assign dataGroup_lo_hi_1166 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1167;
  assign dataGroup_lo_hi_1167 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1168;
  assign dataGroup_lo_hi_1168 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1169;
  assign dataGroup_lo_hi_1169 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1170;
  assign dataGroup_lo_hi_1170 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1171;
  assign dataGroup_lo_hi_1171 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1172;
  assign dataGroup_lo_hi_1172 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1173;
  assign dataGroup_lo_hi_1173 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1174;
  assign dataGroup_lo_hi_1174 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1175;
  assign dataGroup_lo_hi_1175 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1176;
  assign dataGroup_lo_hi_1176 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1177;
  assign dataGroup_lo_hi_1177 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1178;
  assign dataGroup_lo_hi_1178 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1179;
  assign dataGroup_lo_hi_1179 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1180;
  assign dataGroup_lo_hi_1180 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1181;
  assign dataGroup_lo_hi_1181 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1182;
  assign dataGroup_lo_hi_1182 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1183;
  assign dataGroup_lo_hi_1183 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1184;
  assign dataGroup_lo_hi_1184 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1185;
  assign dataGroup_lo_hi_1185 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1186;
  assign dataGroup_lo_hi_1186 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1187;
  assign dataGroup_lo_hi_1187 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1188;
  assign dataGroup_lo_hi_1188 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1189;
  assign dataGroup_lo_hi_1189 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1190;
  assign dataGroup_lo_hi_1190 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1191;
  assign dataGroup_lo_hi_1191 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1192;
  assign dataGroup_lo_hi_1192 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1193;
  assign dataGroup_lo_hi_1193 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1194;
  assign dataGroup_lo_hi_1194 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1195;
  assign dataGroup_lo_hi_1195 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1196;
  assign dataGroup_lo_hi_1196 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1197;
  assign dataGroup_lo_hi_1197 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1198;
  assign dataGroup_lo_hi_1198 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1199;
  assign dataGroup_lo_hi_1199 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1200;
  assign dataGroup_lo_hi_1200 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1201;
  assign dataGroup_lo_hi_1201 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1202;
  assign dataGroup_lo_hi_1202 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1203;
  assign dataGroup_lo_hi_1203 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1204;
  assign dataGroup_lo_hi_1204 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1205;
  assign dataGroup_lo_hi_1205 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1206;
  assign dataGroup_lo_hi_1206 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1207;
  assign dataGroup_lo_hi_1207 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1208;
  assign dataGroup_lo_hi_1208 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1209;
  assign dataGroup_lo_hi_1209 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1210;
  assign dataGroup_lo_hi_1210 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1211;
  assign dataGroup_lo_hi_1211 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1212;
  assign dataGroup_lo_hi_1212 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1213;
  assign dataGroup_lo_hi_1213 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1214;
  assign dataGroup_lo_hi_1214 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1215;
  assign dataGroup_lo_hi_1215 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1216;
  assign dataGroup_lo_hi_1216 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1217;
  assign dataGroup_lo_hi_1217 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1218;
  assign dataGroup_lo_hi_1218 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1219;
  assign dataGroup_lo_hi_1219 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1220;
  assign dataGroup_lo_hi_1220 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1221;
  assign dataGroup_lo_hi_1221 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1222;
  assign dataGroup_lo_hi_1222 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1223;
  assign dataGroup_lo_hi_1223 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1224;
  assign dataGroup_lo_hi_1224 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1225;
  assign dataGroup_lo_hi_1225 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1226;
  assign dataGroup_lo_hi_1226 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1227;
  assign dataGroup_lo_hi_1227 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1228;
  assign dataGroup_lo_hi_1228 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1229;
  assign dataGroup_lo_hi_1229 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1230;
  assign dataGroup_lo_hi_1230 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1231;
  assign dataGroup_lo_hi_1231 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1232;
  assign dataGroup_lo_hi_1232 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1233;
  assign dataGroup_lo_hi_1233 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1234;
  assign dataGroup_lo_hi_1234 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1235;
  assign dataGroup_lo_hi_1235 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1236;
  assign dataGroup_lo_hi_1236 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1237;
  assign dataGroup_lo_hi_1237 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1238;
  assign dataGroup_lo_hi_1238 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1239;
  assign dataGroup_lo_hi_1239 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1240;
  assign dataGroup_lo_hi_1240 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1241;
  assign dataGroup_lo_hi_1241 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1242;
  assign dataGroup_lo_hi_1242 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1243;
  assign dataGroup_lo_hi_1243 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1244;
  assign dataGroup_lo_hi_1244 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1245;
  assign dataGroup_lo_hi_1245 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1246;
  assign dataGroup_lo_hi_1246 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1247;
  assign dataGroup_lo_hi_1247 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1248;
  assign dataGroup_lo_hi_1248 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1249;
  assign dataGroup_lo_hi_1249 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1250;
  assign dataGroup_lo_hi_1250 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1251;
  assign dataGroup_lo_hi_1251 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1252;
  assign dataGroup_lo_hi_1252 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1253;
  assign dataGroup_lo_hi_1253 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1254;
  assign dataGroup_lo_hi_1254 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1255;
  assign dataGroup_lo_hi_1255 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1256;
  assign dataGroup_lo_hi_1256 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1257;
  assign dataGroup_lo_hi_1257 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1258;
  assign dataGroup_lo_hi_1258 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1259;
  assign dataGroup_lo_hi_1259 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1260;
  assign dataGroup_lo_hi_1260 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1261;
  assign dataGroup_lo_hi_1261 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1262;
  assign dataGroup_lo_hi_1262 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1263;
  assign dataGroup_lo_hi_1263 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1264;
  assign dataGroup_lo_hi_1264 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1265;
  assign dataGroup_lo_hi_1265 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1266;
  assign dataGroup_lo_hi_1266 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1267;
  assign dataGroup_lo_hi_1267 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1268;
  assign dataGroup_lo_hi_1268 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1269;
  assign dataGroup_lo_hi_1269 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1270;
  assign dataGroup_lo_hi_1270 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1271;
  assign dataGroup_lo_hi_1271 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1272;
  assign dataGroup_lo_hi_1272 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1273;
  assign dataGroup_lo_hi_1273 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1274;
  assign dataGroup_lo_hi_1274 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1275;
  assign dataGroup_lo_hi_1275 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1276;
  assign dataGroup_lo_hi_1276 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1277;
  assign dataGroup_lo_hi_1277 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1278;
  assign dataGroup_lo_hi_1278 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1279;
  assign dataGroup_lo_hi_1279 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1280;
  assign dataGroup_lo_hi_1280 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1281;
  assign dataGroup_lo_hi_1281 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1282;
  assign dataGroup_lo_hi_1282 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1283;
  assign dataGroup_lo_hi_1283 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1284;
  assign dataGroup_lo_hi_1284 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1285;
  assign dataGroup_lo_hi_1285 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1286;
  assign dataGroup_lo_hi_1286 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1287;
  assign dataGroup_lo_hi_1287 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1288;
  assign dataGroup_lo_hi_1288 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1289;
  assign dataGroup_lo_hi_1289 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1290;
  assign dataGroup_lo_hi_1290 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1291;
  assign dataGroup_lo_hi_1291 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1292;
  assign dataGroup_lo_hi_1292 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1293;
  assign dataGroup_lo_hi_1293 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1294;
  assign dataGroup_lo_hi_1294 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1295;
  assign dataGroup_lo_hi_1295 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1296;
  assign dataGroup_lo_hi_1296 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1297;
  assign dataGroup_lo_hi_1297 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1298;
  assign dataGroup_lo_hi_1298 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1299;
  assign dataGroup_lo_hi_1299 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1300;
  assign dataGroup_lo_hi_1300 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1301;
  assign dataGroup_lo_hi_1301 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1302;
  assign dataGroup_lo_hi_1302 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1303;
  assign dataGroup_lo_hi_1303 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1304;
  assign dataGroup_lo_hi_1304 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1305;
  assign dataGroup_lo_hi_1305 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1306;
  assign dataGroup_lo_hi_1306 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1307;
  assign dataGroup_lo_hi_1307 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1308;
  assign dataGroup_lo_hi_1308 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1309;
  assign dataGroup_lo_hi_1309 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1310;
  assign dataGroup_lo_hi_1310 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1311;
  assign dataGroup_lo_hi_1311 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1312;
  assign dataGroup_lo_hi_1312 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1313;
  assign dataGroup_lo_hi_1313 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1314;
  assign dataGroup_lo_hi_1314 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1315;
  assign dataGroup_lo_hi_1315 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1316;
  assign dataGroup_lo_hi_1316 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1317;
  assign dataGroup_lo_hi_1317 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1318;
  assign dataGroup_lo_hi_1318 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1319;
  assign dataGroup_lo_hi_1319 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1320;
  assign dataGroup_lo_hi_1320 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1321;
  assign dataGroup_lo_hi_1321 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1322;
  assign dataGroup_lo_hi_1322 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1323;
  assign dataGroup_lo_hi_1323 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1324;
  assign dataGroup_lo_hi_1324 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1325;
  assign dataGroup_lo_hi_1325 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1326;
  assign dataGroup_lo_hi_1326 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1327;
  assign dataGroup_lo_hi_1327 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1328;
  assign dataGroup_lo_hi_1328 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1329;
  assign dataGroup_lo_hi_1329 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1330;
  assign dataGroup_lo_hi_1330 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1331;
  assign dataGroup_lo_hi_1331 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1332;
  assign dataGroup_lo_hi_1332 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1333;
  assign dataGroup_lo_hi_1333 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1334;
  assign dataGroup_lo_hi_1334 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1335;
  assign dataGroup_lo_hi_1335 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1336;
  assign dataGroup_lo_hi_1336 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1337;
  assign dataGroup_lo_hi_1337 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1338;
  assign dataGroup_lo_hi_1338 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1339;
  assign dataGroup_lo_hi_1339 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1340;
  assign dataGroup_lo_hi_1340 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1341;
  assign dataGroup_lo_hi_1341 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1342;
  assign dataGroup_lo_hi_1342 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1343;
  assign dataGroup_lo_hi_1343 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1344;
  assign dataGroup_lo_hi_1344 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1345;
  assign dataGroup_lo_hi_1345 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1346;
  assign dataGroup_lo_hi_1346 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1347;
  assign dataGroup_lo_hi_1347 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1348;
  assign dataGroup_lo_hi_1348 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1349;
  assign dataGroup_lo_hi_1349 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1350;
  assign dataGroup_lo_hi_1350 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1351;
  assign dataGroup_lo_hi_1351 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1352;
  assign dataGroup_lo_hi_1352 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1353;
  assign dataGroup_lo_hi_1353 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1354;
  assign dataGroup_lo_hi_1354 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1355;
  assign dataGroup_lo_hi_1355 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1356;
  assign dataGroup_lo_hi_1356 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1357;
  assign dataGroup_lo_hi_1357 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1358;
  assign dataGroup_lo_hi_1358 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1359;
  assign dataGroup_lo_hi_1359 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1360;
  assign dataGroup_lo_hi_1360 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1361;
  assign dataGroup_lo_hi_1361 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1362;
  assign dataGroup_lo_hi_1362 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1363;
  assign dataGroup_lo_hi_1363 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1364;
  assign dataGroup_lo_hi_1364 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1365;
  assign dataGroup_lo_hi_1365 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1366;
  assign dataGroup_lo_hi_1366 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1367;
  assign dataGroup_lo_hi_1367 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1368;
  assign dataGroup_lo_hi_1368 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1369;
  assign dataGroup_lo_hi_1369 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1370;
  assign dataGroup_lo_hi_1370 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1371;
  assign dataGroup_lo_hi_1371 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1372;
  assign dataGroup_lo_hi_1372 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1373;
  assign dataGroup_lo_hi_1373 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1374;
  assign dataGroup_lo_hi_1374 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1375;
  assign dataGroup_lo_hi_1375 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1376;
  assign dataGroup_lo_hi_1376 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1377;
  assign dataGroup_lo_hi_1377 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1378;
  assign dataGroup_lo_hi_1378 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1379;
  assign dataGroup_lo_hi_1379 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1380;
  assign dataGroup_lo_hi_1380 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1381;
  assign dataGroup_lo_hi_1381 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1382;
  assign dataGroup_lo_hi_1382 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1383;
  assign dataGroup_lo_hi_1383 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1384;
  assign dataGroup_lo_hi_1384 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1385;
  assign dataGroup_lo_hi_1385 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1386;
  assign dataGroup_lo_hi_1386 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1387;
  assign dataGroup_lo_hi_1387 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1388;
  assign dataGroup_lo_hi_1388 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1389;
  assign dataGroup_lo_hi_1389 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1390;
  assign dataGroup_lo_hi_1390 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1391;
  assign dataGroup_lo_hi_1391 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1392;
  assign dataGroup_lo_hi_1392 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1393;
  assign dataGroup_lo_hi_1393 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1394;
  assign dataGroup_lo_hi_1394 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1395;
  assign dataGroup_lo_hi_1395 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1396;
  assign dataGroup_lo_hi_1396 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1397;
  assign dataGroup_lo_hi_1397 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1398;
  assign dataGroup_lo_hi_1398 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1399;
  assign dataGroup_lo_hi_1399 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1400;
  assign dataGroup_lo_hi_1400 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1401;
  assign dataGroup_lo_hi_1401 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1402;
  assign dataGroup_lo_hi_1402 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1403;
  assign dataGroup_lo_hi_1403 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1404;
  assign dataGroup_lo_hi_1404 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1405;
  assign dataGroup_lo_hi_1405 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1406;
  assign dataGroup_lo_hi_1406 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1407;
  assign dataGroup_lo_hi_1407 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1408;
  assign dataGroup_lo_hi_1408 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1409;
  assign dataGroup_lo_hi_1409 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1410;
  assign dataGroup_lo_hi_1410 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1411;
  assign dataGroup_lo_hi_1411 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1412;
  assign dataGroup_lo_hi_1412 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1413;
  assign dataGroup_lo_hi_1413 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1414;
  assign dataGroup_lo_hi_1414 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1415;
  assign dataGroup_lo_hi_1415 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1416;
  assign dataGroup_lo_hi_1416 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1417;
  assign dataGroup_lo_hi_1417 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1418;
  assign dataGroup_lo_hi_1418 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1419;
  assign dataGroup_lo_hi_1419 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1420;
  assign dataGroup_lo_hi_1420 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1421;
  assign dataGroup_lo_hi_1421 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1422;
  assign dataGroup_lo_hi_1422 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1423;
  assign dataGroup_lo_hi_1423 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1424;
  assign dataGroup_lo_hi_1424 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1425;
  assign dataGroup_lo_hi_1425 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1426;
  assign dataGroup_lo_hi_1426 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1427;
  assign dataGroup_lo_hi_1427 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1428;
  assign dataGroup_lo_hi_1428 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1429;
  assign dataGroup_lo_hi_1429 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1430;
  assign dataGroup_lo_hi_1430 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1431;
  assign dataGroup_lo_hi_1431 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1432;
  assign dataGroup_lo_hi_1432 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1433;
  assign dataGroup_lo_hi_1433 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1434;
  assign dataGroup_lo_hi_1434 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1435;
  assign dataGroup_lo_hi_1435 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1436;
  assign dataGroup_lo_hi_1436 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1437;
  assign dataGroup_lo_hi_1437 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1438;
  assign dataGroup_lo_hi_1438 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1439;
  assign dataGroup_lo_hi_1439 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1440;
  assign dataGroup_lo_hi_1440 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1441;
  assign dataGroup_lo_hi_1441 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1442;
  assign dataGroup_lo_hi_1442 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1443;
  assign dataGroup_lo_hi_1443 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1444;
  assign dataGroup_lo_hi_1444 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1445;
  assign dataGroup_lo_hi_1445 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1446;
  assign dataGroup_lo_hi_1446 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1447;
  assign dataGroup_lo_hi_1447 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1448;
  assign dataGroup_lo_hi_1448 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1449;
  assign dataGroup_lo_hi_1449 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1450;
  assign dataGroup_lo_hi_1450 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1451;
  assign dataGroup_lo_hi_1451 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1452;
  assign dataGroup_lo_hi_1452 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1453;
  assign dataGroup_lo_hi_1453 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1454;
  assign dataGroup_lo_hi_1454 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1455;
  assign dataGroup_lo_hi_1455 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1456;
  assign dataGroup_lo_hi_1456 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1457;
  assign dataGroup_lo_hi_1457 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1458;
  assign dataGroup_lo_hi_1458 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1459;
  assign dataGroup_lo_hi_1459 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1460;
  assign dataGroup_lo_hi_1460 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1461;
  assign dataGroup_lo_hi_1461 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1462;
  assign dataGroup_lo_hi_1462 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1463;
  assign dataGroup_lo_hi_1463 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1464;
  assign dataGroup_lo_hi_1464 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1465;
  assign dataGroup_lo_hi_1465 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1466;
  assign dataGroup_lo_hi_1466 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1467;
  assign dataGroup_lo_hi_1467 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1468;
  assign dataGroup_lo_hi_1468 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1469;
  assign dataGroup_lo_hi_1469 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1470;
  assign dataGroup_lo_hi_1470 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1471;
  assign dataGroup_lo_hi_1471 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1472;
  assign dataGroup_lo_hi_1472 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1473;
  assign dataGroup_lo_hi_1473 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1474;
  assign dataGroup_lo_hi_1474 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1475;
  assign dataGroup_lo_hi_1475 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1476;
  assign dataGroup_lo_hi_1476 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1477;
  assign dataGroup_lo_hi_1477 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1478;
  assign dataGroup_lo_hi_1478 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1479;
  assign dataGroup_lo_hi_1479 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1480;
  assign dataGroup_lo_hi_1480 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1481;
  assign dataGroup_lo_hi_1481 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1482;
  assign dataGroup_lo_hi_1482 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1483;
  assign dataGroup_lo_hi_1483 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1484;
  assign dataGroup_lo_hi_1484 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1485;
  assign dataGroup_lo_hi_1485 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1486;
  assign dataGroup_lo_hi_1486 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1487;
  assign dataGroup_lo_hi_1487 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1488;
  assign dataGroup_lo_hi_1488 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1489;
  assign dataGroup_lo_hi_1489 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1490;
  assign dataGroup_lo_hi_1490 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1491;
  assign dataGroup_lo_hi_1491 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1492;
  assign dataGroup_lo_hi_1492 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1493;
  assign dataGroup_lo_hi_1493 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1494;
  assign dataGroup_lo_hi_1494 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1495;
  assign dataGroup_lo_hi_1495 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1496;
  assign dataGroup_lo_hi_1496 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1497;
  assign dataGroup_lo_hi_1497 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1498;
  assign dataGroup_lo_hi_1498 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1499;
  assign dataGroup_lo_hi_1499 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1500;
  assign dataGroup_lo_hi_1500 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1501;
  assign dataGroup_lo_hi_1501 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1502;
  assign dataGroup_lo_hi_1502 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1503;
  assign dataGroup_lo_hi_1503 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1504;
  assign dataGroup_lo_hi_1504 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1505;
  assign dataGroup_lo_hi_1505 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1506;
  assign dataGroup_lo_hi_1506 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1507;
  assign dataGroup_lo_hi_1507 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1508;
  assign dataGroup_lo_hi_1508 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1509;
  assign dataGroup_lo_hi_1509 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1510;
  assign dataGroup_lo_hi_1510 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1511;
  assign dataGroup_lo_hi_1511 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1512;
  assign dataGroup_lo_hi_1512 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1513;
  assign dataGroup_lo_hi_1513 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1514;
  assign dataGroup_lo_hi_1514 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1515;
  assign dataGroup_lo_hi_1515 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1516;
  assign dataGroup_lo_hi_1516 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1517;
  assign dataGroup_lo_hi_1517 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1518;
  assign dataGroup_lo_hi_1518 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1519;
  assign dataGroup_lo_hi_1519 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1520;
  assign dataGroup_lo_hi_1520 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1521;
  assign dataGroup_lo_hi_1521 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1522;
  assign dataGroup_lo_hi_1522 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1523;
  assign dataGroup_lo_hi_1523 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1524;
  assign dataGroup_lo_hi_1524 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1525;
  assign dataGroup_lo_hi_1525 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1526;
  assign dataGroup_lo_hi_1526 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1527;
  assign dataGroup_lo_hi_1527 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1528;
  assign dataGroup_lo_hi_1528 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1529;
  assign dataGroup_lo_hi_1529 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1530;
  assign dataGroup_lo_hi_1530 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1531;
  assign dataGroup_lo_hi_1531 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1532;
  assign dataGroup_lo_hi_1532 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1533;
  assign dataGroup_lo_hi_1533 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1534;
  assign dataGroup_lo_hi_1534 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1535;
  assign dataGroup_lo_hi_1535 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1536;
  assign dataGroup_lo_hi_1536 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1537;
  assign dataGroup_lo_hi_1537 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1538;
  assign dataGroup_lo_hi_1538 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1539;
  assign dataGroup_lo_hi_1539 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1540;
  assign dataGroup_lo_hi_1540 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1541;
  assign dataGroup_lo_hi_1541 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1542;
  assign dataGroup_lo_hi_1542 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1543;
  assign dataGroup_lo_hi_1543 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1544;
  assign dataGroup_lo_hi_1544 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1545;
  assign dataGroup_lo_hi_1545 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1546;
  assign dataGroup_lo_hi_1546 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1547;
  assign dataGroup_lo_hi_1547 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1548;
  assign dataGroup_lo_hi_1548 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1549;
  assign dataGroup_lo_hi_1549 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1550;
  assign dataGroup_lo_hi_1550 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1551;
  assign dataGroup_lo_hi_1551 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1552;
  assign dataGroup_lo_hi_1552 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1553;
  assign dataGroup_lo_hi_1553 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1554;
  assign dataGroup_lo_hi_1554 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1555;
  assign dataGroup_lo_hi_1555 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1556;
  assign dataGroup_lo_hi_1556 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1557;
  assign dataGroup_lo_hi_1557 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1558;
  assign dataGroup_lo_hi_1558 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1559;
  assign dataGroup_lo_hi_1559 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1560;
  assign dataGroup_lo_hi_1560 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1561;
  assign dataGroup_lo_hi_1561 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1562;
  assign dataGroup_lo_hi_1562 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1563;
  assign dataGroup_lo_hi_1563 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1564;
  assign dataGroup_lo_hi_1564 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1565;
  assign dataGroup_lo_hi_1565 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1566;
  assign dataGroup_lo_hi_1566 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1567;
  assign dataGroup_lo_hi_1567 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1568;
  assign dataGroup_lo_hi_1568 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1569;
  assign dataGroup_lo_hi_1569 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1570;
  assign dataGroup_lo_hi_1570 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1571;
  assign dataGroup_lo_hi_1571 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1572;
  assign dataGroup_lo_hi_1572 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1573;
  assign dataGroup_lo_hi_1573 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1574;
  assign dataGroup_lo_hi_1574 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1575;
  assign dataGroup_lo_hi_1575 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1576;
  assign dataGroup_lo_hi_1576 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1577;
  assign dataGroup_lo_hi_1577 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1578;
  assign dataGroup_lo_hi_1578 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1579;
  assign dataGroup_lo_hi_1579 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1580;
  assign dataGroup_lo_hi_1580 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1581;
  assign dataGroup_lo_hi_1581 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1582;
  assign dataGroup_lo_hi_1582 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1583;
  assign dataGroup_lo_hi_1583 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1584;
  assign dataGroup_lo_hi_1584 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1585;
  assign dataGroup_lo_hi_1585 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1586;
  assign dataGroup_lo_hi_1586 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1587;
  assign dataGroup_lo_hi_1587 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1588;
  assign dataGroup_lo_hi_1588 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1589;
  assign dataGroup_lo_hi_1589 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1590;
  assign dataGroup_lo_hi_1590 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1591;
  assign dataGroup_lo_hi_1591 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1592;
  assign dataGroup_lo_hi_1592 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1593;
  assign dataGroup_lo_hi_1593 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1594;
  assign dataGroup_lo_hi_1594 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1595;
  assign dataGroup_lo_hi_1595 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1596;
  assign dataGroup_lo_hi_1596 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1597;
  assign dataGroup_lo_hi_1597 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1598;
  assign dataGroup_lo_hi_1598 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1599;
  assign dataGroup_lo_hi_1599 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1600;
  assign dataGroup_lo_hi_1600 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1601;
  assign dataGroup_lo_hi_1601 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1602;
  assign dataGroup_lo_hi_1602 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1603;
  assign dataGroup_lo_hi_1603 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1604;
  assign dataGroup_lo_hi_1604 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1605;
  assign dataGroup_lo_hi_1605 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1606;
  assign dataGroup_lo_hi_1606 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1607;
  assign dataGroup_lo_hi_1607 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1608;
  assign dataGroup_lo_hi_1608 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1609;
  assign dataGroup_lo_hi_1609 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1610;
  assign dataGroup_lo_hi_1610 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1611;
  assign dataGroup_lo_hi_1611 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1612;
  assign dataGroup_lo_hi_1612 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1613;
  assign dataGroup_lo_hi_1613 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1614;
  assign dataGroup_lo_hi_1614 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1615;
  assign dataGroup_lo_hi_1615 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1616;
  assign dataGroup_lo_hi_1616 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1617;
  assign dataGroup_lo_hi_1617 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1618;
  assign dataGroup_lo_hi_1618 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1619;
  assign dataGroup_lo_hi_1619 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1620;
  assign dataGroup_lo_hi_1620 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1621;
  assign dataGroup_lo_hi_1621 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1622;
  assign dataGroup_lo_hi_1622 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1623;
  assign dataGroup_lo_hi_1623 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1624;
  assign dataGroup_lo_hi_1624 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1625;
  assign dataGroup_lo_hi_1625 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1626;
  assign dataGroup_lo_hi_1626 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1627;
  assign dataGroup_lo_hi_1627 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1628;
  assign dataGroup_lo_hi_1628 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1629;
  assign dataGroup_lo_hi_1629 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1630;
  assign dataGroup_lo_hi_1630 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1631;
  assign dataGroup_lo_hi_1631 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1632;
  assign dataGroup_lo_hi_1632 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1633;
  assign dataGroup_lo_hi_1633 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1634;
  assign dataGroup_lo_hi_1634 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1635;
  assign dataGroup_lo_hi_1635 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1636;
  assign dataGroup_lo_hi_1636 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1637;
  assign dataGroup_lo_hi_1637 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1638;
  assign dataGroup_lo_hi_1638 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1639;
  assign dataGroup_lo_hi_1639 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1640;
  assign dataGroup_lo_hi_1640 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1641;
  assign dataGroup_lo_hi_1641 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1642;
  assign dataGroup_lo_hi_1642 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1643;
  assign dataGroup_lo_hi_1643 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1644;
  assign dataGroup_lo_hi_1644 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1645;
  assign dataGroup_lo_hi_1645 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1646;
  assign dataGroup_lo_hi_1646 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1647;
  assign dataGroup_lo_hi_1647 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1648;
  assign dataGroup_lo_hi_1648 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1649;
  assign dataGroup_lo_hi_1649 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1650;
  assign dataGroup_lo_hi_1650 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1651;
  assign dataGroup_lo_hi_1651 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1652;
  assign dataGroup_lo_hi_1652 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1653;
  assign dataGroup_lo_hi_1653 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1654;
  assign dataGroup_lo_hi_1654 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1655;
  assign dataGroup_lo_hi_1655 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1656;
  assign dataGroup_lo_hi_1656 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1657;
  assign dataGroup_lo_hi_1657 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1658;
  assign dataGroup_lo_hi_1658 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1659;
  assign dataGroup_lo_hi_1659 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1660;
  assign dataGroup_lo_hi_1660 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1661;
  assign dataGroup_lo_hi_1661 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1662;
  assign dataGroup_lo_hi_1662 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1663;
  assign dataGroup_lo_hi_1663 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1664;
  assign dataGroup_lo_hi_1664 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1665;
  assign dataGroup_lo_hi_1665 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1666;
  assign dataGroup_lo_hi_1666 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1667;
  assign dataGroup_lo_hi_1667 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1668;
  assign dataGroup_lo_hi_1668 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1669;
  assign dataGroup_lo_hi_1669 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1670;
  assign dataGroup_lo_hi_1670 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1671;
  assign dataGroup_lo_hi_1671 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1672;
  assign dataGroup_lo_hi_1672 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1673;
  assign dataGroup_lo_hi_1673 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1674;
  assign dataGroup_lo_hi_1674 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1675;
  assign dataGroup_lo_hi_1675 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1676;
  assign dataGroup_lo_hi_1676 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1677;
  assign dataGroup_lo_hi_1677 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1678;
  assign dataGroup_lo_hi_1678 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1679;
  assign dataGroup_lo_hi_1679 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1680;
  assign dataGroup_lo_hi_1680 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1681;
  assign dataGroup_lo_hi_1681 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1682;
  assign dataGroup_lo_hi_1682 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1683;
  assign dataGroup_lo_hi_1683 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1684;
  assign dataGroup_lo_hi_1684 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1685;
  assign dataGroup_lo_hi_1685 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1686;
  assign dataGroup_lo_hi_1686 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1687;
  assign dataGroup_lo_hi_1687 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1688;
  assign dataGroup_lo_hi_1688 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1689;
  assign dataGroup_lo_hi_1689 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1690;
  assign dataGroup_lo_hi_1690 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1691;
  assign dataGroup_lo_hi_1691 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1692;
  assign dataGroup_lo_hi_1692 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1693;
  assign dataGroup_lo_hi_1693 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1694;
  assign dataGroup_lo_hi_1694 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1695;
  assign dataGroup_lo_hi_1695 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1696;
  assign dataGroup_lo_hi_1696 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1697;
  assign dataGroup_lo_hi_1697 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1698;
  assign dataGroup_lo_hi_1698 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1699;
  assign dataGroup_lo_hi_1699 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1700;
  assign dataGroup_lo_hi_1700 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1701;
  assign dataGroup_lo_hi_1701 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1702;
  assign dataGroup_lo_hi_1702 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1703;
  assign dataGroup_lo_hi_1703 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1704;
  assign dataGroup_lo_hi_1704 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1705;
  assign dataGroup_lo_hi_1705 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1706;
  assign dataGroup_lo_hi_1706 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1707;
  assign dataGroup_lo_hi_1707 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1708;
  assign dataGroup_lo_hi_1708 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1709;
  assign dataGroup_lo_hi_1709 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1710;
  assign dataGroup_lo_hi_1710 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1711;
  assign dataGroup_lo_hi_1711 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1712;
  assign dataGroup_lo_hi_1712 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1713;
  assign dataGroup_lo_hi_1713 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1714;
  assign dataGroup_lo_hi_1714 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1715;
  assign dataGroup_lo_hi_1715 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1716;
  assign dataGroup_lo_hi_1716 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1717;
  assign dataGroup_lo_hi_1717 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1718;
  assign dataGroup_lo_hi_1718 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1719;
  assign dataGroup_lo_hi_1719 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1720;
  assign dataGroup_lo_hi_1720 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1721;
  assign dataGroup_lo_hi_1721 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1722;
  assign dataGroup_lo_hi_1722 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1723;
  assign dataGroup_lo_hi_1723 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1724;
  assign dataGroup_lo_hi_1724 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1725;
  assign dataGroup_lo_hi_1725 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1726;
  assign dataGroup_lo_hi_1726 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1727;
  assign dataGroup_lo_hi_1727 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1728;
  assign dataGroup_lo_hi_1728 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1729;
  assign dataGroup_lo_hi_1729 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1730;
  assign dataGroup_lo_hi_1730 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1731;
  assign dataGroup_lo_hi_1731 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1732;
  assign dataGroup_lo_hi_1732 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1733;
  assign dataGroup_lo_hi_1733 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1734;
  assign dataGroup_lo_hi_1734 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1735;
  assign dataGroup_lo_hi_1735 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1736;
  assign dataGroup_lo_hi_1736 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1737;
  assign dataGroup_lo_hi_1737 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1738;
  assign dataGroup_lo_hi_1738 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1739;
  assign dataGroup_lo_hi_1739 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1740;
  assign dataGroup_lo_hi_1740 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1741;
  assign dataGroup_lo_hi_1741 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1742;
  assign dataGroup_lo_hi_1742 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1743;
  assign dataGroup_lo_hi_1743 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1744;
  assign dataGroup_lo_hi_1744 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1745;
  assign dataGroup_lo_hi_1745 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1746;
  assign dataGroup_lo_hi_1746 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1747;
  assign dataGroup_lo_hi_1747 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1748;
  assign dataGroup_lo_hi_1748 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1749;
  assign dataGroup_lo_hi_1749 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1750;
  assign dataGroup_lo_hi_1750 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1751;
  assign dataGroup_lo_hi_1751 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1752;
  assign dataGroup_lo_hi_1752 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1753;
  assign dataGroup_lo_hi_1753 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1754;
  assign dataGroup_lo_hi_1754 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1755;
  assign dataGroup_lo_hi_1755 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1756;
  assign dataGroup_lo_hi_1756 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1757;
  assign dataGroup_lo_hi_1757 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1758;
  assign dataGroup_lo_hi_1758 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1759;
  assign dataGroup_lo_hi_1759 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1760;
  assign dataGroup_lo_hi_1760 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1761;
  assign dataGroup_lo_hi_1761 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1762;
  assign dataGroup_lo_hi_1762 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1763;
  assign dataGroup_lo_hi_1763 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1764;
  assign dataGroup_lo_hi_1764 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1765;
  assign dataGroup_lo_hi_1765 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1766;
  assign dataGroup_lo_hi_1766 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1767;
  assign dataGroup_lo_hi_1767 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1768;
  assign dataGroup_lo_hi_1768 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1769;
  assign dataGroup_lo_hi_1769 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1770;
  assign dataGroup_lo_hi_1770 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1771;
  assign dataGroup_lo_hi_1771 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1772;
  assign dataGroup_lo_hi_1772 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1773;
  assign dataGroup_lo_hi_1773 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1774;
  assign dataGroup_lo_hi_1774 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1775;
  assign dataGroup_lo_hi_1775 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1776;
  assign dataGroup_lo_hi_1776 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1777;
  assign dataGroup_lo_hi_1777 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1778;
  assign dataGroup_lo_hi_1778 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1779;
  assign dataGroup_lo_hi_1779 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1780;
  assign dataGroup_lo_hi_1780 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1781;
  assign dataGroup_lo_hi_1781 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1782;
  assign dataGroup_lo_hi_1782 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1783;
  assign dataGroup_lo_hi_1783 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1784;
  assign dataGroup_lo_hi_1784 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1785;
  assign dataGroup_lo_hi_1785 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1786;
  assign dataGroup_lo_hi_1786 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1787;
  assign dataGroup_lo_hi_1787 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1788;
  assign dataGroup_lo_hi_1788 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1789;
  assign dataGroup_lo_hi_1789 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1790;
  assign dataGroup_lo_hi_1790 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1791;
  assign dataGroup_lo_hi_1791 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1792;
  assign dataGroup_lo_hi_1792 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1793;
  assign dataGroup_lo_hi_1793 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1794;
  assign dataGroup_lo_hi_1794 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1795;
  assign dataGroup_lo_hi_1795 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1796;
  assign dataGroup_lo_hi_1796 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1797;
  assign dataGroup_lo_hi_1797 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1798;
  assign dataGroup_lo_hi_1798 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1799;
  assign dataGroup_lo_hi_1799 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1800;
  assign dataGroup_lo_hi_1800 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1801;
  assign dataGroup_lo_hi_1801 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1802;
  assign dataGroup_lo_hi_1802 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1803;
  assign dataGroup_lo_hi_1803 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1804;
  assign dataGroup_lo_hi_1804 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1805;
  assign dataGroup_lo_hi_1805 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1806;
  assign dataGroup_lo_hi_1806 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1807;
  assign dataGroup_lo_hi_1807 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1808;
  assign dataGroup_lo_hi_1808 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1809;
  assign dataGroup_lo_hi_1809 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1810;
  assign dataGroup_lo_hi_1810 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1811;
  assign dataGroup_lo_hi_1811 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1812;
  assign dataGroup_lo_hi_1812 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1813;
  assign dataGroup_lo_hi_1813 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1814;
  assign dataGroup_lo_hi_1814 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1815;
  assign dataGroup_lo_hi_1815 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1816;
  assign dataGroup_lo_hi_1816 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1817;
  assign dataGroup_lo_hi_1817 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1818;
  assign dataGroup_lo_hi_1818 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1819;
  assign dataGroup_lo_hi_1819 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1820;
  assign dataGroup_lo_hi_1820 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1821;
  assign dataGroup_lo_hi_1821 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1822;
  assign dataGroup_lo_hi_1822 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1823;
  assign dataGroup_lo_hi_1823 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1824;
  assign dataGroup_lo_hi_1824 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1825;
  assign dataGroup_lo_hi_1825 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1826;
  assign dataGroup_lo_hi_1826 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1827;
  assign dataGroup_lo_hi_1827 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1828;
  assign dataGroup_lo_hi_1828 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1829;
  assign dataGroup_lo_hi_1829 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1830;
  assign dataGroup_lo_hi_1830 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1831;
  assign dataGroup_lo_hi_1831 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1832;
  assign dataGroup_lo_hi_1832 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1833;
  assign dataGroup_lo_hi_1833 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1834;
  assign dataGroup_lo_hi_1834 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1835;
  assign dataGroup_lo_hi_1835 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1836;
  assign dataGroup_lo_hi_1836 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1837;
  assign dataGroup_lo_hi_1837 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1838;
  assign dataGroup_lo_hi_1838 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1839;
  assign dataGroup_lo_hi_1839 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1840;
  assign dataGroup_lo_hi_1840 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1841;
  assign dataGroup_lo_hi_1841 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1842;
  assign dataGroup_lo_hi_1842 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1843;
  assign dataGroup_lo_hi_1843 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1844;
  assign dataGroup_lo_hi_1844 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1845;
  assign dataGroup_lo_hi_1845 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1846;
  assign dataGroup_lo_hi_1846 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1847;
  assign dataGroup_lo_hi_1847 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1848;
  assign dataGroup_lo_hi_1848 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1849;
  assign dataGroup_lo_hi_1849 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1850;
  assign dataGroup_lo_hi_1850 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1851;
  assign dataGroup_lo_hi_1851 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1852;
  assign dataGroup_lo_hi_1852 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1853;
  assign dataGroup_lo_hi_1853 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1854;
  assign dataGroup_lo_hi_1854 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1855;
  assign dataGroup_lo_hi_1855 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1856;
  assign dataGroup_lo_hi_1856 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1857;
  assign dataGroup_lo_hi_1857 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1858;
  assign dataGroup_lo_hi_1858 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1859;
  assign dataGroup_lo_hi_1859 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1860;
  assign dataGroup_lo_hi_1860 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1861;
  assign dataGroup_lo_hi_1861 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1862;
  assign dataGroup_lo_hi_1862 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1863;
  assign dataGroup_lo_hi_1863 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1864;
  assign dataGroup_lo_hi_1864 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1865;
  assign dataGroup_lo_hi_1865 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1866;
  assign dataGroup_lo_hi_1866 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1867;
  assign dataGroup_lo_hi_1867 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1868;
  assign dataGroup_lo_hi_1868 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1869;
  assign dataGroup_lo_hi_1869 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1870;
  assign dataGroup_lo_hi_1870 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1871;
  assign dataGroup_lo_hi_1871 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1872;
  assign dataGroup_lo_hi_1872 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1873;
  assign dataGroup_lo_hi_1873 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1874;
  assign dataGroup_lo_hi_1874 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1875;
  assign dataGroup_lo_hi_1875 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1876;
  assign dataGroup_lo_hi_1876 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1877;
  assign dataGroup_lo_hi_1877 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1878;
  assign dataGroup_lo_hi_1878 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1879;
  assign dataGroup_lo_hi_1879 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1880;
  assign dataGroup_lo_hi_1880 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1881;
  assign dataGroup_lo_hi_1881 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1882;
  assign dataGroup_lo_hi_1882 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1883;
  assign dataGroup_lo_hi_1883 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1884;
  assign dataGroup_lo_hi_1884 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1885;
  assign dataGroup_lo_hi_1885 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1886;
  assign dataGroup_lo_hi_1886 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1887;
  assign dataGroup_lo_hi_1887 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1888;
  assign dataGroup_lo_hi_1888 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1889;
  assign dataGroup_lo_hi_1889 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1890;
  assign dataGroup_lo_hi_1890 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1891;
  assign dataGroup_lo_hi_1891 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1892;
  assign dataGroup_lo_hi_1892 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1893;
  assign dataGroup_lo_hi_1893 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1894;
  assign dataGroup_lo_hi_1894 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1895;
  assign dataGroup_lo_hi_1895 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1896;
  assign dataGroup_lo_hi_1896 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1897;
  assign dataGroup_lo_hi_1897 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1898;
  assign dataGroup_lo_hi_1898 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1899;
  assign dataGroup_lo_hi_1899 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1900;
  assign dataGroup_lo_hi_1900 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1901;
  assign dataGroup_lo_hi_1901 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1902;
  assign dataGroup_lo_hi_1902 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1903;
  assign dataGroup_lo_hi_1903 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1904;
  assign dataGroup_lo_hi_1904 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1905;
  assign dataGroup_lo_hi_1905 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1906;
  assign dataGroup_lo_hi_1906 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1907;
  assign dataGroup_lo_hi_1907 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1908;
  assign dataGroup_lo_hi_1908 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1909;
  assign dataGroup_lo_hi_1909 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1910;
  assign dataGroup_lo_hi_1910 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1911;
  assign dataGroup_lo_hi_1911 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1912;
  assign dataGroup_lo_hi_1912 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1913;
  assign dataGroup_lo_hi_1913 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1914;
  assign dataGroup_lo_hi_1914 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1915;
  assign dataGroup_lo_hi_1915 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1916;
  assign dataGroup_lo_hi_1916 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1917;
  assign dataGroup_lo_hi_1917 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1918;
  assign dataGroup_lo_hi_1918 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1919;
  assign dataGroup_lo_hi_1919 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1920;
  assign dataGroup_lo_hi_1920 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1921;
  assign dataGroup_lo_hi_1921 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1922;
  assign dataGroup_lo_hi_1922 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1923;
  assign dataGroup_lo_hi_1923 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1924;
  assign dataGroup_lo_hi_1924 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1925;
  assign dataGroup_lo_hi_1925 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1926;
  assign dataGroup_lo_hi_1926 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1927;
  assign dataGroup_lo_hi_1927 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1928;
  assign dataGroup_lo_hi_1928 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1929;
  assign dataGroup_lo_hi_1929 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1930;
  assign dataGroup_lo_hi_1930 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1931;
  assign dataGroup_lo_hi_1931 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1932;
  assign dataGroup_lo_hi_1932 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1933;
  assign dataGroup_lo_hi_1933 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1934;
  assign dataGroup_lo_hi_1934 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1935;
  assign dataGroup_lo_hi_1935 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1936;
  assign dataGroup_lo_hi_1936 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1937;
  assign dataGroup_lo_hi_1937 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1938;
  assign dataGroup_lo_hi_1938 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1939;
  assign dataGroup_lo_hi_1939 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1940;
  assign dataGroup_lo_hi_1940 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1941;
  assign dataGroup_lo_hi_1941 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1942;
  assign dataGroup_lo_hi_1942 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1943;
  assign dataGroup_lo_hi_1943 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1944;
  assign dataGroup_lo_hi_1944 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1945;
  assign dataGroup_lo_hi_1945 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1946;
  assign dataGroup_lo_hi_1946 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1947;
  assign dataGroup_lo_hi_1947 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1948;
  assign dataGroup_lo_hi_1948 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1949;
  assign dataGroup_lo_hi_1949 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1950;
  assign dataGroup_lo_hi_1950 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1951;
  assign dataGroup_lo_hi_1951 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1952;
  assign dataGroup_lo_hi_1952 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1953;
  assign dataGroup_lo_hi_1953 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1954;
  assign dataGroup_lo_hi_1954 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1955;
  assign dataGroup_lo_hi_1955 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1956;
  assign dataGroup_lo_hi_1956 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1957;
  assign dataGroup_lo_hi_1957 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1958;
  assign dataGroup_lo_hi_1958 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1959;
  assign dataGroup_lo_hi_1959 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1960;
  assign dataGroup_lo_hi_1960 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1961;
  assign dataGroup_lo_hi_1961 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1962;
  assign dataGroup_lo_hi_1962 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1963;
  assign dataGroup_lo_hi_1963 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1964;
  assign dataGroup_lo_hi_1964 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1965;
  assign dataGroup_lo_hi_1965 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1966;
  assign dataGroup_lo_hi_1966 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1967;
  assign dataGroup_lo_hi_1967 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1968;
  assign dataGroup_lo_hi_1968 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1969;
  assign dataGroup_lo_hi_1969 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1970;
  assign dataGroup_lo_hi_1970 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1971;
  assign dataGroup_lo_hi_1971 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1972;
  assign dataGroup_lo_hi_1972 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1973;
  assign dataGroup_lo_hi_1973 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1974;
  assign dataGroup_lo_hi_1974 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1975;
  assign dataGroup_lo_hi_1975 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1976;
  assign dataGroup_lo_hi_1976 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1977;
  assign dataGroup_lo_hi_1977 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1978;
  assign dataGroup_lo_hi_1978 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1979;
  assign dataGroup_lo_hi_1979 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1980;
  assign dataGroup_lo_hi_1980 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1981;
  assign dataGroup_lo_hi_1981 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1982;
  assign dataGroup_lo_hi_1982 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1983;
  assign dataGroup_lo_hi_1983 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1984;
  assign dataGroup_lo_hi_1984 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1985;
  assign dataGroup_lo_hi_1985 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1986;
  assign dataGroup_lo_hi_1986 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1987;
  assign dataGroup_lo_hi_1987 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1988;
  assign dataGroup_lo_hi_1988 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1989;
  assign dataGroup_lo_hi_1989 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1990;
  assign dataGroup_lo_hi_1990 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1991;
  assign dataGroup_lo_hi_1991 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1992;
  assign dataGroup_lo_hi_1992 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1993;
  assign dataGroup_lo_hi_1993 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1994;
  assign dataGroup_lo_hi_1994 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1995;
  assign dataGroup_lo_hi_1995 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1996;
  assign dataGroup_lo_hi_1996 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1997;
  assign dataGroup_lo_hi_1997 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1998;
  assign dataGroup_lo_hi_1998 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_1999;
  assign dataGroup_lo_hi_1999 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2000;
  assign dataGroup_lo_hi_2000 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2001;
  assign dataGroup_lo_hi_2001 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2002;
  assign dataGroup_lo_hi_2002 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2003;
  assign dataGroup_lo_hi_2003 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2004;
  assign dataGroup_lo_hi_2004 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2005;
  assign dataGroup_lo_hi_2005 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2006;
  assign dataGroup_lo_hi_2006 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2007;
  assign dataGroup_lo_hi_2007 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2008;
  assign dataGroup_lo_hi_2008 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2009;
  assign dataGroup_lo_hi_2009 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2010;
  assign dataGroup_lo_hi_2010 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2011;
  assign dataGroup_lo_hi_2011 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2012;
  assign dataGroup_lo_hi_2012 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2013;
  assign dataGroup_lo_hi_2013 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2014;
  assign dataGroup_lo_hi_2014 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2015;
  assign dataGroup_lo_hi_2015 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2016;
  assign dataGroup_lo_hi_2016 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2017;
  assign dataGroup_lo_hi_2017 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2018;
  assign dataGroup_lo_hi_2018 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2019;
  assign dataGroup_lo_hi_2019 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2020;
  assign dataGroup_lo_hi_2020 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2021;
  assign dataGroup_lo_hi_2021 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2022;
  assign dataGroup_lo_hi_2022 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2023;
  assign dataGroup_lo_hi_2023 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2024;
  assign dataGroup_lo_hi_2024 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2025;
  assign dataGroup_lo_hi_2025 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2026;
  assign dataGroup_lo_hi_2026 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2027;
  assign dataGroup_lo_hi_2027 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2028;
  assign dataGroup_lo_hi_2028 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2029;
  assign dataGroup_lo_hi_2029 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2030;
  assign dataGroup_lo_hi_2030 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2031;
  assign dataGroup_lo_hi_2031 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2032;
  assign dataGroup_lo_hi_2032 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2033;
  assign dataGroup_lo_hi_2033 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2034;
  assign dataGroup_lo_hi_2034 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2035;
  assign dataGroup_lo_hi_2035 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2036;
  assign dataGroup_lo_hi_2036 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2037;
  assign dataGroup_lo_hi_2037 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2038;
  assign dataGroup_lo_hi_2038 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2039;
  assign dataGroup_lo_hi_2039 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2040;
  assign dataGroup_lo_hi_2040 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2041;
  assign dataGroup_lo_hi_2041 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2042;
  assign dataGroup_lo_hi_2042 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2043;
  assign dataGroup_lo_hi_2043 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2044;
  assign dataGroup_lo_hi_2044 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2045;
  assign dataGroup_lo_hi_2045 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2046;
  assign dataGroup_lo_hi_2046 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2047;
  assign dataGroup_lo_hi_2047 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2048;
  assign dataGroup_lo_hi_2048 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2049;
  assign dataGroup_lo_hi_2049 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2050;
  assign dataGroup_lo_hi_2050 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2051;
  assign dataGroup_lo_hi_2051 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2052;
  assign dataGroup_lo_hi_2052 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2053;
  assign dataGroup_lo_hi_2053 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2054;
  assign dataGroup_lo_hi_2054 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2055;
  assign dataGroup_lo_hi_2055 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2056;
  assign dataGroup_lo_hi_2056 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2057;
  assign dataGroup_lo_hi_2057 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2058;
  assign dataGroup_lo_hi_2058 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2059;
  assign dataGroup_lo_hi_2059 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2060;
  assign dataGroup_lo_hi_2060 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2061;
  assign dataGroup_lo_hi_2061 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2062;
  assign dataGroup_lo_hi_2062 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2063;
  assign dataGroup_lo_hi_2063 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2064;
  assign dataGroup_lo_hi_2064 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2065;
  assign dataGroup_lo_hi_2065 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2066;
  assign dataGroup_lo_hi_2066 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2067;
  assign dataGroup_lo_hi_2067 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2068;
  assign dataGroup_lo_hi_2068 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2069;
  assign dataGroup_lo_hi_2069 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2070;
  assign dataGroup_lo_hi_2070 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2071;
  assign dataGroup_lo_hi_2071 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2072;
  assign dataGroup_lo_hi_2072 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2073;
  assign dataGroup_lo_hi_2073 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2074;
  assign dataGroup_lo_hi_2074 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2075;
  assign dataGroup_lo_hi_2075 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2076;
  assign dataGroup_lo_hi_2076 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2077;
  assign dataGroup_lo_hi_2077 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2078;
  assign dataGroup_lo_hi_2078 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2079;
  assign dataGroup_lo_hi_2079 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2080;
  assign dataGroup_lo_hi_2080 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2081;
  assign dataGroup_lo_hi_2081 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2082;
  assign dataGroup_lo_hi_2082 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2083;
  assign dataGroup_lo_hi_2083 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2084;
  assign dataGroup_lo_hi_2084 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2085;
  assign dataGroup_lo_hi_2085 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2086;
  assign dataGroup_lo_hi_2086 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2087;
  assign dataGroup_lo_hi_2087 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2088;
  assign dataGroup_lo_hi_2088 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2089;
  assign dataGroup_lo_hi_2089 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2090;
  assign dataGroup_lo_hi_2090 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2091;
  assign dataGroup_lo_hi_2091 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2092;
  assign dataGroup_lo_hi_2092 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2093;
  assign dataGroup_lo_hi_2093 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2094;
  assign dataGroup_lo_hi_2094 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2095;
  assign dataGroup_lo_hi_2095 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2096;
  assign dataGroup_lo_hi_2096 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2097;
  assign dataGroup_lo_hi_2097 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2098;
  assign dataGroup_lo_hi_2098 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2099;
  assign dataGroup_lo_hi_2099 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2100;
  assign dataGroup_lo_hi_2100 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2101;
  assign dataGroup_lo_hi_2101 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2102;
  assign dataGroup_lo_hi_2102 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2103;
  assign dataGroup_lo_hi_2103 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2104;
  assign dataGroup_lo_hi_2104 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2105;
  assign dataGroup_lo_hi_2105 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2106;
  assign dataGroup_lo_hi_2106 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2107;
  assign dataGroup_lo_hi_2107 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2108;
  assign dataGroup_lo_hi_2108 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2109;
  assign dataGroup_lo_hi_2109 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2110;
  assign dataGroup_lo_hi_2110 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2111;
  assign dataGroup_lo_hi_2111 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2112;
  assign dataGroup_lo_hi_2112 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2113;
  assign dataGroup_lo_hi_2113 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2114;
  assign dataGroup_lo_hi_2114 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2115;
  assign dataGroup_lo_hi_2115 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2116;
  assign dataGroup_lo_hi_2116 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2117;
  assign dataGroup_lo_hi_2117 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2118;
  assign dataGroup_lo_hi_2118 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2119;
  assign dataGroup_lo_hi_2119 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2120;
  assign dataGroup_lo_hi_2120 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2121;
  assign dataGroup_lo_hi_2121 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2122;
  assign dataGroup_lo_hi_2122 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2123;
  assign dataGroup_lo_hi_2123 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2124;
  assign dataGroup_lo_hi_2124 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2125;
  assign dataGroup_lo_hi_2125 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2126;
  assign dataGroup_lo_hi_2126 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2127;
  assign dataGroup_lo_hi_2127 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2128;
  assign dataGroup_lo_hi_2128 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2129;
  assign dataGroup_lo_hi_2129 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2130;
  assign dataGroup_lo_hi_2130 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2131;
  assign dataGroup_lo_hi_2131 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2132;
  assign dataGroup_lo_hi_2132 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2133;
  assign dataGroup_lo_hi_2133 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2134;
  assign dataGroup_lo_hi_2134 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2135;
  assign dataGroup_lo_hi_2135 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2136;
  assign dataGroup_lo_hi_2136 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2137;
  assign dataGroup_lo_hi_2137 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2138;
  assign dataGroup_lo_hi_2138 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2139;
  assign dataGroup_lo_hi_2139 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2140;
  assign dataGroup_lo_hi_2140 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2141;
  assign dataGroup_lo_hi_2141 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2142;
  assign dataGroup_lo_hi_2142 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2143;
  assign dataGroup_lo_hi_2143 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2144;
  assign dataGroup_lo_hi_2144 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2145;
  assign dataGroup_lo_hi_2145 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2146;
  assign dataGroup_lo_hi_2146 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2147;
  assign dataGroup_lo_hi_2147 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2148;
  assign dataGroup_lo_hi_2148 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2149;
  assign dataGroup_lo_hi_2149 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2150;
  assign dataGroup_lo_hi_2150 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2151;
  assign dataGroup_lo_hi_2151 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2152;
  assign dataGroup_lo_hi_2152 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2153;
  assign dataGroup_lo_hi_2153 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2154;
  assign dataGroup_lo_hi_2154 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2155;
  assign dataGroup_lo_hi_2155 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2156;
  assign dataGroup_lo_hi_2156 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2157;
  assign dataGroup_lo_hi_2157 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2158;
  assign dataGroup_lo_hi_2158 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2159;
  assign dataGroup_lo_hi_2159 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2160;
  assign dataGroup_lo_hi_2160 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2161;
  assign dataGroup_lo_hi_2161 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2162;
  assign dataGroup_lo_hi_2162 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2163;
  assign dataGroup_lo_hi_2163 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2164;
  assign dataGroup_lo_hi_2164 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2165;
  assign dataGroup_lo_hi_2165 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2166;
  assign dataGroup_lo_hi_2166 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2167;
  assign dataGroup_lo_hi_2167 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2168;
  assign dataGroup_lo_hi_2168 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2169;
  assign dataGroup_lo_hi_2169 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2170;
  assign dataGroup_lo_hi_2170 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2171;
  assign dataGroup_lo_hi_2171 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2172;
  assign dataGroup_lo_hi_2172 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2173;
  assign dataGroup_lo_hi_2173 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2174;
  assign dataGroup_lo_hi_2174 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2175;
  assign dataGroup_lo_hi_2175 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2176;
  assign dataGroup_lo_hi_2176 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2177;
  assign dataGroup_lo_hi_2177 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2178;
  assign dataGroup_lo_hi_2178 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2179;
  assign dataGroup_lo_hi_2179 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2180;
  assign dataGroup_lo_hi_2180 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2181;
  assign dataGroup_lo_hi_2181 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2182;
  assign dataGroup_lo_hi_2182 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2183;
  assign dataGroup_lo_hi_2183 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2184;
  assign dataGroup_lo_hi_2184 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2185;
  assign dataGroup_lo_hi_2185 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2186;
  assign dataGroup_lo_hi_2186 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2187;
  assign dataGroup_lo_hi_2187 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2188;
  assign dataGroup_lo_hi_2188 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2189;
  assign dataGroup_lo_hi_2189 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2190;
  assign dataGroup_lo_hi_2190 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2191;
  assign dataGroup_lo_hi_2191 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2192;
  assign dataGroup_lo_hi_2192 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2193;
  assign dataGroup_lo_hi_2193 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2194;
  assign dataGroup_lo_hi_2194 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2195;
  assign dataGroup_lo_hi_2195 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2196;
  assign dataGroup_lo_hi_2196 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2197;
  assign dataGroup_lo_hi_2197 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2198;
  assign dataGroup_lo_hi_2198 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2199;
  assign dataGroup_lo_hi_2199 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2200;
  assign dataGroup_lo_hi_2200 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2201;
  assign dataGroup_lo_hi_2201 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2202;
  assign dataGroup_lo_hi_2202 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2203;
  assign dataGroup_lo_hi_2203 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2204;
  assign dataGroup_lo_hi_2204 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2205;
  assign dataGroup_lo_hi_2205 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2206;
  assign dataGroup_lo_hi_2206 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2207;
  assign dataGroup_lo_hi_2207 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2208;
  assign dataGroup_lo_hi_2208 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2209;
  assign dataGroup_lo_hi_2209 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2210;
  assign dataGroup_lo_hi_2210 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2211;
  assign dataGroup_lo_hi_2211 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2212;
  assign dataGroup_lo_hi_2212 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2213;
  assign dataGroup_lo_hi_2213 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2214;
  assign dataGroup_lo_hi_2214 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2215;
  assign dataGroup_lo_hi_2215 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2216;
  assign dataGroup_lo_hi_2216 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2217;
  assign dataGroup_lo_hi_2217 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2218;
  assign dataGroup_lo_hi_2218 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2219;
  assign dataGroup_lo_hi_2219 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2220;
  assign dataGroup_lo_hi_2220 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2221;
  assign dataGroup_lo_hi_2221 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2222;
  assign dataGroup_lo_hi_2222 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2223;
  assign dataGroup_lo_hi_2223 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2224;
  assign dataGroup_lo_hi_2224 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2225;
  assign dataGroup_lo_hi_2225 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2226;
  assign dataGroup_lo_hi_2226 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2227;
  assign dataGroup_lo_hi_2227 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2228;
  assign dataGroup_lo_hi_2228 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2229;
  assign dataGroup_lo_hi_2229 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2230;
  assign dataGroup_lo_hi_2230 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2231;
  assign dataGroup_lo_hi_2231 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2232;
  assign dataGroup_lo_hi_2232 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2233;
  assign dataGroup_lo_hi_2233 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2234;
  assign dataGroup_lo_hi_2234 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2235;
  assign dataGroup_lo_hi_2235 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2236;
  assign dataGroup_lo_hi_2236 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2237;
  assign dataGroup_lo_hi_2237 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2238;
  assign dataGroup_lo_hi_2238 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2239;
  assign dataGroup_lo_hi_2239 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2240;
  assign dataGroup_lo_hi_2240 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2241;
  assign dataGroup_lo_hi_2241 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2242;
  assign dataGroup_lo_hi_2242 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2243;
  assign dataGroup_lo_hi_2243 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2244;
  assign dataGroup_lo_hi_2244 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2245;
  assign dataGroup_lo_hi_2245 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2246;
  assign dataGroup_lo_hi_2246 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2247;
  assign dataGroup_lo_hi_2247 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2248;
  assign dataGroup_lo_hi_2248 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2249;
  assign dataGroup_lo_hi_2249 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2250;
  assign dataGroup_lo_hi_2250 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2251;
  assign dataGroup_lo_hi_2251 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2252;
  assign dataGroup_lo_hi_2252 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2253;
  assign dataGroup_lo_hi_2253 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2254;
  assign dataGroup_lo_hi_2254 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2255;
  assign dataGroup_lo_hi_2255 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2256;
  assign dataGroup_lo_hi_2256 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2257;
  assign dataGroup_lo_hi_2257 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2258;
  assign dataGroup_lo_hi_2258 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2259;
  assign dataGroup_lo_hi_2259 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2260;
  assign dataGroup_lo_hi_2260 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2261;
  assign dataGroup_lo_hi_2261 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2262;
  assign dataGroup_lo_hi_2262 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2263;
  assign dataGroup_lo_hi_2263 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2264;
  assign dataGroup_lo_hi_2264 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2265;
  assign dataGroup_lo_hi_2265 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2266;
  assign dataGroup_lo_hi_2266 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2267;
  assign dataGroup_lo_hi_2267 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2268;
  assign dataGroup_lo_hi_2268 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2269;
  assign dataGroup_lo_hi_2269 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2270;
  assign dataGroup_lo_hi_2270 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2271;
  assign dataGroup_lo_hi_2271 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2272;
  assign dataGroup_lo_hi_2272 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2273;
  assign dataGroup_lo_hi_2273 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2274;
  assign dataGroup_lo_hi_2274 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2275;
  assign dataGroup_lo_hi_2275 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2276;
  assign dataGroup_lo_hi_2276 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2277;
  assign dataGroup_lo_hi_2277 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2278;
  assign dataGroup_lo_hi_2278 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2279;
  assign dataGroup_lo_hi_2279 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2280;
  assign dataGroup_lo_hi_2280 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2281;
  assign dataGroup_lo_hi_2281 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2282;
  assign dataGroup_lo_hi_2282 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2283;
  assign dataGroup_lo_hi_2283 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2284;
  assign dataGroup_lo_hi_2284 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2285;
  assign dataGroup_lo_hi_2285 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2286;
  assign dataGroup_lo_hi_2286 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2287;
  assign dataGroup_lo_hi_2287 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2288;
  assign dataGroup_lo_hi_2288 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2289;
  assign dataGroup_lo_hi_2289 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2290;
  assign dataGroup_lo_hi_2290 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2291;
  assign dataGroup_lo_hi_2291 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2292;
  assign dataGroup_lo_hi_2292 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2293;
  assign dataGroup_lo_hi_2293 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2294;
  assign dataGroup_lo_hi_2294 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2295;
  assign dataGroup_lo_hi_2295 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2296;
  assign dataGroup_lo_hi_2296 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2297;
  assign dataGroup_lo_hi_2297 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2298;
  assign dataGroup_lo_hi_2298 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2299;
  assign dataGroup_lo_hi_2299 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2300;
  assign dataGroup_lo_hi_2300 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2301;
  assign dataGroup_lo_hi_2301 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2302;
  assign dataGroup_lo_hi_2302 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2303;
  assign dataGroup_lo_hi_2303 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2304;
  assign dataGroup_lo_hi_2304 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2305;
  assign dataGroup_lo_hi_2305 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2306;
  assign dataGroup_lo_hi_2306 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2307;
  assign dataGroup_lo_hi_2307 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2308;
  assign dataGroup_lo_hi_2308 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2309;
  assign dataGroup_lo_hi_2309 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2310;
  assign dataGroup_lo_hi_2310 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2311;
  assign dataGroup_lo_hi_2311 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2312;
  assign dataGroup_lo_hi_2312 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2313;
  assign dataGroup_lo_hi_2313 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2314;
  assign dataGroup_lo_hi_2314 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2315;
  assign dataGroup_lo_hi_2315 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2316;
  assign dataGroup_lo_hi_2316 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2317;
  assign dataGroup_lo_hi_2317 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2318;
  assign dataGroup_lo_hi_2318 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2319;
  assign dataGroup_lo_hi_2319 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2320;
  assign dataGroup_lo_hi_2320 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2321;
  assign dataGroup_lo_hi_2321 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2322;
  assign dataGroup_lo_hi_2322 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2323;
  assign dataGroup_lo_hi_2323 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2324;
  assign dataGroup_lo_hi_2324 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2325;
  assign dataGroup_lo_hi_2325 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2326;
  assign dataGroup_lo_hi_2326 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2327;
  assign dataGroup_lo_hi_2327 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2328;
  assign dataGroup_lo_hi_2328 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2329;
  assign dataGroup_lo_hi_2329 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2330;
  assign dataGroup_lo_hi_2330 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2331;
  assign dataGroup_lo_hi_2331 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2332;
  assign dataGroup_lo_hi_2332 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2333;
  assign dataGroup_lo_hi_2333 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2334;
  assign dataGroup_lo_hi_2334 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2335;
  assign dataGroup_lo_hi_2335 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2336;
  assign dataGroup_lo_hi_2336 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2337;
  assign dataGroup_lo_hi_2337 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2338;
  assign dataGroup_lo_hi_2338 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2339;
  assign dataGroup_lo_hi_2339 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2340;
  assign dataGroup_lo_hi_2340 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2341;
  assign dataGroup_lo_hi_2341 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2342;
  assign dataGroup_lo_hi_2342 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2343;
  assign dataGroup_lo_hi_2343 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2344;
  assign dataGroup_lo_hi_2344 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2345;
  assign dataGroup_lo_hi_2345 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2346;
  assign dataGroup_lo_hi_2346 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2347;
  assign dataGroup_lo_hi_2347 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2348;
  assign dataGroup_lo_hi_2348 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2349;
  assign dataGroup_lo_hi_2349 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2350;
  assign dataGroup_lo_hi_2350 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2351;
  assign dataGroup_lo_hi_2351 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2352;
  assign dataGroup_lo_hi_2352 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2353;
  assign dataGroup_lo_hi_2353 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2354;
  assign dataGroup_lo_hi_2354 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2355;
  assign dataGroup_lo_hi_2355 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2356;
  assign dataGroup_lo_hi_2356 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2357;
  assign dataGroup_lo_hi_2357 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2358;
  assign dataGroup_lo_hi_2358 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2359;
  assign dataGroup_lo_hi_2359 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2360;
  assign dataGroup_lo_hi_2360 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2361;
  assign dataGroup_lo_hi_2361 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2362;
  assign dataGroup_lo_hi_2362 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2363;
  assign dataGroup_lo_hi_2363 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2364;
  assign dataGroup_lo_hi_2364 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2365;
  assign dataGroup_lo_hi_2365 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2366;
  assign dataGroup_lo_hi_2366 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2367;
  assign dataGroup_lo_hi_2367 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2368;
  assign dataGroup_lo_hi_2368 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2369;
  assign dataGroup_lo_hi_2369 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2370;
  assign dataGroup_lo_hi_2370 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2371;
  assign dataGroup_lo_hi_2371 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2372;
  assign dataGroup_lo_hi_2372 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2373;
  assign dataGroup_lo_hi_2373 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2374;
  assign dataGroup_lo_hi_2374 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2375;
  assign dataGroup_lo_hi_2375 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2376;
  assign dataGroup_lo_hi_2376 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2377;
  assign dataGroup_lo_hi_2377 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2378;
  assign dataGroup_lo_hi_2378 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2379;
  assign dataGroup_lo_hi_2379 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2380;
  assign dataGroup_lo_hi_2380 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2381;
  assign dataGroup_lo_hi_2381 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2382;
  assign dataGroup_lo_hi_2382 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2383;
  assign dataGroup_lo_hi_2383 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2384;
  assign dataGroup_lo_hi_2384 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2385;
  assign dataGroup_lo_hi_2385 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2386;
  assign dataGroup_lo_hi_2386 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2387;
  assign dataGroup_lo_hi_2387 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2388;
  assign dataGroup_lo_hi_2388 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2389;
  assign dataGroup_lo_hi_2389 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2390;
  assign dataGroup_lo_hi_2390 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2391;
  assign dataGroup_lo_hi_2391 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2392;
  assign dataGroup_lo_hi_2392 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2393;
  assign dataGroup_lo_hi_2393 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2394;
  assign dataGroup_lo_hi_2394 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2395;
  assign dataGroup_lo_hi_2395 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2396;
  assign dataGroup_lo_hi_2396 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2397;
  assign dataGroup_lo_hi_2397 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2398;
  assign dataGroup_lo_hi_2398 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2399;
  assign dataGroup_lo_hi_2399 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2400;
  assign dataGroup_lo_hi_2400 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2401;
  assign dataGroup_lo_hi_2401 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2402;
  assign dataGroup_lo_hi_2402 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2403;
  assign dataGroup_lo_hi_2403 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2404;
  assign dataGroup_lo_hi_2404 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2405;
  assign dataGroup_lo_hi_2405 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2406;
  assign dataGroup_lo_hi_2406 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2407;
  assign dataGroup_lo_hi_2407 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2408;
  assign dataGroup_lo_hi_2408 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2409;
  assign dataGroup_lo_hi_2409 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2410;
  assign dataGroup_lo_hi_2410 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2411;
  assign dataGroup_lo_hi_2411 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2412;
  assign dataGroup_lo_hi_2412 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2413;
  assign dataGroup_lo_hi_2413 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2414;
  assign dataGroup_lo_hi_2414 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2415;
  assign dataGroup_lo_hi_2415 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2416;
  assign dataGroup_lo_hi_2416 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2417;
  assign dataGroup_lo_hi_2417 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2418;
  assign dataGroup_lo_hi_2418 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2419;
  assign dataGroup_lo_hi_2419 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2420;
  assign dataGroup_lo_hi_2420 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2421;
  assign dataGroup_lo_hi_2421 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2422;
  assign dataGroup_lo_hi_2422 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2423;
  assign dataGroup_lo_hi_2423 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2424;
  assign dataGroup_lo_hi_2424 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2425;
  assign dataGroup_lo_hi_2425 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2426;
  assign dataGroup_lo_hi_2426 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2427;
  assign dataGroup_lo_hi_2427 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2428;
  assign dataGroup_lo_hi_2428 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2429;
  assign dataGroup_lo_hi_2429 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2430;
  assign dataGroup_lo_hi_2430 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2431;
  assign dataGroup_lo_hi_2431 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2432;
  assign dataGroup_lo_hi_2432 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2433;
  assign dataGroup_lo_hi_2433 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2434;
  assign dataGroup_lo_hi_2434 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2435;
  assign dataGroup_lo_hi_2435 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2436;
  assign dataGroup_lo_hi_2436 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2437;
  assign dataGroup_lo_hi_2437 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2438;
  assign dataGroup_lo_hi_2438 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2439;
  assign dataGroup_lo_hi_2439 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2440;
  assign dataGroup_lo_hi_2440 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2441;
  assign dataGroup_lo_hi_2441 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2442;
  assign dataGroup_lo_hi_2442 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2443;
  assign dataGroup_lo_hi_2443 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2444;
  assign dataGroup_lo_hi_2444 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2445;
  assign dataGroup_lo_hi_2445 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2446;
  assign dataGroup_lo_hi_2446 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2447;
  assign dataGroup_lo_hi_2447 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2448;
  assign dataGroup_lo_hi_2448 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2449;
  assign dataGroup_lo_hi_2449 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2450;
  assign dataGroup_lo_hi_2450 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2451;
  assign dataGroup_lo_hi_2451 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2452;
  assign dataGroup_lo_hi_2452 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2453;
  assign dataGroup_lo_hi_2453 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2454;
  assign dataGroup_lo_hi_2454 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2455;
  assign dataGroup_lo_hi_2455 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2456;
  assign dataGroup_lo_hi_2456 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2457;
  assign dataGroup_lo_hi_2457 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2458;
  assign dataGroup_lo_hi_2458 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2459;
  assign dataGroup_lo_hi_2459 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2460;
  assign dataGroup_lo_hi_2460 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2461;
  assign dataGroup_lo_hi_2461 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2462;
  assign dataGroup_lo_hi_2462 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2463;
  assign dataGroup_lo_hi_2463 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2464;
  assign dataGroup_lo_hi_2464 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2465;
  assign dataGroup_lo_hi_2465 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2466;
  assign dataGroup_lo_hi_2466 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2467;
  assign dataGroup_lo_hi_2467 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2468;
  assign dataGroup_lo_hi_2468 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2469;
  assign dataGroup_lo_hi_2469 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2470;
  assign dataGroup_lo_hi_2470 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2471;
  assign dataGroup_lo_hi_2471 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2472;
  assign dataGroup_lo_hi_2472 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2473;
  assign dataGroup_lo_hi_2473 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2474;
  assign dataGroup_lo_hi_2474 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2475;
  assign dataGroup_lo_hi_2475 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2476;
  assign dataGroup_lo_hi_2476 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2477;
  assign dataGroup_lo_hi_2477 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2478;
  assign dataGroup_lo_hi_2478 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2479;
  assign dataGroup_lo_hi_2479 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2480;
  assign dataGroup_lo_hi_2480 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2481;
  assign dataGroup_lo_hi_2481 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2482;
  assign dataGroup_lo_hi_2482 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2483;
  assign dataGroup_lo_hi_2483 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2484;
  assign dataGroup_lo_hi_2484 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2485;
  assign dataGroup_lo_hi_2485 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2486;
  assign dataGroup_lo_hi_2486 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2487;
  assign dataGroup_lo_hi_2487 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2488;
  assign dataGroup_lo_hi_2488 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2489;
  assign dataGroup_lo_hi_2489 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2490;
  assign dataGroup_lo_hi_2490 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2491;
  assign dataGroup_lo_hi_2491 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2492;
  assign dataGroup_lo_hi_2492 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2493;
  assign dataGroup_lo_hi_2493 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2494;
  assign dataGroup_lo_hi_2494 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2495;
  assign dataGroup_lo_hi_2495 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2496;
  assign dataGroup_lo_hi_2496 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2497;
  assign dataGroup_lo_hi_2497 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2498;
  assign dataGroup_lo_hi_2498 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2499;
  assign dataGroup_lo_hi_2499 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2500;
  assign dataGroup_lo_hi_2500 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2501;
  assign dataGroup_lo_hi_2501 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2502;
  assign dataGroup_lo_hi_2502 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2503;
  assign dataGroup_lo_hi_2503 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2504;
  assign dataGroup_lo_hi_2504 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2505;
  assign dataGroup_lo_hi_2505 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2506;
  assign dataGroup_lo_hi_2506 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2507;
  assign dataGroup_lo_hi_2507 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2508;
  assign dataGroup_lo_hi_2508 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2509;
  assign dataGroup_lo_hi_2509 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2510;
  assign dataGroup_lo_hi_2510 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2511;
  assign dataGroup_lo_hi_2511 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2512;
  assign dataGroup_lo_hi_2512 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2513;
  assign dataGroup_lo_hi_2513 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2514;
  assign dataGroup_lo_hi_2514 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2515;
  assign dataGroup_lo_hi_2515 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2516;
  assign dataGroup_lo_hi_2516 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2517;
  assign dataGroup_lo_hi_2517 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2518;
  assign dataGroup_lo_hi_2518 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2519;
  assign dataGroup_lo_hi_2519 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2520;
  assign dataGroup_lo_hi_2520 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2521;
  assign dataGroup_lo_hi_2521 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2522;
  assign dataGroup_lo_hi_2522 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2523;
  assign dataGroup_lo_hi_2523 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2524;
  assign dataGroup_lo_hi_2524 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2525;
  assign dataGroup_lo_hi_2525 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2526;
  assign dataGroup_lo_hi_2526 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2527;
  assign dataGroup_lo_hi_2527 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2528;
  assign dataGroup_lo_hi_2528 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2529;
  assign dataGroup_lo_hi_2529 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2530;
  assign dataGroup_lo_hi_2530 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2531;
  assign dataGroup_lo_hi_2531 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2532;
  assign dataGroup_lo_hi_2532 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2533;
  assign dataGroup_lo_hi_2533 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2534;
  assign dataGroup_lo_hi_2534 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2535;
  assign dataGroup_lo_hi_2535 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2536;
  assign dataGroup_lo_hi_2536 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2537;
  assign dataGroup_lo_hi_2537 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2538;
  assign dataGroup_lo_hi_2538 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2539;
  assign dataGroup_lo_hi_2539 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2540;
  assign dataGroup_lo_hi_2540 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2541;
  assign dataGroup_lo_hi_2541 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2542;
  assign dataGroup_lo_hi_2542 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2543;
  assign dataGroup_lo_hi_2543 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2544;
  assign dataGroup_lo_hi_2544 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2545;
  assign dataGroup_lo_hi_2545 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2546;
  assign dataGroup_lo_hi_2546 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2547;
  assign dataGroup_lo_hi_2547 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2548;
  assign dataGroup_lo_hi_2548 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2549;
  assign dataGroup_lo_hi_2549 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2550;
  assign dataGroup_lo_hi_2550 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2551;
  assign dataGroup_lo_hi_2551 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2552;
  assign dataGroup_lo_hi_2552 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2553;
  assign dataGroup_lo_hi_2553 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2554;
  assign dataGroup_lo_hi_2554 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2555;
  assign dataGroup_lo_hi_2555 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2556;
  assign dataGroup_lo_hi_2556 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2557;
  assign dataGroup_lo_hi_2557 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2558;
  assign dataGroup_lo_hi_2558 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2559;
  assign dataGroup_lo_hi_2559 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2560;
  assign dataGroup_lo_hi_2560 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2561;
  assign dataGroup_lo_hi_2561 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2562;
  assign dataGroup_lo_hi_2562 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2563;
  assign dataGroup_lo_hi_2563 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2564;
  assign dataGroup_lo_hi_2564 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2565;
  assign dataGroup_lo_hi_2565 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2566;
  assign dataGroup_lo_hi_2566 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2567;
  assign dataGroup_lo_hi_2567 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2568;
  assign dataGroup_lo_hi_2568 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2569;
  assign dataGroup_lo_hi_2569 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2570;
  assign dataGroup_lo_hi_2570 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2571;
  assign dataGroup_lo_hi_2571 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2572;
  assign dataGroup_lo_hi_2572 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2573;
  assign dataGroup_lo_hi_2573 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2574;
  assign dataGroup_lo_hi_2574 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2575;
  assign dataGroup_lo_hi_2575 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2576;
  assign dataGroup_lo_hi_2576 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2577;
  assign dataGroup_lo_hi_2577 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2578;
  assign dataGroup_lo_hi_2578 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2579;
  assign dataGroup_lo_hi_2579 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2580;
  assign dataGroup_lo_hi_2580 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2581;
  assign dataGroup_lo_hi_2581 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2582;
  assign dataGroup_lo_hi_2582 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2583;
  assign dataGroup_lo_hi_2583 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2584;
  assign dataGroup_lo_hi_2584 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2585;
  assign dataGroup_lo_hi_2585 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2586;
  assign dataGroup_lo_hi_2586 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2587;
  assign dataGroup_lo_hi_2587 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2588;
  assign dataGroup_lo_hi_2588 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2589;
  assign dataGroup_lo_hi_2589 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2590;
  assign dataGroup_lo_hi_2590 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2591;
  assign dataGroup_lo_hi_2591 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2592;
  assign dataGroup_lo_hi_2592 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2593;
  assign dataGroup_lo_hi_2593 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2594;
  assign dataGroup_lo_hi_2594 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2595;
  assign dataGroup_lo_hi_2595 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2596;
  assign dataGroup_lo_hi_2596 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2597;
  assign dataGroup_lo_hi_2597 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2598;
  assign dataGroup_lo_hi_2598 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2599;
  assign dataGroup_lo_hi_2599 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2600;
  assign dataGroup_lo_hi_2600 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2601;
  assign dataGroup_lo_hi_2601 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2602;
  assign dataGroup_lo_hi_2602 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2603;
  assign dataGroup_lo_hi_2603 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2604;
  assign dataGroup_lo_hi_2604 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2605;
  assign dataGroup_lo_hi_2605 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2606;
  assign dataGroup_lo_hi_2606 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2607;
  assign dataGroup_lo_hi_2607 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2608;
  assign dataGroup_lo_hi_2608 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2609;
  assign dataGroup_lo_hi_2609 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2610;
  assign dataGroup_lo_hi_2610 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2611;
  assign dataGroup_lo_hi_2611 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2612;
  assign dataGroup_lo_hi_2612 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2613;
  assign dataGroup_lo_hi_2613 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2614;
  assign dataGroup_lo_hi_2614 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2615;
  assign dataGroup_lo_hi_2615 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2616;
  assign dataGroup_lo_hi_2616 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2617;
  assign dataGroup_lo_hi_2617 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2618;
  assign dataGroup_lo_hi_2618 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2619;
  assign dataGroup_lo_hi_2619 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2620;
  assign dataGroup_lo_hi_2620 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2621;
  assign dataGroup_lo_hi_2621 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2622;
  assign dataGroup_lo_hi_2622 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2623;
  assign dataGroup_lo_hi_2623 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2624;
  assign dataGroup_lo_hi_2624 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2625;
  assign dataGroup_lo_hi_2625 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2626;
  assign dataGroup_lo_hi_2626 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2627;
  assign dataGroup_lo_hi_2627 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2628;
  assign dataGroup_lo_hi_2628 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2629;
  assign dataGroup_lo_hi_2629 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2630;
  assign dataGroup_lo_hi_2630 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2631;
  assign dataGroup_lo_hi_2631 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2632;
  assign dataGroup_lo_hi_2632 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2633;
  assign dataGroup_lo_hi_2633 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2634;
  assign dataGroup_lo_hi_2634 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2635;
  assign dataGroup_lo_hi_2635 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2636;
  assign dataGroup_lo_hi_2636 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2637;
  assign dataGroup_lo_hi_2637 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2638;
  assign dataGroup_lo_hi_2638 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2639;
  assign dataGroup_lo_hi_2639 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2640;
  assign dataGroup_lo_hi_2640 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2641;
  assign dataGroup_lo_hi_2641 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2642;
  assign dataGroup_lo_hi_2642 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2643;
  assign dataGroup_lo_hi_2643 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2644;
  assign dataGroup_lo_hi_2644 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2645;
  assign dataGroup_lo_hi_2645 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2646;
  assign dataGroup_lo_hi_2646 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2647;
  assign dataGroup_lo_hi_2647 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2648;
  assign dataGroup_lo_hi_2648 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2649;
  assign dataGroup_lo_hi_2649 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2650;
  assign dataGroup_lo_hi_2650 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2651;
  assign dataGroup_lo_hi_2651 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2652;
  assign dataGroup_lo_hi_2652 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2653;
  assign dataGroup_lo_hi_2653 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2654;
  assign dataGroup_lo_hi_2654 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2655;
  assign dataGroup_lo_hi_2655 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2656;
  assign dataGroup_lo_hi_2656 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2657;
  assign dataGroup_lo_hi_2657 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2658;
  assign dataGroup_lo_hi_2658 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2659;
  assign dataGroup_lo_hi_2659 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2660;
  assign dataGroup_lo_hi_2660 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2661;
  assign dataGroup_lo_hi_2661 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2662;
  assign dataGroup_lo_hi_2662 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2663;
  assign dataGroup_lo_hi_2663 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2664;
  assign dataGroup_lo_hi_2664 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2665;
  assign dataGroup_lo_hi_2665 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2666;
  assign dataGroup_lo_hi_2666 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2667;
  assign dataGroup_lo_hi_2667 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2668;
  assign dataGroup_lo_hi_2668 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2669;
  assign dataGroup_lo_hi_2669 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2670;
  assign dataGroup_lo_hi_2670 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2671;
  assign dataGroup_lo_hi_2671 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2672;
  assign dataGroup_lo_hi_2672 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2673;
  assign dataGroup_lo_hi_2673 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2674;
  assign dataGroup_lo_hi_2674 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2675;
  assign dataGroup_lo_hi_2675 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2676;
  assign dataGroup_lo_hi_2676 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2677;
  assign dataGroup_lo_hi_2677 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2678;
  assign dataGroup_lo_hi_2678 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2679;
  assign dataGroup_lo_hi_2679 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2680;
  assign dataGroup_lo_hi_2680 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2681;
  assign dataGroup_lo_hi_2681 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2682;
  assign dataGroup_lo_hi_2682 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2683;
  assign dataGroup_lo_hi_2683 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2684;
  assign dataGroup_lo_hi_2684 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2685;
  assign dataGroup_lo_hi_2685 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2686;
  assign dataGroup_lo_hi_2686 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2687;
  assign dataGroup_lo_hi_2687 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2688;
  assign dataGroup_lo_hi_2688 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2689;
  assign dataGroup_lo_hi_2689 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2690;
  assign dataGroup_lo_hi_2690 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2691;
  assign dataGroup_lo_hi_2691 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2692;
  assign dataGroup_lo_hi_2692 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2693;
  assign dataGroup_lo_hi_2693 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2694;
  assign dataGroup_lo_hi_2694 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2695;
  assign dataGroup_lo_hi_2695 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2696;
  assign dataGroup_lo_hi_2696 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2697;
  assign dataGroup_lo_hi_2697 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2698;
  assign dataGroup_lo_hi_2698 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2699;
  assign dataGroup_lo_hi_2699 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2700;
  assign dataGroup_lo_hi_2700 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2701;
  assign dataGroup_lo_hi_2701 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2702;
  assign dataGroup_lo_hi_2702 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2703;
  assign dataGroup_lo_hi_2703 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2704;
  assign dataGroup_lo_hi_2704 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2705;
  assign dataGroup_lo_hi_2705 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2706;
  assign dataGroup_lo_hi_2706 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2707;
  assign dataGroup_lo_hi_2707 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2708;
  assign dataGroup_lo_hi_2708 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2709;
  assign dataGroup_lo_hi_2709 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2710;
  assign dataGroup_lo_hi_2710 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2711;
  assign dataGroup_lo_hi_2711 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2712;
  assign dataGroup_lo_hi_2712 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2713;
  assign dataGroup_lo_hi_2713 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2714;
  assign dataGroup_lo_hi_2714 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2715;
  assign dataGroup_lo_hi_2715 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2716;
  assign dataGroup_lo_hi_2716 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2717;
  assign dataGroup_lo_hi_2717 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2718;
  assign dataGroup_lo_hi_2718 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2719;
  assign dataGroup_lo_hi_2719 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2720;
  assign dataGroup_lo_hi_2720 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2721;
  assign dataGroup_lo_hi_2721 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2722;
  assign dataGroup_lo_hi_2722 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2723;
  assign dataGroup_lo_hi_2723 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2724;
  assign dataGroup_lo_hi_2724 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2725;
  assign dataGroup_lo_hi_2725 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2726;
  assign dataGroup_lo_hi_2726 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2727;
  assign dataGroup_lo_hi_2727 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2728;
  assign dataGroup_lo_hi_2728 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2729;
  assign dataGroup_lo_hi_2729 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2730;
  assign dataGroup_lo_hi_2730 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2731;
  assign dataGroup_lo_hi_2731 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2732;
  assign dataGroup_lo_hi_2732 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2733;
  assign dataGroup_lo_hi_2733 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2734;
  assign dataGroup_lo_hi_2734 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2735;
  assign dataGroup_lo_hi_2735 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2736;
  assign dataGroup_lo_hi_2736 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2737;
  assign dataGroup_lo_hi_2737 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2738;
  assign dataGroup_lo_hi_2738 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2739;
  assign dataGroup_lo_hi_2739 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2740;
  assign dataGroup_lo_hi_2740 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2741;
  assign dataGroup_lo_hi_2741 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2742;
  assign dataGroup_lo_hi_2742 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2743;
  assign dataGroup_lo_hi_2743 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2744;
  assign dataGroup_lo_hi_2744 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2745;
  assign dataGroup_lo_hi_2745 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2746;
  assign dataGroup_lo_hi_2746 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2747;
  assign dataGroup_lo_hi_2747 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2748;
  assign dataGroup_lo_hi_2748 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2749;
  assign dataGroup_lo_hi_2749 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2750;
  assign dataGroup_lo_hi_2750 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2751;
  assign dataGroup_lo_hi_2751 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2752;
  assign dataGroup_lo_hi_2752 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2753;
  assign dataGroup_lo_hi_2753 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2754;
  assign dataGroup_lo_hi_2754 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2755;
  assign dataGroup_lo_hi_2755 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2756;
  assign dataGroup_lo_hi_2756 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2757;
  assign dataGroup_lo_hi_2757 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2758;
  assign dataGroup_lo_hi_2758 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2759;
  assign dataGroup_lo_hi_2759 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2760;
  assign dataGroup_lo_hi_2760 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2761;
  assign dataGroup_lo_hi_2761 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2762;
  assign dataGroup_lo_hi_2762 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2763;
  assign dataGroup_lo_hi_2763 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2764;
  assign dataGroup_lo_hi_2764 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2765;
  assign dataGroup_lo_hi_2765 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2766;
  assign dataGroup_lo_hi_2766 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2767;
  assign dataGroup_lo_hi_2767 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2768;
  assign dataGroup_lo_hi_2768 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2769;
  assign dataGroup_lo_hi_2769 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2770;
  assign dataGroup_lo_hi_2770 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2771;
  assign dataGroup_lo_hi_2771 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2772;
  assign dataGroup_lo_hi_2772 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2773;
  assign dataGroup_lo_hi_2773 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2774;
  assign dataGroup_lo_hi_2774 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2775;
  assign dataGroup_lo_hi_2775 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2776;
  assign dataGroup_lo_hi_2776 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2777;
  assign dataGroup_lo_hi_2777 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2778;
  assign dataGroup_lo_hi_2778 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2779;
  assign dataGroup_lo_hi_2779 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2780;
  assign dataGroup_lo_hi_2780 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2781;
  assign dataGroup_lo_hi_2781 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2782;
  assign dataGroup_lo_hi_2782 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2783;
  assign dataGroup_lo_hi_2783 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2784;
  assign dataGroup_lo_hi_2784 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2785;
  assign dataGroup_lo_hi_2785 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2786;
  assign dataGroup_lo_hi_2786 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2787;
  assign dataGroup_lo_hi_2787 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2788;
  assign dataGroup_lo_hi_2788 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2789;
  assign dataGroup_lo_hi_2789 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2790;
  assign dataGroup_lo_hi_2790 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2791;
  assign dataGroup_lo_hi_2791 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2792;
  assign dataGroup_lo_hi_2792 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2793;
  assign dataGroup_lo_hi_2793 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2794;
  assign dataGroup_lo_hi_2794 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2795;
  assign dataGroup_lo_hi_2795 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2796;
  assign dataGroup_lo_hi_2796 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2797;
  assign dataGroup_lo_hi_2797 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2798;
  assign dataGroup_lo_hi_2798 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2799;
  assign dataGroup_lo_hi_2799 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2800;
  assign dataGroup_lo_hi_2800 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2801;
  assign dataGroup_lo_hi_2801 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2802;
  assign dataGroup_lo_hi_2802 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2803;
  assign dataGroup_lo_hi_2803 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2804;
  assign dataGroup_lo_hi_2804 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2805;
  assign dataGroup_lo_hi_2805 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2806;
  assign dataGroup_lo_hi_2806 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2807;
  assign dataGroup_lo_hi_2807 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2808;
  assign dataGroup_lo_hi_2808 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2809;
  assign dataGroup_lo_hi_2809 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2810;
  assign dataGroup_lo_hi_2810 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2811;
  assign dataGroup_lo_hi_2811 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2812;
  assign dataGroup_lo_hi_2812 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2813;
  assign dataGroup_lo_hi_2813 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2814;
  assign dataGroup_lo_hi_2814 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2815;
  assign dataGroup_lo_hi_2815 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2816;
  assign dataGroup_lo_hi_2816 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2817;
  assign dataGroup_lo_hi_2817 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2818;
  assign dataGroup_lo_hi_2818 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2819;
  assign dataGroup_lo_hi_2819 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2820;
  assign dataGroup_lo_hi_2820 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2821;
  assign dataGroup_lo_hi_2821 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2822;
  assign dataGroup_lo_hi_2822 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2823;
  assign dataGroup_lo_hi_2823 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2824;
  assign dataGroup_lo_hi_2824 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2825;
  assign dataGroup_lo_hi_2825 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2826;
  assign dataGroup_lo_hi_2826 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2827;
  assign dataGroup_lo_hi_2827 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2828;
  assign dataGroup_lo_hi_2828 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2829;
  assign dataGroup_lo_hi_2829 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2830;
  assign dataGroup_lo_hi_2830 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2831;
  assign dataGroup_lo_hi_2831 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2832;
  assign dataGroup_lo_hi_2832 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2833;
  assign dataGroup_lo_hi_2833 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2834;
  assign dataGroup_lo_hi_2834 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2835;
  assign dataGroup_lo_hi_2835 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2836;
  assign dataGroup_lo_hi_2836 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2837;
  assign dataGroup_lo_hi_2837 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2838;
  assign dataGroup_lo_hi_2838 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2839;
  assign dataGroup_lo_hi_2839 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2840;
  assign dataGroup_lo_hi_2840 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2841;
  assign dataGroup_lo_hi_2841 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2842;
  assign dataGroup_lo_hi_2842 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2843;
  assign dataGroup_lo_hi_2843 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2844;
  assign dataGroup_lo_hi_2844 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2845;
  assign dataGroup_lo_hi_2845 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2846;
  assign dataGroup_lo_hi_2846 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2847;
  assign dataGroup_lo_hi_2847 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2848;
  assign dataGroup_lo_hi_2848 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2849;
  assign dataGroup_lo_hi_2849 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2850;
  assign dataGroup_lo_hi_2850 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2851;
  assign dataGroup_lo_hi_2851 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2852;
  assign dataGroup_lo_hi_2852 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2853;
  assign dataGroup_lo_hi_2853 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2854;
  assign dataGroup_lo_hi_2854 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2855;
  assign dataGroup_lo_hi_2855 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2856;
  assign dataGroup_lo_hi_2856 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2857;
  assign dataGroup_lo_hi_2857 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2858;
  assign dataGroup_lo_hi_2858 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2859;
  assign dataGroup_lo_hi_2859 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2860;
  assign dataGroup_lo_hi_2860 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2861;
  assign dataGroup_lo_hi_2861 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2862;
  assign dataGroup_lo_hi_2862 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2863;
  assign dataGroup_lo_hi_2863 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2864;
  assign dataGroup_lo_hi_2864 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2865;
  assign dataGroup_lo_hi_2865 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2866;
  assign dataGroup_lo_hi_2866 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2867;
  assign dataGroup_lo_hi_2867 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2868;
  assign dataGroup_lo_hi_2868 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2869;
  assign dataGroup_lo_hi_2869 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2870;
  assign dataGroup_lo_hi_2870 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2871;
  assign dataGroup_lo_hi_2871 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2872;
  assign dataGroup_lo_hi_2872 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2873;
  assign dataGroup_lo_hi_2873 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2874;
  assign dataGroup_lo_hi_2874 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2875;
  assign dataGroup_lo_hi_2875 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2876;
  assign dataGroup_lo_hi_2876 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2877;
  assign dataGroup_lo_hi_2877 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2878;
  assign dataGroup_lo_hi_2878 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2879;
  assign dataGroup_lo_hi_2879 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2880;
  assign dataGroup_lo_hi_2880 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2881;
  assign dataGroup_lo_hi_2881 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2882;
  assign dataGroup_lo_hi_2882 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2883;
  assign dataGroup_lo_hi_2883 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2884;
  assign dataGroup_lo_hi_2884 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2885;
  assign dataGroup_lo_hi_2885 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2886;
  assign dataGroup_lo_hi_2886 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2887;
  assign dataGroup_lo_hi_2887 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2888;
  assign dataGroup_lo_hi_2888 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2889;
  assign dataGroup_lo_hi_2889 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2890;
  assign dataGroup_lo_hi_2890 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2891;
  assign dataGroup_lo_hi_2891 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2892;
  assign dataGroup_lo_hi_2892 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2893;
  assign dataGroup_lo_hi_2893 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2894;
  assign dataGroup_lo_hi_2894 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2895;
  assign dataGroup_lo_hi_2895 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2896;
  assign dataGroup_lo_hi_2896 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2897;
  assign dataGroup_lo_hi_2897 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2898;
  assign dataGroup_lo_hi_2898 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2899;
  assign dataGroup_lo_hi_2899 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2900;
  assign dataGroup_lo_hi_2900 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2901;
  assign dataGroup_lo_hi_2901 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2902;
  assign dataGroup_lo_hi_2902 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2903;
  assign dataGroup_lo_hi_2903 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2904;
  assign dataGroup_lo_hi_2904 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2905;
  assign dataGroup_lo_hi_2905 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2906;
  assign dataGroup_lo_hi_2906 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2907;
  assign dataGroup_lo_hi_2907 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2908;
  assign dataGroup_lo_hi_2908 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2909;
  assign dataGroup_lo_hi_2909 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2910;
  assign dataGroup_lo_hi_2910 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2911;
  assign dataGroup_lo_hi_2911 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2912;
  assign dataGroup_lo_hi_2912 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2913;
  assign dataGroup_lo_hi_2913 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2914;
  assign dataGroup_lo_hi_2914 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2915;
  assign dataGroup_lo_hi_2915 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2916;
  assign dataGroup_lo_hi_2916 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2917;
  assign dataGroup_lo_hi_2917 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2918;
  assign dataGroup_lo_hi_2918 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2919;
  assign dataGroup_lo_hi_2919 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2920;
  assign dataGroup_lo_hi_2920 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2921;
  assign dataGroup_lo_hi_2921 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2922;
  assign dataGroup_lo_hi_2922 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2923;
  assign dataGroup_lo_hi_2923 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2924;
  assign dataGroup_lo_hi_2924 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2925;
  assign dataGroup_lo_hi_2925 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2926;
  assign dataGroup_lo_hi_2926 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2927;
  assign dataGroup_lo_hi_2927 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2928;
  assign dataGroup_lo_hi_2928 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2929;
  assign dataGroup_lo_hi_2929 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2930;
  assign dataGroup_lo_hi_2930 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2931;
  assign dataGroup_lo_hi_2931 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2932;
  assign dataGroup_lo_hi_2932 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2933;
  assign dataGroup_lo_hi_2933 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2934;
  assign dataGroup_lo_hi_2934 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2935;
  assign dataGroup_lo_hi_2935 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2936;
  assign dataGroup_lo_hi_2936 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2937;
  assign dataGroup_lo_hi_2937 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2938;
  assign dataGroup_lo_hi_2938 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2939;
  assign dataGroup_lo_hi_2939 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2940;
  assign dataGroup_lo_hi_2940 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2941;
  assign dataGroup_lo_hi_2941 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2942;
  assign dataGroup_lo_hi_2942 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2943;
  assign dataGroup_lo_hi_2943 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2944;
  assign dataGroup_lo_hi_2944 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2945;
  assign dataGroup_lo_hi_2945 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2946;
  assign dataGroup_lo_hi_2946 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2947;
  assign dataGroup_lo_hi_2947 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2948;
  assign dataGroup_lo_hi_2948 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2949;
  assign dataGroup_lo_hi_2949 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2950;
  assign dataGroup_lo_hi_2950 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2951;
  assign dataGroup_lo_hi_2951 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2952;
  assign dataGroup_lo_hi_2952 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2953;
  assign dataGroup_lo_hi_2953 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2954;
  assign dataGroup_lo_hi_2954 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2955;
  assign dataGroup_lo_hi_2955 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2956;
  assign dataGroup_lo_hi_2956 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2957;
  assign dataGroup_lo_hi_2957 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2958;
  assign dataGroup_lo_hi_2958 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2959;
  assign dataGroup_lo_hi_2959 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2960;
  assign dataGroup_lo_hi_2960 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2961;
  assign dataGroup_lo_hi_2961 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2962;
  assign dataGroup_lo_hi_2962 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2963;
  assign dataGroup_lo_hi_2963 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2964;
  assign dataGroup_lo_hi_2964 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2965;
  assign dataGroup_lo_hi_2965 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2966;
  assign dataGroup_lo_hi_2966 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2967;
  assign dataGroup_lo_hi_2967 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2968;
  assign dataGroup_lo_hi_2968 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2969;
  assign dataGroup_lo_hi_2969 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2970;
  assign dataGroup_lo_hi_2970 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2971;
  assign dataGroup_lo_hi_2971 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2972;
  assign dataGroup_lo_hi_2972 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2973;
  assign dataGroup_lo_hi_2973 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2974;
  assign dataGroup_lo_hi_2974 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2975;
  assign dataGroup_lo_hi_2975 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2976;
  assign dataGroup_lo_hi_2976 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2977;
  assign dataGroup_lo_hi_2977 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2978;
  assign dataGroup_lo_hi_2978 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2979;
  assign dataGroup_lo_hi_2979 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2980;
  assign dataGroup_lo_hi_2980 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2981;
  assign dataGroup_lo_hi_2981 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2982;
  assign dataGroup_lo_hi_2982 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2983;
  assign dataGroup_lo_hi_2983 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2984;
  assign dataGroup_lo_hi_2984 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2985;
  assign dataGroup_lo_hi_2985 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2986;
  assign dataGroup_lo_hi_2986 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2987;
  assign dataGroup_lo_hi_2987 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2988;
  assign dataGroup_lo_hi_2988 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2989;
  assign dataGroup_lo_hi_2989 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2990;
  assign dataGroup_lo_hi_2990 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2991;
  assign dataGroup_lo_hi_2991 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2992;
  assign dataGroup_lo_hi_2992 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2993;
  assign dataGroup_lo_hi_2993 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2994;
  assign dataGroup_lo_hi_2994 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2995;
  assign dataGroup_lo_hi_2995 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2996;
  assign dataGroup_lo_hi_2996 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2997;
  assign dataGroup_lo_hi_2997 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2998;
  assign dataGroup_lo_hi_2998 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_2999;
  assign dataGroup_lo_hi_2999 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3000;
  assign dataGroup_lo_hi_3000 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3001;
  assign dataGroup_lo_hi_3001 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3002;
  assign dataGroup_lo_hi_3002 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3003;
  assign dataGroup_lo_hi_3003 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3004;
  assign dataGroup_lo_hi_3004 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3005;
  assign dataGroup_lo_hi_3005 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3006;
  assign dataGroup_lo_hi_3006 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3007;
  assign dataGroup_lo_hi_3007 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3008;
  assign dataGroup_lo_hi_3008 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3009;
  assign dataGroup_lo_hi_3009 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3010;
  assign dataGroup_lo_hi_3010 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3011;
  assign dataGroup_lo_hi_3011 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3012;
  assign dataGroup_lo_hi_3012 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3013;
  assign dataGroup_lo_hi_3013 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3014;
  assign dataGroup_lo_hi_3014 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3015;
  assign dataGroup_lo_hi_3015 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3016;
  assign dataGroup_lo_hi_3016 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3017;
  assign dataGroup_lo_hi_3017 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3018;
  assign dataGroup_lo_hi_3018 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3019;
  assign dataGroup_lo_hi_3019 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3020;
  assign dataGroup_lo_hi_3020 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3021;
  assign dataGroup_lo_hi_3021 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3022;
  assign dataGroup_lo_hi_3022 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3023;
  assign dataGroup_lo_hi_3023 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3024;
  assign dataGroup_lo_hi_3024 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3025;
  assign dataGroup_lo_hi_3025 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3026;
  assign dataGroup_lo_hi_3026 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3027;
  assign dataGroup_lo_hi_3027 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3028;
  assign dataGroup_lo_hi_3028 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3029;
  assign dataGroup_lo_hi_3029 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3030;
  assign dataGroup_lo_hi_3030 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3031;
  assign dataGroup_lo_hi_3031 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3032;
  assign dataGroup_lo_hi_3032 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3033;
  assign dataGroup_lo_hi_3033 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3034;
  assign dataGroup_lo_hi_3034 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3035;
  assign dataGroup_lo_hi_3035 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3036;
  assign dataGroup_lo_hi_3036 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3037;
  assign dataGroup_lo_hi_3037 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3038;
  assign dataGroup_lo_hi_3038 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3039;
  assign dataGroup_lo_hi_3039 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3040;
  assign dataGroup_lo_hi_3040 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3041;
  assign dataGroup_lo_hi_3041 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3042;
  assign dataGroup_lo_hi_3042 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3043;
  assign dataGroup_lo_hi_3043 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3044;
  assign dataGroup_lo_hi_3044 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3045;
  assign dataGroup_lo_hi_3045 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3046;
  assign dataGroup_lo_hi_3046 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3047;
  assign dataGroup_lo_hi_3047 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3048;
  assign dataGroup_lo_hi_3048 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3049;
  assign dataGroup_lo_hi_3049 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3050;
  assign dataGroup_lo_hi_3050 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3051;
  assign dataGroup_lo_hi_3051 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3052;
  assign dataGroup_lo_hi_3052 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3053;
  assign dataGroup_lo_hi_3053 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3054;
  assign dataGroup_lo_hi_3054 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3055;
  assign dataGroup_lo_hi_3055 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3056;
  assign dataGroup_lo_hi_3056 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3057;
  assign dataGroup_lo_hi_3057 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3058;
  assign dataGroup_lo_hi_3058 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3059;
  assign dataGroup_lo_hi_3059 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3060;
  assign dataGroup_lo_hi_3060 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3061;
  assign dataGroup_lo_hi_3061 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3062;
  assign dataGroup_lo_hi_3062 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3063;
  assign dataGroup_lo_hi_3063 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3064;
  assign dataGroup_lo_hi_3064 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3065;
  assign dataGroup_lo_hi_3065 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3066;
  assign dataGroup_lo_hi_3066 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3067;
  assign dataGroup_lo_hi_3067 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3068;
  assign dataGroup_lo_hi_3068 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3069;
  assign dataGroup_lo_hi_3069 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3070;
  assign dataGroup_lo_hi_3070 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3071;
  assign dataGroup_lo_hi_3071 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3072;
  assign dataGroup_lo_hi_3072 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3073;
  assign dataGroup_lo_hi_3073 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3074;
  assign dataGroup_lo_hi_3074 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3075;
  assign dataGroup_lo_hi_3075 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3076;
  assign dataGroup_lo_hi_3076 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3077;
  assign dataGroup_lo_hi_3077 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3078;
  assign dataGroup_lo_hi_3078 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3079;
  assign dataGroup_lo_hi_3079 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3080;
  assign dataGroup_lo_hi_3080 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3081;
  assign dataGroup_lo_hi_3081 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3082;
  assign dataGroup_lo_hi_3082 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3083;
  assign dataGroup_lo_hi_3083 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3084;
  assign dataGroup_lo_hi_3084 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3085;
  assign dataGroup_lo_hi_3085 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3086;
  assign dataGroup_lo_hi_3086 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3087;
  assign dataGroup_lo_hi_3087 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3088;
  assign dataGroup_lo_hi_3088 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3089;
  assign dataGroup_lo_hi_3089 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3090;
  assign dataGroup_lo_hi_3090 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3091;
  assign dataGroup_lo_hi_3091 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3092;
  assign dataGroup_lo_hi_3092 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3093;
  assign dataGroup_lo_hi_3093 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3094;
  assign dataGroup_lo_hi_3094 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3095;
  assign dataGroup_lo_hi_3095 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3096;
  assign dataGroup_lo_hi_3096 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3097;
  assign dataGroup_lo_hi_3097 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3098;
  assign dataGroup_lo_hi_3098 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3099;
  assign dataGroup_lo_hi_3099 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3100;
  assign dataGroup_lo_hi_3100 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3101;
  assign dataGroup_lo_hi_3101 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3102;
  assign dataGroup_lo_hi_3102 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3103;
  assign dataGroup_lo_hi_3103 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3104;
  assign dataGroup_lo_hi_3104 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3105;
  assign dataGroup_lo_hi_3105 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3106;
  assign dataGroup_lo_hi_3106 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3107;
  assign dataGroup_lo_hi_3107 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3108;
  assign dataGroup_lo_hi_3108 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3109;
  assign dataGroup_lo_hi_3109 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3110;
  assign dataGroup_lo_hi_3110 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3111;
  assign dataGroup_lo_hi_3111 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3112;
  assign dataGroup_lo_hi_3112 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3113;
  assign dataGroup_lo_hi_3113 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3114;
  assign dataGroup_lo_hi_3114 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3115;
  assign dataGroup_lo_hi_3115 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3116;
  assign dataGroup_lo_hi_3116 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3117;
  assign dataGroup_lo_hi_3117 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3118;
  assign dataGroup_lo_hi_3118 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3119;
  assign dataGroup_lo_hi_3119 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3120;
  assign dataGroup_lo_hi_3120 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3121;
  assign dataGroup_lo_hi_3121 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3122;
  assign dataGroup_lo_hi_3122 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3123;
  assign dataGroup_lo_hi_3123 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3124;
  assign dataGroup_lo_hi_3124 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3125;
  assign dataGroup_lo_hi_3125 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3126;
  assign dataGroup_lo_hi_3126 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3127;
  assign dataGroup_lo_hi_3127 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3128;
  assign dataGroup_lo_hi_3128 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3129;
  assign dataGroup_lo_hi_3129 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3130;
  assign dataGroup_lo_hi_3130 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3131;
  assign dataGroup_lo_hi_3131 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3132;
  assign dataGroup_lo_hi_3132 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3133;
  assign dataGroup_lo_hi_3133 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3134;
  assign dataGroup_lo_hi_3134 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3135;
  assign dataGroup_lo_hi_3135 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3136;
  assign dataGroup_lo_hi_3136 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3137;
  assign dataGroup_lo_hi_3137 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3138;
  assign dataGroup_lo_hi_3138 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3139;
  assign dataGroup_lo_hi_3139 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3140;
  assign dataGroup_lo_hi_3140 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3141;
  assign dataGroup_lo_hi_3141 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3142;
  assign dataGroup_lo_hi_3142 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3143;
  assign dataGroup_lo_hi_3143 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3144;
  assign dataGroup_lo_hi_3144 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3145;
  assign dataGroup_lo_hi_3145 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3146;
  assign dataGroup_lo_hi_3146 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3147;
  assign dataGroup_lo_hi_3147 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3148;
  assign dataGroup_lo_hi_3148 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3149;
  assign dataGroup_lo_hi_3149 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3150;
  assign dataGroup_lo_hi_3150 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3151;
  assign dataGroup_lo_hi_3151 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3152;
  assign dataGroup_lo_hi_3152 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3153;
  assign dataGroup_lo_hi_3153 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3154;
  assign dataGroup_lo_hi_3154 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3155;
  assign dataGroup_lo_hi_3155 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3156;
  assign dataGroup_lo_hi_3156 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3157;
  assign dataGroup_lo_hi_3157 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3158;
  assign dataGroup_lo_hi_3158 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3159;
  assign dataGroup_lo_hi_3159 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3160;
  assign dataGroup_lo_hi_3160 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3161;
  assign dataGroup_lo_hi_3161 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3162;
  assign dataGroup_lo_hi_3162 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3163;
  assign dataGroup_lo_hi_3163 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3164;
  assign dataGroup_lo_hi_3164 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3165;
  assign dataGroup_lo_hi_3165 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3166;
  assign dataGroup_lo_hi_3166 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3167;
  assign dataGroup_lo_hi_3167 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3168;
  assign dataGroup_lo_hi_3168 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3169;
  assign dataGroup_lo_hi_3169 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3170;
  assign dataGroup_lo_hi_3170 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3171;
  assign dataGroup_lo_hi_3171 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3172;
  assign dataGroup_lo_hi_3172 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3173;
  assign dataGroup_lo_hi_3173 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3174;
  assign dataGroup_lo_hi_3174 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3175;
  assign dataGroup_lo_hi_3175 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3176;
  assign dataGroup_lo_hi_3176 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3177;
  assign dataGroup_lo_hi_3177 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3178;
  assign dataGroup_lo_hi_3178 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3179;
  assign dataGroup_lo_hi_3179 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3180;
  assign dataGroup_lo_hi_3180 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3181;
  assign dataGroup_lo_hi_3181 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3182;
  assign dataGroup_lo_hi_3182 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3183;
  assign dataGroup_lo_hi_3183 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3184;
  assign dataGroup_lo_hi_3184 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3185;
  assign dataGroup_lo_hi_3185 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3186;
  assign dataGroup_lo_hi_3186 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3187;
  assign dataGroup_lo_hi_3187 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3188;
  assign dataGroup_lo_hi_3188 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3189;
  assign dataGroup_lo_hi_3189 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3190;
  assign dataGroup_lo_hi_3190 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3191;
  assign dataGroup_lo_hi_3191 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3192;
  assign dataGroup_lo_hi_3192 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3193;
  assign dataGroup_lo_hi_3193 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3194;
  assign dataGroup_lo_hi_3194 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3195;
  assign dataGroup_lo_hi_3195 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3196;
  assign dataGroup_lo_hi_3196 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3197;
  assign dataGroup_lo_hi_3197 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3198;
  assign dataGroup_lo_hi_3198 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3199;
  assign dataGroup_lo_hi_3199 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3200;
  assign dataGroup_lo_hi_3200 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3201;
  assign dataGroup_lo_hi_3201 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3202;
  assign dataGroup_lo_hi_3202 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3203;
  assign dataGroup_lo_hi_3203 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3204;
  assign dataGroup_lo_hi_3204 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3205;
  assign dataGroup_lo_hi_3205 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3206;
  assign dataGroup_lo_hi_3206 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3207;
  assign dataGroup_lo_hi_3207 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3208;
  assign dataGroup_lo_hi_3208 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3209;
  assign dataGroup_lo_hi_3209 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3210;
  assign dataGroup_lo_hi_3210 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3211;
  assign dataGroup_lo_hi_3211 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3212;
  assign dataGroup_lo_hi_3212 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3213;
  assign dataGroup_lo_hi_3213 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3214;
  assign dataGroup_lo_hi_3214 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3215;
  assign dataGroup_lo_hi_3215 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3216;
  assign dataGroup_lo_hi_3216 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3217;
  assign dataGroup_lo_hi_3217 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3218;
  assign dataGroup_lo_hi_3218 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3219;
  assign dataGroup_lo_hi_3219 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3220;
  assign dataGroup_lo_hi_3220 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3221;
  assign dataGroup_lo_hi_3221 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3222;
  assign dataGroup_lo_hi_3222 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3223;
  assign dataGroup_lo_hi_3223 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3224;
  assign dataGroup_lo_hi_3224 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3225;
  assign dataGroup_lo_hi_3225 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3226;
  assign dataGroup_lo_hi_3226 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3227;
  assign dataGroup_lo_hi_3227 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3228;
  assign dataGroup_lo_hi_3228 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3229;
  assign dataGroup_lo_hi_3229 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3230;
  assign dataGroup_lo_hi_3230 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3231;
  assign dataGroup_lo_hi_3231 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3232;
  assign dataGroup_lo_hi_3232 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3233;
  assign dataGroup_lo_hi_3233 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3234;
  assign dataGroup_lo_hi_3234 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3235;
  assign dataGroup_lo_hi_3235 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3236;
  assign dataGroup_lo_hi_3236 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3237;
  assign dataGroup_lo_hi_3237 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3238;
  assign dataGroup_lo_hi_3238 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3239;
  assign dataGroup_lo_hi_3239 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3240;
  assign dataGroup_lo_hi_3240 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3241;
  assign dataGroup_lo_hi_3241 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3242;
  assign dataGroup_lo_hi_3242 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3243;
  assign dataGroup_lo_hi_3243 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3244;
  assign dataGroup_lo_hi_3244 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3245;
  assign dataGroup_lo_hi_3245 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3246;
  assign dataGroup_lo_hi_3246 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3247;
  assign dataGroup_lo_hi_3247 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3248;
  assign dataGroup_lo_hi_3248 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3249;
  assign dataGroup_lo_hi_3249 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3250;
  assign dataGroup_lo_hi_3250 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3251;
  assign dataGroup_lo_hi_3251 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3252;
  assign dataGroup_lo_hi_3252 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3253;
  assign dataGroup_lo_hi_3253 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3254;
  assign dataGroup_lo_hi_3254 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3255;
  assign dataGroup_lo_hi_3255 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3256;
  assign dataGroup_lo_hi_3256 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3257;
  assign dataGroup_lo_hi_3257 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3258;
  assign dataGroup_lo_hi_3258 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3259;
  assign dataGroup_lo_hi_3259 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3260;
  assign dataGroup_lo_hi_3260 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3261;
  assign dataGroup_lo_hi_3261 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3262;
  assign dataGroup_lo_hi_3262 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3263;
  assign dataGroup_lo_hi_3263 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3264;
  assign dataGroup_lo_hi_3264 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3265;
  assign dataGroup_lo_hi_3265 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3266;
  assign dataGroup_lo_hi_3266 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3267;
  assign dataGroup_lo_hi_3267 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3268;
  assign dataGroup_lo_hi_3268 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3269;
  assign dataGroup_lo_hi_3269 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3270;
  assign dataGroup_lo_hi_3270 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3271;
  assign dataGroup_lo_hi_3271 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3272;
  assign dataGroup_lo_hi_3272 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3273;
  assign dataGroup_lo_hi_3273 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3274;
  assign dataGroup_lo_hi_3274 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3275;
  assign dataGroup_lo_hi_3275 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3276;
  assign dataGroup_lo_hi_3276 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3277;
  assign dataGroup_lo_hi_3277 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3278;
  assign dataGroup_lo_hi_3278 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3279;
  assign dataGroup_lo_hi_3279 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3280;
  assign dataGroup_lo_hi_3280 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3281;
  assign dataGroup_lo_hi_3281 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3282;
  assign dataGroup_lo_hi_3282 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3283;
  assign dataGroup_lo_hi_3283 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3284;
  assign dataGroup_lo_hi_3284 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3285;
  assign dataGroup_lo_hi_3285 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3286;
  assign dataGroup_lo_hi_3286 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3287;
  assign dataGroup_lo_hi_3287 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3288;
  assign dataGroup_lo_hi_3288 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3289;
  assign dataGroup_lo_hi_3289 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3290;
  assign dataGroup_lo_hi_3290 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3291;
  assign dataGroup_lo_hi_3291 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3292;
  assign dataGroup_lo_hi_3292 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3293;
  assign dataGroup_lo_hi_3293 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3294;
  assign dataGroup_lo_hi_3294 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3295;
  assign dataGroup_lo_hi_3295 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3296;
  assign dataGroup_lo_hi_3296 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3297;
  assign dataGroup_lo_hi_3297 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3298;
  assign dataGroup_lo_hi_3298 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3299;
  assign dataGroup_lo_hi_3299 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3300;
  assign dataGroup_lo_hi_3300 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3301;
  assign dataGroup_lo_hi_3301 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3302;
  assign dataGroup_lo_hi_3302 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3303;
  assign dataGroup_lo_hi_3303 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3304;
  assign dataGroup_lo_hi_3304 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3305;
  assign dataGroup_lo_hi_3305 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3306;
  assign dataGroup_lo_hi_3306 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3307;
  assign dataGroup_lo_hi_3307 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3308;
  assign dataGroup_lo_hi_3308 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3309;
  assign dataGroup_lo_hi_3309 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3310;
  assign dataGroup_lo_hi_3310 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3311;
  assign dataGroup_lo_hi_3311 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3312;
  assign dataGroup_lo_hi_3312 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3313;
  assign dataGroup_lo_hi_3313 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3314;
  assign dataGroup_lo_hi_3314 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3315;
  assign dataGroup_lo_hi_3315 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3316;
  assign dataGroup_lo_hi_3316 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3317;
  assign dataGroup_lo_hi_3317 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3318;
  assign dataGroup_lo_hi_3318 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3319;
  assign dataGroup_lo_hi_3319 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3320;
  assign dataGroup_lo_hi_3320 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3321;
  assign dataGroup_lo_hi_3321 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3322;
  assign dataGroup_lo_hi_3322 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3323;
  assign dataGroup_lo_hi_3323 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3324;
  assign dataGroup_lo_hi_3324 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3325;
  assign dataGroup_lo_hi_3325 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3326;
  assign dataGroup_lo_hi_3326 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3327;
  assign dataGroup_lo_hi_3327 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3328;
  assign dataGroup_lo_hi_3328 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3329;
  assign dataGroup_lo_hi_3329 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3330;
  assign dataGroup_lo_hi_3330 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3331;
  assign dataGroup_lo_hi_3331 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3332;
  assign dataGroup_lo_hi_3332 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3333;
  assign dataGroup_lo_hi_3333 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3334;
  assign dataGroup_lo_hi_3334 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3335;
  assign dataGroup_lo_hi_3335 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3336;
  assign dataGroup_lo_hi_3336 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3337;
  assign dataGroup_lo_hi_3337 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3338;
  assign dataGroup_lo_hi_3338 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3339;
  assign dataGroup_lo_hi_3339 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3340;
  assign dataGroup_lo_hi_3340 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3341;
  assign dataGroup_lo_hi_3341 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3342;
  assign dataGroup_lo_hi_3342 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3343;
  assign dataGroup_lo_hi_3343 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3344;
  assign dataGroup_lo_hi_3344 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3345;
  assign dataGroup_lo_hi_3345 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3346;
  assign dataGroup_lo_hi_3346 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3347;
  assign dataGroup_lo_hi_3347 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3348;
  assign dataGroup_lo_hi_3348 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3349;
  assign dataGroup_lo_hi_3349 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3350;
  assign dataGroup_lo_hi_3350 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3351;
  assign dataGroup_lo_hi_3351 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3352;
  assign dataGroup_lo_hi_3352 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3353;
  assign dataGroup_lo_hi_3353 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3354;
  assign dataGroup_lo_hi_3354 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3355;
  assign dataGroup_lo_hi_3355 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3356;
  assign dataGroup_lo_hi_3356 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3357;
  assign dataGroup_lo_hi_3357 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3358;
  assign dataGroup_lo_hi_3358 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3359;
  assign dataGroup_lo_hi_3359 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3360;
  assign dataGroup_lo_hi_3360 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3361;
  assign dataGroup_lo_hi_3361 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3362;
  assign dataGroup_lo_hi_3362 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3363;
  assign dataGroup_lo_hi_3363 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3364;
  assign dataGroup_lo_hi_3364 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3365;
  assign dataGroup_lo_hi_3365 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3366;
  assign dataGroup_lo_hi_3366 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3367;
  assign dataGroup_lo_hi_3367 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3368;
  assign dataGroup_lo_hi_3368 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3369;
  assign dataGroup_lo_hi_3369 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3370;
  assign dataGroup_lo_hi_3370 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3371;
  assign dataGroup_lo_hi_3371 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3372;
  assign dataGroup_lo_hi_3372 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3373;
  assign dataGroup_lo_hi_3373 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3374;
  assign dataGroup_lo_hi_3374 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3375;
  assign dataGroup_lo_hi_3375 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3376;
  assign dataGroup_lo_hi_3376 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3377;
  assign dataGroup_lo_hi_3377 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3378;
  assign dataGroup_lo_hi_3378 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3379;
  assign dataGroup_lo_hi_3379 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3380;
  assign dataGroup_lo_hi_3380 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3381;
  assign dataGroup_lo_hi_3381 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3382;
  assign dataGroup_lo_hi_3382 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3383;
  assign dataGroup_lo_hi_3383 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3384;
  assign dataGroup_lo_hi_3384 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3385;
  assign dataGroup_lo_hi_3385 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3386;
  assign dataGroup_lo_hi_3386 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3387;
  assign dataGroup_lo_hi_3387 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3388;
  assign dataGroup_lo_hi_3388 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3389;
  assign dataGroup_lo_hi_3389 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3390;
  assign dataGroup_lo_hi_3390 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3391;
  assign dataGroup_lo_hi_3391 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3392;
  assign dataGroup_lo_hi_3392 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3393;
  assign dataGroup_lo_hi_3393 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3394;
  assign dataGroup_lo_hi_3394 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3395;
  assign dataGroup_lo_hi_3395 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3396;
  assign dataGroup_lo_hi_3396 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3397;
  assign dataGroup_lo_hi_3397 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3398;
  assign dataGroup_lo_hi_3398 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3399;
  assign dataGroup_lo_hi_3399 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3400;
  assign dataGroup_lo_hi_3400 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3401;
  assign dataGroup_lo_hi_3401 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3402;
  assign dataGroup_lo_hi_3402 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3403;
  assign dataGroup_lo_hi_3403 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3404;
  assign dataGroup_lo_hi_3404 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3405;
  assign dataGroup_lo_hi_3405 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3406;
  assign dataGroup_lo_hi_3406 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3407;
  assign dataGroup_lo_hi_3407 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3408;
  assign dataGroup_lo_hi_3408 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3409;
  assign dataGroup_lo_hi_3409 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3410;
  assign dataGroup_lo_hi_3410 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3411;
  assign dataGroup_lo_hi_3411 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3412;
  assign dataGroup_lo_hi_3412 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3413;
  assign dataGroup_lo_hi_3413 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3414;
  assign dataGroup_lo_hi_3414 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3415;
  assign dataGroup_lo_hi_3415 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3416;
  assign dataGroup_lo_hi_3416 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3417;
  assign dataGroup_lo_hi_3417 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3418;
  assign dataGroup_lo_hi_3418 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3419;
  assign dataGroup_lo_hi_3419 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3420;
  assign dataGroup_lo_hi_3420 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3421;
  assign dataGroup_lo_hi_3421 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3422;
  assign dataGroup_lo_hi_3422 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3423;
  assign dataGroup_lo_hi_3423 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3424;
  assign dataGroup_lo_hi_3424 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3425;
  assign dataGroup_lo_hi_3425 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3426;
  assign dataGroup_lo_hi_3426 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3427;
  assign dataGroup_lo_hi_3427 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3428;
  assign dataGroup_lo_hi_3428 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3429;
  assign dataGroup_lo_hi_3429 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3430;
  assign dataGroup_lo_hi_3430 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3431;
  assign dataGroup_lo_hi_3431 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3432;
  assign dataGroup_lo_hi_3432 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3433;
  assign dataGroup_lo_hi_3433 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3434;
  assign dataGroup_lo_hi_3434 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3435;
  assign dataGroup_lo_hi_3435 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3436;
  assign dataGroup_lo_hi_3436 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3437;
  assign dataGroup_lo_hi_3437 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3438;
  assign dataGroup_lo_hi_3438 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3439;
  assign dataGroup_lo_hi_3439 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3440;
  assign dataGroup_lo_hi_3440 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3441;
  assign dataGroup_lo_hi_3441 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3442;
  assign dataGroup_lo_hi_3442 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3443;
  assign dataGroup_lo_hi_3443 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3444;
  assign dataGroup_lo_hi_3444 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3445;
  assign dataGroup_lo_hi_3445 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3446;
  assign dataGroup_lo_hi_3446 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3447;
  assign dataGroup_lo_hi_3447 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3448;
  assign dataGroup_lo_hi_3448 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3449;
  assign dataGroup_lo_hi_3449 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3450;
  assign dataGroup_lo_hi_3450 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3451;
  assign dataGroup_lo_hi_3451 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3452;
  assign dataGroup_lo_hi_3452 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3453;
  assign dataGroup_lo_hi_3453 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3454;
  assign dataGroup_lo_hi_3454 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3455;
  assign dataGroup_lo_hi_3455 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3456;
  assign dataGroup_lo_hi_3456 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3457;
  assign dataGroup_lo_hi_3457 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3458;
  assign dataGroup_lo_hi_3458 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3459;
  assign dataGroup_lo_hi_3459 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3460;
  assign dataGroup_lo_hi_3460 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3461;
  assign dataGroup_lo_hi_3461 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3462;
  assign dataGroup_lo_hi_3462 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3463;
  assign dataGroup_lo_hi_3463 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3464;
  assign dataGroup_lo_hi_3464 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3465;
  assign dataGroup_lo_hi_3465 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3466;
  assign dataGroup_lo_hi_3466 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3467;
  assign dataGroup_lo_hi_3467 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3468;
  assign dataGroup_lo_hi_3468 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3469;
  assign dataGroup_lo_hi_3469 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3470;
  assign dataGroup_lo_hi_3470 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3471;
  assign dataGroup_lo_hi_3471 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3472;
  assign dataGroup_lo_hi_3472 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3473;
  assign dataGroup_lo_hi_3473 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3474;
  assign dataGroup_lo_hi_3474 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3475;
  assign dataGroup_lo_hi_3475 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3476;
  assign dataGroup_lo_hi_3476 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3477;
  assign dataGroup_lo_hi_3477 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3478;
  assign dataGroup_lo_hi_3478 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3479;
  assign dataGroup_lo_hi_3479 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3480;
  assign dataGroup_lo_hi_3480 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3481;
  assign dataGroup_lo_hi_3481 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3482;
  assign dataGroup_lo_hi_3482 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3483;
  assign dataGroup_lo_hi_3483 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3484;
  assign dataGroup_lo_hi_3484 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3485;
  assign dataGroup_lo_hi_3485 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3486;
  assign dataGroup_lo_hi_3486 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3487;
  assign dataGroup_lo_hi_3487 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3488;
  assign dataGroup_lo_hi_3488 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3489;
  assign dataGroup_lo_hi_3489 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3490;
  assign dataGroup_lo_hi_3490 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3491;
  assign dataGroup_lo_hi_3491 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3492;
  assign dataGroup_lo_hi_3492 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3493;
  assign dataGroup_lo_hi_3493 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3494;
  assign dataGroup_lo_hi_3494 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3495;
  assign dataGroup_lo_hi_3495 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3496;
  assign dataGroup_lo_hi_3496 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3497;
  assign dataGroup_lo_hi_3497 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3498;
  assign dataGroup_lo_hi_3498 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3499;
  assign dataGroup_lo_hi_3499 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3500;
  assign dataGroup_lo_hi_3500 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3501;
  assign dataGroup_lo_hi_3501 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3502;
  assign dataGroup_lo_hi_3502 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3503;
  assign dataGroup_lo_hi_3503 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3504;
  assign dataGroup_lo_hi_3504 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3505;
  assign dataGroup_lo_hi_3505 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3506;
  assign dataGroup_lo_hi_3506 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3507;
  assign dataGroup_lo_hi_3507 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3508;
  assign dataGroup_lo_hi_3508 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3509;
  assign dataGroup_lo_hi_3509 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3510;
  assign dataGroup_lo_hi_3510 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3511;
  assign dataGroup_lo_hi_3511 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3512;
  assign dataGroup_lo_hi_3512 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3513;
  assign dataGroup_lo_hi_3513 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3514;
  assign dataGroup_lo_hi_3514 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3515;
  assign dataGroup_lo_hi_3515 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3516;
  assign dataGroup_lo_hi_3516 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3517;
  assign dataGroup_lo_hi_3517 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3518;
  assign dataGroup_lo_hi_3518 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3519;
  assign dataGroup_lo_hi_3519 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3520;
  assign dataGroup_lo_hi_3520 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3521;
  assign dataGroup_lo_hi_3521 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3522;
  assign dataGroup_lo_hi_3522 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3523;
  assign dataGroup_lo_hi_3523 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3524;
  assign dataGroup_lo_hi_3524 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3525;
  assign dataGroup_lo_hi_3525 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3526;
  assign dataGroup_lo_hi_3526 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3527;
  assign dataGroup_lo_hi_3527 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3528;
  assign dataGroup_lo_hi_3528 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3529;
  assign dataGroup_lo_hi_3529 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3530;
  assign dataGroup_lo_hi_3530 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3531;
  assign dataGroup_lo_hi_3531 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3532;
  assign dataGroup_lo_hi_3532 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3533;
  assign dataGroup_lo_hi_3533 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3534;
  assign dataGroup_lo_hi_3534 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3535;
  assign dataGroup_lo_hi_3535 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3536;
  assign dataGroup_lo_hi_3536 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3537;
  assign dataGroup_lo_hi_3537 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3538;
  assign dataGroup_lo_hi_3538 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3539;
  assign dataGroup_lo_hi_3539 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3540;
  assign dataGroup_lo_hi_3540 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3541;
  assign dataGroup_lo_hi_3541 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3542;
  assign dataGroup_lo_hi_3542 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3543;
  assign dataGroup_lo_hi_3543 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3544;
  assign dataGroup_lo_hi_3544 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3545;
  assign dataGroup_lo_hi_3545 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3546;
  assign dataGroup_lo_hi_3546 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3547;
  assign dataGroup_lo_hi_3547 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3548;
  assign dataGroup_lo_hi_3548 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3549;
  assign dataGroup_lo_hi_3549 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3550;
  assign dataGroup_lo_hi_3550 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3551;
  assign dataGroup_lo_hi_3551 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3552;
  assign dataGroup_lo_hi_3552 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3553;
  assign dataGroup_lo_hi_3553 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3554;
  assign dataGroup_lo_hi_3554 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3555;
  assign dataGroup_lo_hi_3555 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3556;
  assign dataGroup_lo_hi_3556 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3557;
  assign dataGroup_lo_hi_3557 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3558;
  assign dataGroup_lo_hi_3558 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3559;
  assign dataGroup_lo_hi_3559 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3560;
  assign dataGroup_lo_hi_3560 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3561;
  assign dataGroup_lo_hi_3561 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3562;
  assign dataGroup_lo_hi_3562 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3563;
  assign dataGroup_lo_hi_3563 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3564;
  assign dataGroup_lo_hi_3564 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3565;
  assign dataGroup_lo_hi_3565 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3566;
  assign dataGroup_lo_hi_3566 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3567;
  assign dataGroup_lo_hi_3567 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3568;
  assign dataGroup_lo_hi_3568 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3569;
  assign dataGroup_lo_hi_3569 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3570;
  assign dataGroup_lo_hi_3570 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3571;
  assign dataGroup_lo_hi_3571 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3572;
  assign dataGroup_lo_hi_3572 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3573;
  assign dataGroup_lo_hi_3573 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3574;
  assign dataGroup_lo_hi_3574 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3575;
  assign dataGroup_lo_hi_3575 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3576;
  assign dataGroup_lo_hi_3576 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3577;
  assign dataGroup_lo_hi_3577 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3578;
  assign dataGroup_lo_hi_3578 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3579;
  assign dataGroup_lo_hi_3579 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3580;
  assign dataGroup_lo_hi_3580 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3581;
  assign dataGroup_lo_hi_3581 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3582;
  assign dataGroup_lo_hi_3582 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3583;
  assign dataGroup_lo_hi_3583 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3584;
  assign dataGroup_lo_hi_3584 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3585;
  assign dataGroup_lo_hi_3585 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3586;
  assign dataGroup_lo_hi_3586 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3587;
  assign dataGroup_lo_hi_3587 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3588;
  assign dataGroup_lo_hi_3588 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3589;
  assign dataGroup_lo_hi_3589 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3590;
  assign dataGroup_lo_hi_3590 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3591;
  assign dataGroup_lo_hi_3591 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3592;
  assign dataGroup_lo_hi_3592 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3593;
  assign dataGroup_lo_hi_3593 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3594;
  assign dataGroup_lo_hi_3594 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3595;
  assign dataGroup_lo_hi_3595 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3596;
  assign dataGroup_lo_hi_3596 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3597;
  assign dataGroup_lo_hi_3597 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3598;
  assign dataGroup_lo_hi_3598 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3599;
  assign dataGroup_lo_hi_3599 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3600;
  assign dataGroup_lo_hi_3600 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3601;
  assign dataGroup_lo_hi_3601 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3602;
  assign dataGroup_lo_hi_3602 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3603;
  assign dataGroup_lo_hi_3603 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3604;
  assign dataGroup_lo_hi_3604 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3605;
  assign dataGroup_lo_hi_3605 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3606;
  assign dataGroup_lo_hi_3606 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3607;
  assign dataGroup_lo_hi_3607 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3608;
  assign dataGroup_lo_hi_3608 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3609;
  assign dataGroup_lo_hi_3609 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3610;
  assign dataGroup_lo_hi_3610 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3611;
  assign dataGroup_lo_hi_3611 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3612;
  assign dataGroup_lo_hi_3612 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3613;
  assign dataGroup_lo_hi_3613 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3614;
  assign dataGroup_lo_hi_3614 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3615;
  assign dataGroup_lo_hi_3615 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3616;
  assign dataGroup_lo_hi_3616 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3617;
  assign dataGroup_lo_hi_3617 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3618;
  assign dataGroup_lo_hi_3618 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3619;
  assign dataGroup_lo_hi_3619 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3620;
  assign dataGroup_lo_hi_3620 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3621;
  assign dataGroup_lo_hi_3621 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3622;
  assign dataGroup_lo_hi_3622 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3623;
  assign dataGroup_lo_hi_3623 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3624;
  assign dataGroup_lo_hi_3624 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3625;
  assign dataGroup_lo_hi_3625 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3626;
  assign dataGroup_lo_hi_3626 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3627;
  assign dataGroup_lo_hi_3627 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3628;
  assign dataGroup_lo_hi_3628 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3629;
  assign dataGroup_lo_hi_3629 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3630;
  assign dataGroup_lo_hi_3630 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3631;
  assign dataGroup_lo_hi_3631 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3632;
  assign dataGroup_lo_hi_3632 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3633;
  assign dataGroup_lo_hi_3633 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3634;
  assign dataGroup_lo_hi_3634 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3635;
  assign dataGroup_lo_hi_3635 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3636;
  assign dataGroup_lo_hi_3636 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3637;
  assign dataGroup_lo_hi_3637 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3638;
  assign dataGroup_lo_hi_3638 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3639;
  assign dataGroup_lo_hi_3639 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3640;
  assign dataGroup_lo_hi_3640 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3641;
  assign dataGroup_lo_hi_3641 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3642;
  assign dataGroup_lo_hi_3642 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3643;
  assign dataGroup_lo_hi_3643 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3644;
  assign dataGroup_lo_hi_3644 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3645;
  assign dataGroup_lo_hi_3645 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3646;
  assign dataGroup_lo_hi_3646 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3647;
  assign dataGroup_lo_hi_3647 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3648;
  assign dataGroup_lo_hi_3648 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3649;
  assign dataGroup_lo_hi_3649 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3650;
  assign dataGroup_lo_hi_3650 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3651;
  assign dataGroup_lo_hi_3651 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3652;
  assign dataGroup_lo_hi_3652 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3653;
  assign dataGroup_lo_hi_3653 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3654;
  assign dataGroup_lo_hi_3654 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3655;
  assign dataGroup_lo_hi_3655 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3656;
  assign dataGroup_lo_hi_3656 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3657;
  assign dataGroup_lo_hi_3657 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3658;
  assign dataGroup_lo_hi_3658 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3659;
  assign dataGroup_lo_hi_3659 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3660;
  assign dataGroup_lo_hi_3660 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3661;
  assign dataGroup_lo_hi_3661 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3662;
  assign dataGroup_lo_hi_3662 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3663;
  assign dataGroup_lo_hi_3663 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3664;
  assign dataGroup_lo_hi_3664 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3665;
  assign dataGroup_lo_hi_3665 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3666;
  assign dataGroup_lo_hi_3666 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3667;
  assign dataGroup_lo_hi_3667 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3668;
  assign dataGroup_lo_hi_3668 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3669;
  assign dataGroup_lo_hi_3669 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3670;
  assign dataGroup_lo_hi_3670 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3671;
  assign dataGroup_lo_hi_3671 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3672;
  assign dataGroup_lo_hi_3672 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3673;
  assign dataGroup_lo_hi_3673 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3674;
  assign dataGroup_lo_hi_3674 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3675;
  assign dataGroup_lo_hi_3675 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3676;
  assign dataGroup_lo_hi_3676 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3677;
  assign dataGroup_lo_hi_3677 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3678;
  assign dataGroup_lo_hi_3678 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3679;
  assign dataGroup_lo_hi_3679 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3680;
  assign dataGroup_lo_hi_3680 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3681;
  assign dataGroup_lo_hi_3681 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3682;
  assign dataGroup_lo_hi_3682 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3683;
  assign dataGroup_lo_hi_3683 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3684;
  assign dataGroup_lo_hi_3684 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3685;
  assign dataGroup_lo_hi_3685 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3686;
  assign dataGroup_lo_hi_3686 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3687;
  assign dataGroup_lo_hi_3687 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3688;
  assign dataGroup_lo_hi_3688 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3689;
  assign dataGroup_lo_hi_3689 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3690;
  assign dataGroup_lo_hi_3690 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3691;
  assign dataGroup_lo_hi_3691 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3692;
  assign dataGroup_lo_hi_3692 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3693;
  assign dataGroup_lo_hi_3693 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3694;
  assign dataGroup_lo_hi_3694 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3695;
  assign dataGroup_lo_hi_3695 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3696;
  assign dataGroup_lo_hi_3696 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3697;
  assign dataGroup_lo_hi_3697 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3698;
  assign dataGroup_lo_hi_3698 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3699;
  assign dataGroup_lo_hi_3699 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3700;
  assign dataGroup_lo_hi_3700 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3701;
  assign dataGroup_lo_hi_3701 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3702;
  assign dataGroup_lo_hi_3702 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3703;
  assign dataGroup_lo_hi_3703 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3704;
  assign dataGroup_lo_hi_3704 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3705;
  assign dataGroup_lo_hi_3705 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3706;
  assign dataGroup_lo_hi_3706 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3707;
  assign dataGroup_lo_hi_3707 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3708;
  assign dataGroup_lo_hi_3708 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3709;
  assign dataGroup_lo_hi_3709 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3710;
  assign dataGroup_lo_hi_3710 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3711;
  assign dataGroup_lo_hi_3711 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3712;
  assign dataGroup_lo_hi_3712 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3713;
  assign dataGroup_lo_hi_3713 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3714;
  assign dataGroup_lo_hi_3714 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3715;
  assign dataGroup_lo_hi_3715 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3716;
  assign dataGroup_lo_hi_3716 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3717;
  assign dataGroup_lo_hi_3717 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3718;
  assign dataGroup_lo_hi_3718 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3719;
  assign dataGroup_lo_hi_3719 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3720;
  assign dataGroup_lo_hi_3720 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3721;
  assign dataGroup_lo_hi_3721 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3722;
  assign dataGroup_lo_hi_3722 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3723;
  assign dataGroup_lo_hi_3723 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3724;
  assign dataGroup_lo_hi_3724 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3725;
  assign dataGroup_lo_hi_3725 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3726;
  assign dataGroup_lo_hi_3726 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3727;
  assign dataGroup_lo_hi_3727 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3728;
  assign dataGroup_lo_hi_3728 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3729;
  assign dataGroup_lo_hi_3729 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3730;
  assign dataGroup_lo_hi_3730 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3731;
  assign dataGroup_lo_hi_3731 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3732;
  assign dataGroup_lo_hi_3732 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3733;
  assign dataGroup_lo_hi_3733 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3734;
  assign dataGroup_lo_hi_3734 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3735;
  assign dataGroup_lo_hi_3735 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3736;
  assign dataGroup_lo_hi_3736 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3737;
  assign dataGroup_lo_hi_3737 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3738;
  assign dataGroup_lo_hi_3738 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3739;
  assign dataGroup_lo_hi_3739 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3740;
  assign dataGroup_lo_hi_3740 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3741;
  assign dataGroup_lo_hi_3741 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3742;
  assign dataGroup_lo_hi_3742 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3743;
  assign dataGroup_lo_hi_3743 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3744;
  assign dataGroup_lo_hi_3744 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3745;
  assign dataGroup_lo_hi_3745 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3746;
  assign dataGroup_lo_hi_3746 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3747;
  assign dataGroup_lo_hi_3747 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3748;
  assign dataGroup_lo_hi_3748 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3749;
  assign dataGroup_lo_hi_3749 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3750;
  assign dataGroup_lo_hi_3750 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3751;
  assign dataGroup_lo_hi_3751 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3752;
  assign dataGroup_lo_hi_3752 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3753;
  assign dataGroup_lo_hi_3753 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3754;
  assign dataGroup_lo_hi_3754 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3755;
  assign dataGroup_lo_hi_3755 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3756;
  assign dataGroup_lo_hi_3756 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3757;
  assign dataGroup_lo_hi_3757 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3758;
  assign dataGroup_lo_hi_3758 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3759;
  assign dataGroup_lo_hi_3759 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3760;
  assign dataGroup_lo_hi_3760 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3761;
  assign dataGroup_lo_hi_3761 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3762;
  assign dataGroup_lo_hi_3762 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3763;
  assign dataGroup_lo_hi_3763 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3764;
  assign dataGroup_lo_hi_3764 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3765;
  assign dataGroup_lo_hi_3765 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3766;
  assign dataGroup_lo_hi_3766 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3767;
  assign dataGroup_lo_hi_3767 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3768;
  assign dataGroup_lo_hi_3768 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3769;
  assign dataGroup_lo_hi_3769 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3770;
  assign dataGroup_lo_hi_3770 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3771;
  assign dataGroup_lo_hi_3771 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3772;
  assign dataGroup_lo_hi_3772 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3773;
  assign dataGroup_lo_hi_3773 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3774;
  assign dataGroup_lo_hi_3774 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3775;
  assign dataGroup_lo_hi_3775 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3776;
  assign dataGroup_lo_hi_3776 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3777;
  assign dataGroup_lo_hi_3777 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3778;
  assign dataGroup_lo_hi_3778 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3779;
  assign dataGroup_lo_hi_3779 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3780;
  assign dataGroup_lo_hi_3780 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3781;
  assign dataGroup_lo_hi_3781 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3782;
  assign dataGroup_lo_hi_3782 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3783;
  assign dataGroup_lo_hi_3783 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3784;
  assign dataGroup_lo_hi_3784 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3785;
  assign dataGroup_lo_hi_3785 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3786;
  assign dataGroup_lo_hi_3786 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3787;
  assign dataGroup_lo_hi_3787 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3788;
  assign dataGroup_lo_hi_3788 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3789;
  assign dataGroup_lo_hi_3789 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3790;
  assign dataGroup_lo_hi_3790 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3791;
  assign dataGroup_lo_hi_3791 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3792;
  assign dataGroup_lo_hi_3792 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3793;
  assign dataGroup_lo_hi_3793 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3794;
  assign dataGroup_lo_hi_3794 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3795;
  assign dataGroup_lo_hi_3795 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3796;
  assign dataGroup_lo_hi_3796 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3797;
  assign dataGroup_lo_hi_3797 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3798;
  assign dataGroup_lo_hi_3798 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3799;
  assign dataGroup_lo_hi_3799 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3800;
  assign dataGroup_lo_hi_3800 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3801;
  assign dataGroup_lo_hi_3801 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3802;
  assign dataGroup_lo_hi_3802 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3803;
  assign dataGroup_lo_hi_3803 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3804;
  assign dataGroup_lo_hi_3804 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3805;
  assign dataGroup_lo_hi_3805 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3806;
  assign dataGroup_lo_hi_3806 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3807;
  assign dataGroup_lo_hi_3807 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3808;
  assign dataGroup_lo_hi_3808 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3809;
  assign dataGroup_lo_hi_3809 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3810;
  assign dataGroup_lo_hi_3810 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3811;
  assign dataGroup_lo_hi_3811 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3812;
  assign dataGroup_lo_hi_3812 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3813;
  assign dataGroup_lo_hi_3813 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3814;
  assign dataGroup_lo_hi_3814 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3815;
  assign dataGroup_lo_hi_3815 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3816;
  assign dataGroup_lo_hi_3816 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3817;
  assign dataGroup_lo_hi_3817 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3818;
  assign dataGroup_lo_hi_3818 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3819;
  assign dataGroup_lo_hi_3819 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3820;
  assign dataGroup_lo_hi_3820 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3821;
  assign dataGroup_lo_hi_3821 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3822;
  assign dataGroup_lo_hi_3822 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3823;
  assign dataGroup_lo_hi_3823 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3824;
  assign dataGroup_lo_hi_3824 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3825;
  assign dataGroup_lo_hi_3825 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3826;
  assign dataGroup_lo_hi_3826 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3827;
  assign dataGroup_lo_hi_3827 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3828;
  assign dataGroup_lo_hi_3828 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3829;
  assign dataGroup_lo_hi_3829 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3830;
  assign dataGroup_lo_hi_3830 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3831;
  assign dataGroup_lo_hi_3831 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3832;
  assign dataGroup_lo_hi_3832 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3833;
  assign dataGroup_lo_hi_3833 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3834;
  assign dataGroup_lo_hi_3834 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3835;
  assign dataGroup_lo_hi_3835 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3836;
  assign dataGroup_lo_hi_3836 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3837;
  assign dataGroup_lo_hi_3837 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3838;
  assign dataGroup_lo_hi_3838 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3839;
  assign dataGroup_lo_hi_3839 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3840;
  assign dataGroup_lo_hi_3840 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3841;
  assign dataGroup_lo_hi_3841 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3842;
  assign dataGroup_lo_hi_3842 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3843;
  assign dataGroup_lo_hi_3843 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3844;
  assign dataGroup_lo_hi_3844 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3845;
  assign dataGroup_lo_hi_3845 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3846;
  assign dataGroup_lo_hi_3846 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3847;
  assign dataGroup_lo_hi_3847 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3848;
  assign dataGroup_lo_hi_3848 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3849;
  assign dataGroup_lo_hi_3849 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3850;
  assign dataGroup_lo_hi_3850 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3851;
  assign dataGroup_lo_hi_3851 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3852;
  assign dataGroup_lo_hi_3852 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3853;
  assign dataGroup_lo_hi_3853 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3854;
  assign dataGroup_lo_hi_3854 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3855;
  assign dataGroup_lo_hi_3855 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3856;
  assign dataGroup_lo_hi_3856 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3857;
  assign dataGroup_lo_hi_3857 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3858;
  assign dataGroup_lo_hi_3858 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3859;
  assign dataGroup_lo_hi_3859 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3860;
  assign dataGroup_lo_hi_3860 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3861;
  assign dataGroup_lo_hi_3861 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3862;
  assign dataGroup_lo_hi_3862 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3863;
  assign dataGroup_lo_hi_3863 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3864;
  assign dataGroup_lo_hi_3864 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3865;
  assign dataGroup_lo_hi_3865 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3866;
  assign dataGroup_lo_hi_3866 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3867;
  assign dataGroup_lo_hi_3867 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3868;
  assign dataGroup_lo_hi_3868 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3869;
  assign dataGroup_lo_hi_3869 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3870;
  assign dataGroup_lo_hi_3870 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3871;
  assign dataGroup_lo_hi_3871 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3872;
  assign dataGroup_lo_hi_3872 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3873;
  assign dataGroup_lo_hi_3873 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3874;
  assign dataGroup_lo_hi_3874 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3875;
  assign dataGroup_lo_hi_3875 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3876;
  assign dataGroup_lo_hi_3876 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3877;
  assign dataGroup_lo_hi_3877 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3878;
  assign dataGroup_lo_hi_3878 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3879;
  assign dataGroup_lo_hi_3879 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3880;
  assign dataGroup_lo_hi_3880 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3881;
  assign dataGroup_lo_hi_3881 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3882;
  assign dataGroup_lo_hi_3882 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3883;
  assign dataGroup_lo_hi_3883 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3884;
  assign dataGroup_lo_hi_3884 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3885;
  assign dataGroup_lo_hi_3885 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3886;
  assign dataGroup_lo_hi_3886 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3887;
  assign dataGroup_lo_hi_3887 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3888;
  assign dataGroup_lo_hi_3888 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3889;
  assign dataGroup_lo_hi_3889 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3890;
  assign dataGroup_lo_hi_3890 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3891;
  assign dataGroup_lo_hi_3891 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3892;
  assign dataGroup_lo_hi_3892 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3893;
  assign dataGroup_lo_hi_3893 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3894;
  assign dataGroup_lo_hi_3894 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3895;
  assign dataGroup_lo_hi_3895 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3896;
  assign dataGroup_lo_hi_3896 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3897;
  assign dataGroup_lo_hi_3897 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3898;
  assign dataGroup_lo_hi_3898 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3899;
  assign dataGroup_lo_hi_3899 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3900;
  assign dataGroup_lo_hi_3900 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3901;
  assign dataGroup_lo_hi_3901 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3902;
  assign dataGroup_lo_hi_3902 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3903;
  assign dataGroup_lo_hi_3903 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3904;
  assign dataGroup_lo_hi_3904 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3905;
  assign dataGroup_lo_hi_3905 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3906;
  assign dataGroup_lo_hi_3906 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3907;
  assign dataGroup_lo_hi_3907 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3908;
  assign dataGroup_lo_hi_3908 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3909;
  assign dataGroup_lo_hi_3909 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3910;
  assign dataGroup_lo_hi_3910 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3911;
  assign dataGroup_lo_hi_3911 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3912;
  assign dataGroup_lo_hi_3912 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3913;
  assign dataGroup_lo_hi_3913 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3914;
  assign dataGroup_lo_hi_3914 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3915;
  assign dataGroup_lo_hi_3915 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3916;
  assign dataGroup_lo_hi_3916 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3917;
  assign dataGroup_lo_hi_3917 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3918;
  assign dataGroup_lo_hi_3918 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3919;
  assign dataGroup_lo_hi_3919 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3920;
  assign dataGroup_lo_hi_3920 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3921;
  assign dataGroup_lo_hi_3921 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3922;
  assign dataGroup_lo_hi_3922 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3923;
  assign dataGroup_lo_hi_3923 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3924;
  assign dataGroup_lo_hi_3924 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3925;
  assign dataGroup_lo_hi_3925 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3926;
  assign dataGroup_lo_hi_3926 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3927;
  assign dataGroup_lo_hi_3927 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3928;
  assign dataGroup_lo_hi_3928 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3929;
  assign dataGroup_lo_hi_3929 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3930;
  assign dataGroup_lo_hi_3930 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3931;
  assign dataGroup_lo_hi_3931 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3932;
  assign dataGroup_lo_hi_3932 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3933;
  assign dataGroup_lo_hi_3933 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3934;
  assign dataGroup_lo_hi_3934 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3935;
  assign dataGroup_lo_hi_3935 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3936;
  assign dataGroup_lo_hi_3936 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3937;
  assign dataGroup_lo_hi_3937 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3938;
  assign dataGroup_lo_hi_3938 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3939;
  assign dataGroup_lo_hi_3939 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3940;
  assign dataGroup_lo_hi_3940 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3941;
  assign dataGroup_lo_hi_3941 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3942;
  assign dataGroup_lo_hi_3942 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3943;
  assign dataGroup_lo_hi_3943 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3944;
  assign dataGroup_lo_hi_3944 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3945;
  assign dataGroup_lo_hi_3945 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3946;
  assign dataGroup_lo_hi_3946 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3947;
  assign dataGroup_lo_hi_3947 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3948;
  assign dataGroup_lo_hi_3948 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3949;
  assign dataGroup_lo_hi_3949 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3950;
  assign dataGroup_lo_hi_3950 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3951;
  assign dataGroup_lo_hi_3951 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3952;
  assign dataGroup_lo_hi_3952 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3953;
  assign dataGroup_lo_hi_3953 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3954;
  assign dataGroup_lo_hi_3954 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3955;
  assign dataGroup_lo_hi_3955 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3956;
  assign dataGroup_lo_hi_3956 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3957;
  assign dataGroup_lo_hi_3957 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3958;
  assign dataGroup_lo_hi_3958 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3959;
  assign dataGroup_lo_hi_3959 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3960;
  assign dataGroup_lo_hi_3960 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3961;
  assign dataGroup_lo_hi_3961 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3962;
  assign dataGroup_lo_hi_3962 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3963;
  assign dataGroup_lo_hi_3963 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3964;
  assign dataGroup_lo_hi_3964 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3965;
  assign dataGroup_lo_hi_3965 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3966;
  assign dataGroup_lo_hi_3966 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3967;
  assign dataGroup_lo_hi_3967 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3968;
  assign dataGroup_lo_hi_3968 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3969;
  assign dataGroup_lo_hi_3969 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3970;
  assign dataGroup_lo_hi_3970 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3971;
  assign dataGroup_lo_hi_3971 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3972;
  assign dataGroup_lo_hi_3972 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3973;
  assign dataGroup_lo_hi_3973 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3974;
  assign dataGroup_lo_hi_3974 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3975;
  assign dataGroup_lo_hi_3975 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3976;
  assign dataGroup_lo_hi_3976 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3977;
  assign dataGroup_lo_hi_3977 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3978;
  assign dataGroup_lo_hi_3978 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3979;
  assign dataGroup_lo_hi_3979 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3980;
  assign dataGroup_lo_hi_3980 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3981;
  assign dataGroup_lo_hi_3981 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3982;
  assign dataGroup_lo_hi_3982 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3983;
  assign dataGroup_lo_hi_3983 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3984;
  assign dataGroup_lo_hi_3984 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3985;
  assign dataGroup_lo_hi_3985 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3986;
  assign dataGroup_lo_hi_3986 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3987;
  assign dataGroup_lo_hi_3987 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3988;
  assign dataGroup_lo_hi_3988 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3989;
  assign dataGroup_lo_hi_3989 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3990;
  assign dataGroup_lo_hi_3990 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3991;
  assign dataGroup_lo_hi_3991 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3992;
  assign dataGroup_lo_hi_3992 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3993;
  assign dataGroup_lo_hi_3993 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3994;
  assign dataGroup_lo_hi_3994 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3995;
  assign dataGroup_lo_hi_3995 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3996;
  assign dataGroup_lo_hi_3996 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3997;
  assign dataGroup_lo_hi_3997 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3998;
  assign dataGroup_lo_hi_3998 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_3999;
  assign dataGroup_lo_hi_3999 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4000;
  assign dataGroup_lo_hi_4000 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4001;
  assign dataGroup_lo_hi_4001 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4002;
  assign dataGroup_lo_hi_4002 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4003;
  assign dataGroup_lo_hi_4003 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4004;
  assign dataGroup_lo_hi_4004 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4005;
  assign dataGroup_lo_hi_4005 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4006;
  assign dataGroup_lo_hi_4006 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4007;
  assign dataGroup_lo_hi_4007 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4008;
  assign dataGroup_lo_hi_4008 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4009;
  assign dataGroup_lo_hi_4009 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4010;
  assign dataGroup_lo_hi_4010 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4011;
  assign dataGroup_lo_hi_4011 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4012;
  assign dataGroup_lo_hi_4012 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4013;
  assign dataGroup_lo_hi_4013 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4014;
  assign dataGroup_lo_hi_4014 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4015;
  assign dataGroup_lo_hi_4015 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4016;
  assign dataGroup_lo_hi_4016 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4017;
  assign dataGroup_lo_hi_4017 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4018;
  assign dataGroup_lo_hi_4018 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4019;
  assign dataGroup_lo_hi_4019 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4020;
  assign dataGroup_lo_hi_4020 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4021;
  assign dataGroup_lo_hi_4021 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4022;
  assign dataGroup_lo_hi_4022 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4023;
  assign dataGroup_lo_hi_4023 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4024;
  assign dataGroup_lo_hi_4024 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4025;
  assign dataGroup_lo_hi_4025 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4026;
  assign dataGroup_lo_hi_4026 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4027;
  assign dataGroup_lo_hi_4027 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4028;
  assign dataGroup_lo_hi_4028 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4029;
  assign dataGroup_lo_hi_4029 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4030;
  assign dataGroup_lo_hi_4030 = _GEN_6;
  wire [1023:0] dataGroup_lo_hi_4031;
  assign dataGroup_lo_hi_4031 = _GEN_6;
  wire [2047:0] dataGroup_lo = {dataGroup_lo_hi, dataGroup_lo_lo};
  wire [1023:0] _GEN_7 = {dataSelect_5, dataSelect_4};
  wire [1023:0] dataGroup_hi_lo;
  assign dataGroup_hi_lo = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1;
  assign dataGroup_hi_lo_1 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2;
  assign dataGroup_hi_lo_2 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3;
  assign dataGroup_hi_lo_3 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4;
  assign dataGroup_hi_lo_4 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_5;
  assign dataGroup_hi_lo_5 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_6;
  assign dataGroup_hi_lo_6 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_7;
  assign dataGroup_hi_lo_7 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_8;
  assign dataGroup_hi_lo_8 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_9;
  assign dataGroup_hi_lo_9 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_10;
  assign dataGroup_hi_lo_10 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_11;
  assign dataGroup_hi_lo_11 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_12;
  assign dataGroup_hi_lo_12 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_13;
  assign dataGroup_hi_lo_13 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_14;
  assign dataGroup_hi_lo_14 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_15;
  assign dataGroup_hi_lo_15 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_16;
  assign dataGroup_hi_lo_16 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_17;
  assign dataGroup_hi_lo_17 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_18;
  assign dataGroup_hi_lo_18 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_19;
  assign dataGroup_hi_lo_19 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_20;
  assign dataGroup_hi_lo_20 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_21;
  assign dataGroup_hi_lo_21 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_22;
  assign dataGroup_hi_lo_22 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_23;
  assign dataGroup_hi_lo_23 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_24;
  assign dataGroup_hi_lo_24 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_25;
  assign dataGroup_hi_lo_25 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_26;
  assign dataGroup_hi_lo_26 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_27;
  assign dataGroup_hi_lo_27 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_28;
  assign dataGroup_hi_lo_28 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_29;
  assign dataGroup_hi_lo_29 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_30;
  assign dataGroup_hi_lo_30 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_31;
  assign dataGroup_hi_lo_31 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_32;
  assign dataGroup_hi_lo_32 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_33;
  assign dataGroup_hi_lo_33 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_34;
  assign dataGroup_hi_lo_34 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_35;
  assign dataGroup_hi_lo_35 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_36;
  assign dataGroup_hi_lo_36 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_37;
  assign dataGroup_hi_lo_37 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_38;
  assign dataGroup_hi_lo_38 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_39;
  assign dataGroup_hi_lo_39 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_40;
  assign dataGroup_hi_lo_40 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_41;
  assign dataGroup_hi_lo_41 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_42;
  assign dataGroup_hi_lo_42 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_43;
  assign dataGroup_hi_lo_43 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_44;
  assign dataGroup_hi_lo_44 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_45;
  assign dataGroup_hi_lo_45 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_46;
  assign dataGroup_hi_lo_46 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_47;
  assign dataGroup_hi_lo_47 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_48;
  assign dataGroup_hi_lo_48 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_49;
  assign dataGroup_hi_lo_49 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_50;
  assign dataGroup_hi_lo_50 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_51;
  assign dataGroup_hi_lo_51 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_52;
  assign dataGroup_hi_lo_52 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_53;
  assign dataGroup_hi_lo_53 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_54;
  assign dataGroup_hi_lo_54 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_55;
  assign dataGroup_hi_lo_55 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_56;
  assign dataGroup_hi_lo_56 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_57;
  assign dataGroup_hi_lo_57 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_58;
  assign dataGroup_hi_lo_58 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_59;
  assign dataGroup_hi_lo_59 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_60;
  assign dataGroup_hi_lo_60 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_61;
  assign dataGroup_hi_lo_61 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_62;
  assign dataGroup_hi_lo_62 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_63;
  assign dataGroup_hi_lo_63 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_64;
  assign dataGroup_hi_lo_64 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_65;
  assign dataGroup_hi_lo_65 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_66;
  assign dataGroup_hi_lo_66 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_67;
  assign dataGroup_hi_lo_67 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_68;
  assign dataGroup_hi_lo_68 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_69;
  assign dataGroup_hi_lo_69 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_70;
  assign dataGroup_hi_lo_70 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_71;
  assign dataGroup_hi_lo_71 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_72;
  assign dataGroup_hi_lo_72 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_73;
  assign dataGroup_hi_lo_73 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_74;
  assign dataGroup_hi_lo_74 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_75;
  assign dataGroup_hi_lo_75 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_76;
  assign dataGroup_hi_lo_76 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_77;
  assign dataGroup_hi_lo_77 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_78;
  assign dataGroup_hi_lo_78 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_79;
  assign dataGroup_hi_lo_79 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_80;
  assign dataGroup_hi_lo_80 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_81;
  assign dataGroup_hi_lo_81 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_82;
  assign dataGroup_hi_lo_82 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_83;
  assign dataGroup_hi_lo_83 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_84;
  assign dataGroup_hi_lo_84 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_85;
  assign dataGroup_hi_lo_85 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_86;
  assign dataGroup_hi_lo_86 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_87;
  assign dataGroup_hi_lo_87 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_88;
  assign dataGroup_hi_lo_88 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_89;
  assign dataGroup_hi_lo_89 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_90;
  assign dataGroup_hi_lo_90 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_91;
  assign dataGroup_hi_lo_91 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_92;
  assign dataGroup_hi_lo_92 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_93;
  assign dataGroup_hi_lo_93 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_94;
  assign dataGroup_hi_lo_94 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_95;
  assign dataGroup_hi_lo_95 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_96;
  assign dataGroup_hi_lo_96 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_97;
  assign dataGroup_hi_lo_97 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_98;
  assign dataGroup_hi_lo_98 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_99;
  assign dataGroup_hi_lo_99 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_100;
  assign dataGroup_hi_lo_100 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_101;
  assign dataGroup_hi_lo_101 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_102;
  assign dataGroup_hi_lo_102 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_103;
  assign dataGroup_hi_lo_103 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_104;
  assign dataGroup_hi_lo_104 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_105;
  assign dataGroup_hi_lo_105 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_106;
  assign dataGroup_hi_lo_106 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_107;
  assign dataGroup_hi_lo_107 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_108;
  assign dataGroup_hi_lo_108 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_109;
  assign dataGroup_hi_lo_109 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_110;
  assign dataGroup_hi_lo_110 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_111;
  assign dataGroup_hi_lo_111 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_112;
  assign dataGroup_hi_lo_112 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_113;
  assign dataGroup_hi_lo_113 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_114;
  assign dataGroup_hi_lo_114 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_115;
  assign dataGroup_hi_lo_115 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_116;
  assign dataGroup_hi_lo_116 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_117;
  assign dataGroup_hi_lo_117 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_118;
  assign dataGroup_hi_lo_118 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_119;
  assign dataGroup_hi_lo_119 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_120;
  assign dataGroup_hi_lo_120 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_121;
  assign dataGroup_hi_lo_121 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_122;
  assign dataGroup_hi_lo_122 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_123;
  assign dataGroup_hi_lo_123 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_124;
  assign dataGroup_hi_lo_124 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_125;
  assign dataGroup_hi_lo_125 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_126;
  assign dataGroup_hi_lo_126 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_127;
  assign dataGroup_hi_lo_127 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_128;
  assign dataGroup_hi_lo_128 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_129;
  assign dataGroup_hi_lo_129 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_130;
  assign dataGroup_hi_lo_130 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_131;
  assign dataGroup_hi_lo_131 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_132;
  assign dataGroup_hi_lo_132 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_133;
  assign dataGroup_hi_lo_133 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_134;
  assign dataGroup_hi_lo_134 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_135;
  assign dataGroup_hi_lo_135 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_136;
  assign dataGroup_hi_lo_136 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_137;
  assign dataGroup_hi_lo_137 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_138;
  assign dataGroup_hi_lo_138 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_139;
  assign dataGroup_hi_lo_139 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_140;
  assign dataGroup_hi_lo_140 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_141;
  assign dataGroup_hi_lo_141 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_142;
  assign dataGroup_hi_lo_142 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_143;
  assign dataGroup_hi_lo_143 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_144;
  assign dataGroup_hi_lo_144 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_145;
  assign dataGroup_hi_lo_145 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_146;
  assign dataGroup_hi_lo_146 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_147;
  assign dataGroup_hi_lo_147 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_148;
  assign dataGroup_hi_lo_148 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_149;
  assign dataGroup_hi_lo_149 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_150;
  assign dataGroup_hi_lo_150 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_151;
  assign dataGroup_hi_lo_151 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_152;
  assign dataGroup_hi_lo_152 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_153;
  assign dataGroup_hi_lo_153 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_154;
  assign dataGroup_hi_lo_154 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_155;
  assign dataGroup_hi_lo_155 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_156;
  assign dataGroup_hi_lo_156 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_157;
  assign dataGroup_hi_lo_157 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_158;
  assign dataGroup_hi_lo_158 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_159;
  assign dataGroup_hi_lo_159 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_160;
  assign dataGroup_hi_lo_160 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_161;
  assign dataGroup_hi_lo_161 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_162;
  assign dataGroup_hi_lo_162 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_163;
  assign dataGroup_hi_lo_163 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_164;
  assign dataGroup_hi_lo_164 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_165;
  assign dataGroup_hi_lo_165 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_166;
  assign dataGroup_hi_lo_166 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_167;
  assign dataGroup_hi_lo_167 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_168;
  assign dataGroup_hi_lo_168 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_169;
  assign dataGroup_hi_lo_169 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_170;
  assign dataGroup_hi_lo_170 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_171;
  assign dataGroup_hi_lo_171 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_172;
  assign dataGroup_hi_lo_172 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_173;
  assign dataGroup_hi_lo_173 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_174;
  assign dataGroup_hi_lo_174 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_175;
  assign dataGroup_hi_lo_175 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_176;
  assign dataGroup_hi_lo_176 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_177;
  assign dataGroup_hi_lo_177 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_178;
  assign dataGroup_hi_lo_178 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_179;
  assign dataGroup_hi_lo_179 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_180;
  assign dataGroup_hi_lo_180 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_181;
  assign dataGroup_hi_lo_181 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_182;
  assign dataGroup_hi_lo_182 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_183;
  assign dataGroup_hi_lo_183 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_184;
  assign dataGroup_hi_lo_184 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_185;
  assign dataGroup_hi_lo_185 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_186;
  assign dataGroup_hi_lo_186 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_187;
  assign dataGroup_hi_lo_187 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_188;
  assign dataGroup_hi_lo_188 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_189;
  assign dataGroup_hi_lo_189 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_190;
  assign dataGroup_hi_lo_190 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_191;
  assign dataGroup_hi_lo_191 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_192;
  assign dataGroup_hi_lo_192 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_193;
  assign dataGroup_hi_lo_193 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_194;
  assign dataGroup_hi_lo_194 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_195;
  assign dataGroup_hi_lo_195 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_196;
  assign dataGroup_hi_lo_196 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_197;
  assign dataGroup_hi_lo_197 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_198;
  assign dataGroup_hi_lo_198 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_199;
  assign dataGroup_hi_lo_199 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_200;
  assign dataGroup_hi_lo_200 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_201;
  assign dataGroup_hi_lo_201 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_202;
  assign dataGroup_hi_lo_202 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_203;
  assign dataGroup_hi_lo_203 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_204;
  assign dataGroup_hi_lo_204 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_205;
  assign dataGroup_hi_lo_205 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_206;
  assign dataGroup_hi_lo_206 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_207;
  assign dataGroup_hi_lo_207 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_208;
  assign dataGroup_hi_lo_208 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_209;
  assign dataGroup_hi_lo_209 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_210;
  assign dataGroup_hi_lo_210 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_211;
  assign dataGroup_hi_lo_211 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_212;
  assign dataGroup_hi_lo_212 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_213;
  assign dataGroup_hi_lo_213 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_214;
  assign dataGroup_hi_lo_214 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_215;
  assign dataGroup_hi_lo_215 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_216;
  assign dataGroup_hi_lo_216 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_217;
  assign dataGroup_hi_lo_217 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_218;
  assign dataGroup_hi_lo_218 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_219;
  assign dataGroup_hi_lo_219 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_220;
  assign dataGroup_hi_lo_220 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_221;
  assign dataGroup_hi_lo_221 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_222;
  assign dataGroup_hi_lo_222 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_223;
  assign dataGroup_hi_lo_223 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_224;
  assign dataGroup_hi_lo_224 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_225;
  assign dataGroup_hi_lo_225 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_226;
  assign dataGroup_hi_lo_226 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_227;
  assign dataGroup_hi_lo_227 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_228;
  assign dataGroup_hi_lo_228 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_229;
  assign dataGroup_hi_lo_229 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_230;
  assign dataGroup_hi_lo_230 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_231;
  assign dataGroup_hi_lo_231 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_232;
  assign dataGroup_hi_lo_232 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_233;
  assign dataGroup_hi_lo_233 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_234;
  assign dataGroup_hi_lo_234 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_235;
  assign dataGroup_hi_lo_235 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_236;
  assign dataGroup_hi_lo_236 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_237;
  assign dataGroup_hi_lo_237 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_238;
  assign dataGroup_hi_lo_238 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_239;
  assign dataGroup_hi_lo_239 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_240;
  assign dataGroup_hi_lo_240 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_241;
  assign dataGroup_hi_lo_241 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_242;
  assign dataGroup_hi_lo_242 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_243;
  assign dataGroup_hi_lo_243 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_244;
  assign dataGroup_hi_lo_244 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_245;
  assign dataGroup_hi_lo_245 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_246;
  assign dataGroup_hi_lo_246 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_247;
  assign dataGroup_hi_lo_247 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_248;
  assign dataGroup_hi_lo_248 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_249;
  assign dataGroup_hi_lo_249 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_250;
  assign dataGroup_hi_lo_250 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_251;
  assign dataGroup_hi_lo_251 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_252;
  assign dataGroup_hi_lo_252 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_253;
  assign dataGroup_hi_lo_253 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_254;
  assign dataGroup_hi_lo_254 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_255;
  assign dataGroup_hi_lo_255 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_256;
  assign dataGroup_hi_lo_256 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_257;
  assign dataGroup_hi_lo_257 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_258;
  assign dataGroup_hi_lo_258 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_259;
  assign dataGroup_hi_lo_259 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_260;
  assign dataGroup_hi_lo_260 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_261;
  assign dataGroup_hi_lo_261 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_262;
  assign dataGroup_hi_lo_262 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_263;
  assign dataGroup_hi_lo_263 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_264;
  assign dataGroup_hi_lo_264 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_265;
  assign dataGroup_hi_lo_265 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_266;
  assign dataGroup_hi_lo_266 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_267;
  assign dataGroup_hi_lo_267 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_268;
  assign dataGroup_hi_lo_268 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_269;
  assign dataGroup_hi_lo_269 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_270;
  assign dataGroup_hi_lo_270 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_271;
  assign dataGroup_hi_lo_271 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_272;
  assign dataGroup_hi_lo_272 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_273;
  assign dataGroup_hi_lo_273 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_274;
  assign dataGroup_hi_lo_274 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_275;
  assign dataGroup_hi_lo_275 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_276;
  assign dataGroup_hi_lo_276 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_277;
  assign dataGroup_hi_lo_277 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_278;
  assign dataGroup_hi_lo_278 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_279;
  assign dataGroup_hi_lo_279 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_280;
  assign dataGroup_hi_lo_280 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_281;
  assign dataGroup_hi_lo_281 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_282;
  assign dataGroup_hi_lo_282 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_283;
  assign dataGroup_hi_lo_283 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_284;
  assign dataGroup_hi_lo_284 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_285;
  assign dataGroup_hi_lo_285 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_286;
  assign dataGroup_hi_lo_286 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_287;
  assign dataGroup_hi_lo_287 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_288;
  assign dataGroup_hi_lo_288 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_289;
  assign dataGroup_hi_lo_289 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_290;
  assign dataGroup_hi_lo_290 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_291;
  assign dataGroup_hi_lo_291 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_292;
  assign dataGroup_hi_lo_292 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_293;
  assign dataGroup_hi_lo_293 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_294;
  assign dataGroup_hi_lo_294 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_295;
  assign dataGroup_hi_lo_295 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_296;
  assign dataGroup_hi_lo_296 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_297;
  assign dataGroup_hi_lo_297 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_298;
  assign dataGroup_hi_lo_298 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_299;
  assign dataGroup_hi_lo_299 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_300;
  assign dataGroup_hi_lo_300 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_301;
  assign dataGroup_hi_lo_301 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_302;
  assign dataGroup_hi_lo_302 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_303;
  assign dataGroup_hi_lo_303 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_304;
  assign dataGroup_hi_lo_304 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_305;
  assign dataGroup_hi_lo_305 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_306;
  assign dataGroup_hi_lo_306 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_307;
  assign dataGroup_hi_lo_307 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_308;
  assign dataGroup_hi_lo_308 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_309;
  assign dataGroup_hi_lo_309 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_310;
  assign dataGroup_hi_lo_310 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_311;
  assign dataGroup_hi_lo_311 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_312;
  assign dataGroup_hi_lo_312 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_313;
  assign dataGroup_hi_lo_313 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_314;
  assign dataGroup_hi_lo_314 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_315;
  assign dataGroup_hi_lo_315 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_316;
  assign dataGroup_hi_lo_316 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_317;
  assign dataGroup_hi_lo_317 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_318;
  assign dataGroup_hi_lo_318 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_319;
  assign dataGroup_hi_lo_319 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_320;
  assign dataGroup_hi_lo_320 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_321;
  assign dataGroup_hi_lo_321 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_322;
  assign dataGroup_hi_lo_322 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_323;
  assign dataGroup_hi_lo_323 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_324;
  assign dataGroup_hi_lo_324 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_325;
  assign dataGroup_hi_lo_325 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_326;
  assign dataGroup_hi_lo_326 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_327;
  assign dataGroup_hi_lo_327 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_328;
  assign dataGroup_hi_lo_328 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_329;
  assign dataGroup_hi_lo_329 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_330;
  assign dataGroup_hi_lo_330 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_331;
  assign dataGroup_hi_lo_331 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_332;
  assign dataGroup_hi_lo_332 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_333;
  assign dataGroup_hi_lo_333 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_334;
  assign dataGroup_hi_lo_334 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_335;
  assign dataGroup_hi_lo_335 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_336;
  assign dataGroup_hi_lo_336 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_337;
  assign dataGroup_hi_lo_337 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_338;
  assign dataGroup_hi_lo_338 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_339;
  assign dataGroup_hi_lo_339 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_340;
  assign dataGroup_hi_lo_340 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_341;
  assign dataGroup_hi_lo_341 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_342;
  assign dataGroup_hi_lo_342 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_343;
  assign dataGroup_hi_lo_343 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_344;
  assign dataGroup_hi_lo_344 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_345;
  assign dataGroup_hi_lo_345 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_346;
  assign dataGroup_hi_lo_346 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_347;
  assign dataGroup_hi_lo_347 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_348;
  assign dataGroup_hi_lo_348 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_349;
  assign dataGroup_hi_lo_349 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_350;
  assign dataGroup_hi_lo_350 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_351;
  assign dataGroup_hi_lo_351 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_352;
  assign dataGroup_hi_lo_352 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_353;
  assign dataGroup_hi_lo_353 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_354;
  assign dataGroup_hi_lo_354 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_355;
  assign dataGroup_hi_lo_355 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_356;
  assign dataGroup_hi_lo_356 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_357;
  assign dataGroup_hi_lo_357 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_358;
  assign dataGroup_hi_lo_358 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_359;
  assign dataGroup_hi_lo_359 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_360;
  assign dataGroup_hi_lo_360 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_361;
  assign dataGroup_hi_lo_361 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_362;
  assign dataGroup_hi_lo_362 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_363;
  assign dataGroup_hi_lo_363 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_364;
  assign dataGroup_hi_lo_364 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_365;
  assign dataGroup_hi_lo_365 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_366;
  assign dataGroup_hi_lo_366 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_367;
  assign dataGroup_hi_lo_367 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_368;
  assign dataGroup_hi_lo_368 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_369;
  assign dataGroup_hi_lo_369 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_370;
  assign dataGroup_hi_lo_370 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_371;
  assign dataGroup_hi_lo_371 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_372;
  assign dataGroup_hi_lo_372 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_373;
  assign dataGroup_hi_lo_373 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_374;
  assign dataGroup_hi_lo_374 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_375;
  assign dataGroup_hi_lo_375 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_376;
  assign dataGroup_hi_lo_376 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_377;
  assign dataGroup_hi_lo_377 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_378;
  assign dataGroup_hi_lo_378 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_379;
  assign dataGroup_hi_lo_379 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_380;
  assign dataGroup_hi_lo_380 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_381;
  assign dataGroup_hi_lo_381 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_382;
  assign dataGroup_hi_lo_382 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_383;
  assign dataGroup_hi_lo_383 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_384;
  assign dataGroup_hi_lo_384 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_385;
  assign dataGroup_hi_lo_385 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_386;
  assign dataGroup_hi_lo_386 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_387;
  assign dataGroup_hi_lo_387 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_388;
  assign dataGroup_hi_lo_388 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_389;
  assign dataGroup_hi_lo_389 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_390;
  assign dataGroup_hi_lo_390 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_391;
  assign dataGroup_hi_lo_391 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_392;
  assign dataGroup_hi_lo_392 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_393;
  assign dataGroup_hi_lo_393 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_394;
  assign dataGroup_hi_lo_394 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_395;
  assign dataGroup_hi_lo_395 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_396;
  assign dataGroup_hi_lo_396 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_397;
  assign dataGroup_hi_lo_397 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_398;
  assign dataGroup_hi_lo_398 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_399;
  assign dataGroup_hi_lo_399 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_400;
  assign dataGroup_hi_lo_400 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_401;
  assign dataGroup_hi_lo_401 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_402;
  assign dataGroup_hi_lo_402 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_403;
  assign dataGroup_hi_lo_403 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_404;
  assign dataGroup_hi_lo_404 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_405;
  assign dataGroup_hi_lo_405 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_406;
  assign dataGroup_hi_lo_406 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_407;
  assign dataGroup_hi_lo_407 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_408;
  assign dataGroup_hi_lo_408 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_409;
  assign dataGroup_hi_lo_409 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_410;
  assign dataGroup_hi_lo_410 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_411;
  assign dataGroup_hi_lo_411 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_412;
  assign dataGroup_hi_lo_412 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_413;
  assign dataGroup_hi_lo_413 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_414;
  assign dataGroup_hi_lo_414 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_415;
  assign dataGroup_hi_lo_415 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_416;
  assign dataGroup_hi_lo_416 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_417;
  assign dataGroup_hi_lo_417 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_418;
  assign dataGroup_hi_lo_418 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_419;
  assign dataGroup_hi_lo_419 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_420;
  assign dataGroup_hi_lo_420 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_421;
  assign dataGroup_hi_lo_421 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_422;
  assign dataGroup_hi_lo_422 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_423;
  assign dataGroup_hi_lo_423 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_424;
  assign dataGroup_hi_lo_424 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_425;
  assign dataGroup_hi_lo_425 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_426;
  assign dataGroup_hi_lo_426 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_427;
  assign dataGroup_hi_lo_427 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_428;
  assign dataGroup_hi_lo_428 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_429;
  assign dataGroup_hi_lo_429 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_430;
  assign dataGroup_hi_lo_430 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_431;
  assign dataGroup_hi_lo_431 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_432;
  assign dataGroup_hi_lo_432 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_433;
  assign dataGroup_hi_lo_433 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_434;
  assign dataGroup_hi_lo_434 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_435;
  assign dataGroup_hi_lo_435 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_436;
  assign dataGroup_hi_lo_436 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_437;
  assign dataGroup_hi_lo_437 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_438;
  assign dataGroup_hi_lo_438 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_439;
  assign dataGroup_hi_lo_439 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_440;
  assign dataGroup_hi_lo_440 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_441;
  assign dataGroup_hi_lo_441 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_442;
  assign dataGroup_hi_lo_442 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_443;
  assign dataGroup_hi_lo_443 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_444;
  assign dataGroup_hi_lo_444 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_445;
  assign dataGroup_hi_lo_445 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_446;
  assign dataGroup_hi_lo_446 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_447;
  assign dataGroup_hi_lo_447 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_448;
  assign dataGroup_hi_lo_448 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_449;
  assign dataGroup_hi_lo_449 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_450;
  assign dataGroup_hi_lo_450 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_451;
  assign dataGroup_hi_lo_451 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_452;
  assign dataGroup_hi_lo_452 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_453;
  assign dataGroup_hi_lo_453 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_454;
  assign dataGroup_hi_lo_454 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_455;
  assign dataGroup_hi_lo_455 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_456;
  assign dataGroup_hi_lo_456 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_457;
  assign dataGroup_hi_lo_457 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_458;
  assign dataGroup_hi_lo_458 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_459;
  assign dataGroup_hi_lo_459 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_460;
  assign dataGroup_hi_lo_460 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_461;
  assign dataGroup_hi_lo_461 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_462;
  assign dataGroup_hi_lo_462 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_463;
  assign dataGroup_hi_lo_463 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_464;
  assign dataGroup_hi_lo_464 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_465;
  assign dataGroup_hi_lo_465 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_466;
  assign dataGroup_hi_lo_466 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_467;
  assign dataGroup_hi_lo_467 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_468;
  assign dataGroup_hi_lo_468 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_469;
  assign dataGroup_hi_lo_469 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_470;
  assign dataGroup_hi_lo_470 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_471;
  assign dataGroup_hi_lo_471 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_472;
  assign dataGroup_hi_lo_472 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_473;
  assign dataGroup_hi_lo_473 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_474;
  assign dataGroup_hi_lo_474 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_475;
  assign dataGroup_hi_lo_475 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_476;
  assign dataGroup_hi_lo_476 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_477;
  assign dataGroup_hi_lo_477 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_478;
  assign dataGroup_hi_lo_478 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_479;
  assign dataGroup_hi_lo_479 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_480;
  assign dataGroup_hi_lo_480 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_481;
  assign dataGroup_hi_lo_481 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_482;
  assign dataGroup_hi_lo_482 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_483;
  assign dataGroup_hi_lo_483 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_484;
  assign dataGroup_hi_lo_484 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_485;
  assign dataGroup_hi_lo_485 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_486;
  assign dataGroup_hi_lo_486 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_487;
  assign dataGroup_hi_lo_487 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_488;
  assign dataGroup_hi_lo_488 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_489;
  assign dataGroup_hi_lo_489 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_490;
  assign dataGroup_hi_lo_490 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_491;
  assign dataGroup_hi_lo_491 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_492;
  assign dataGroup_hi_lo_492 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_493;
  assign dataGroup_hi_lo_493 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_494;
  assign dataGroup_hi_lo_494 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_495;
  assign dataGroup_hi_lo_495 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_496;
  assign dataGroup_hi_lo_496 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_497;
  assign dataGroup_hi_lo_497 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_498;
  assign dataGroup_hi_lo_498 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_499;
  assign dataGroup_hi_lo_499 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_500;
  assign dataGroup_hi_lo_500 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_501;
  assign dataGroup_hi_lo_501 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_502;
  assign dataGroup_hi_lo_502 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_503;
  assign dataGroup_hi_lo_503 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_504;
  assign dataGroup_hi_lo_504 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_505;
  assign dataGroup_hi_lo_505 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_506;
  assign dataGroup_hi_lo_506 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_507;
  assign dataGroup_hi_lo_507 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_508;
  assign dataGroup_hi_lo_508 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_509;
  assign dataGroup_hi_lo_509 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_510;
  assign dataGroup_hi_lo_510 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_511;
  assign dataGroup_hi_lo_511 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_512;
  assign dataGroup_hi_lo_512 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_513;
  assign dataGroup_hi_lo_513 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_514;
  assign dataGroup_hi_lo_514 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_515;
  assign dataGroup_hi_lo_515 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_516;
  assign dataGroup_hi_lo_516 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_517;
  assign dataGroup_hi_lo_517 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_518;
  assign dataGroup_hi_lo_518 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_519;
  assign dataGroup_hi_lo_519 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_520;
  assign dataGroup_hi_lo_520 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_521;
  assign dataGroup_hi_lo_521 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_522;
  assign dataGroup_hi_lo_522 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_523;
  assign dataGroup_hi_lo_523 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_524;
  assign dataGroup_hi_lo_524 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_525;
  assign dataGroup_hi_lo_525 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_526;
  assign dataGroup_hi_lo_526 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_527;
  assign dataGroup_hi_lo_527 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_528;
  assign dataGroup_hi_lo_528 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_529;
  assign dataGroup_hi_lo_529 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_530;
  assign dataGroup_hi_lo_530 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_531;
  assign dataGroup_hi_lo_531 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_532;
  assign dataGroup_hi_lo_532 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_533;
  assign dataGroup_hi_lo_533 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_534;
  assign dataGroup_hi_lo_534 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_535;
  assign dataGroup_hi_lo_535 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_536;
  assign dataGroup_hi_lo_536 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_537;
  assign dataGroup_hi_lo_537 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_538;
  assign dataGroup_hi_lo_538 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_539;
  assign dataGroup_hi_lo_539 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_540;
  assign dataGroup_hi_lo_540 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_541;
  assign dataGroup_hi_lo_541 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_542;
  assign dataGroup_hi_lo_542 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_543;
  assign dataGroup_hi_lo_543 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_544;
  assign dataGroup_hi_lo_544 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_545;
  assign dataGroup_hi_lo_545 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_546;
  assign dataGroup_hi_lo_546 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_547;
  assign dataGroup_hi_lo_547 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_548;
  assign dataGroup_hi_lo_548 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_549;
  assign dataGroup_hi_lo_549 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_550;
  assign dataGroup_hi_lo_550 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_551;
  assign dataGroup_hi_lo_551 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_552;
  assign dataGroup_hi_lo_552 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_553;
  assign dataGroup_hi_lo_553 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_554;
  assign dataGroup_hi_lo_554 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_555;
  assign dataGroup_hi_lo_555 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_556;
  assign dataGroup_hi_lo_556 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_557;
  assign dataGroup_hi_lo_557 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_558;
  assign dataGroup_hi_lo_558 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_559;
  assign dataGroup_hi_lo_559 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_560;
  assign dataGroup_hi_lo_560 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_561;
  assign dataGroup_hi_lo_561 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_562;
  assign dataGroup_hi_lo_562 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_563;
  assign dataGroup_hi_lo_563 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_564;
  assign dataGroup_hi_lo_564 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_565;
  assign dataGroup_hi_lo_565 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_566;
  assign dataGroup_hi_lo_566 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_567;
  assign dataGroup_hi_lo_567 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_568;
  assign dataGroup_hi_lo_568 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_569;
  assign dataGroup_hi_lo_569 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_570;
  assign dataGroup_hi_lo_570 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_571;
  assign dataGroup_hi_lo_571 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_572;
  assign dataGroup_hi_lo_572 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_573;
  assign dataGroup_hi_lo_573 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_574;
  assign dataGroup_hi_lo_574 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_575;
  assign dataGroup_hi_lo_575 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_576;
  assign dataGroup_hi_lo_576 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_577;
  assign dataGroup_hi_lo_577 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_578;
  assign dataGroup_hi_lo_578 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_579;
  assign dataGroup_hi_lo_579 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_580;
  assign dataGroup_hi_lo_580 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_581;
  assign dataGroup_hi_lo_581 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_582;
  assign dataGroup_hi_lo_582 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_583;
  assign dataGroup_hi_lo_583 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_584;
  assign dataGroup_hi_lo_584 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_585;
  assign dataGroup_hi_lo_585 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_586;
  assign dataGroup_hi_lo_586 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_587;
  assign dataGroup_hi_lo_587 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_588;
  assign dataGroup_hi_lo_588 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_589;
  assign dataGroup_hi_lo_589 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_590;
  assign dataGroup_hi_lo_590 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_591;
  assign dataGroup_hi_lo_591 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_592;
  assign dataGroup_hi_lo_592 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_593;
  assign dataGroup_hi_lo_593 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_594;
  assign dataGroup_hi_lo_594 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_595;
  assign dataGroup_hi_lo_595 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_596;
  assign dataGroup_hi_lo_596 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_597;
  assign dataGroup_hi_lo_597 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_598;
  assign dataGroup_hi_lo_598 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_599;
  assign dataGroup_hi_lo_599 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_600;
  assign dataGroup_hi_lo_600 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_601;
  assign dataGroup_hi_lo_601 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_602;
  assign dataGroup_hi_lo_602 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_603;
  assign dataGroup_hi_lo_603 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_604;
  assign dataGroup_hi_lo_604 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_605;
  assign dataGroup_hi_lo_605 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_606;
  assign dataGroup_hi_lo_606 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_607;
  assign dataGroup_hi_lo_607 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_608;
  assign dataGroup_hi_lo_608 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_609;
  assign dataGroup_hi_lo_609 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_610;
  assign dataGroup_hi_lo_610 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_611;
  assign dataGroup_hi_lo_611 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_612;
  assign dataGroup_hi_lo_612 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_613;
  assign dataGroup_hi_lo_613 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_614;
  assign dataGroup_hi_lo_614 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_615;
  assign dataGroup_hi_lo_615 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_616;
  assign dataGroup_hi_lo_616 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_617;
  assign dataGroup_hi_lo_617 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_618;
  assign dataGroup_hi_lo_618 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_619;
  assign dataGroup_hi_lo_619 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_620;
  assign dataGroup_hi_lo_620 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_621;
  assign dataGroup_hi_lo_621 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_622;
  assign dataGroup_hi_lo_622 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_623;
  assign dataGroup_hi_lo_623 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_624;
  assign dataGroup_hi_lo_624 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_625;
  assign dataGroup_hi_lo_625 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_626;
  assign dataGroup_hi_lo_626 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_627;
  assign dataGroup_hi_lo_627 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_628;
  assign dataGroup_hi_lo_628 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_629;
  assign dataGroup_hi_lo_629 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_630;
  assign dataGroup_hi_lo_630 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_631;
  assign dataGroup_hi_lo_631 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_632;
  assign dataGroup_hi_lo_632 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_633;
  assign dataGroup_hi_lo_633 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_634;
  assign dataGroup_hi_lo_634 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_635;
  assign dataGroup_hi_lo_635 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_636;
  assign dataGroup_hi_lo_636 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_637;
  assign dataGroup_hi_lo_637 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_638;
  assign dataGroup_hi_lo_638 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_639;
  assign dataGroup_hi_lo_639 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_640;
  assign dataGroup_hi_lo_640 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_641;
  assign dataGroup_hi_lo_641 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_642;
  assign dataGroup_hi_lo_642 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_643;
  assign dataGroup_hi_lo_643 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_644;
  assign dataGroup_hi_lo_644 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_645;
  assign dataGroup_hi_lo_645 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_646;
  assign dataGroup_hi_lo_646 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_647;
  assign dataGroup_hi_lo_647 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_648;
  assign dataGroup_hi_lo_648 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_649;
  assign dataGroup_hi_lo_649 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_650;
  assign dataGroup_hi_lo_650 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_651;
  assign dataGroup_hi_lo_651 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_652;
  assign dataGroup_hi_lo_652 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_653;
  assign dataGroup_hi_lo_653 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_654;
  assign dataGroup_hi_lo_654 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_655;
  assign dataGroup_hi_lo_655 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_656;
  assign dataGroup_hi_lo_656 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_657;
  assign dataGroup_hi_lo_657 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_658;
  assign dataGroup_hi_lo_658 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_659;
  assign dataGroup_hi_lo_659 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_660;
  assign dataGroup_hi_lo_660 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_661;
  assign dataGroup_hi_lo_661 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_662;
  assign dataGroup_hi_lo_662 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_663;
  assign dataGroup_hi_lo_663 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_664;
  assign dataGroup_hi_lo_664 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_665;
  assign dataGroup_hi_lo_665 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_666;
  assign dataGroup_hi_lo_666 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_667;
  assign dataGroup_hi_lo_667 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_668;
  assign dataGroup_hi_lo_668 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_669;
  assign dataGroup_hi_lo_669 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_670;
  assign dataGroup_hi_lo_670 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_671;
  assign dataGroup_hi_lo_671 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_672;
  assign dataGroup_hi_lo_672 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_673;
  assign dataGroup_hi_lo_673 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_674;
  assign dataGroup_hi_lo_674 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_675;
  assign dataGroup_hi_lo_675 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_676;
  assign dataGroup_hi_lo_676 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_677;
  assign dataGroup_hi_lo_677 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_678;
  assign dataGroup_hi_lo_678 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_679;
  assign dataGroup_hi_lo_679 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_680;
  assign dataGroup_hi_lo_680 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_681;
  assign dataGroup_hi_lo_681 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_682;
  assign dataGroup_hi_lo_682 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_683;
  assign dataGroup_hi_lo_683 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_684;
  assign dataGroup_hi_lo_684 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_685;
  assign dataGroup_hi_lo_685 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_686;
  assign dataGroup_hi_lo_686 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_687;
  assign dataGroup_hi_lo_687 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_688;
  assign dataGroup_hi_lo_688 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_689;
  assign dataGroup_hi_lo_689 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_690;
  assign dataGroup_hi_lo_690 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_691;
  assign dataGroup_hi_lo_691 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_692;
  assign dataGroup_hi_lo_692 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_693;
  assign dataGroup_hi_lo_693 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_694;
  assign dataGroup_hi_lo_694 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_695;
  assign dataGroup_hi_lo_695 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_696;
  assign dataGroup_hi_lo_696 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_697;
  assign dataGroup_hi_lo_697 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_698;
  assign dataGroup_hi_lo_698 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_699;
  assign dataGroup_hi_lo_699 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_700;
  assign dataGroup_hi_lo_700 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_701;
  assign dataGroup_hi_lo_701 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_702;
  assign dataGroup_hi_lo_702 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_703;
  assign dataGroup_hi_lo_703 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_704;
  assign dataGroup_hi_lo_704 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_705;
  assign dataGroup_hi_lo_705 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_706;
  assign dataGroup_hi_lo_706 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_707;
  assign dataGroup_hi_lo_707 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_708;
  assign dataGroup_hi_lo_708 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_709;
  assign dataGroup_hi_lo_709 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_710;
  assign dataGroup_hi_lo_710 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_711;
  assign dataGroup_hi_lo_711 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_712;
  assign dataGroup_hi_lo_712 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_713;
  assign dataGroup_hi_lo_713 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_714;
  assign dataGroup_hi_lo_714 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_715;
  assign dataGroup_hi_lo_715 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_716;
  assign dataGroup_hi_lo_716 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_717;
  assign dataGroup_hi_lo_717 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_718;
  assign dataGroup_hi_lo_718 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_719;
  assign dataGroup_hi_lo_719 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_720;
  assign dataGroup_hi_lo_720 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_721;
  assign dataGroup_hi_lo_721 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_722;
  assign dataGroup_hi_lo_722 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_723;
  assign dataGroup_hi_lo_723 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_724;
  assign dataGroup_hi_lo_724 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_725;
  assign dataGroup_hi_lo_725 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_726;
  assign dataGroup_hi_lo_726 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_727;
  assign dataGroup_hi_lo_727 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_728;
  assign dataGroup_hi_lo_728 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_729;
  assign dataGroup_hi_lo_729 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_730;
  assign dataGroup_hi_lo_730 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_731;
  assign dataGroup_hi_lo_731 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_732;
  assign dataGroup_hi_lo_732 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_733;
  assign dataGroup_hi_lo_733 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_734;
  assign dataGroup_hi_lo_734 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_735;
  assign dataGroup_hi_lo_735 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_736;
  assign dataGroup_hi_lo_736 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_737;
  assign dataGroup_hi_lo_737 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_738;
  assign dataGroup_hi_lo_738 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_739;
  assign dataGroup_hi_lo_739 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_740;
  assign dataGroup_hi_lo_740 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_741;
  assign dataGroup_hi_lo_741 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_742;
  assign dataGroup_hi_lo_742 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_743;
  assign dataGroup_hi_lo_743 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_744;
  assign dataGroup_hi_lo_744 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_745;
  assign dataGroup_hi_lo_745 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_746;
  assign dataGroup_hi_lo_746 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_747;
  assign dataGroup_hi_lo_747 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_748;
  assign dataGroup_hi_lo_748 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_749;
  assign dataGroup_hi_lo_749 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_750;
  assign dataGroup_hi_lo_750 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_751;
  assign dataGroup_hi_lo_751 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_752;
  assign dataGroup_hi_lo_752 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_753;
  assign dataGroup_hi_lo_753 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_754;
  assign dataGroup_hi_lo_754 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_755;
  assign dataGroup_hi_lo_755 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_756;
  assign dataGroup_hi_lo_756 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_757;
  assign dataGroup_hi_lo_757 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_758;
  assign dataGroup_hi_lo_758 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_759;
  assign dataGroup_hi_lo_759 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_760;
  assign dataGroup_hi_lo_760 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_761;
  assign dataGroup_hi_lo_761 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_762;
  assign dataGroup_hi_lo_762 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_763;
  assign dataGroup_hi_lo_763 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_764;
  assign dataGroup_hi_lo_764 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_765;
  assign dataGroup_hi_lo_765 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_766;
  assign dataGroup_hi_lo_766 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_767;
  assign dataGroup_hi_lo_767 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_768;
  assign dataGroup_hi_lo_768 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_769;
  assign dataGroup_hi_lo_769 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_770;
  assign dataGroup_hi_lo_770 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_771;
  assign dataGroup_hi_lo_771 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_772;
  assign dataGroup_hi_lo_772 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_773;
  assign dataGroup_hi_lo_773 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_774;
  assign dataGroup_hi_lo_774 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_775;
  assign dataGroup_hi_lo_775 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_776;
  assign dataGroup_hi_lo_776 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_777;
  assign dataGroup_hi_lo_777 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_778;
  assign dataGroup_hi_lo_778 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_779;
  assign dataGroup_hi_lo_779 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_780;
  assign dataGroup_hi_lo_780 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_781;
  assign dataGroup_hi_lo_781 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_782;
  assign dataGroup_hi_lo_782 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_783;
  assign dataGroup_hi_lo_783 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_784;
  assign dataGroup_hi_lo_784 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_785;
  assign dataGroup_hi_lo_785 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_786;
  assign dataGroup_hi_lo_786 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_787;
  assign dataGroup_hi_lo_787 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_788;
  assign dataGroup_hi_lo_788 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_789;
  assign dataGroup_hi_lo_789 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_790;
  assign dataGroup_hi_lo_790 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_791;
  assign dataGroup_hi_lo_791 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_792;
  assign dataGroup_hi_lo_792 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_793;
  assign dataGroup_hi_lo_793 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_794;
  assign dataGroup_hi_lo_794 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_795;
  assign dataGroup_hi_lo_795 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_796;
  assign dataGroup_hi_lo_796 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_797;
  assign dataGroup_hi_lo_797 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_798;
  assign dataGroup_hi_lo_798 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_799;
  assign dataGroup_hi_lo_799 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_800;
  assign dataGroup_hi_lo_800 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_801;
  assign dataGroup_hi_lo_801 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_802;
  assign dataGroup_hi_lo_802 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_803;
  assign dataGroup_hi_lo_803 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_804;
  assign dataGroup_hi_lo_804 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_805;
  assign dataGroup_hi_lo_805 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_806;
  assign dataGroup_hi_lo_806 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_807;
  assign dataGroup_hi_lo_807 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_808;
  assign dataGroup_hi_lo_808 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_809;
  assign dataGroup_hi_lo_809 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_810;
  assign dataGroup_hi_lo_810 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_811;
  assign dataGroup_hi_lo_811 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_812;
  assign dataGroup_hi_lo_812 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_813;
  assign dataGroup_hi_lo_813 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_814;
  assign dataGroup_hi_lo_814 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_815;
  assign dataGroup_hi_lo_815 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_816;
  assign dataGroup_hi_lo_816 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_817;
  assign dataGroup_hi_lo_817 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_818;
  assign dataGroup_hi_lo_818 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_819;
  assign dataGroup_hi_lo_819 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_820;
  assign dataGroup_hi_lo_820 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_821;
  assign dataGroup_hi_lo_821 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_822;
  assign dataGroup_hi_lo_822 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_823;
  assign dataGroup_hi_lo_823 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_824;
  assign dataGroup_hi_lo_824 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_825;
  assign dataGroup_hi_lo_825 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_826;
  assign dataGroup_hi_lo_826 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_827;
  assign dataGroup_hi_lo_827 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_828;
  assign dataGroup_hi_lo_828 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_829;
  assign dataGroup_hi_lo_829 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_830;
  assign dataGroup_hi_lo_830 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_831;
  assign dataGroup_hi_lo_831 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_832;
  assign dataGroup_hi_lo_832 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_833;
  assign dataGroup_hi_lo_833 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_834;
  assign dataGroup_hi_lo_834 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_835;
  assign dataGroup_hi_lo_835 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_836;
  assign dataGroup_hi_lo_836 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_837;
  assign dataGroup_hi_lo_837 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_838;
  assign dataGroup_hi_lo_838 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_839;
  assign dataGroup_hi_lo_839 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_840;
  assign dataGroup_hi_lo_840 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_841;
  assign dataGroup_hi_lo_841 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_842;
  assign dataGroup_hi_lo_842 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_843;
  assign dataGroup_hi_lo_843 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_844;
  assign dataGroup_hi_lo_844 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_845;
  assign dataGroup_hi_lo_845 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_846;
  assign dataGroup_hi_lo_846 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_847;
  assign dataGroup_hi_lo_847 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_848;
  assign dataGroup_hi_lo_848 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_849;
  assign dataGroup_hi_lo_849 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_850;
  assign dataGroup_hi_lo_850 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_851;
  assign dataGroup_hi_lo_851 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_852;
  assign dataGroup_hi_lo_852 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_853;
  assign dataGroup_hi_lo_853 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_854;
  assign dataGroup_hi_lo_854 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_855;
  assign dataGroup_hi_lo_855 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_856;
  assign dataGroup_hi_lo_856 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_857;
  assign dataGroup_hi_lo_857 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_858;
  assign dataGroup_hi_lo_858 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_859;
  assign dataGroup_hi_lo_859 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_860;
  assign dataGroup_hi_lo_860 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_861;
  assign dataGroup_hi_lo_861 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_862;
  assign dataGroup_hi_lo_862 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_863;
  assign dataGroup_hi_lo_863 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_864;
  assign dataGroup_hi_lo_864 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_865;
  assign dataGroup_hi_lo_865 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_866;
  assign dataGroup_hi_lo_866 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_867;
  assign dataGroup_hi_lo_867 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_868;
  assign dataGroup_hi_lo_868 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_869;
  assign dataGroup_hi_lo_869 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_870;
  assign dataGroup_hi_lo_870 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_871;
  assign dataGroup_hi_lo_871 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_872;
  assign dataGroup_hi_lo_872 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_873;
  assign dataGroup_hi_lo_873 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_874;
  assign dataGroup_hi_lo_874 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_875;
  assign dataGroup_hi_lo_875 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_876;
  assign dataGroup_hi_lo_876 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_877;
  assign dataGroup_hi_lo_877 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_878;
  assign dataGroup_hi_lo_878 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_879;
  assign dataGroup_hi_lo_879 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_880;
  assign dataGroup_hi_lo_880 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_881;
  assign dataGroup_hi_lo_881 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_882;
  assign dataGroup_hi_lo_882 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_883;
  assign dataGroup_hi_lo_883 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_884;
  assign dataGroup_hi_lo_884 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_885;
  assign dataGroup_hi_lo_885 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_886;
  assign dataGroup_hi_lo_886 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_887;
  assign dataGroup_hi_lo_887 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_888;
  assign dataGroup_hi_lo_888 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_889;
  assign dataGroup_hi_lo_889 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_890;
  assign dataGroup_hi_lo_890 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_891;
  assign dataGroup_hi_lo_891 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_892;
  assign dataGroup_hi_lo_892 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_893;
  assign dataGroup_hi_lo_893 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_894;
  assign dataGroup_hi_lo_894 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_895;
  assign dataGroup_hi_lo_895 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_896;
  assign dataGroup_hi_lo_896 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_897;
  assign dataGroup_hi_lo_897 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_898;
  assign dataGroup_hi_lo_898 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_899;
  assign dataGroup_hi_lo_899 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_900;
  assign dataGroup_hi_lo_900 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_901;
  assign dataGroup_hi_lo_901 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_902;
  assign dataGroup_hi_lo_902 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_903;
  assign dataGroup_hi_lo_903 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_904;
  assign dataGroup_hi_lo_904 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_905;
  assign dataGroup_hi_lo_905 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_906;
  assign dataGroup_hi_lo_906 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_907;
  assign dataGroup_hi_lo_907 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_908;
  assign dataGroup_hi_lo_908 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_909;
  assign dataGroup_hi_lo_909 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_910;
  assign dataGroup_hi_lo_910 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_911;
  assign dataGroup_hi_lo_911 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_912;
  assign dataGroup_hi_lo_912 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_913;
  assign dataGroup_hi_lo_913 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_914;
  assign dataGroup_hi_lo_914 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_915;
  assign dataGroup_hi_lo_915 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_916;
  assign dataGroup_hi_lo_916 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_917;
  assign dataGroup_hi_lo_917 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_918;
  assign dataGroup_hi_lo_918 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_919;
  assign dataGroup_hi_lo_919 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_920;
  assign dataGroup_hi_lo_920 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_921;
  assign dataGroup_hi_lo_921 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_922;
  assign dataGroup_hi_lo_922 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_923;
  assign dataGroup_hi_lo_923 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_924;
  assign dataGroup_hi_lo_924 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_925;
  assign dataGroup_hi_lo_925 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_926;
  assign dataGroup_hi_lo_926 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_927;
  assign dataGroup_hi_lo_927 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_928;
  assign dataGroup_hi_lo_928 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_929;
  assign dataGroup_hi_lo_929 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_930;
  assign dataGroup_hi_lo_930 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_931;
  assign dataGroup_hi_lo_931 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_932;
  assign dataGroup_hi_lo_932 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_933;
  assign dataGroup_hi_lo_933 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_934;
  assign dataGroup_hi_lo_934 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_935;
  assign dataGroup_hi_lo_935 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_936;
  assign dataGroup_hi_lo_936 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_937;
  assign dataGroup_hi_lo_937 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_938;
  assign dataGroup_hi_lo_938 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_939;
  assign dataGroup_hi_lo_939 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_940;
  assign dataGroup_hi_lo_940 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_941;
  assign dataGroup_hi_lo_941 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_942;
  assign dataGroup_hi_lo_942 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_943;
  assign dataGroup_hi_lo_943 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_944;
  assign dataGroup_hi_lo_944 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_945;
  assign dataGroup_hi_lo_945 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_946;
  assign dataGroup_hi_lo_946 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_947;
  assign dataGroup_hi_lo_947 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_948;
  assign dataGroup_hi_lo_948 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_949;
  assign dataGroup_hi_lo_949 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_950;
  assign dataGroup_hi_lo_950 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_951;
  assign dataGroup_hi_lo_951 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_952;
  assign dataGroup_hi_lo_952 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_953;
  assign dataGroup_hi_lo_953 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_954;
  assign dataGroup_hi_lo_954 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_955;
  assign dataGroup_hi_lo_955 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_956;
  assign dataGroup_hi_lo_956 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_957;
  assign dataGroup_hi_lo_957 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_958;
  assign dataGroup_hi_lo_958 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_959;
  assign dataGroup_hi_lo_959 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_960;
  assign dataGroup_hi_lo_960 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_961;
  assign dataGroup_hi_lo_961 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_962;
  assign dataGroup_hi_lo_962 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_963;
  assign dataGroup_hi_lo_963 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_964;
  assign dataGroup_hi_lo_964 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_965;
  assign dataGroup_hi_lo_965 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_966;
  assign dataGroup_hi_lo_966 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_967;
  assign dataGroup_hi_lo_967 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_968;
  assign dataGroup_hi_lo_968 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_969;
  assign dataGroup_hi_lo_969 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_970;
  assign dataGroup_hi_lo_970 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_971;
  assign dataGroup_hi_lo_971 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_972;
  assign dataGroup_hi_lo_972 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_973;
  assign dataGroup_hi_lo_973 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_974;
  assign dataGroup_hi_lo_974 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_975;
  assign dataGroup_hi_lo_975 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_976;
  assign dataGroup_hi_lo_976 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_977;
  assign dataGroup_hi_lo_977 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_978;
  assign dataGroup_hi_lo_978 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_979;
  assign dataGroup_hi_lo_979 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_980;
  assign dataGroup_hi_lo_980 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_981;
  assign dataGroup_hi_lo_981 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_982;
  assign dataGroup_hi_lo_982 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_983;
  assign dataGroup_hi_lo_983 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_984;
  assign dataGroup_hi_lo_984 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_985;
  assign dataGroup_hi_lo_985 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_986;
  assign dataGroup_hi_lo_986 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_987;
  assign dataGroup_hi_lo_987 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_988;
  assign dataGroup_hi_lo_988 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_989;
  assign dataGroup_hi_lo_989 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_990;
  assign dataGroup_hi_lo_990 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_991;
  assign dataGroup_hi_lo_991 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_992;
  assign dataGroup_hi_lo_992 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_993;
  assign dataGroup_hi_lo_993 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_994;
  assign dataGroup_hi_lo_994 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_995;
  assign dataGroup_hi_lo_995 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_996;
  assign dataGroup_hi_lo_996 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_997;
  assign dataGroup_hi_lo_997 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_998;
  assign dataGroup_hi_lo_998 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_999;
  assign dataGroup_hi_lo_999 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1000;
  assign dataGroup_hi_lo_1000 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1001;
  assign dataGroup_hi_lo_1001 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1002;
  assign dataGroup_hi_lo_1002 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1003;
  assign dataGroup_hi_lo_1003 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1004;
  assign dataGroup_hi_lo_1004 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1005;
  assign dataGroup_hi_lo_1005 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1006;
  assign dataGroup_hi_lo_1006 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1007;
  assign dataGroup_hi_lo_1007 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1008;
  assign dataGroup_hi_lo_1008 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1009;
  assign dataGroup_hi_lo_1009 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1010;
  assign dataGroup_hi_lo_1010 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1011;
  assign dataGroup_hi_lo_1011 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1012;
  assign dataGroup_hi_lo_1012 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1013;
  assign dataGroup_hi_lo_1013 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1014;
  assign dataGroup_hi_lo_1014 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1015;
  assign dataGroup_hi_lo_1015 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1016;
  assign dataGroup_hi_lo_1016 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1017;
  assign dataGroup_hi_lo_1017 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1018;
  assign dataGroup_hi_lo_1018 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1019;
  assign dataGroup_hi_lo_1019 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1020;
  assign dataGroup_hi_lo_1020 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1021;
  assign dataGroup_hi_lo_1021 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1022;
  assign dataGroup_hi_lo_1022 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1023;
  assign dataGroup_hi_lo_1023 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1024;
  assign dataGroup_hi_lo_1024 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1025;
  assign dataGroup_hi_lo_1025 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1026;
  assign dataGroup_hi_lo_1026 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1027;
  assign dataGroup_hi_lo_1027 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1028;
  assign dataGroup_hi_lo_1028 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1029;
  assign dataGroup_hi_lo_1029 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1030;
  assign dataGroup_hi_lo_1030 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1031;
  assign dataGroup_hi_lo_1031 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1032;
  assign dataGroup_hi_lo_1032 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1033;
  assign dataGroup_hi_lo_1033 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1034;
  assign dataGroup_hi_lo_1034 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1035;
  assign dataGroup_hi_lo_1035 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1036;
  assign dataGroup_hi_lo_1036 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1037;
  assign dataGroup_hi_lo_1037 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1038;
  assign dataGroup_hi_lo_1038 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1039;
  assign dataGroup_hi_lo_1039 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1040;
  assign dataGroup_hi_lo_1040 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1041;
  assign dataGroup_hi_lo_1041 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1042;
  assign dataGroup_hi_lo_1042 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1043;
  assign dataGroup_hi_lo_1043 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1044;
  assign dataGroup_hi_lo_1044 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1045;
  assign dataGroup_hi_lo_1045 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1046;
  assign dataGroup_hi_lo_1046 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1047;
  assign dataGroup_hi_lo_1047 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1048;
  assign dataGroup_hi_lo_1048 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1049;
  assign dataGroup_hi_lo_1049 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1050;
  assign dataGroup_hi_lo_1050 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1051;
  assign dataGroup_hi_lo_1051 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1052;
  assign dataGroup_hi_lo_1052 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1053;
  assign dataGroup_hi_lo_1053 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1054;
  assign dataGroup_hi_lo_1054 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1055;
  assign dataGroup_hi_lo_1055 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1056;
  assign dataGroup_hi_lo_1056 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1057;
  assign dataGroup_hi_lo_1057 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1058;
  assign dataGroup_hi_lo_1058 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1059;
  assign dataGroup_hi_lo_1059 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1060;
  assign dataGroup_hi_lo_1060 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1061;
  assign dataGroup_hi_lo_1061 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1062;
  assign dataGroup_hi_lo_1062 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1063;
  assign dataGroup_hi_lo_1063 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1064;
  assign dataGroup_hi_lo_1064 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1065;
  assign dataGroup_hi_lo_1065 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1066;
  assign dataGroup_hi_lo_1066 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1067;
  assign dataGroup_hi_lo_1067 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1068;
  assign dataGroup_hi_lo_1068 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1069;
  assign dataGroup_hi_lo_1069 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1070;
  assign dataGroup_hi_lo_1070 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1071;
  assign dataGroup_hi_lo_1071 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1072;
  assign dataGroup_hi_lo_1072 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1073;
  assign dataGroup_hi_lo_1073 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1074;
  assign dataGroup_hi_lo_1074 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1075;
  assign dataGroup_hi_lo_1075 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1076;
  assign dataGroup_hi_lo_1076 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1077;
  assign dataGroup_hi_lo_1077 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1078;
  assign dataGroup_hi_lo_1078 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1079;
  assign dataGroup_hi_lo_1079 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1080;
  assign dataGroup_hi_lo_1080 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1081;
  assign dataGroup_hi_lo_1081 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1082;
  assign dataGroup_hi_lo_1082 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1083;
  assign dataGroup_hi_lo_1083 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1084;
  assign dataGroup_hi_lo_1084 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1085;
  assign dataGroup_hi_lo_1085 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1086;
  assign dataGroup_hi_lo_1086 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1087;
  assign dataGroup_hi_lo_1087 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1088;
  assign dataGroup_hi_lo_1088 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1089;
  assign dataGroup_hi_lo_1089 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1090;
  assign dataGroup_hi_lo_1090 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1091;
  assign dataGroup_hi_lo_1091 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1092;
  assign dataGroup_hi_lo_1092 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1093;
  assign dataGroup_hi_lo_1093 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1094;
  assign dataGroup_hi_lo_1094 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1095;
  assign dataGroup_hi_lo_1095 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1096;
  assign dataGroup_hi_lo_1096 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1097;
  assign dataGroup_hi_lo_1097 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1098;
  assign dataGroup_hi_lo_1098 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1099;
  assign dataGroup_hi_lo_1099 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1100;
  assign dataGroup_hi_lo_1100 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1101;
  assign dataGroup_hi_lo_1101 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1102;
  assign dataGroup_hi_lo_1102 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1103;
  assign dataGroup_hi_lo_1103 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1104;
  assign dataGroup_hi_lo_1104 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1105;
  assign dataGroup_hi_lo_1105 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1106;
  assign dataGroup_hi_lo_1106 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1107;
  assign dataGroup_hi_lo_1107 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1108;
  assign dataGroup_hi_lo_1108 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1109;
  assign dataGroup_hi_lo_1109 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1110;
  assign dataGroup_hi_lo_1110 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1111;
  assign dataGroup_hi_lo_1111 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1112;
  assign dataGroup_hi_lo_1112 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1113;
  assign dataGroup_hi_lo_1113 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1114;
  assign dataGroup_hi_lo_1114 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1115;
  assign dataGroup_hi_lo_1115 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1116;
  assign dataGroup_hi_lo_1116 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1117;
  assign dataGroup_hi_lo_1117 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1118;
  assign dataGroup_hi_lo_1118 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1119;
  assign dataGroup_hi_lo_1119 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1120;
  assign dataGroup_hi_lo_1120 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1121;
  assign dataGroup_hi_lo_1121 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1122;
  assign dataGroup_hi_lo_1122 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1123;
  assign dataGroup_hi_lo_1123 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1124;
  assign dataGroup_hi_lo_1124 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1125;
  assign dataGroup_hi_lo_1125 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1126;
  assign dataGroup_hi_lo_1126 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1127;
  assign dataGroup_hi_lo_1127 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1128;
  assign dataGroup_hi_lo_1128 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1129;
  assign dataGroup_hi_lo_1129 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1130;
  assign dataGroup_hi_lo_1130 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1131;
  assign dataGroup_hi_lo_1131 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1132;
  assign dataGroup_hi_lo_1132 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1133;
  assign dataGroup_hi_lo_1133 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1134;
  assign dataGroup_hi_lo_1134 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1135;
  assign dataGroup_hi_lo_1135 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1136;
  assign dataGroup_hi_lo_1136 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1137;
  assign dataGroup_hi_lo_1137 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1138;
  assign dataGroup_hi_lo_1138 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1139;
  assign dataGroup_hi_lo_1139 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1140;
  assign dataGroup_hi_lo_1140 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1141;
  assign dataGroup_hi_lo_1141 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1142;
  assign dataGroup_hi_lo_1142 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1143;
  assign dataGroup_hi_lo_1143 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1144;
  assign dataGroup_hi_lo_1144 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1145;
  assign dataGroup_hi_lo_1145 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1146;
  assign dataGroup_hi_lo_1146 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1147;
  assign dataGroup_hi_lo_1147 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1148;
  assign dataGroup_hi_lo_1148 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1149;
  assign dataGroup_hi_lo_1149 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1150;
  assign dataGroup_hi_lo_1150 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1151;
  assign dataGroup_hi_lo_1151 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1152;
  assign dataGroup_hi_lo_1152 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1153;
  assign dataGroup_hi_lo_1153 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1154;
  assign dataGroup_hi_lo_1154 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1155;
  assign dataGroup_hi_lo_1155 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1156;
  assign dataGroup_hi_lo_1156 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1157;
  assign dataGroup_hi_lo_1157 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1158;
  assign dataGroup_hi_lo_1158 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1159;
  assign dataGroup_hi_lo_1159 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1160;
  assign dataGroup_hi_lo_1160 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1161;
  assign dataGroup_hi_lo_1161 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1162;
  assign dataGroup_hi_lo_1162 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1163;
  assign dataGroup_hi_lo_1163 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1164;
  assign dataGroup_hi_lo_1164 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1165;
  assign dataGroup_hi_lo_1165 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1166;
  assign dataGroup_hi_lo_1166 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1167;
  assign dataGroup_hi_lo_1167 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1168;
  assign dataGroup_hi_lo_1168 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1169;
  assign dataGroup_hi_lo_1169 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1170;
  assign dataGroup_hi_lo_1170 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1171;
  assign dataGroup_hi_lo_1171 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1172;
  assign dataGroup_hi_lo_1172 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1173;
  assign dataGroup_hi_lo_1173 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1174;
  assign dataGroup_hi_lo_1174 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1175;
  assign dataGroup_hi_lo_1175 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1176;
  assign dataGroup_hi_lo_1176 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1177;
  assign dataGroup_hi_lo_1177 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1178;
  assign dataGroup_hi_lo_1178 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1179;
  assign dataGroup_hi_lo_1179 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1180;
  assign dataGroup_hi_lo_1180 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1181;
  assign dataGroup_hi_lo_1181 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1182;
  assign dataGroup_hi_lo_1182 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1183;
  assign dataGroup_hi_lo_1183 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1184;
  assign dataGroup_hi_lo_1184 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1185;
  assign dataGroup_hi_lo_1185 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1186;
  assign dataGroup_hi_lo_1186 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1187;
  assign dataGroup_hi_lo_1187 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1188;
  assign dataGroup_hi_lo_1188 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1189;
  assign dataGroup_hi_lo_1189 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1190;
  assign dataGroup_hi_lo_1190 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1191;
  assign dataGroup_hi_lo_1191 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1192;
  assign dataGroup_hi_lo_1192 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1193;
  assign dataGroup_hi_lo_1193 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1194;
  assign dataGroup_hi_lo_1194 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1195;
  assign dataGroup_hi_lo_1195 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1196;
  assign dataGroup_hi_lo_1196 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1197;
  assign dataGroup_hi_lo_1197 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1198;
  assign dataGroup_hi_lo_1198 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1199;
  assign dataGroup_hi_lo_1199 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1200;
  assign dataGroup_hi_lo_1200 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1201;
  assign dataGroup_hi_lo_1201 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1202;
  assign dataGroup_hi_lo_1202 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1203;
  assign dataGroup_hi_lo_1203 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1204;
  assign dataGroup_hi_lo_1204 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1205;
  assign dataGroup_hi_lo_1205 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1206;
  assign dataGroup_hi_lo_1206 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1207;
  assign dataGroup_hi_lo_1207 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1208;
  assign dataGroup_hi_lo_1208 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1209;
  assign dataGroup_hi_lo_1209 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1210;
  assign dataGroup_hi_lo_1210 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1211;
  assign dataGroup_hi_lo_1211 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1212;
  assign dataGroup_hi_lo_1212 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1213;
  assign dataGroup_hi_lo_1213 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1214;
  assign dataGroup_hi_lo_1214 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1215;
  assign dataGroup_hi_lo_1215 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1216;
  assign dataGroup_hi_lo_1216 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1217;
  assign dataGroup_hi_lo_1217 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1218;
  assign dataGroup_hi_lo_1218 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1219;
  assign dataGroup_hi_lo_1219 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1220;
  assign dataGroup_hi_lo_1220 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1221;
  assign dataGroup_hi_lo_1221 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1222;
  assign dataGroup_hi_lo_1222 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1223;
  assign dataGroup_hi_lo_1223 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1224;
  assign dataGroup_hi_lo_1224 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1225;
  assign dataGroup_hi_lo_1225 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1226;
  assign dataGroup_hi_lo_1226 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1227;
  assign dataGroup_hi_lo_1227 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1228;
  assign dataGroup_hi_lo_1228 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1229;
  assign dataGroup_hi_lo_1229 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1230;
  assign dataGroup_hi_lo_1230 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1231;
  assign dataGroup_hi_lo_1231 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1232;
  assign dataGroup_hi_lo_1232 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1233;
  assign dataGroup_hi_lo_1233 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1234;
  assign dataGroup_hi_lo_1234 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1235;
  assign dataGroup_hi_lo_1235 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1236;
  assign dataGroup_hi_lo_1236 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1237;
  assign dataGroup_hi_lo_1237 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1238;
  assign dataGroup_hi_lo_1238 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1239;
  assign dataGroup_hi_lo_1239 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1240;
  assign dataGroup_hi_lo_1240 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1241;
  assign dataGroup_hi_lo_1241 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1242;
  assign dataGroup_hi_lo_1242 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1243;
  assign dataGroup_hi_lo_1243 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1244;
  assign dataGroup_hi_lo_1244 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1245;
  assign dataGroup_hi_lo_1245 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1246;
  assign dataGroup_hi_lo_1246 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1247;
  assign dataGroup_hi_lo_1247 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1248;
  assign dataGroup_hi_lo_1248 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1249;
  assign dataGroup_hi_lo_1249 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1250;
  assign dataGroup_hi_lo_1250 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1251;
  assign dataGroup_hi_lo_1251 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1252;
  assign dataGroup_hi_lo_1252 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1253;
  assign dataGroup_hi_lo_1253 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1254;
  assign dataGroup_hi_lo_1254 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1255;
  assign dataGroup_hi_lo_1255 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1256;
  assign dataGroup_hi_lo_1256 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1257;
  assign dataGroup_hi_lo_1257 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1258;
  assign dataGroup_hi_lo_1258 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1259;
  assign dataGroup_hi_lo_1259 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1260;
  assign dataGroup_hi_lo_1260 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1261;
  assign dataGroup_hi_lo_1261 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1262;
  assign dataGroup_hi_lo_1262 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1263;
  assign dataGroup_hi_lo_1263 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1264;
  assign dataGroup_hi_lo_1264 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1265;
  assign dataGroup_hi_lo_1265 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1266;
  assign dataGroup_hi_lo_1266 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1267;
  assign dataGroup_hi_lo_1267 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1268;
  assign dataGroup_hi_lo_1268 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1269;
  assign dataGroup_hi_lo_1269 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1270;
  assign dataGroup_hi_lo_1270 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1271;
  assign dataGroup_hi_lo_1271 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1272;
  assign dataGroup_hi_lo_1272 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1273;
  assign dataGroup_hi_lo_1273 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1274;
  assign dataGroup_hi_lo_1274 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1275;
  assign dataGroup_hi_lo_1275 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1276;
  assign dataGroup_hi_lo_1276 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1277;
  assign dataGroup_hi_lo_1277 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1278;
  assign dataGroup_hi_lo_1278 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1279;
  assign dataGroup_hi_lo_1279 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1280;
  assign dataGroup_hi_lo_1280 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1281;
  assign dataGroup_hi_lo_1281 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1282;
  assign dataGroup_hi_lo_1282 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1283;
  assign dataGroup_hi_lo_1283 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1284;
  assign dataGroup_hi_lo_1284 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1285;
  assign dataGroup_hi_lo_1285 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1286;
  assign dataGroup_hi_lo_1286 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1287;
  assign dataGroup_hi_lo_1287 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1288;
  assign dataGroup_hi_lo_1288 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1289;
  assign dataGroup_hi_lo_1289 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1290;
  assign dataGroup_hi_lo_1290 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1291;
  assign dataGroup_hi_lo_1291 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1292;
  assign dataGroup_hi_lo_1292 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1293;
  assign dataGroup_hi_lo_1293 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1294;
  assign dataGroup_hi_lo_1294 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1295;
  assign dataGroup_hi_lo_1295 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1296;
  assign dataGroup_hi_lo_1296 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1297;
  assign dataGroup_hi_lo_1297 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1298;
  assign dataGroup_hi_lo_1298 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1299;
  assign dataGroup_hi_lo_1299 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1300;
  assign dataGroup_hi_lo_1300 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1301;
  assign dataGroup_hi_lo_1301 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1302;
  assign dataGroup_hi_lo_1302 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1303;
  assign dataGroup_hi_lo_1303 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1304;
  assign dataGroup_hi_lo_1304 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1305;
  assign dataGroup_hi_lo_1305 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1306;
  assign dataGroup_hi_lo_1306 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1307;
  assign dataGroup_hi_lo_1307 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1308;
  assign dataGroup_hi_lo_1308 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1309;
  assign dataGroup_hi_lo_1309 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1310;
  assign dataGroup_hi_lo_1310 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1311;
  assign dataGroup_hi_lo_1311 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1312;
  assign dataGroup_hi_lo_1312 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1313;
  assign dataGroup_hi_lo_1313 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1314;
  assign dataGroup_hi_lo_1314 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1315;
  assign dataGroup_hi_lo_1315 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1316;
  assign dataGroup_hi_lo_1316 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1317;
  assign dataGroup_hi_lo_1317 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1318;
  assign dataGroup_hi_lo_1318 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1319;
  assign dataGroup_hi_lo_1319 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1320;
  assign dataGroup_hi_lo_1320 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1321;
  assign dataGroup_hi_lo_1321 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1322;
  assign dataGroup_hi_lo_1322 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1323;
  assign dataGroup_hi_lo_1323 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1324;
  assign dataGroup_hi_lo_1324 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1325;
  assign dataGroup_hi_lo_1325 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1326;
  assign dataGroup_hi_lo_1326 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1327;
  assign dataGroup_hi_lo_1327 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1328;
  assign dataGroup_hi_lo_1328 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1329;
  assign dataGroup_hi_lo_1329 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1330;
  assign dataGroup_hi_lo_1330 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1331;
  assign dataGroup_hi_lo_1331 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1332;
  assign dataGroup_hi_lo_1332 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1333;
  assign dataGroup_hi_lo_1333 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1334;
  assign dataGroup_hi_lo_1334 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1335;
  assign dataGroup_hi_lo_1335 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1336;
  assign dataGroup_hi_lo_1336 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1337;
  assign dataGroup_hi_lo_1337 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1338;
  assign dataGroup_hi_lo_1338 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1339;
  assign dataGroup_hi_lo_1339 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1340;
  assign dataGroup_hi_lo_1340 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1341;
  assign dataGroup_hi_lo_1341 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1342;
  assign dataGroup_hi_lo_1342 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1343;
  assign dataGroup_hi_lo_1343 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1344;
  assign dataGroup_hi_lo_1344 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1345;
  assign dataGroup_hi_lo_1345 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1346;
  assign dataGroup_hi_lo_1346 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1347;
  assign dataGroup_hi_lo_1347 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1348;
  assign dataGroup_hi_lo_1348 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1349;
  assign dataGroup_hi_lo_1349 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1350;
  assign dataGroup_hi_lo_1350 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1351;
  assign dataGroup_hi_lo_1351 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1352;
  assign dataGroup_hi_lo_1352 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1353;
  assign dataGroup_hi_lo_1353 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1354;
  assign dataGroup_hi_lo_1354 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1355;
  assign dataGroup_hi_lo_1355 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1356;
  assign dataGroup_hi_lo_1356 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1357;
  assign dataGroup_hi_lo_1357 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1358;
  assign dataGroup_hi_lo_1358 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1359;
  assign dataGroup_hi_lo_1359 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1360;
  assign dataGroup_hi_lo_1360 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1361;
  assign dataGroup_hi_lo_1361 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1362;
  assign dataGroup_hi_lo_1362 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1363;
  assign dataGroup_hi_lo_1363 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1364;
  assign dataGroup_hi_lo_1364 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1365;
  assign dataGroup_hi_lo_1365 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1366;
  assign dataGroup_hi_lo_1366 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1367;
  assign dataGroup_hi_lo_1367 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1368;
  assign dataGroup_hi_lo_1368 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1369;
  assign dataGroup_hi_lo_1369 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1370;
  assign dataGroup_hi_lo_1370 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1371;
  assign dataGroup_hi_lo_1371 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1372;
  assign dataGroup_hi_lo_1372 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1373;
  assign dataGroup_hi_lo_1373 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1374;
  assign dataGroup_hi_lo_1374 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1375;
  assign dataGroup_hi_lo_1375 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1376;
  assign dataGroup_hi_lo_1376 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1377;
  assign dataGroup_hi_lo_1377 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1378;
  assign dataGroup_hi_lo_1378 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1379;
  assign dataGroup_hi_lo_1379 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1380;
  assign dataGroup_hi_lo_1380 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1381;
  assign dataGroup_hi_lo_1381 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1382;
  assign dataGroup_hi_lo_1382 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1383;
  assign dataGroup_hi_lo_1383 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1384;
  assign dataGroup_hi_lo_1384 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1385;
  assign dataGroup_hi_lo_1385 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1386;
  assign dataGroup_hi_lo_1386 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1387;
  assign dataGroup_hi_lo_1387 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1388;
  assign dataGroup_hi_lo_1388 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1389;
  assign dataGroup_hi_lo_1389 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1390;
  assign dataGroup_hi_lo_1390 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1391;
  assign dataGroup_hi_lo_1391 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1392;
  assign dataGroup_hi_lo_1392 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1393;
  assign dataGroup_hi_lo_1393 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1394;
  assign dataGroup_hi_lo_1394 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1395;
  assign dataGroup_hi_lo_1395 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1396;
  assign dataGroup_hi_lo_1396 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1397;
  assign dataGroup_hi_lo_1397 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1398;
  assign dataGroup_hi_lo_1398 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1399;
  assign dataGroup_hi_lo_1399 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1400;
  assign dataGroup_hi_lo_1400 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1401;
  assign dataGroup_hi_lo_1401 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1402;
  assign dataGroup_hi_lo_1402 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1403;
  assign dataGroup_hi_lo_1403 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1404;
  assign dataGroup_hi_lo_1404 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1405;
  assign dataGroup_hi_lo_1405 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1406;
  assign dataGroup_hi_lo_1406 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1407;
  assign dataGroup_hi_lo_1407 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1408;
  assign dataGroup_hi_lo_1408 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1409;
  assign dataGroup_hi_lo_1409 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1410;
  assign dataGroup_hi_lo_1410 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1411;
  assign dataGroup_hi_lo_1411 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1412;
  assign dataGroup_hi_lo_1412 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1413;
  assign dataGroup_hi_lo_1413 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1414;
  assign dataGroup_hi_lo_1414 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1415;
  assign dataGroup_hi_lo_1415 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1416;
  assign dataGroup_hi_lo_1416 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1417;
  assign dataGroup_hi_lo_1417 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1418;
  assign dataGroup_hi_lo_1418 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1419;
  assign dataGroup_hi_lo_1419 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1420;
  assign dataGroup_hi_lo_1420 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1421;
  assign dataGroup_hi_lo_1421 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1422;
  assign dataGroup_hi_lo_1422 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1423;
  assign dataGroup_hi_lo_1423 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1424;
  assign dataGroup_hi_lo_1424 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1425;
  assign dataGroup_hi_lo_1425 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1426;
  assign dataGroup_hi_lo_1426 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1427;
  assign dataGroup_hi_lo_1427 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1428;
  assign dataGroup_hi_lo_1428 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1429;
  assign dataGroup_hi_lo_1429 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1430;
  assign dataGroup_hi_lo_1430 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1431;
  assign dataGroup_hi_lo_1431 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1432;
  assign dataGroup_hi_lo_1432 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1433;
  assign dataGroup_hi_lo_1433 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1434;
  assign dataGroup_hi_lo_1434 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1435;
  assign dataGroup_hi_lo_1435 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1436;
  assign dataGroup_hi_lo_1436 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1437;
  assign dataGroup_hi_lo_1437 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1438;
  assign dataGroup_hi_lo_1438 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1439;
  assign dataGroup_hi_lo_1439 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1440;
  assign dataGroup_hi_lo_1440 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1441;
  assign dataGroup_hi_lo_1441 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1442;
  assign dataGroup_hi_lo_1442 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1443;
  assign dataGroup_hi_lo_1443 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1444;
  assign dataGroup_hi_lo_1444 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1445;
  assign dataGroup_hi_lo_1445 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1446;
  assign dataGroup_hi_lo_1446 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1447;
  assign dataGroup_hi_lo_1447 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1448;
  assign dataGroup_hi_lo_1448 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1449;
  assign dataGroup_hi_lo_1449 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1450;
  assign dataGroup_hi_lo_1450 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1451;
  assign dataGroup_hi_lo_1451 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1452;
  assign dataGroup_hi_lo_1452 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1453;
  assign dataGroup_hi_lo_1453 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1454;
  assign dataGroup_hi_lo_1454 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1455;
  assign dataGroup_hi_lo_1455 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1456;
  assign dataGroup_hi_lo_1456 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1457;
  assign dataGroup_hi_lo_1457 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1458;
  assign dataGroup_hi_lo_1458 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1459;
  assign dataGroup_hi_lo_1459 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1460;
  assign dataGroup_hi_lo_1460 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1461;
  assign dataGroup_hi_lo_1461 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1462;
  assign dataGroup_hi_lo_1462 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1463;
  assign dataGroup_hi_lo_1463 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1464;
  assign dataGroup_hi_lo_1464 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1465;
  assign dataGroup_hi_lo_1465 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1466;
  assign dataGroup_hi_lo_1466 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1467;
  assign dataGroup_hi_lo_1467 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1468;
  assign dataGroup_hi_lo_1468 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1469;
  assign dataGroup_hi_lo_1469 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1470;
  assign dataGroup_hi_lo_1470 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1471;
  assign dataGroup_hi_lo_1471 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1472;
  assign dataGroup_hi_lo_1472 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1473;
  assign dataGroup_hi_lo_1473 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1474;
  assign dataGroup_hi_lo_1474 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1475;
  assign dataGroup_hi_lo_1475 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1476;
  assign dataGroup_hi_lo_1476 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1477;
  assign dataGroup_hi_lo_1477 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1478;
  assign dataGroup_hi_lo_1478 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1479;
  assign dataGroup_hi_lo_1479 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1480;
  assign dataGroup_hi_lo_1480 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1481;
  assign dataGroup_hi_lo_1481 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1482;
  assign dataGroup_hi_lo_1482 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1483;
  assign dataGroup_hi_lo_1483 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1484;
  assign dataGroup_hi_lo_1484 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1485;
  assign dataGroup_hi_lo_1485 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1486;
  assign dataGroup_hi_lo_1486 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1487;
  assign dataGroup_hi_lo_1487 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1488;
  assign dataGroup_hi_lo_1488 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1489;
  assign dataGroup_hi_lo_1489 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1490;
  assign dataGroup_hi_lo_1490 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1491;
  assign dataGroup_hi_lo_1491 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1492;
  assign dataGroup_hi_lo_1492 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1493;
  assign dataGroup_hi_lo_1493 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1494;
  assign dataGroup_hi_lo_1494 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1495;
  assign dataGroup_hi_lo_1495 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1496;
  assign dataGroup_hi_lo_1496 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1497;
  assign dataGroup_hi_lo_1497 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1498;
  assign dataGroup_hi_lo_1498 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1499;
  assign dataGroup_hi_lo_1499 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1500;
  assign dataGroup_hi_lo_1500 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1501;
  assign dataGroup_hi_lo_1501 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1502;
  assign dataGroup_hi_lo_1502 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1503;
  assign dataGroup_hi_lo_1503 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1504;
  assign dataGroup_hi_lo_1504 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1505;
  assign dataGroup_hi_lo_1505 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1506;
  assign dataGroup_hi_lo_1506 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1507;
  assign dataGroup_hi_lo_1507 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1508;
  assign dataGroup_hi_lo_1508 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1509;
  assign dataGroup_hi_lo_1509 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1510;
  assign dataGroup_hi_lo_1510 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1511;
  assign dataGroup_hi_lo_1511 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1512;
  assign dataGroup_hi_lo_1512 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1513;
  assign dataGroup_hi_lo_1513 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1514;
  assign dataGroup_hi_lo_1514 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1515;
  assign dataGroup_hi_lo_1515 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1516;
  assign dataGroup_hi_lo_1516 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1517;
  assign dataGroup_hi_lo_1517 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1518;
  assign dataGroup_hi_lo_1518 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1519;
  assign dataGroup_hi_lo_1519 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1520;
  assign dataGroup_hi_lo_1520 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1521;
  assign dataGroup_hi_lo_1521 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1522;
  assign dataGroup_hi_lo_1522 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1523;
  assign dataGroup_hi_lo_1523 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1524;
  assign dataGroup_hi_lo_1524 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1525;
  assign dataGroup_hi_lo_1525 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1526;
  assign dataGroup_hi_lo_1526 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1527;
  assign dataGroup_hi_lo_1527 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1528;
  assign dataGroup_hi_lo_1528 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1529;
  assign dataGroup_hi_lo_1529 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1530;
  assign dataGroup_hi_lo_1530 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1531;
  assign dataGroup_hi_lo_1531 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1532;
  assign dataGroup_hi_lo_1532 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1533;
  assign dataGroup_hi_lo_1533 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1534;
  assign dataGroup_hi_lo_1534 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1535;
  assign dataGroup_hi_lo_1535 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1536;
  assign dataGroup_hi_lo_1536 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1537;
  assign dataGroup_hi_lo_1537 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1538;
  assign dataGroup_hi_lo_1538 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1539;
  assign dataGroup_hi_lo_1539 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1540;
  assign dataGroup_hi_lo_1540 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1541;
  assign dataGroup_hi_lo_1541 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1542;
  assign dataGroup_hi_lo_1542 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1543;
  assign dataGroup_hi_lo_1543 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1544;
  assign dataGroup_hi_lo_1544 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1545;
  assign dataGroup_hi_lo_1545 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1546;
  assign dataGroup_hi_lo_1546 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1547;
  assign dataGroup_hi_lo_1547 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1548;
  assign dataGroup_hi_lo_1548 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1549;
  assign dataGroup_hi_lo_1549 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1550;
  assign dataGroup_hi_lo_1550 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1551;
  assign dataGroup_hi_lo_1551 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1552;
  assign dataGroup_hi_lo_1552 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1553;
  assign dataGroup_hi_lo_1553 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1554;
  assign dataGroup_hi_lo_1554 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1555;
  assign dataGroup_hi_lo_1555 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1556;
  assign dataGroup_hi_lo_1556 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1557;
  assign dataGroup_hi_lo_1557 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1558;
  assign dataGroup_hi_lo_1558 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1559;
  assign dataGroup_hi_lo_1559 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1560;
  assign dataGroup_hi_lo_1560 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1561;
  assign dataGroup_hi_lo_1561 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1562;
  assign dataGroup_hi_lo_1562 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1563;
  assign dataGroup_hi_lo_1563 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1564;
  assign dataGroup_hi_lo_1564 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1565;
  assign dataGroup_hi_lo_1565 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1566;
  assign dataGroup_hi_lo_1566 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1567;
  assign dataGroup_hi_lo_1567 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1568;
  assign dataGroup_hi_lo_1568 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1569;
  assign dataGroup_hi_lo_1569 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1570;
  assign dataGroup_hi_lo_1570 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1571;
  assign dataGroup_hi_lo_1571 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1572;
  assign dataGroup_hi_lo_1572 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1573;
  assign dataGroup_hi_lo_1573 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1574;
  assign dataGroup_hi_lo_1574 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1575;
  assign dataGroup_hi_lo_1575 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1576;
  assign dataGroup_hi_lo_1576 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1577;
  assign dataGroup_hi_lo_1577 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1578;
  assign dataGroup_hi_lo_1578 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1579;
  assign dataGroup_hi_lo_1579 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1580;
  assign dataGroup_hi_lo_1580 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1581;
  assign dataGroup_hi_lo_1581 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1582;
  assign dataGroup_hi_lo_1582 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1583;
  assign dataGroup_hi_lo_1583 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1584;
  assign dataGroup_hi_lo_1584 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1585;
  assign dataGroup_hi_lo_1585 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1586;
  assign dataGroup_hi_lo_1586 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1587;
  assign dataGroup_hi_lo_1587 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1588;
  assign dataGroup_hi_lo_1588 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1589;
  assign dataGroup_hi_lo_1589 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1590;
  assign dataGroup_hi_lo_1590 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1591;
  assign dataGroup_hi_lo_1591 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1592;
  assign dataGroup_hi_lo_1592 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1593;
  assign dataGroup_hi_lo_1593 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1594;
  assign dataGroup_hi_lo_1594 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1595;
  assign dataGroup_hi_lo_1595 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1596;
  assign dataGroup_hi_lo_1596 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1597;
  assign dataGroup_hi_lo_1597 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1598;
  assign dataGroup_hi_lo_1598 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1599;
  assign dataGroup_hi_lo_1599 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1600;
  assign dataGroup_hi_lo_1600 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1601;
  assign dataGroup_hi_lo_1601 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1602;
  assign dataGroup_hi_lo_1602 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1603;
  assign dataGroup_hi_lo_1603 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1604;
  assign dataGroup_hi_lo_1604 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1605;
  assign dataGroup_hi_lo_1605 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1606;
  assign dataGroup_hi_lo_1606 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1607;
  assign dataGroup_hi_lo_1607 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1608;
  assign dataGroup_hi_lo_1608 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1609;
  assign dataGroup_hi_lo_1609 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1610;
  assign dataGroup_hi_lo_1610 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1611;
  assign dataGroup_hi_lo_1611 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1612;
  assign dataGroup_hi_lo_1612 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1613;
  assign dataGroup_hi_lo_1613 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1614;
  assign dataGroup_hi_lo_1614 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1615;
  assign dataGroup_hi_lo_1615 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1616;
  assign dataGroup_hi_lo_1616 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1617;
  assign dataGroup_hi_lo_1617 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1618;
  assign dataGroup_hi_lo_1618 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1619;
  assign dataGroup_hi_lo_1619 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1620;
  assign dataGroup_hi_lo_1620 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1621;
  assign dataGroup_hi_lo_1621 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1622;
  assign dataGroup_hi_lo_1622 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1623;
  assign dataGroup_hi_lo_1623 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1624;
  assign dataGroup_hi_lo_1624 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1625;
  assign dataGroup_hi_lo_1625 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1626;
  assign dataGroup_hi_lo_1626 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1627;
  assign dataGroup_hi_lo_1627 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1628;
  assign dataGroup_hi_lo_1628 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1629;
  assign dataGroup_hi_lo_1629 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1630;
  assign dataGroup_hi_lo_1630 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1631;
  assign dataGroup_hi_lo_1631 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1632;
  assign dataGroup_hi_lo_1632 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1633;
  assign dataGroup_hi_lo_1633 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1634;
  assign dataGroup_hi_lo_1634 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1635;
  assign dataGroup_hi_lo_1635 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1636;
  assign dataGroup_hi_lo_1636 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1637;
  assign dataGroup_hi_lo_1637 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1638;
  assign dataGroup_hi_lo_1638 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1639;
  assign dataGroup_hi_lo_1639 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1640;
  assign dataGroup_hi_lo_1640 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1641;
  assign dataGroup_hi_lo_1641 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1642;
  assign dataGroup_hi_lo_1642 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1643;
  assign dataGroup_hi_lo_1643 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1644;
  assign dataGroup_hi_lo_1644 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1645;
  assign dataGroup_hi_lo_1645 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1646;
  assign dataGroup_hi_lo_1646 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1647;
  assign dataGroup_hi_lo_1647 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1648;
  assign dataGroup_hi_lo_1648 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1649;
  assign dataGroup_hi_lo_1649 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1650;
  assign dataGroup_hi_lo_1650 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1651;
  assign dataGroup_hi_lo_1651 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1652;
  assign dataGroup_hi_lo_1652 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1653;
  assign dataGroup_hi_lo_1653 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1654;
  assign dataGroup_hi_lo_1654 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1655;
  assign dataGroup_hi_lo_1655 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1656;
  assign dataGroup_hi_lo_1656 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1657;
  assign dataGroup_hi_lo_1657 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1658;
  assign dataGroup_hi_lo_1658 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1659;
  assign dataGroup_hi_lo_1659 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1660;
  assign dataGroup_hi_lo_1660 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1661;
  assign dataGroup_hi_lo_1661 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1662;
  assign dataGroup_hi_lo_1662 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1663;
  assign dataGroup_hi_lo_1663 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1664;
  assign dataGroup_hi_lo_1664 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1665;
  assign dataGroup_hi_lo_1665 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1666;
  assign dataGroup_hi_lo_1666 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1667;
  assign dataGroup_hi_lo_1667 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1668;
  assign dataGroup_hi_lo_1668 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1669;
  assign dataGroup_hi_lo_1669 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1670;
  assign dataGroup_hi_lo_1670 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1671;
  assign dataGroup_hi_lo_1671 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1672;
  assign dataGroup_hi_lo_1672 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1673;
  assign dataGroup_hi_lo_1673 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1674;
  assign dataGroup_hi_lo_1674 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1675;
  assign dataGroup_hi_lo_1675 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1676;
  assign dataGroup_hi_lo_1676 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1677;
  assign dataGroup_hi_lo_1677 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1678;
  assign dataGroup_hi_lo_1678 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1679;
  assign dataGroup_hi_lo_1679 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1680;
  assign dataGroup_hi_lo_1680 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1681;
  assign dataGroup_hi_lo_1681 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1682;
  assign dataGroup_hi_lo_1682 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1683;
  assign dataGroup_hi_lo_1683 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1684;
  assign dataGroup_hi_lo_1684 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1685;
  assign dataGroup_hi_lo_1685 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1686;
  assign dataGroup_hi_lo_1686 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1687;
  assign dataGroup_hi_lo_1687 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1688;
  assign dataGroup_hi_lo_1688 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1689;
  assign dataGroup_hi_lo_1689 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1690;
  assign dataGroup_hi_lo_1690 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1691;
  assign dataGroup_hi_lo_1691 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1692;
  assign dataGroup_hi_lo_1692 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1693;
  assign dataGroup_hi_lo_1693 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1694;
  assign dataGroup_hi_lo_1694 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1695;
  assign dataGroup_hi_lo_1695 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1696;
  assign dataGroup_hi_lo_1696 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1697;
  assign dataGroup_hi_lo_1697 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1698;
  assign dataGroup_hi_lo_1698 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1699;
  assign dataGroup_hi_lo_1699 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1700;
  assign dataGroup_hi_lo_1700 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1701;
  assign dataGroup_hi_lo_1701 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1702;
  assign dataGroup_hi_lo_1702 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1703;
  assign dataGroup_hi_lo_1703 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1704;
  assign dataGroup_hi_lo_1704 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1705;
  assign dataGroup_hi_lo_1705 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1706;
  assign dataGroup_hi_lo_1706 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1707;
  assign dataGroup_hi_lo_1707 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1708;
  assign dataGroup_hi_lo_1708 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1709;
  assign dataGroup_hi_lo_1709 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1710;
  assign dataGroup_hi_lo_1710 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1711;
  assign dataGroup_hi_lo_1711 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1712;
  assign dataGroup_hi_lo_1712 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1713;
  assign dataGroup_hi_lo_1713 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1714;
  assign dataGroup_hi_lo_1714 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1715;
  assign dataGroup_hi_lo_1715 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1716;
  assign dataGroup_hi_lo_1716 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1717;
  assign dataGroup_hi_lo_1717 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1718;
  assign dataGroup_hi_lo_1718 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1719;
  assign dataGroup_hi_lo_1719 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1720;
  assign dataGroup_hi_lo_1720 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1721;
  assign dataGroup_hi_lo_1721 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1722;
  assign dataGroup_hi_lo_1722 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1723;
  assign dataGroup_hi_lo_1723 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1724;
  assign dataGroup_hi_lo_1724 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1725;
  assign dataGroup_hi_lo_1725 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1726;
  assign dataGroup_hi_lo_1726 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1727;
  assign dataGroup_hi_lo_1727 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1728;
  assign dataGroup_hi_lo_1728 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1729;
  assign dataGroup_hi_lo_1729 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1730;
  assign dataGroup_hi_lo_1730 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1731;
  assign dataGroup_hi_lo_1731 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1732;
  assign dataGroup_hi_lo_1732 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1733;
  assign dataGroup_hi_lo_1733 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1734;
  assign dataGroup_hi_lo_1734 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1735;
  assign dataGroup_hi_lo_1735 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1736;
  assign dataGroup_hi_lo_1736 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1737;
  assign dataGroup_hi_lo_1737 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1738;
  assign dataGroup_hi_lo_1738 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1739;
  assign dataGroup_hi_lo_1739 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1740;
  assign dataGroup_hi_lo_1740 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1741;
  assign dataGroup_hi_lo_1741 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1742;
  assign dataGroup_hi_lo_1742 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1743;
  assign dataGroup_hi_lo_1743 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1744;
  assign dataGroup_hi_lo_1744 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1745;
  assign dataGroup_hi_lo_1745 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1746;
  assign dataGroup_hi_lo_1746 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1747;
  assign dataGroup_hi_lo_1747 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1748;
  assign dataGroup_hi_lo_1748 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1749;
  assign dataGroup_hi_lo_1749 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1750;
  assign dataGroup_hi_lo_1750 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1751;
  assign dataGroup_hi_lo_1751 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1752;
  assign dataGroup_hi_lo_1752 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1753;
  assign dataGroup_hi_lo_1753 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1754;
  assign dataGroup_hi_lo_1754 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1755;
  assign dataGroup_hi_lo_1755 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1756;
  assign dataGroup_hi_lo_1756 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1757;
  assign dataGroup_hi_lo_1757 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1758;
  assign dataGroup_hi_lo_1758 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1759;
  assign dataGroup_hi_lo_1759 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1760;
  assign dataGroup_hi_lo_1760 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1761;
  assign dataGroup_hi_lo_1761 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1762;
  assign dataGroup_hi_lo_1762 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1763;
  assign dataGroup_hi_lo_1763 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1764;
  assign dataGroup_hi_lo_1764 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1765;
  assign dataGroup_hi_lo_1765 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1766;
  assign dataGroup_hi_lo_1766 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1767;
  assign dataGroup_hi_lo_1767 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1768;
  assign dataGroup_hi_lo_1768 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1769;
  assign dataGroup_hi_lo_1769 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1770;
  assign dataGroup_hi_lo_1770 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1771;
  assign dataGroup_hi_lo_1771 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1772;
  assign dataGroup_hi_lo_1772 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1773;
  assign dataGroup_hi_lo_1773 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1774;
  assign dataGroup_hi_lo_1774 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1775;
  assign dataGroup_hi_lo_1775 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1776;
  assign dataGroup_hi_lo_1776 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1777;
  assign dataGroup_hi_lo_1777 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1778;
  assign dataGroup_hi_lo_1778 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1779;
  assign dataGroup_hi_lo_1779 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1780;
  assign dataGroup_hi_lo_1780 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1781;
  assign dataGroup_hi_lo_1781 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1782;
  assign dataGroup_hi_lo_1782 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1783;
  assign dataGroup_hi_lo_1783 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1784;
  assign dataGroup_hi_lo_1784 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1785;
  assign dataGroup_hi_lo_1785 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1786;
  assign dataGroup_hi_lo_1786 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1787;
  assign dataGroup_hi_lo_1787 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1788;
  assign dataGroup_hi_lo_1788 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1789;
  assign dataGroup_hi_lo_1789 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1790;
  assign dataGroup_hi_lo_1790 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1791;
  assign dataGroup_hi_lo_1791 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1792;
  assign dataGroup_hi_lo_1792 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1793;
  assign dataGroup_hi_lo_1793 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1794;
  assign dataGroup_hi_lo_1794 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1795;
  assign dataGroup_hi_lo_1795 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1796;
  assign dataGroup_hi_lo_1796 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1797;
  assign dataGroup_hi_lo_1797 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1798;
  assign dataGroup_hi_lo_1798 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1799;
  assign dataGroup_hi_lo_1799 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1800;
  assign dataGroup_hi_lo_1800 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1801;
  assign dataGroup_hi_lo_1801 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1802;
  assign dataGroup_hi_lo_1802 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1803;
  assign dataGroup_hi_lo_1803 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1804;
  assign dataGroup_hi_lo_1804 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1805;
  assign dataGroup_hi_lo_1805 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1806;
  assign dataGroup_hi_lo_1806 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1807;
  assign dataGroup_hi_lo_1807 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1808;
  assign dataGroup_hi_lo_1808 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1809;
  assign dataGroup_hi_lo_1809 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1810;
  assign dataGroup_hi_lo_1810 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1811;
  assign dataGroup_hi_lo_1811 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1812;
  assign dataGroup_hi_lo_1812 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1813;
  assign dataGroup_hi_lo_1813 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1814;
  assign dataGroup_hi_lo_1814 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1815;
  assign dataGroup_hi_lo_1815 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1816;
  assign dataGroup_hi_lo_1816 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1817;
  assign dataGroup_hi_lo_1817 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1818;
  assign dataGroup_hi_lo_1818 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1819;
  assign dataGroup_hi_lo_1819 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1820;
  assign dataGroup_hi_lo_1820 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1821;
  assign dataGroup_hi_lo_1821 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1822;
  assign dataGroup_hi_lo_1822 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1823;
  assign dataGroup_hi_lo_1823 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1824;
  assign dataGroup_hi_lo_1824 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1825;
  assign dataGroup_hi_lo_1825 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1826;
  assign dataGroup_hi_lo_1826 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1827;
  assign dataGroup_hi_lo_1827 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1828;
  assign dataGroup_hi_lo_1828 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1829;
  assign dataGroup_hi_lo_1829 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1830;
  assign dataGroup_hi_lo_1830 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1831;
  assign dataGroup_hi_lo_1831 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1832;
  assign dataGroup_hi_lo_1832 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1833;
  assign dataGroup_hi_lo_1833 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1834;
  assign dataGroup_hi_lo_1834 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1835;
  assign dataGroup_hi_lo_1835 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1836;
  assign dataGroup_hi_lo_1836 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1837;
  assign dataGroup_hi_lo_1837 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1838;
  assign dataGroup_hi_lo_1838 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1839;
  assign dataGroup_hi_lo_1839 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1840;
  assign dataGroup_hi_lo_1840 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1841;
  assign dataGroup_hi_lo_1841 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1842;
  assign dataGroup_hi_lo_1842 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1843;
  assign dataGroup_hi_lo_1843 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1844;
  assign dataGroup_hi_lo_1844 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1845;
  assign dataGroup_hi_lo_1845 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1846;
  assign dataGroup_hi_lo_1846 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1847;
  assign dataGroup_hi_lo_1847 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1848;
  assign dataGroup_hi_lo_1848 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1849;
  assign dataGroup_hi_lo_1849 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1850;
  assign dataGroup_hi_lo_1850 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1851;
  assign dataGroup_hi_lo_1851 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1852;
  assign dataGroup_hi_lo_1852 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1853;
  assign dataGroup_hi_lo_1853 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1854;
  assign dataGroup_hi_lo_1854 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1855;
  assign dataGroup_hi_lo_1855 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1856;
  assign dataGroup_hi_lo_1856 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1857;
  assign dataGroup_hi_lo_1857 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1858;
  assign dataGroup_hi_lo_1858 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1859;
  assign dataGroup_hi_lo_1859 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1860;
  assign dataGroup_hi_lo_1860 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1861;
  assign dataGroup_hi_lo_1861 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1862;
  assign dataGroup_hi_lo_1862 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1863;
  assign dataGroup_hi_lo_1863 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1864;
  assign dataGroup_hi_lo_1864 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1865;
  assign dataGroup_hi_lo_1865 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1866;
  assign dataGroup_hi_lo_1866 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1867;
  assign dataGroup_hi_lo_1867 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1868;
  assign dataGroup_hi_lo_1868 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1869;
  assign dataGroup_hi_lo_1869 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1870;
  assign dataGroup_hi_lo_1870 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1871;
  assign dataGroup_hi_lo_1871 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1872;
  assign dataGroup_hi_lo_1872 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1873;
  assign dataGroup_hi_lo_1873 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1874;
  assign dataGroup_hi_lo_1874 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1875;
  assign dataGroup_hi_lo_1875 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1876;
  assign dataGroup_hi_lo_1876 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1877;
  assign dataGroup_hi_lo_1877 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1878;
  assign dataGroup_hi_lo_1878 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1879;
  assign dataGroup_hi_lo_1879 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1880;
  assign dataGroup_hi_lo_1880 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1881;
  assign dataGroup_hi_lo_1881 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1882;
  assign dataGroup_hi_lo_1882 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1883;
  assign dataGroup_hi_lo_1883 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1884;
  assign dataGroup_hi_lo_1884 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1885;
  assign dataGroup_hi_lo_1885 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1886;
  assign dataGroup_hi_lo_1886 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1887;
  assign dataGroup_hi_lo_1887 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1888;
  assign dataGroup_hi_lo_1888 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1889;
  assign dataGroup_hi_lo_1889 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1890;
  assign dataGroup_hi_lo_1890 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1891;
  assign dataGroup_hi_lo_1891 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1892;
  assign dataGroup_hi_lo_1892 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1893;
  assign dataGroup_hi_lo_1893 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1894;
  assign dataGroup_hi_lo_1894 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1895;
  assign dataGroup_hi_lo_1895 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1896;
  assign dataGroup_hi_lo_1896 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1897;
  assign dataGroup_hi_lo_1897 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1898;
  assign dataGroup_hi_lo_1898 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1899;
  assign dataGroup_hi_lo_1899 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1900;
  assign dataGroup_hi_lo_1900 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1901;
  assign dataGroup_hi_lo_1901 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1902;
  assign dataGroup_hi_lo_1902 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1903;
  assign dataGroup_hi_lo_1903 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1904;
  assign dataGroup_hi_lo_1904 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1905;
  assign dataGroup_hi_lo_1905 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1906;
  assign dataGroup_hi_lo_1906 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1907;
  assign dataGroup_hi_lo_1907 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1908;
  assign dataGroup_hi_lo_1908 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1909;
  assign dataGroup_hi_lo_1909 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1910;
  assign dataGroup_hi_lo_1910 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1911;
  assign dataGroup_hi_lo_1911 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1912;
  assign dataGroup_hi_lo_1912 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1913;
  assign dataGroup_hi_lo_1913 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1914;
  assign dataGroup_hi_lo_1914 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1915;
  assign dataGroup_hi_lo_1915 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1916;
  assign dataGroup_hi_lo_1916 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1917;
  assign dataGroup_hi_lo_1917 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1918;
  assign dataGroup_hi_lo_1918 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1919;
  assign dataGroup_hi_lo_1919 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1920;
  assign dataGroup_hi_lo_1920 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1921;
  assign dataGroup_hi_lo_1921 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1922;
  assign dataGroup_hi_lo_1922 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1923;
  assign dataGroup_hi_lo_1923 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1924;
  assign dataGroup_hi_lo_1924 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1925;
  assign dataGroup_hi_lo_1925 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1926;
  assign dataGroup_hi_lo_1926 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1927;
  assign dataGroup_hi_lo_1927 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1928;
  assign dataGroup_hi_lo_1928 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1929;
  assign dataGroup_hi_lo_1929 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1930;
  assign dataGroup_hi_lo_1930 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1931;
  assign dataGroup_hi_lo_1931 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1932;
  assign dataGroup_hi_lo_1932 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1933;
  assign dataGroup_hi_lo_1933 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1934;
  assign dataGroup_hi_lo_1934 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1935;
  assign dataGroup_hi_lo_1935 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1936;
  assign dataGroup_hi_lo_1936 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1937;
  assign dataGroup_hi_lo_1937 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1938;
  assign dataGroup_hi_lo_1938 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1939;
  assign dataGroup_hi_lo_1939 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1940;
  assign dataGroup_hi_lo_1940 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1941;
  assign dataGroup_hi_lo_1941 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1942;
  assign dataGroup_hi_lo_1942 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1943;
  assign dataGroup_hi_lo_1943 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1944;
  assign dataGroup_hi_lo_1944 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1945;
  assign dataGroup_hi_lo_1945 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1946;
  assign dataGroup_hi_lo_1946 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1947;
  assign dataGroup_hi_lo_1947 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1948;
  assign dataGroup_hi_lo_1948 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1949;
  assign dataGroup_hi_lo_1949 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1950;
  assign dataGroup_hi_lo_1950 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1951;
  assign dataGroup_hi_lo_1951 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1952;
  assign dataGroup_hi_lo_1952 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1953;
  assign dataGroup_hi_lo_1953 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1954;
  assign dataGroup_hi_lo_1954 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1955;
  assign dataGroup_hi_lo_1955 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1956;
  assign dataGroup_hi_lo_1956 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1957;
  assign dataGroup_hi_lo_1957 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1958;
  assign dataGroup_hi_lo_1958 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1959;
  assign dataGroup_hi_lo_1959 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1960;
  assign dataGroup_hi_lo_1960 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1961;
  assign dataGroup_hi_lo_1961 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1962;
  assign dataGroup_hi_lo_1962 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1963;
  assign dataGroup_hi_lo_1963 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1964;
  assign dataGroup_hi_lo_1964 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1965;
  assign dataGroup_hi_lo_1965 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1966;
  assign dataGroup_hi_lo_1966 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1967;
  assign dataGroup_hi_lo_1967 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1968;
  assign dataGroup_hi_lo_1968 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1969;
  assign dataGroup_hi_lo_1969 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1970;
  assign dataGroup_hi_lo_1970 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1971;
  assign dataGroup_hi_lo_1971 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1972;
  assign dataGroup_hi_lo_1972 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1973;
  assign dataGroup_hi_lo_1973 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1974;
  assign dataGroup_hi_lo_1974 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1975;
  assign dataGroup_hi_lo_1975 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1976;
  assign dataGroup_hi_lo_1976 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1977;
  assign dataGroup_hi_lo_1977 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1978;
  assign dataGroup_hi_lo_1978 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1979;
  assign dataGroup_hi_lo_1979 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1980;
  assign dataGroup_hi_lo_1980 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1981;
  assign dataGroup_hi_lo_1981 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1982;
  assign dataGroup_hi_lo_1982 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1983;
  assign dataGroup_hi_lo_1983 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1984;
  assign dataGroup_hi_lo_1984 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1985;
  assign dataGroup_hi_lo_1985 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1986;
  assign dataGroup_hi_lo_1986 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1987;
  assign dataGroup_hi_lo_1987 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1988;
  assign dataGroup_hi_lo_1988 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1989;
  assign dataGroup_hi_lo_1989 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1990;
  assign dataGroup_hi_lo_1990 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1991;
  assign dataGroup_hi_lo_1991 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1992;
  assign dataGroup_hi_lo_1992 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1993;
  assign dataGroup_hi_lo_1993 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1994;
  assign dataGroup_hi_lo_1994 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1995;
  assign dataGroup_hi_lo_1995 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1996;
  assign dataGroup_hi_lo_1996 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1997;
  assign dataGroup_hi_lo_1997 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1998;
  assign dataGroup_hi_lo_1998 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_1999;
  assign dataGroup_hi_lo_1999 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2000;
  assign dataGroup_hi_lo_2000 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2001;
  assign dataGroup_hi_lo_2001 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2002;
  assign dataGroup_hi_lo_2002 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2003;
  assign dataGroup_hi_lo_2003 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2004;
  assign dataGroup_hi_lo_2004 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2005;
  assign dataGroup_hi_lo_2005 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2006;
  assign dataGroup_hi_lo_2006 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2007;
  assign dataGroup_hi_lo_2007 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2008;
  assign dataGroup_hi_lo_2008 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2009;
  assign dataGroup_hi_lo_2009 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2010;
  assign dataGroup_hi_lo_2010 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2011;
  assign dataGroup_hi_lo_2011 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2012;
  assign dataGroup_hi_lo_2012 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2013;
  assign dataGroup_hi_lo_2013 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2014;
  assign dataGroup_hi_lo_2014 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2015;
  assign dataGroup_hi_lo_2015 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2016;
  assign dataGroup_hi_lo_2016 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2017;
  assign dataGroup_hi_lo_2017 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2018;
  assign dataGroup_hi_lo_2018 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2019;
  assign dataGroup_hi_lo_2019 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2020;
  assign dataGroup_hi_lo_2020 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2021;
  assign dataGroup_hi_lo_2021 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2022;
  assign dataGroup_hi_lo_2022 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2023;
  assign dataGroup_hi_lo_2023 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2024;
  assign dataGroup_hi_lo_2024 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2025;
  assign dataGroup_hi_lo_2025 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2026;
  assign dataGroup_hi_lo_2026 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2027;
  assign dataGroup_hi_lo_2027 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2028;
  assign dataGroup_hi_lo_2028 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2029;
  assign dataGroup_hi_lo_2029 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2030;
  assign dataGroup_hi_lo_2030 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2031;
  assign dataGroup_hi_lo_2031 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2032;
  assign dataGroup_hi_lo_2032 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2033;
  assign dataGroup_hi_lo_2033 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2034;
  assign dataGroup_hi_lo_2034 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2035;
  assign dataGroup_hi_lo_2035 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2036;
  assign dataGroup_hi_lo_2036 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2037;
  assign dataGroup_hi_lo_2037 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2038;
  assign dataGroup_hi_lo_2038 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2039;
  assign dataGroup_hi_lo_2039 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2040;
  assign dataGroup_hi_lo_2040 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2041;
  assign dataGroup_hi_lo_2041 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2042;
  assign dataGroup_hi_lo_2042 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2043;
  assign dataGroup_hi_lo_2043 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2044;
  assign dataGroup_hi_lo_2044 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2045;
  assign dataGroup_hi_lo_2045 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2046;
  assign dataGroup_hi_lo_2046 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2047;
  assign dataGroup_hi_lo_2047 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2048;
  assign dataGroup_hi_lo_2048 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2049;
  assign dataGroup_hi_lo_2049 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2050;
  assign dataGroup_hi_lo_2050 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2051;
  assign dataGroup_hi_lo_2051 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2052;
  assign dataGroup_hi_lo_2052 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2053;
  assign dataGroup_hi_lo_2053 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2054;
  assign dataGroup_hi_lo_2054 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2055;
  assign dataGroup_hi_lo_2055 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2056;
  assign dataGroup_hi_lo_2056 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2057;
  assign dataGroup_hi_lo_2057 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2058;
  assign dataGroup_hi_lo_2058 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2059;
  assign dataGroup_hi_lo_2059 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2060;
  assign dataGroup_hi_lo_2060 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2061;
  assign dataGroup_hi_lo_2061 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2062;
  assign dataGroup_hi_lo_2062 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2063;
  assign dataGroup_hi_lo_2063 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2064;
  assign dataGroup_hi_lo_2064 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2065;
  assign dataGroup_hi_lo_2065 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2066;
  assign dataGroup_hi_lo_2066 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2067;
  assign dataGroup_hi_lo_2067 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2068;
  assign dataGroup_hi_lo_2068 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2069;
  assign dataGroup_hi_lo_2069 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2070;
  assign dataGroup_hi_lo_2070 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2071;
  assign dataGroup_hi_lo_2071 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2072;
  assign dataGroup_hi_lo_2072 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2073;
  assign dataGroup_hi_lo_2073 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2074;
  assign dataGroup_hi_lo_2074 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2075;
  assign dataGroup_hi_lo_2075 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2076;
  assign dataGroup_hi_lo_2076 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2077;
  assign dataGroup_hi_lo_2077 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2078;
  assign dataGroup_hi_lo_2078 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2079;
  assign dataGroup_hi_lo_2079 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2080;
  assign dataGroup_hi_lo_2080 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2081;
  assign dataGroup_hi_lo_2081 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2082;
  assign dataGroup_hi_lo_2082 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2083;
  assign dataGroup_hi_lo_2083 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2084;
  assign dataGroup_hi_lo_2084 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2085;
  assign dataGroup_hi_lo_2085 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2086;
  assign dataGroup_hi_lo_2086 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2087;
  assign dataGroup_hi_lo_2087 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2088;
  assign dataGroup_hi_lo_2088 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2089;
  assign dataGroup_hi_lo_2089 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2090;
  assign dataGroup_hi_lo_2090 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2091;
  assign dataGroup_hi_lo_2091 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2092;
  assign dataGroup_hi_lo_2092 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2093;
  assign dataGroup_hi_lo_2093 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2094;
  assign dataGroup_hi_lo_2094 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2095;
  assign dataGroup_hi_lo_2095 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2096;
  assign dataGroup_hi_lo_2096 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2097;
  assign dataGroup_hi_lo_2097 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2098;
  assign dataGroup_hi_lo_2098 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2099;
  assign dataGroup_hi_lo_2099 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2100;
  assign dataGroup_hi_lo_2100 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2101;
  assign dataGroup_hi_lo_2101 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2102;
  assign dataGroup_hi_lo_2102 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2103;
  assign dataGroup_hi_lo_2103 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2104;
  assign dataGroup_hi_lo_2104 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2105;
  assign dataGroup_hi_lo_2105 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2106;
  assign dataGroup_hi_lo_2106 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2107;
  assign dataGroup_hi_lo_2107 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2108;
  assign dataGroup_hi_lo_2108 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2109;
  assign dataGroup_hi_lo_2109 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2110;
  assign dataGroup_hi_lo_2110 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2111;
  assign dataGroup_hi_lo_2111 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2112;
  assign dataGroup_hi_lo_2112 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2113;
  assign dataGroup_hi_lo_2113 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2114;
  assign dataGroup_hi_lo_2114 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2115;
  assign dataGroup_hi_lo_2115 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2116;
  assign dataGroup_hi_lo_2116 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2117;
  assign dataGroup_hi_lo_2117 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2118;
  assign dataGroup_hi_lo_2118 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2119;
  assign dataGroup_hi_lo_2119 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2120;
  assign dataGroup_hi_lo_2120 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2121;
  assign dataGroup_hi_lo_2121 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2122;
  assign dataGroup_hi_lo_2122 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2123;
  assign dataGroup_hi_lo_2123 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2124;
  assign dataGroup_hi_lo_2124 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2125;
  assign dataGroup_hi_lo_2125 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2126;
  assign dataGroup_hi_lo_2126 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2127;
  assign dataGroup_hi_lo_2127 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2128;
  assign dataGroup_hi_lo_2128 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2129;
  assign dataGroup_hi_lo_2129 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2130;
  assign dataGroup_hi_lo_2130 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2131;
  assign dataGroup_hi_lo_2131 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2132;
  assign dataGroup_hi_lo_2132 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2133;
  assign dataGroup_hi_lo_2133 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2134;
  assign dataGroup_hi_lo_2134 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2135;
  assign dataGroup_hi_lo_2135 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2136;
  assign dataGroup_hi_lo_2136 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2137;
  assign dataGroup_hi_lo_2137 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2138;
  assign dataGroup_hi_lo_2138 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2139;
  assign dataGroup_hi_lo_2139 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2140;
  assign dataGroup_hi_lo_2140 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2141;
  assign dataGroup_hi_lo_2141 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2142;
  assign dataGroup_hi_lo_2142 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2143;
  assign dataGroup_hi_lo_2143 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2144;
  assign dataGroup_hi_lo_2144 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2145;
  assign dataGroup_hi_lo_2145 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2146;
  assign dataGroup_hi_lo_2146 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2147;
  assign dataGroup_hi_lo_2147 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2148;
  assign dataGroup_hi_lo_2148 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2149;
  assign dataGroup_hi_lo_2149 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2150;
  assign dataGroup_hi_lo_2150 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2151;
  assign dataGroup_hi_lo_2151 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2152;
  assign dataGroup_hi_lo_2152 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2153;
  assign dataGroup_hi_lo_2153 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2154;
  assign dataGroup_hi_lo_2154 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2155;
  assign dataGroup_hi_lo_2155 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2156;
  assign dataGroup_hi_lo_2156 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2157;
  assign dataGroup_hi_lo_2157 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2158;
  assign dataGroup_hi_lo_2158 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2159;
  assign dataGroup_hi_lo_2159 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2160;
  assign dataGroup_hi_lo_2160 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2161;
  assign dataGroup_hi_lo_2161 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2162;
  assign dataGroup_hi_lo_2162 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2163;
  assign dataGroup_hi_lo_2163 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2164;
  assign dataGroup_hi_lo_2164 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2165;
  assign dataGroup_hi_lo_2165 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2166;
  assign dataGroup_hi_lo_2166 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2167;
  assign dataGroup_hi_lo_2167 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2168;
  assign dataGroup_hi_lo_2168 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2169;
  assign dataGroup_hi_lo_2169 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2170;
  assign dataGroup_hi_lo_2170 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2171;
  assign dataGroup_hi_lo_2171 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2172;
  assign dataGroup_hi_lo_2172 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2173;
  assign dataGroup_hi_lo_2173 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2174;
  assign dataGroup_hi_lo_2174 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2175;
  assign dataGroup_hi_lo_2175 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2176;
  assign dataGroup_hi_lo_2176 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2177;
  assign dataGroup_hi_lo_2177 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2178;
  assign dataGroup_hi_lo_2178 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2179;
  assign dataGroup_hi_lo_2179 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2180;
  assign dataGroup_hi_lo_2180 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2181;
  assign dataGroup_hi_lo_2181 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2182;
  assign dataGroup_hi_lo_2182 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2183;
  assign dataGroup_hi_lo_2183 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2184;
  assign dataGroup_hi_lo_2184 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2185;
  assign dataGroup_hi_lo_2185 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2186;
  assign dataGroup_hi_lo_2186 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2187;
  assign dataGroup_hi_lo_2187 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2188;
  assign dataGroup_hi_lo_2188 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2189;
  assign dataGroup_hi_lo_2189 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2190;
  assign dataGroup_hi_lo_2190 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2191;
  assign dataGroup_hi_lo_2191 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2192;
  assign dataGroup_hi_lo_2192 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2193;
  assign dataGroup_hi_lo_2193 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2194;
  assign dataGroup_hi_lo_2194 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2195;
  assign dataGroup_hi_lo_2195 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2196;
  assign dataGroup_hi_lo_2196 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2197;
  assign dataGroup_hi_lo_2197 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2198;
  assign dataGroup_hi_lo_2198 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2199;
  assign dataGroup_hi_lo_2199 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2200;
  assign dataGroup_hi_lo_2200 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2201;
  assign dataGroup_hi_lo_2201 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2202;
  assign dataGroup_hi_lo_2202 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2203;
  assign dataGroup_hi_lo_2203 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2204;
  assign dataGroup_hi_lo_2204 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2205;
  assign dataGroup_hi_lo_2205 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2206;
  assign dataGroup_hi_lo_2206 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2207;
  assign dataGroup_hi_lo_2207 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2208;
  assign dataGroup_hi_lo_2208 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2209;
  assign dataGroup_hi_lo_2209 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2210;
  assign dataGroup_hi_lo_2210 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2211;
  assign dataGroup_hi_lo_2211 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2212;
  assign dataGroup_hi_lo_2212 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2213;
  assign dataGroup_hi_lo_2213 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2214;
  assign dataGroup_hi_lo_2214 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2215;
  assign dataGroup_hi_lo_2215 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2216;
  assign dataGroup_hi_lo_2216 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2217;
  assign dataGroup_hi_lo_2217 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2218;
  assign dataGroup_hi_lo_2218 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2219;
  assign dataGroup_hi_lo_2219 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2220;
  assign dataGroup_hi_lo_2220 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2221;
  assign dataGroup_hi_lo_2221 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2222;
  assign dataGroup_hi_lo_2222 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2223;
  assign dataGroup_hi_lo_2223 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2224;
  assign dataGroup_hi_lo_2224 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2225;
  assign dataGroup_hi_lo_2225 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2226;
  assign dataGroup_hi_lo_2226 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2227;
  assign dataGroup_hi_lo_2227 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2228;
  assign dataGroup_hi_lo_2228 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2229;
  assign dataGroup_hi_lo_2229 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2230;
  assign dataGroup_hi_lo_2230 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2231;
  assign dataGroup_hi_lo_2231 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2232;
  assign dataGroup_hi_lo_2232 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2233;
  assign dataGroup_hi_lo_2233 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2234;
  assign dataGroup_hi_lo_2234 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2235;
  assign dataGroup_hi_lo_2235 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2236;
  assign dataGroup_hi_lo_2236 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2237;
  assign dataGroup_hi_lo_2237 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2238;
  assign dataGroup_hi_lo_2238 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2239;
  assign dataGroup_hi_lo_2239 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2240;
  assign dataGroup_hi_lo_2240 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2241;
  assign dataGroup_hi_lo_2241 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2242;
  assign dataGroup_hi_lo_2242 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2243;
  assign dataGroup_hi_lo_2243 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2244;
  assign dataGroup_hi_lo_2244 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2245;
  assign dataGroup_hi_lo_2245 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2246;
  assign dataGroup_hi_lo_2246 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2247;
  assign dataGroup_hi_lo_2247 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2248;
  assign dataGroup_hi_lo_2248 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2249;
  assign dataGroup_hi_lo_2249 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2250;
  assign dataGroup_hi_lo_2250 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2251;
  assign dataGroup_hi_lo_2251 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2252;
  assign dataGroup_hi_lo_2252 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2253;
  assign dataGroup_hi_lo_2253 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2254;
  assign dataGroup_hi_lo_2254 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2255;
  assign dataGroup_hi_lo_2255 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2256;
  assign dataGroup_hi_lo_2256 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2257;
  assign dataGroup_hi_lo_2257 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2258;
  assign dataGroup_hi_lo_2258 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2259;
  assign dataGroup_hi_lo_2259 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2260;
  assign dataGroup_hi_lo_2260 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2261;
  assign dataGroup_hi_lo_2261 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2262;
  assign dataGroup_hi_lo_2262 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2263;
  assign dataGroup_hi_lo_2263 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2264;
  assign dataGroup_hi_lo_2264 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2265;
  assign dataGroup_hi_lo_2265 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2266;
  assign dataGroup_hi_lo_2266 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2267;
  assign dataGroup_hi_lo_2267 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2268;
  assign dataGroup_hi_lo_2268 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2269;
  assign dataGroup_hi_lo_2269 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2270;
  assign dataGroup_hi_lo_2270 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2271;
  assign dataGroup_hi_lo_2271 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2272;
  assign dataGroup_hi_lo_2272 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2273;
  assign dataGroup_hi_lo_2273 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2274;
  assign dataGroup_hi_lo_2274 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2275;
  assign dataGroup_hi_lo_2275 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2276;
  assign dataGroup_hi_lo_2276 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2277;
  assign dataGroup_hi_lo_2277 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2278;
  assign dataGroup_hi_lo_2278 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2279;
  assign dataGroup_hi_lo_2279 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2280;
  assign dataGroup_hi_lo_2280 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2281;
  assign dataGroup_hi_lo_2281 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2282;
  assign dataGroup_hi_lo_2282 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2283;
  assign dataGroup_hi_lo_2283 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2284;
  assign dataGroup_hi_lo_2284 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2285;
  assign dataGroup_hi_lo_2285 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2286;
  assign dataGroup_hi_lo_2286 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2287;
  assign dataGroup_hi_lo_2287 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2288;
  assign dataGroup_hi_lo_2288 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2289;
  assign dataGroup_hi_lo_2289 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2290;
  assign dataGroup_hi_lo_2290 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2291;
  assign dataGroup_hi_lo_2291 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2292;
  assign dataGroup_hi_lo_2292 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2293;
  assign dataGroup_hi_lo_2293 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2294;
  assign dataGroup_hi_lo_2294 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2295;
  assign dataGroup_hi_lo_2295 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2296;
  assign dataGroup_hi_lo_2296 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2297;
  assign dataGroup_hi_lo_2297 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2298;
  assign dataGroup_hi_lo_2298 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2299;
  assign dataGroup_hi_lo_2299 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2300;
  assign dataGroup_hi_lo_2300 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2301;
  assign dataGroup_hi_lo_2301 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2302;
  assign dataGroup_hi_lo_2302 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2303;
  assign dataGroup_hi_lo_2303 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2304;
  assign dataGroup_hi_lo_2304 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2305;
  assign dataGroup_hi_lo_2305 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2306;
  assign dataGroup_hi_lo_2306 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2307;
  assign dataGroup_hi_lo_2307 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2308;
  assign dataGroup_hi_lo_2308 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2309;
  assign dataGroup_hi_lo_2309 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2310;
  assign dataGroup_hi_lo_2310 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2311;
  assign dataGroup_hi_lo_2311 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2312;
  assign dataGroup_hi_lo_2312 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2313;
  assign dataGroup_hi_lo_2313 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2314;
  assign dataGroup_hi_lo_2314 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2315;
  assign dataGroup_hi_lo_2315 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2316;
  assign dataGroup_hi_lo_2316 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2317;
  assign dataGroup_hi_lo_2317 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2318;
  assign dataGroup_hi_lo_2318 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2319;
  assign dataGroup_hi_lo_2319 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2320;
  assign dataGroup_hi_lo_2320 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2321;
  assign dataGroup_hi_lo_2321 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2322;
  assign dataGroup_hi_lo_2322 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2323;
  assign dataGroup_hi_lo_2323 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2324;
  assign dataGroup_hi_lo_2324 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2325;
  assign dataGroup_hi_lo_2325 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2326;
  assign dataGroup_hi_lo_2326 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2327;
  assign dataGroup_hi_lo_2327 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2328;
  assign dataGroup_hi_lo_2328 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2329;
  assign dataGroup_hi_lo_2329 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2330;
  assign dataGroup_hi_lo_2330 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2331;
  assign dataGroup_hi_lo_2331 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2332;
  assign dataGroup_hi_lo_2332 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2333;
  assign dataGroup_hi_lo_2333 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2334;
  assign dataGroup_hi_lo_2334 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2335;
  assign dataGroup_hi_lo_2335 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2336;
  assign dataGroup_hi_lo_2336 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2337;
  assign dataGroup_hi_lo_2337 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2338;
  assign dataGroup_hi_lo_2338 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2339;
  assign dataGroup_hi_lo_2339 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2340;
  assign dataGroup_hi_lo_2340 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2341;
  assign dataGroup_hi_lo_2341 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2342;
  assign dataGroup_hi_lo_2342 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2343;
  assign dataGroup_hi_lo_2343 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2344;
  assign dataGroup_hi_lo_2344 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2345;
  assign dataGroup_hi_lo_2345 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2346;
  assign dataGroup_hi_lo_2346 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2347;
  assign dataGroup_hi_lo_2347 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2348;
  assign dataGroup_hi_lo_2348 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2349;
  assign dataGroup_hi_lo_2349 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2350;
  assign dataGroup_hi_lo_2350 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2351;
  assign dataGroup_hi_lo_2351 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2352;
  assign dataGroup_hi_lo_2352 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2353;
  assign dataGroup_hi_lo_2353 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2354;
  assign dataGroup_hi_lo_2354 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2355;
  assign dataGroup_hi_lo_2355 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2356;
  assign dataGroup_hi_lo_2356 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2357;
  assign dataGroup_hi_lo_2357 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2358;
  assign dataGroup_hi_lo_2358 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2359;
  assign dataGroup_hi_lo_2359 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2360;
  assign dataGroup_hi_lo_2360 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2361;
  assign dataGroup_hi_lo_2361 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2362;
  assign dataGroup_hi_lo_2362 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2363;
  assign dataGroup_hi_lo_2363 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2364;
  assign dataGroup_hi_lo_2364 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2365;
  assign dataGroup_hi_lo_2365 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2366;
  assign dataGroup_hi_lo_2366 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2367;
  assign dataGroup_hi_lo_2367 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2368;
  assign dataGroup_hi_lo_2368 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2369;
  assign dataGroup_hi_lo_2369 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2370;
  assign dataGroup_hi_lo_2370 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2371;
  assign dataGroup_hi_lo_2371 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2372;
  assign dataGroup_hi_lo_2372 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2373;
  assign dataGroup_hi_lo_2373 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2374;
  assign dataGroup_hi_lo_2374 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2375;
  assign dataGroup_hi_lo_2375 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2376;
  assign dataGroup_hi_lo_2376 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2377;
  assign dataGroup_hi_lo_2377 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2378;
  assign dataGroup_hi_lo_2378 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2379;
  assign dataGroup_hi_lo_2379 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2380;
  assign dataGroup_hi_lo_2380 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2381;
  assign dataGroup_hi_lo_2381 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2382;
  assign dataGroup_hi_lo_2382 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2383;
  assign dataGroup_hi_lo_2383 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2384;
  assign dataGroup_hi_lo_2384 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2385;
  assign dataGroup_hi_lo_2385 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2386;
  assign dataGroup_hi_lo_2386 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2387;
  assign dataGroup_hi_lo_2387 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2388;
  assign dataGroup_hi_lo_2388 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2389;
  assign dataGroup_hi_lo_2389 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2390;
  assign dataGroup_hi_lo_2390 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2391;
  assign dataGroup_hi_lo_2391 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2392;
  assign dataGroup_hi_lo_2392 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2393;
  assign dataGroup_hi_lo_2393 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2394;
  assign dataGroup_hi_lo_2394 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2395;
  assign dataGroup_hi_lo_2395 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2396;
  assign dataGroup_hi_lo_2396 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2397;
  assign dataGroup_hi_lo_2397 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2398;
  assign dataGroup_hi_lo_2398 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2399;
  assign dataGroup_hi_lo_2399 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2400;
  assign dataGroup_hi_lo_2400 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2401;
  assign dataGroup_hi_lo_2401 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2402;
  assign dataGroup_hi_lo_2402 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2403;
  assign dataGroup_hi_lo_2403 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2404;
  assign dataGroup_hi_lo_2404 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2405;
  assign dataGroup_hi_lo_2405 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2406;
  assign dataGroup_hi_lo_2406 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2407;
  assign dataGroup_hi_lo_2407 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2408;
  assign dataGroup_hi_lo_2408 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2409;
  assign dataGroup_hi_lo_2409 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2410;
  assign dataGroup_hi_lo_2410 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2411;
  assign dataGroup_hi_lo_2411 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2412;
  assign dataGroup_hi_lo_2412 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2413;
  assign dataGroup_hi_lo_2413 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2414;
  assign dataGroup_hi_lo_2414 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2415;
  assign dataGroup_hi_lo_2415 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2416;
  assign dataGroup_hi_lo_2416 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2417;
  assign dataGroup_hi_lo_2417 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2418;
  assign dataGroup_hi_lo_2418 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2419;
  assign dataGroup_hi_lo_2419 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2420;
  assign dataGroup_hi_lo_2420 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2421;
  assign dataGroup_hi_lo_2421 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2422;
  assign dataGroup_hi_lo_2422 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2423;
  assign dataGroup_hi_lo_2423 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2424;
  assign dataGroup_hi_lo_2424 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2425;
  assign dataGroup_hi_lo_2425 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2426;
  assign dataGroup_hi_lo_2426 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2427;
  assign dataGroup_hi_lo_2427 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2428;
  assign dataGroup_hi_lo_2428 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2429;
  assign dataGroup_hi_lo_2429 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2430;
  assign dataGroup_hi_lo_2430 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2431;
  assign dataGroup_hi_lo_2431 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2432;
  assign dataGroup_hi_lo_2432 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2433;
  assign dataGroup_hi_lo_2433 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2434;
  assign dataGroup_hi_lo_2434 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2435;
  assign dataGroup_hi_lo_2435 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2436;
  assign dataGroup_hi_lo_2436 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2437;
  assign dataGroup_hi_lo_2437 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2438;
  assign dataGroup_hi_lo_2438 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2439;
  assign dataGroup_hi_lo_2439 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2440;
  assign dataGroup_hi_lo_2440 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2441;
  assign dataGroup_hi_lo_2441 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2442;
  assign dataGroup_hi_lo_2442 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2443;
  assign dataGroup_hi_lo_2443 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2444;
  assign dataGroup_hi_lo_2444 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2445;
  assign dataGroup_hi_lo_2445 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2446;
  assign dataGroup_hi_lo_2446 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2447;
  assign dataGroup_hi_lo_2447 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2448;
  assign dataGroup_hi_lo_2448 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2449;
  assign dataGroup_hi_lo_2449 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2450;
  assign dataGroup_hi_lo_2450 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2451;
  assign dataGroup_hi_lo_2451 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2452;
  assign dataGroup_hi_lo_2452 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2453;
  assign dataGroup_hi_lo_2453 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2454;
  assign dataGroup_hi_lo_2454 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2455;
  assign dataGroup_hi_lo_2455 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2456;
  assign dataGroup_hi_lo_2456 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2457;
  assign dataGroup_hi_lo_2457 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2458;
  assign dataGroup_hi_lo_2458 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2459;
  assign dataGroup_hi_lo_2459 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2460;
  assign dataGroup_hi_lo_2460 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2461;
  assign dataGroup_hi_lo_2461 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2462;
  assign dataGroup_hi_lo_2462 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2463;
  assign dataGroup_hi_lo_2463 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2464;
  assign dataGroup_hi_lo_2464 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2465;
  assign dataGroup_hi_lo_2465 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2466;
  assign dataGroup_hi_lo_2466 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2467;
  assign dataGroup_hi_lo_2467 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2468;
  assign dataGroup_hi_lo_2468 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2469;
  assign dataGroup_hi_lo_2469 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2470;
  assign dataGroup_hi_lo_2470 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2471;
  assign dataGroup_hi_lo_2471 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2472;
  assign dataGroup_hi_lo_2472 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2473;
  assign dataGroup_hi_lo_2473 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2474;
  assign dataGroup_hi_lo_2474 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2475;
  assign dataGroup_hi_lo_2475 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2476;
  assign dataGroup_hi_lo_2476 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2477;
  assign dataGroup_hi_lo_2477 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2478;
  assign dataGroup_hi_lo_2478 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2479;
  assign dataGroup_hi_lo_2479 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2480;
  assign dataGroup_hi_lo_2480 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2481;
  assign dataGroup_hi_lo_2481 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2482;
  assign dataGroup_hi_lo_2482 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2483;
  assign dataGroup_hi_lo_2483 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2484;
  assign dataGroup_hi_lo_2484 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2485;
  assign dataGroup_hi_lo_2485 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2486;
  assign dataGroup_hi_lo_2486 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2487;
  assign dataGroup_hi_lo_2487 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2488;
  assign dataGroup_hi_lo_2488 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2489;
  assign dataGroup_hi_lo_2489 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2490;
  assign dataGroup_hi_lo_2490 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2491;
  assign dataGroup_hi_lo_2491 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2492;
  assign dataGroup_hi_lo_2492 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2493;
  assign dataGroup_hi_lo_2493 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2494;
  assign dataGroup_hi_lo_2494 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2495;
  assign dataGroup_hi_lo_2495 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2496;
  assign dataGroup_hi_lo_2496 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2497;
  assign dataGroup_hi_lo_2497 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2498;
  assign dataGroup_hi_lo_2498 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2499;
  assign dataGroup_hi_lo_2499 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2500;
  assign dataGroup_hi_lo_2500 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2501;
  assign dataGroup_hi_lo_2501 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2502;
  assign dataGroup_hi_lo_2502 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2503;
  assign dataGroup_hi_lo_2503 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2504;
  assign dataGroup_hi_lo_2504 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2505;
  assign dataGroup_hi_lo_2505 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2506;
  assign dataGroup_hi_lo_2506 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2507;
  assign dataGroup_hi_lo_2507 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2508;
  assign dataGroup_hi_lo_2508 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2509;
  assign dataGroup_hi_lo_2509 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2510;
  assign dataGroup_hi_lo_2510 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2511;
  assign dataGroup_hi_lo_2511 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2512;
  assign dataGroup_hi_lo_2512 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2513;
  assign dataGroup_hi_lo_2513 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2514;
  assign dataGroup_hi_lo_2514 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2515;
  assign dataGroup_hi_lo_2515 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2516;
  assign dataGroup_hi_lo_2516 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2517;
  assign dataGroup_hi_lo_2517 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2518;
  assign dataGroup_hi_lo_2518 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2519;
  assign dataGroup_hi_lo_2519 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2520;
  assign dataGroup_hi_lo_2520 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2521;
  assign dataGroup_hi_lo_2521 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2522;
  assign dataGroup_hi_lo_2522 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2523;
  assign dataGroup_hi_lo_2523 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2524;
  assign dataGroup_hi_lo_2524 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2525;
  assign dataGroup_hi_lo_2525 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2526;
  assign dataGroup_hi_lo_2526 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2527;
  assign dataGroup_hi_lo_2527 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2528;
  assign dataGroup_hi_lo_2528 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2529;
  assign dataGroup_hi_lo_2529 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2530;
  assign dataGroup_hi_lo_2530 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2531;
  assign dataGroup_hi_lo_2531 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2532;
  assign dataGroup_hi_lo_2532 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2533;
  assign dataGroup_hi_lo_2533 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2534;
  assign dataGroup_hi_lo_2534 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2535;
  assign dataGroup_hi_lo_2535 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2536;
  assign dataGroup_hi_lo_2536 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2537;
  assign dataGroup_hi_lo_2537 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2538;
  assign dataGroup_hi_lo_2538 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2539;
  assign dataGroup_hi_lo_2539 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2540;
  assign dataGroup_hi_lo_2540 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2541;
  assign dataGroup_hi_lo_2541 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2542;
  assign dataGroup_hi_lo_2542 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2543;
  assign dataGroup_hi_lo_2543 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2544;
  assign dataGroup_hi_lo_2544 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2545;
  assign dataGroup_hi_lo_2545 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2546;
  assign dataGroup_hi_lo_2546 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2547;
  assign dataGroup_hi_lo_2547 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2548;
  assign dataGroup_hi_lo_2548 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2549;
  assign dataGroup_hi_lo_2549 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2550;
  assign dataGroup_hi_lo_2550 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2551;
  assign dataGroup_hi_lo_2551 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2552;
  assign dataGroup_hi_lo_2552 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2553;
  assign dataGroup_hi_lo_2553 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2554;
  assign dataGroup_hi_lo_2554 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2555;
  assign dataGroup_hi_lo_2555 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2556;
  assign dataGroup_hi_lo_2556 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2557;
  assign dataGroup_hi_lo_2557 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2558;
  assign dataGroup_hi_lo_2558 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2559;
  assign dataGroup_hi_lo_2559 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2560;
  assign dataGroup_hi_lo_2560 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2561;
  assign dataGroup_hi_lo_2561 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2562;
  assign dataGroup_hi_lo_2562 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2563;
  assign dataGroup_hi_lo_2563 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2564;
  assign dataGroup_hi_lo_2564 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2565;
  assign dataGroup_hi_lo_2565 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2566;
  assign dataGroup_hi_lo_2566 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2567;
  assign dataGroup_hi_lo_2567 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2568;
  assign dataGroup_hi_lo_2568 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2569;
  assign dataGroup_hi_lo_2569 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2570;
  assign dataGroup_hi_lo_2570 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2571;
  assign dataGroup_hi_lo_2571 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2572;
  assign dataGroup_hi_lo_2572 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2573;
  assign dataGroup_hi_lo_2573 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2574;
  assign dataGroup_hi_lo_2574 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2575;
  assign dataGroup_hi_lo_2575 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2576;
  assign dataGroup_hi_lo_2576 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2577;
  assign dataGroup_hi_lo_2577 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2578;
  assign dataGroup_hi_lo_2578 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2579;
  assign dataGroup_hi_lo_2579 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2580;
  assign dataGroup_hi_lo_2580 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2581;
  assign dataGroup_hi_lo_2581 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2582;
  assign dataGroup_hi_lo_2582 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2583;
  assign dataGroup_hi_lo_2583 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2584;
  assign dataGroup_hi_lo_2584 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2585;
  assign dataGroup_hi_lo_2585 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2586;
  assign dataGroup_hi_lo_2586 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2587;
  assign dataGroup_hi_lo_2587 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2588;
  assign dataGroup_hi_lo_2588 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2589;
  assign dataGroup_hi_lo_2589 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2590;
  assign dataGroup_hi_lo_2590 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2591;
  assign dataGroup_hi_lo_2591 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2592;
  assign dataGroup_hi_lo_2592 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2593;
  assign dataGroup_hi_lo_2593 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2594;
  assign dataGroup_hi_lo_2594 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2595;
  assign dataGroup_hi_lo_2595 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2596;
  assign dataGroup_hi_lo_2596 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2597;
  assign dataGroup_hi_lo_2597 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2598;
  assign dataGroup_hi_lo_2598 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2599;
  assign dataGroup_hi_lo_2599 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2600;
  assign dataGroup_hi_lo_2600 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2601;
  assign dataGroup_hi_lo_2601 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2602;
  assign dataGroup_hi_lo_2602 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2603;
  assign dataGroup_hi_lo_2603 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2604;
  assign dataGroup_hi_lo_2604 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2605;
  assign dataGroup_hi_lo_2605 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2606;
  assign dataGroup_hi_lo_2606 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2607;
  assign dataGroup_hi_lo_2607 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2608;
  assign dataGroup_hi_lo_2608 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2609;
  assign dataGroup_hi_lo_2609 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2610;
  assign dataGroup_hi_lo_2610 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2611;
  assign dataGroup_hi_lo_2611 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2612;
  assign dataGroup_hi_lo_2612 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2613;
  assign dataGroup_hi_lo_2613 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2614;
  assign dataGroup_hi_lo_2614 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2615;
  assign dataGroup_hi_lo_2615 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2616;
  assign dataGroup_hi_lo_2616 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2617;
  assign dataGroup_hi_lo_2617 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2618;
  assign dataGroup_hi_lo_2618 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2619;
  assign dataGroup_hi_lo_2619 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2620;
  assign dataGroup_hi_lo_2620 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2621;
  assign dataGroup_hi_lo_2621 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2622;
  assign dataGroup_hi_lo_2622 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2623;
  assign dataGroup_hi_lo_2623 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2624;
  assign dataGroup_hi_lo_2624 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2625;
  assign dataGroup_hi_lo_2625 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2626;
  assign dataGroup_hi_lo_2626 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2627;
  assign dataGroup_hi_lo_2627 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2628;
  assign dataGroup_hi_lo_2628 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2629;
  assign dataGroup_hi_lo_2629 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2630;
  assign dataGroup_hi_lo_2630 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2631;
  assign dataGroup_hi_lo_2631 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2632;
  assign dataGroup_hi_lo_2632 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2633;
  assign dataGroup_hi_lo_2633 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2634;
  assign dataGroup_hi_lo_2634 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2635;
  assign dataGroup_hi_lo_2635 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2636;
  assign dataGroup_hi_lo_2636 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2637;
  assign dataGroup_hi_lo_2637 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2638;
  assign dataGroup_hi_lo_2638 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2639;
  assign dataGroup_hi_lo_2639 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2640;
  assign dataGroup_hi_lo_2640 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2641;
  assign dataGroup_hi_lo_2641 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2642;
  assign dataGroup_hi_lo_2642 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2643;
  assign dataGroup_hi_lo_2643 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2644;
  assign dataGroup_hi_lo_2644 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2645;
  assign dataGroup_hi_lo_2645 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2646;
  assign dataGroup_hi_lo_2646 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2647;
  assign dataGroup_hi_lo_2647 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2648;
  assign dataGroup_hi_lo_2648 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2649;
  assign dataGroup_hi_lo_2649 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2650;
  assign dataGroup_hi_lo_2650 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2651;
  assign dataGroup_hi_lo_2651 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2652;
  assign dataGroup_hi_lo_2652 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2653;
  assign dataGroup_hi_lo_2653 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2654;
  assign dataGroup_hi_lo_2654 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2655;
  assign dataGroup_hi_lo_2655 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2656;
  assign dataGroup_hi_lo_2656 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2657;
  assign dataGroup_hi_lo_2657 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2658;
  assign dataGroup_hi_lo_2658 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2659;
  assign dataGroup_hi_lo_2659 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2660;
  assign dataGroup_hi_lo_2660 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2661;
  assign dataGroup_hi_lo_2661 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2662;
  assign dataGroup_hi_lo_2662 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2663;
  assign dataGroup_hi_lo_2663 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2664;
  assign dataGroup_hi_lo_2664 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2665;
  assign dataGroup_hi_lo_2665 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2666;
  assign dataGroup_hi_lo_2666 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2667;
  assign dataGroup_hi_lo_2667 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2668;
  assign dataGroup_hi_lo_2668 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2669;
  assign dataGroup_hi_lo_2669 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2670;
  assign dataGroup_hi_lo_2670 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2671;
  assign dataGroup_hi_lo_2671 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2672;
  assign dataGroup_hi_lo_2672 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2673;
  assign dataGroup_hi_lo_2673 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2674;
  assign dataGroup_hi_lo_2674 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2675;
  assign dataGroup_hi_lo_2675 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2676;
  assign dataGroup_hi_lo_2676 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2677;
  assign dataGroup_hi_lo_2677 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2678;
  assign dataGroup_hi_lo_2678 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2679;
  assign dataGroup_hi_lo_2679 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2680;
  assign dataGroup_hi_lo_2680 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2681;
  assign dataGroup_hi_lo_2681 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2682;
  assign dataGroup_hi_lo_2682 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2683;
  assign dataGroup_hi_lo_2683 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2684;
  assign dataGroup_hi_lo_2684 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2685;
  assign dataGroup_hi_lo_2685 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2686;
  assign dataGroup_hi_lo_2686 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2687;
  assign dataGroup_hi_lo_2687 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2688;
  assign dataGroup_hi_lo_2688 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2689;
  assign dataGroup_hi_lo_2689 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2690;
  assign dataGroup_hi_lo_2690 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2691;
  assign dataGroup_hi_lo_2691 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2692;
  assign dataGroup_hi_lo_2692 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2693;
  assign dataGroup_hi_lo_2693 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2694;
  assign dataGroup_hi_lo_2694 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2695;
  assign dataGroup_hi_lo_2695 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2696;
  assign dataGroup_hi_lo_2696 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2697;
  assign dataGroup_hi_lo_2697 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2698;
  assign dataGroup_hi_lo_2698 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2699;
  assign dataGroup_hi_lo_2699 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2700;
  assign dataGroup_hi_lo_2700 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2701;
  assign dataGroup_hi_lo_2701 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2702;
  assign dataGroup_hi_lo_2702 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2703;
  assign dataGroup_hi_lo_2703 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2704;
  assign dataGroup_hi_lo_2704 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2705;
  assign dataGroup_hi_lo_2705 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2706;
  assign dataGroup_hi_lo_2706 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2707;
  assign dataGroup_hi_lo_2707 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2708;
  assign dataGroup_hi_lo_2708 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2709;
  assign dataGroup_hi_lo_2709 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2710;
  assign dataGroup_hi_lo_2710 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2711;
  assign dataGroup_hi_lo_2711 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2712;
  assign dataGroup_hi_lo_2712 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2713;
  assign dataGroup_hi_lo_2713 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2714;
  assign dataGroup_hi_lo_2714 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2715;
  assign dataGroup_hi_lo_2715 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2716;
  assign dataGroup_hi_lo_2716 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2717;
  assign dataGroup_hi_lo_2717 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2718;
  assign dataGroup_hi_lo_2718 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2719;
  assign dataGroup_hi_lo_2719 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2720;
  assign dataGroup_hi_lo_2720 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2721;
  assign dataGroup_hi_lo_2721 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2722;
  assign dataGroup_hi_lo_2722 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2723;
  assign dataGroup_hi_lo_2723 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2724;
  assign dataGroup_hi_lo_2724 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2725;
  assign dataGroup_hi_lo_2725 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2726;
  assign dataGroup_hi_lo_2726 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2727;
  assign dataGroup_hi_lo_2727 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2728;
  assign dataGroup_hi_lo_2728 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2729;
  assign dataGroup_hi_lo_2729 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2730;
  assign dataGroup_hi_lo_2730 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2731;
  assign dataGroup_hi_lo_2731 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2732;
  assign dataGroup_hi_lo_2732 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2733;
  assign dataGroup_hi_lo_2733 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2734;
  assign dataGroup_hi_lo_2734 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2735;
  assign dataGroup_hi_lo_2735 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2736;
  assign dataGroup_hi_lo_2736 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2737;
  assign dataGroup_hi_lo_2737 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2738;
  assign dataGroup_hi_lo_2738 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2739;
  assign dataGroup_hi_lo_2739 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2740;
  assign dataGroup_hi_lo_2740 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2741;
  assign dataGroup_hi_lo_2741 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2742;
  assign dataGroup_hi_lo_2742 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2743;
  assign dataGroup_hi_lo_2743 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2744;
  assign dataGroup_hi_lo_2744 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2745;
  assign dataGroup_hi_lo_2745 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2746;
  assign dataGroup_hi_lo_2746 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2747;
  assign dataGroup_hi_lo_2747 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2748;
  assign dataGroup_hi_lo_2748 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2749;
  assign dataGroup_hi_lo_2749 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2750;
  assign dataGroup_hi_lo_2750 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2751;
  assign dataGroup_hi_lo_2751 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2752;
  assign dataGroup_hi_lo_2752 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2753;
  assign dataGroup_hi_lo_2753 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2754;
  assign dataGroup_hi_lo_2754 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2755;
  assign dataGroup_hi_lo_2755 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2756;
  assign dataGroup_hi_lo_2756 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2757;
  assign dataGroup_hi_lo_2757 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2758;
  assign dataGroup_hi_lo_2758 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2759;
  assign dataGroup_hi_lo_2759 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2760;
  assign dataGroup_hi_lo_2760 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2761;
  assign dataGroup_hi_lo_2761 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2762;
  assign dataGroup_hi_lo_2762 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2763;
  assign dataGroup_hi_lo_2763 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2764;
  assign dataGroup_hi_lo_2764 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2765;
  assign dataGroup_hi_lo_2765 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2766;
  assign dataGroup_hi_lo_2766 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2767;
  assign dataGroup_hi_lo_2767 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2768;
  assign dataGroup_hi_lo_2768 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2769;
  assign dataGroup_hi_lo_2769 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2770;
  assign dataGroup_hi_lo_2770 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2771;
  assign dataGroup_hi_lo_2771 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2772;
  assign dataGroup_hi_lo_2772 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2773;
  assign dataGroup_hi_lo_2773 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2774;
  assign dataGroup_hi_lo_2774 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2775;
  assign dataGroup_hi_lo_2775 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2776;
  assign dataGroup_hi_lo_2776 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2777;
  assign dataGroup_hi_lo_2777 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2778;
  assign dataGroup_hi_lo_2778 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2779;
  assign dataGroup_hi_lo_2779 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2780;
  assign dataGroup_hi_lo_2780 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2781;
  assign dataGroup_hi_lo_2781 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2782;
  assign dataGroup_hi_lo_2782 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2783;
  assign dataGroup_hi_lo_2783 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2784;
  assign dataGroup_hi_lo_2784 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2785;
  assign dataGroup_hi_lo_2785 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2786;
  assign dataGroup_hi_lo_2786 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2787;
  assign dataGroup_hi_lo_2787 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2788;
  assign dataGroup_hi_lo_2788 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2789;
  assign dataGroup_hi_lo_2789 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2790;
  assign dataGroup_hi_lo_2790 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2791;
  assign dataGroup_hi_lo_2791 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2792;
  assign dataGroup_hi_lo_2792 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2793;
  assign dataGroup_hi_lo_2793 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2794;
  assign dataGroup_hi_lo_2794 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2795;
  assign dataGroup_hi_lo_2795 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2796;
  assign dataGroup_hi_lo_2796 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2797;
  assign dataGroup_hi_lo_2797 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2798;
  assign dataGroup_hi_lo_2798 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2799;
  assign dataGroup_hi_lo_2799 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2800;
  assign dataGroup_hi_lo_2800 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2801;
  assign dataGroup_hi_lo_2801 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2802;
  assign dataGroup_hi_lo_2802 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2803;
  assign dataGroup_hi_lo_2803 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2804;
  assign dataGroup_hi_lo_2804 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2805;
  assign dataGroup_hi_lo_2805 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2806;
  assign dataGroup_hi_lo_2806 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2807;
  assign dataGroup_hi_lo_2807 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2808;
  assign dataGroup_hi_lo_2808 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2809;
  assign dataGroup_hi_lo_2809 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2810;
  assign dataGroup_hi_lo_2810 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2811;
  assign dataGroup_hi_lo_2811 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2812;
  assign dataGroup_hi_lo_2812 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2813;
  assign dataGroup_hi_lo_2813 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2814;
  assign dataGroup_hi_lo_2814 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2815;
  assign dataGroup_hi_lo_2815 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2816;
  assign dataGroup_hi_lo_2816 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2817;
  assign dataGroup_hi_lo_2817 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2818;
  assign dataGroup_hi_lo_2818 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2819;
  assign dataGroup_hi_lo_2819 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2820;
  assign dataGroup_hi_lo_2820 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2821;
  assign dataGroup_hi_lo_2821 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2822;
  assign dataGroup_hi_lo_2822 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2823;
  assign dataGroup_hi_lo_2823 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2824;
  assign dataGroup_hi_lo_2824 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2825;
  assign dataGroup_hi_lo_2825 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2826;
  assign dataGroup_hi_lo_2826 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2827;
  assign dataGroup_hi_lo_2827 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2828;
  assign dataGroup_hi_lo_2828 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2829;
  assign dataGroup_hi_lo_2829 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2830;
  assign dataGroup_hi_lo_2830 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2831;
  assign dataGroup_hi_lo_2831 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2832;
  assign dataGroup_hi_lo_2832 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2833;
  assign dataGroup_hi_lo_2833 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2834;
  assign dataGroup_hi_lo_2834 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2835;
  assign dataGroup_hi_lo_2835 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2836;
  assign dataGroup_hi_lo_2836 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2837;
  assign dataGroup_hi_lo_2837 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2838;
  assign dataGroup_hi_lo_2838 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2839;
  assign dataGroup_hi_lo_2839 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2840;
  assign dataGroup_hi_lo_2840 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2841;
  assign dataGroup_hi_lo_2841 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2842;
  assign dataGroup_hi_lo_2842 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2843;
  assign dataGroup_hi_lo_2843 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2844;
  assign dataGroup_hi_lo_2844 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2845;
  assign dataGroup_hi_lo_2845 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2846;
  assign dataGroup_hi_lo_2846 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2847;
  assign dataGroup_hi_lo_2847 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2848;
  assign dataGroup_hi_lo_2848 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2849;
  assign dataGroup_hi_lo_2849 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2850;
  assign dataGroup_hi_lo_2850 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2851;
  assign dataGroup_hi_lo_2851 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2852;
  assign dataGroup_hi_lo_2852 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2853;
  assign dataGroup_hi_lo_2853 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2854;
  assign dataGroup_hi_lo_2854 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2855;
  assign dataGroup_hi_lo_2855 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2856;
  assign dataGroup_hi_lo_2856 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2857;
  assign dataGroup_hi_lo_2857 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2858;
  assign dataGroup_hi_lo_2858 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2859;
  assign dataGroup_hi_lo_2859 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2860;
  assign dataGroup_hi_lo_2860 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2861;
  assign dataGroup_hi_lo_2861 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2862;
  assign dataGroup_hi_lo_2862 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2863;
  assign dataGroup_hi_lo_2863 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2864;
  assign dataGroup_hi_lo_2864 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2865;
  assign dataGroup_hi_lo_2865 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2866;
  assign dataGroup_hi_lo_2866 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2867;
  assign dataGroup_hi_lo_2867 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2868;
  assign dataGroup_hi_lo_2868 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2869;
  assign dataGroup_hi_lo_2869 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2870;
  assign dataGroup_hi_lo_2870 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2871;
  assign dataGroup_hi_lo_2871 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2872;
  assign dataGroup_hi_lo_2872 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2873;
  assign dataGroup_hi_lo_2873 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2874;
  assign dataGroup_hi_lo_2874 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2875;
  assign dataGroup_hi_lo_2875 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2876;
  assign dataGroup_hi_lo_2876 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2877;
  assign dataGroup_hi_lo_2877 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2878;
  assign dataGroup_hi_lo_2878 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2879;
  assign dataGroup_hi_lo_2879 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2880;
  assign dataGroup_hi_lo_2880 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2881;
  assign dataGroup_hi_lo_2881 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2882;
  assign dataGroup_hi_lo_2882 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2883;
  assign dataGroup_hi_lo_2883 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2884;
  assign dataGroup_hi_lo_2884 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2885;
  assign dataGroup_hi_lo_2885 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2886;
  assign dataGroup_hi_lo_2886 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2887;
  assign dataGroup_hi_lo_2887 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2888;
  assign dataGroup_hi_lo_2888 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2889;
  assign dataGroup_hi_lo_2889 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2890;
  assign dataGroup_hi_lo_2890 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2891;
  assign dataGroup_hi_lo_2891 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2892;
  assign dataGroup_hi_lo_2892 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2893;
  assign dataGroup_hi_lo_2893 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2894;
  assign dataGroup_hi_lo_2894 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2895;
  assign dataGroup_hi_lo_2895 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2896;
  assign dataGroup_hi_lo_2896 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2897;
  assign dataGroup_hi_lo_2897 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2898;
  assign dataGroup_hi_lo_2898 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2899;
  assign dataGroup_hi_lo_2899 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2900;
  assign dataGroup_hi_lo_2900 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2901;
  assign dataGroup_hi_lo_2901 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2902;
  assign dataGroup_hi_lo_2902 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2903;
  assign dataGroup_hi_lo_2903 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2904;
  assign dataGroup_hi_lo_2904 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2905;
  assign dataGroup_hi_lo_2905 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2906;
  assign dataGroup_hi_lo_2906 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2907;
  assign dataGroup_hi_lo_2907 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2908;
  assign dataGroup_hi_lo_2908 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2909;
  assign dataGroup_hi_lo_2909 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2910;
  assign dataGroup_hi_lo_2910 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2911;
  assign dataGroup_hi_lo_2911 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2912;
  assign dataGroup_hi_lo_2912 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2913;
  assign dataGroup_hi_lo_2913 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2914;
  assign dataGroup_hi_lo_2914 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2915;
  assign dataGroup_hi_lo_2915 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2916;
  assign dataGroup_hi_lo_2916 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2917;
  assign dataGroup_hi_lo_2917 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2918;
  assign dataGroup_hi_lo_2918 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2919;
  assign dataGroup_hi_lo_2919 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2920;
  assign dataGroup_hi_lo_2920 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2921;
  assign dataGroup_hi_lo_2921 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2922;
  assign dataGroup_hi_lo_2922 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2923;
  assign dataGroup_hi_lo_2923 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2924;
  assign dataGroup_hi_lo_2924 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2925;
  assign dataGroup_hi_lo_2925 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2926;
  assign dataGroup_hi_lo_2926 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2927;
  assign dataGroup_hi_lo_2927 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2928;
  assign dataGroup_hi_lo_2928 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2929;
  assign dataGroup_hi_lo_2929 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2930;
  assign dataGroup_hi_lo_2930 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2931;
  assign dataGroup_hi_lo_2931 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2932;
  assign dataGroup_hi_lo_2932 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2933;
  assign dataGroup_hi_lo_2933 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2934;
  assign dataGroup_hi_lo_2934 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2935;
  assign dataGroup_hi_lo_2935 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2936;
  assign dataGroup_hi_lo_2936 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2937;
  assign dataGroup_hi_lo_2937 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2938;
  assign dataGroup_hi_lo_2938 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2939;
  assign dataGroup_hi_lo_2939 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2940;
  assign dataGroup_hi_lo_2940 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2941;
  assign dataGroup_hi_lo_2941 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2942;
  assign dataGroup_hi_lo_2942 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2943;
  assign dataGroup_hi_lo_2943 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2944;
  assign dataGroup_hi_lo_2944 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2945;
  assign dataGroup_hi_lo_2945 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2946;
  assign dataGroup_hi_lo_2946 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2947;
  assign dataGroup_hi_lo_2947 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2948;
  assign dataGroup_hi_lo_2948 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2949;
  assign dataGroup_hi_lo_2949 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2950;
  assign dataGroup_hi_lo_2950 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2951;
  assign dataGroup_hi_lo_2951 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2952;
  assign dataGroup_hi_lo_2952 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2953;
  assign dataGroup_hi_lo_2953 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2954;
  assign dataGroup_hi_lo_2954 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2955;
  assign dataGroup_hi_lo_2955 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2956;
  assign dataGroup_hi_lo_2956 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2957;
  assign dataGroup_hi_lo_2957 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2958;
  assign dataGroup_hi_lo_2958 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2959;
  assign dataGroup_hi_lo_2959 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2960;
  assign dataGroup_hi_lo_2960 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2961;
  assign dataGroup_hi_lo_2961 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2962;
  assign dataGroup_hi_lo_2962 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2963;
  assign dataGroup_hi_lo_2963 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2964;
  assign dataGroup_hi_lo_2964 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2965;
  assign dataGroup_hi_lo_2965 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2966;
  assign dataGroup_hi_lo_2966 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2967;
  assign dataGroup_hi_lo_2967 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2968;
  assign dataGroup_hi_lo_2968 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2969;
  assign dataGroup_hi_lo_2969 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2970;
  assign dataGroup_hi_lo_2970 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2971;
  assign dataGroup_hi_lo_2971 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2972;
  assign dataGroup_hi_lo_2972 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2973;
  assign dataGroup_hi_lo_2973 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2974;
  assign dataGroup_hi_lo_2974 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2975;
  assign dataGroup_hi_lo_2975 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2976;
  assign dataGroup_hi_lo_2976 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2977;
  assign dataGroup_hi_lo_2977 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2978;
  assign dataGroup_hi_lo_2978 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2979;
  assign dataGroup_hi_lo_2979 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2980;
  assign dataGroup_hi_lo_2980 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2981;
  assign dataGroup_hi_lo_2981 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2982;
  assign dataGroup_hi_lo_2982 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2983;
  assign dataGroup_hi_lo_2983 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2984;
  assign dataGroup_hi_lo_2984 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2985;
  assign dataGroup_hi_lo_2985 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2986;
  assign dataGroup_hi_lo_2986 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2987;
  assign dataGroup_hi_lo_2987 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2988;
  assign dataGroup_hi_lo_2988 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2989;
  assign dataGroup_hi_lo_2989 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2990;
  assign dataGroup_hi_lo_2990 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2991;
  assign dataGroup_hi_lo_2991 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2992;
  assign dataGroup_hi_lo_2992 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2993;
  assign dataGroup_hi_lo_2993 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2994;
  assign dataGroup_hi_lo_2994 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2995;
  assign dataGroup_hi_lo_2995 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2996;
  assign dataGroup_hi_lo_2996 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2997;
  assign dataGroup_hi_lo_2997 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2998;
  assign dataGroup_hi_lo_2998 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_2999;
  assign dataGroup_hi_lo_2999 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3000;
  assign dataGroup_hi_lo_3000 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3001;
  assign dataGroup_hi_lo_3001 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3002;
  assign dataGroup_hi_lo_3002 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3003;
  assign dataGroup_hi_lo_3003 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3004;
  assign dataGroup_hi_lo_3004 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3005;
  assign dataGroup_hi_lo_3005 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3006;
  assign dataGroup_hi_lo_3006 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3007;
  assign dataGroup_hi_lo_3007 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3008;
  assign dataGroup_hi_lo_3008 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3009;
  assign dataGroup_hi_lo_3009 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3010;
  assign dataGroup_hi_lo_3010 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3011;
  assign dataGroup_hi_lo_3011 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3012;
  assign dataGroup_hi_lo_3012 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3013;
  assign dataGroup_hi_lo_3013 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3014;
  assign dataGroup_hi_lo_3014 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3015;
  assign dataGroup_hi_lo_3015 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3016;
  assign dataGroup_hi_lo_3016 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3017;
  assign dataGroup_hi_lo_3017 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3018;
  assign dataGroup_hi_lo_3018 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3019;
  assign dataGroup_hi_lo_3019 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3020;
  assign dataGroup_hi_lo_3020 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3021;
  assign dataGroup_hi_lo_3021 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3022;
  assign dataGroup_hi_lo_3022 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3023;
  assign dataGroup_hi_lo_3023 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3024;
  assign dataGroup_hi_lo_3024 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3025;
  assign dataGroup_hi_lo_3025 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3026;
  assign dataGroup_hi_lo_3026 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3027;
  assign dataGroup_hi_lo_3027 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3028;
  assign dataGroup_hi_lo_3028 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3029;
  assign dataGroup_hi_lo_3029 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3030;
  assign dataGroup_hi_lo_3030 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3031;
  assign dataGroup_hi_lo_3031 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3032;
  assign dataGroup_hi_lo_3032 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3033;
  assign dataGroup_hi_lo_3033 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3034;
  assign dataGroup_hi_lo_3034 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3035;
  assign dataGroup_hi_lo_3035 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3036;
  assign dataGroup_hi_lo_3036 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3037;
  assign dataGroup_hi_lo_3037 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3038;
  assign dataGroup_hi_lo_3038 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3039;
  assign dataGroup_hi_lo_3039 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3040;
  assign dataGroup_hi_lo_3040 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3041;
  assign dataGroup_hi_lo_3041 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3042;
  assign dataGroup_hi_lo_3042 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3043;
  assign dataGroup_hi_lo_3043 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3044;
  assign dataGroup_hi_lo_3044 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3045;
  assign dataGroup_hi_lo_3045 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3046;
  assign dataGroup_hi_lo_3046 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3047;
  assign dataGroup_hi_lo_3047 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3048;
  assign dataGroup_hi_lo_3048 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3049;
  assign dataGroup_hi_lo_3049 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3050;
  assign dataGroup_hi_lo_3050 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3051;
  assign dataGroup_hi_lo_3051 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3052;
  assign dataGroup_hi_lo_3052 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3053;
  assign dataGroup_hi_lo_3053 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3054;
  assign dataGroup_hi_lo_3054 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3055;
  assign dataGroup_hi_lo_3055 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3056;
  assign dataGroup_hi_lo_3056 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3057;
  assign dataGroup_hi_lo_3057 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3058;
  assign dataGroup_hi_lo_3058 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3059;
  assign dataGroup_hi_lo_3059 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3060;
  assign dataGroup_hi_lo_3060 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3061;
  assign dataGroup_hi_lo_3061 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3062;
  assign dataGroup_hi_lo_3062 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3063;
  assign dataGroup_hi_lo_3063 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3064;
  assign dataGroup_hi_lo_3064 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3065;
  assign dataGroup_hi_lo_3065 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3066;
  assign dataGroup_hi_lo_3066 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3067;
  assign dataGroup_hi_lo_3067 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3068;
  assign dataGroup_hi_lo_3068 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3069;
  assign dataGroup_hi_lo_3069 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3070;
  assign dataGroup_hi_lo_3070 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3071;
  assign dataGroup_hi_lo_3071 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3072;
  assign dataGroup_hi_lo_3072 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3073;
  assign dataGroup_hi_lo_3073 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3074;
  assign dataGroup_hi_lo_3074 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3075;
  assign dataGroup_hi_lo_3075 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3076;
  assign dataGroup_hi_lo_3076 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3077;
  assign dataGroup_hi_lo_3077 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3078;
  assign dataGroup_hi_lo_3078 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3079;
  assign dataGroup_hi_lo_3079 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3080;
  assign dataGroup_hi_lo_3080 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3081;
  assign dataGroup_hi_lo_3081 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3082;
  assign dataGroup_hi_lo_3082 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3083;
  assign dataGroup_hi_lo_3083 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3084;
  assign dataGroup_hi_lo_3084 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3085;
  assign dataGroup_hi_lo_3085 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3086;
  assign dataGroup_hi_lo_3086 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3087;
  assign dataGroup_hi_lo_3087 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3088;
  assign dataGroup_hi_lo_3088 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3089;
  assign dataGroup_hi_lo_3089 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3090;
  assign dataGroup_hi_lo_3090 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3091;
  assign dataGroup_hi_lo_3091 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3092;
  assign dataGroup_hi_lo_3092 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3093;
  assign dataGroup_hi_lo_3093 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3094;
  assign dataGroup_hi_lo_3094 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3095;
  assign dataGroup_hi_lo_3095 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3096;
  assign dataGroup_hi_lo_3096 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3097;
  assign dataGroup_hi_lo_3097 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3098;
  assign dataGroup_hi_lo_3098 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3099;
  assign dataGroup_hi_lo_3099 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3100;
  assign dataGroup_hi_lo_3100 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3101;
  assign dataGroup_hi_lo_3101 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3102;
  assign dataGroup_hi_lo_3102 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3103;
  assign dataGroup_hi_lo_3103 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3104;
  assign dataGroup_hi_lo_3104 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3105;
  assign dataGroup_hi_lo_3105 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3106;
  assign dataGroup_hi_lo_3106 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3107;
  assign dataGroup_hi_lo_3107 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3108;
  assign dataGroup_hi_lo_3108 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3109;
  assign dataGroup_hi_lo_3109 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3110;
  assign dataGroup_hi_lo_3110 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3111;
  assign dataGroup_hi_lo_3111 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3112;
  assign dataGroup_hi_lo_3112 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3113;
  assign dataGroup_hi_lo_3113 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3114;
  assign dataGroup_hi_lo_3114 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3115;
  assign dataGroup_hi_lo_3115 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3116;
  assign dataGroup_hi_lo_3116 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3117;
  assign dataGroup_hi_lo_3117 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3118;
  assign dataGroup_hi_lo_3118 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3119;
  assign dataGroup_hi_lo_3119 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3120;
  assign dataGroup_hi_lo_3120 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3121;
  assign dataGroup_hi_lo_3121 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3122;
  assign dataGroup_hi_lo_3122 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3123;
  assign dataGroup_hi_lo_3123 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3124;
  assign dataGroup_hi_lo_3124 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3125;
  assign dataGroup_hi_lo_3125 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3126;
  assign dataGroup_hi_lo_3126 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3127;
  assign dataGroup_hi_lo_3127 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3128;
  assign dataGroup_hi_lo_3128 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3129;
  assign dataGroup_hi_lo_3129 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3130;
  assign dataGroup_hi_lo_3130 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3131;
  assign dataGroup_hi_lo_3131 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3132;
  assign dataGroup_hi_lo_3132 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3133;
  assign dataGroup_hi_lo_3133 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3134;
  assign dataGroup_hi_lo_3134 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3135;
  assign dataGroup_hi_lo_3135 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3136;
  assign dataGroup_hi_lo_3136 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3137;
  assign dataGroup_hi_lo_3137 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3138;
  assign dataGroup_hi_lo_3138 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3139;
  assign dataGroup_hi_lo_3139 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3140;
  assign dataGroup_hi_lo_3140 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3141;
  assign dataGroup_hi_lo_3141 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3142;
  assign dataGroup_hi_lo_3142 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3143;
  assign dataGroup_hi_lo_3143 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3144;
  assign dataGroup_hi_lo_3144 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3145;
  assign dataGroup_hi_lo_3145 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3146;
  assign dataGroup_hi_lo_3146 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3147;
  assign dataGroup_hi_lo_3147 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3148;
  assign dataGroup_hi_lo_3148 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3149;
  assign dataGroup_hi_lo_3149 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3150;
  assign dataGroup_hi_lo_3150 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3151;
  assign dataGroup_hi_lo_3151 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3152;
  assign dataGroup_hi_lo_3152 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3153;
  assign dataGroup_hi_lo_3153 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3154;
  assign dataGroup_hi_lo_3154 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3155;
  assign dataGroup_hi_lo_3155 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3156;
  assign dataGroup_hi_lo_3156 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3157;
  assign dataGroup_hi_lo_3157 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3158;
  assign dataGroup_hi_lo_3158 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3159;
  assign dataGroup_hi_lo_3159 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3160;
  assign dataGroup_hi_lo_3160 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3161;
  assign dataGroup_hi_lo_3161 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3162;
  assign dataGroup_hi_lo_3162 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3163;
  assign dataGroup_hi_lo_3163 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3164;
  assign dataGroup_hi_lo_3164 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3165;
  assign dataGroup_hi_lo_3165 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3166;
  assign dataGroup_hi_lo_3166 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3167;
  assign dataGroup_hi_lo_3167 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3168;
  assign dataGroup_hi_lo_3168 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3169;
  assign dataGroup_hi_lo_3169 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3170;
  assign dataGroup_hi_lo_3170 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3171;
  assign dataGroup_hi_lo_3171 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3172;
  assign dataGroup_hi_lo_3172 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3173;
  assign dataGroup_hi_lo_3173 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3174;
  assign dataGroup_hi_lo_3174 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3175;
  assign dataGroup_hi_lo_3175 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3176;
  assign dataGroup_hi_lo_3176 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3177;
  assign dataGroup_hi_lo_3177 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3178;
  assign dataGroup_hi_lo_3178 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3179;
  assign dataGroup_hi_lo_3179 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3180;
  assign dataGroup_hi_lo_3180 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3181;
  assign dataGroup_hi_lo_3181 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3182;
  assign dataGroup_hi_lo_3182 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3183;
  assign dataGroup_hi_lo_3183 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3184;
  assign dataGroup_hi_lo_3184 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3185;
  assign dataGroup_hi_lo_3185 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3186;
  assign dataGroup_hi_lo_3186 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3187;
  assign dataGroup_hi_lo_3187 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3188;
  assign dataGroup_hi_lo_3188 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3189;
  assign dataGroup_hi_lo_3189 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3190;
  assign dataGroup_hi_lo_3190 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3191;
  assign dataGroup_hi_lo_3191 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3192;
  assign dataGroup_hi_lo_3192 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3193;
  assign dataGroup_hi_lo_3193 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3194;
  assign dataGroup_hi_lo_3194 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3195;
  assign dataGroup_hi_lo_3195 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3196;
  assign dataGroup_hi_lo_3196 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3197;
  assign dataGroup_hi_lo_3197 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3198;
  assign dataGroup_hi_lo_3198 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3199;
  assign dataGroup_hi_lo_3199 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3200;
  assign dataGroup_hi_lo_3200 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3201;
  assign dataGroup_hi_lo_3201 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3202;
  assign dataGroup_hi_lo_3202 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3203;
  assign dataGroup_hi_lo_3203 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3204;
  assign dataGroup_hi_lo_3204 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3205;
  assign dataGroup_hi_lo_3205 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3206;
  assign dataGroup_hi_lo_3206 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3207;
  assign dataGroup_hi_lo_3207 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3208;
  assign dataGroup_hi_lo_3208 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3209;
  assign dataGroup_hi_lo_3209 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3210;
  assign dataGroup_hi_lo_3210 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3211;
  assign dataGroup_hi_lo_3211 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3212;
  assign dataGroup_hi_lo_3212 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3213;
  assign dataGroup_hi_lo_3213 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3214;
  assign dataGroup_hi_lo_3214 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3215;
  assign dataGroup_hi_lo_3215 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3216;
  assign dataGroup_hi_lo_3216 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3217;
  assign dataGroup_hi_lo_3217 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3218;
  assign dataGroup_hi_lo_3218 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3219;
  assign dataGroup_hi_lo_3219 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3220;
  assign dataGroup_hi_lo_3220 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3221;
  assign dataGroup_hi_lo_3221 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3222;
  assign dataGroup_hi_lo_3222 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3223;
  assign dataGroup_hi_lo_3223 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3224;
  assign dataGroup_hi_lo_3224 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3225;
  assign dataGroup_hi_lo_3225 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3226;
  assign dataGroup_hi_lo_3226 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3227;
  assign dataGroup_hi_lo_3227 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3228;
  assign dataGroup_hi_lo_3228 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3229;
  assign dataGroup_hi_lo_3229 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3230;
  assign dataGroup_hi_lo_3230 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3231;
  assign dataGroup_hi_lo_3231 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3232;
  assign dataGroup_hi_lo_3232 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3233;
  assign dataGroup_hi_lo_3233 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3234;
  assign dataGroup_hi_lo_3234 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3235;
  assign dataGroup_hi_lo_3235 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3236;
  assign dataGroup_hi_lo_3236 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3237;
  assign dataGroup_hi_lo_3237 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3238;
  assign dataGroup_hi_lo_3238 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3239;
  assign dataGroup_hi_lo_3239 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3240;
  assign dataGroup_hi_lo_3240 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3241;
  assign dataGroup_hi_lo_3241 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3242;
  assign dataGroup_hi_lo_3242 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3243;
  assign dataGroup_hi_lo_3243 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3244;
  assign dataGroup_hi_lo_3244 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3245;
  assign dataGroup_hi_lo_3245 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3246;
  assign dataGroup_hi_lo_3246 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3247;
  assign dataGroup_hi_lo_3247 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3248;
  assign dataGroup_hi_lo_3248 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3249;
  assign dataGroup_hi_lo_3249 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3250;
  assign dataGroup_hi_lo_3250 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3251;
  assign dataGroup_hi_lo_3251 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3252;
  assign dataGroup_hi_lo_3252 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3253;
  assign dataGroup_hi_lo_3253 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3254;
  assign dataGroup_hi_lo_3254 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3255;
  assign dataGroup_hi_lo_3255 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3256;
  assign dataGroup_hi_lo_3256 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3257;
  assign dataGroup_hi_lo_3257 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3258;
  assign dataGroup_hi_lo_3258 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3259;
  assign dataGroup_hi_lo_3259 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3260;
  assign dataGroup_hi_lo_3260 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3261;
  assign dataGroup_hi_lo_3261 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3262;
  assign dataGroup_hi_lo_3262 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3263;
  assign dataGroup_hi_lo_3263 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3264;
  assign dataGroup_hi_lo_3264 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3265;
  assign dataGroup_hi_lo_3265 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3266;
  assign dataGroup_hi_lo_3266 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3267;
  assign dataGroup_hi_lo_3267 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3268;
  assign dataGroup_hi_lo_3268 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3269;
  assign dataGroup_hi_lo_3269 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3270;
  assign dataGroup_hi_lo_3270 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3271;
  assign dataGroup_hi_lo_3271 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3272;
  assign dataGroup_hi_lo_3272 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3273;
  assign dataGroup_hi_lo_3273 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3274;
  assign dataGroup_hi_lo_3274 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3275;
  assign dataGroup_hi_lo_3275 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3276;
  assign dataGroup_hi_lo_3276 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3277;
  assign dataGroup_hi_lo_3277 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3278;
  assign dataGroup_hi_lo_3278 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3279;
  assign dataGroup_hi_lo_3279 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3280;
  assign dataGroup_hi_lo_3280 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3281;
  assign dataGroup_hi_lo_3281 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3282;
  assign dataGroup_hi_lo_3282 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3283;
  assign dataGroup_hi_lo_3283 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3284;
  assign dataGroup_hi_lo_3284 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3285;
  assign dataGroup_hi_lo_3285 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3286;
  assign dataGroup_hi_lo_3286 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3287;
  assign dataGroup_hi_lo_3287 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3288;
  assign dataGroup_hi_lo_3288 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3289;
  assign dataGroup_hi_lo_3289 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3290;
  assign dataGroup_hi_lo_3290 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3291;
  assign dataGroup_hi_lo_3291 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3292;
  assign dataGroup_hi_lo_3292 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3293;
  assign dataGroup_hi_lo_3293 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3294;
  assign dataGroup_hi_lo_3294 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3295;
  assign dataGroup_hi_lo_3295 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3296;
  assign dataGroup_hi_lo_3296 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3297;
  assign dataGroup_hi_lo_3297 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3298;
  assign dataGroup_hi_lo_3298 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3299;
  assign dataGroup_hi_lo_3299 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3300;
  assign dataGroup_hi_lo_3300 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3301;
  assign dataGroup_hi_lo_3301 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3302;
  assign dataGroup_hi_lo_3302 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3303;
  assign dataGroup_hi_lo_3303 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3304;
  assign dataGroup_hi_lo_3304 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3305;
  assign dataGroup_hi_lo_3305 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3306;
  assign dataGroup_hi_lo_3306 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3307;
  assign dataGroup_hi_lo_3307 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3308;
  assign dataGroup_hi_lo_3308 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3309;
  assign dataGroup_hi_lo_3309 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3310;
  assign dataGroup_hi_lo_3310 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3311;
  assign dataGroup_hi_lo_3311 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3312;
  assign dataGroup_hi_lo_3312 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3313;
  assign dataGroup_hi_lo_3313 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3314;
  assign dataGroup_hi_lo_3314 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3315;
  assign dataGroup_hi_lo_3315 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3316;
  assign dataGroup_hi_lo_3316 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3317;
  assign dataGroup_hi_lo_3317 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3318;
  assign dataGroup_hi_lo_3318 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3319;
  assign dataGroup_hi_lo_3319 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3320;
  assign dataGroup_hi_lo_3320 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3321;
  assign dataGroup_hi_lo_3321 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3322;
  assign dataGroup_hi_lo_3322 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3323;
  assign dataGroup_hi_lo_3323 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3324;
  assign dataGroup_hi_lo_3324 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3325;
  assign dataGroup_hi_lo_3325 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3326;
  assign dataGroup_hi_lo_3326 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3327;
  assign dataGroup_hi_lo_3327 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3328;
  assign dataGroup_hi_lo_3328 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3329;
  assign dataGroup_hi_lo_3329 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3330;
  assign dataGroup_hi_lo_3330 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3331;
  assign dataGroup_hi_lo_3331 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3332;
  assign dataGroup_hi_lo_3332 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3333;
  assign dataGroup_hi_lo_3333 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3334;
  assign dataGroup_hi_lo_3334 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3335;
  assign dataGroup_hi_lo_3335 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3336;
  assign dataGroup_hi_lo_3336 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3337;
  assign dataGroup_hi_lo_3337 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3338;
  assign dataGroup_hi_lo_3338 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3339;
  assign dataGroup_hi_lo_3339 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3340;
  assign dataGroup_hi_lo_3340 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3341;
  assign dataGroup_hi_lo_3341 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3342;
  assign dataGroup_hi_lo_3342 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3343;
  assign dataGroup_hi_lo_3343 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3344;
  assign dataGroup_hi_lo_3344 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3345;
  assign dataGroup_hi_lo_3345 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3346;
  assign dataGroup_hi_lo_3346 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3347;
  assign dataGroup_hi_lo_3347 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3348;
  assign dataGroup_hi_lo_3348 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3349;
  assign dataGroup_hi_lo_3349 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3350;
  assign dataGroup_hi_lo_3350 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3351;
  assign dataGroup_hi_lo_3351 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3352;
  assign dataGroup_hi_lo_3352 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3353;
  assign dataGroup_hi_lo_3353 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3354;
  assign dataGroup_hi_lo_3354 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3355;
  assign dataGroup_hi_lo_3355 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3356;
  assign dataGroup_hi_lo_3356 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3357;
  assign dataGroup_hi_lo_3357 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3358;
  assign dataGroup_hi_lo_3358 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3359;
  assign dataGroup_hi_lo_3359 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3360;
  assign dataGroup_hi_lo_3360 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3361;
  assign dataGroup_hi_lo_3361 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3362;
  assign dataGroup_hi_lo_3362 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3363;
  assign dataGroup_hi_lo_3363 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3364;
  assign dataGroup_hi_lo_3364 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3365;
  assign dataGroup_hi_lo_3365 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3366;
  assign dataGroup_hi_lo_3366 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3367;
  assign dataGroup_hi_lo_3367 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3368;
  assign dataGroup_hi_lo_3368 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3369;
  assign dataGroup_hi_lo_3369 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3370;
  assign dataGroup_hi_lo_3370 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3371;
  assign dataGroup_hi_lo_3371 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3372;
  assign dataGroup_hi_lo_3372 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3373;
  assign dataGroup_hi_lo_3373 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3374;
  assign dataGroup_hi_lo_3374 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3375;
  assign dataGroup_hi_lo_3375 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3376;
  assign dataGroup_hi_lo_3376 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3377;
  assign dataGroup_hi_lo_3377 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3378;
  assign dataGroup_hi_lo_3378 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3379;
  assign dataGroup_hi_lo_3379 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3380;
  assign dataGroup_hi_lo_3380 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3381;
  assign dataGroup_hi_lo_3381 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3382;
  assign dataGroup_hi_lo_3382 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3383;
  assign dataGroup_hi_lo_3383 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3384;
  assign dataGroup_hi_lo_3384 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3385;
  assign dataGroup_hi_lo_3385 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3386;
  assign dataGroup_hi_lo_3386 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3387;
  assign dataGroup_hi_lo_3387 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3388;
  assign dataGroup_hi_lo_3388 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3389;
  assign dataGroup_hi_lo_3389 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3390;
  assign dataGroup_hi_lo_3390 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3391;
  assign dataGroup_hi_lo_3391 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3392;
  assign dataGroup_hi_lo_3392 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3393;
  assign dataGroup_hi_lo_3393 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3394;
  assign dataGroup_hi_lo_3394 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3395;
  assign dataGroup_hi_lo_3395 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3396;
  assign dataGroup_hi_lo_3396 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3397;
  assign dataGroup_hi_lo_3397 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3398;
  assign dataGroup_hi_lo_3398 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3399;
  assign dataGroup_hi_lo_3399 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3400;
  assign dataGroup_hi_lo_3400 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3401;
  assign dataGroup_hi_lo_3401 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3402;
  assign dataGroup_hi_lo_3402 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3403;
  assign dataGroup_hi_lo_3403 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3404;
  assign dataGroup_hi_lo_3404 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3405;
  assign dataGroup_hi_lo_3405 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3406;
  assign dataGroup_hi_lo_3406 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3407;
  assign dataGroup_hi_lo_3407 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3408;
  assign dataGroup_hi_lo_3408 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3409;
  assign dataGroup_hi_lo_3409 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3410;
  assign dataGroup_hi_lo_3410 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3411;
  assign dataGroup_hi_lo_3411 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3412;
  assign dataGroup_hi_lo_3412 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3413;
  assign dataGroup_hi_lo_3413 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3414;
  assign dataGroup_hi_lo_3414 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3415;
  assign dataGroup_hi_lo_3415 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3416;
  assign dataGroup_hi_lo_3416 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3417;
  assign dataGroup_hi_lo_3417 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3418;
  assign dataGroup_hi_lo_3418 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3419;
  assign dataGroup_hi_lo_3419 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3420;
  assign dataGroup_hi_lo_3420 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3421;
  assign dataGroup_hi_lo_3421 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3422;
  assign dataGroup_hi_lo_3422 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3423;
  assign dataGroup_hi_lo_3423 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3424;
  assign dataGroup_hi_lo_3424 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3425;
  assign dataGroup_hi_lo_3425 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3426;
  assign dataGroup_hi_lo_3426 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3427;
  assign dataGroup_hi_lo_3427 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3428;
  assign dataGroup_hi_lo_3428 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3429;
  assign dataGroup_hi_lo_3429 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3430;
  assign dataGroup_hi_lo_3430 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3431;
  assign dataGroup_hi_lo_3431 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3432;
  assign dataGroup_hi_lo_3432 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3433;
  assign dataGroup_hi_lo_3433 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3434;
  assign dataGroup_hi_lo_3434 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3435;
  assign dataGroup_hi_lo_3435 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3436;
  assign dataGroup_hi_lo_3436 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3437;
  assign dataGroup_hi_lo_3437 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3438;
  assign dataGroup_hi_lo_3438 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3439;
  assign dataGroup_hi_lo_3439 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3440;
  assign dataGroup_hi_lo_3440 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3441;
  assign dataGroup_hi_lo_3441 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3442;
  assign dataGroup_hi_lo_3442 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3443;
  assign dataGroup_hi_lo_3443 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3444;
  assign dataGroup_hi_lo_3444 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3445;
  assign dataGroup_hi_lo_3445 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3446;
  assign dataGroup_hi_lo_3446 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3447;
  assign dataGroup_hi_lo_3447 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3448;
  assign dataGroup_hi_lo_3448 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3449;
  assign dataGroup_hi_lo_3449 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3450;
  assign dataGroup_hi_lo_3450 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3451;
  assign dataGroup_hi_lo_3451 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3452;
  assign dataGroup_hi_lo_3452 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3453;
  assign dataGroup_hi_lo_3453 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3454;
  assign dataGroup_hi_lo_3454 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3455;
  assign dataGroup_hi_lo_3455 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3456;
  assign dataGroup_hi_lo_3456 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3457;
  assign dataGroup_hi_lo_3457 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3458;
  assign dataGroup_hi_lo_3458 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3459;
  assign dataGroup_hi_lo_3459 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3460;
  assign dataGroup_hi_lo_3460 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3461;
  assign dataGroup_hi_lo_3461 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3462;
  assign dataGroup_hi_lo_3462 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3463;
  assign dataGroup_hi_lo_3463 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3464;
  assign dataGroup_hi_lo_3464 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3465;
  assign dataGroup_hi_lo_3465 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3466;
  assign dataGroup_hi_lo_3466 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3467;
  assign dataGroup_hi_lo_3467 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3468;
  assign dataGroup_hi_lo_3468 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3469;
  assign dataGroup_hi_lo_3469 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3470;
  assign dataGroup_hi_lo_3470 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3471;
  assign dataGroup_hi_lo_3471 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3472;
  assign dataGroup_hi_lo_3472 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3473;
  assign dataGroup_hi_lo_3473 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3474;
  assign dataGroup_hi_lo_3474 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3475;
  assign dataGroup_hi_lo_3475 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3476;
  assign dataGroup_hi_lo_3476 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3477;
  assign dataGroup_hi_lo_3477 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3478;
  assign dataGroup_hi_lo_3478 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3479;
  assign dataGroup_hi_lo_3479 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3480;
  assign dataGroup_hi_lo_3480 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3481;
  assign dataGroup_hi_lo_3481 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3482;
  assign dataGroup_hi_lo_3482 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3483;
  assign dataGroup_hi_lo_3483 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3484;
  assign dataGroup_hi_lo_3484 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3485;
  assign dataGroup_hi_lo_3485 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3486;
  assign dataGroup_hi_lo_3486 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3487;
  assign dataGroup_hi_lo_3487 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3488;
  assign dataGroup_hi_lo_3488 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3489;
  assign dataGroup_hi_lo_3489 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3490;
  assign dataGroup_hi_lo_3490 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3491;
  assign dataGroup_hi_lo_3491 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3492;
  assign dataGroup_hi_lo_3492 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3493;
  assign dataGroup_hi_lo_3493 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3494;
  assign dataGroup_hi_lo_3494 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3495;
  assign dataGroup_hi_lo_3495 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3496;
  assign dataGroup_hi_lo_3496 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3497;
  assign dataGroup_hi_lo_3497 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3498;
  assign dataGroup_hi_lo_3498 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3499;
  assign dataGroup_hi_lo_3499 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3500;
  assign dataGroup_hi_lo_3500 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3501;
  assign dataGroup_hi_lo_3501 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3502;
  assign dataGroup_hi_lo_3502 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3503;
  assign dataGroup_hi_lo_3503 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3504;
  assign dataGroup_hi_lo_3504 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3505;
  assign dataGroup_hi_lo_3505 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3506;
  assign dataGroup_hi_lo_3506 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3507;
  assign dataGroup_hi_lo_3507 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3508;
  assign dataGroup_hi_lo_3508 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3509;
  assign dataGroup_hi_lo_3509 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3510;
  assign dataGroup_hi_lo_3510 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3511;
  assign dataGroup_hi_lo_3511 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3512;
  assign dataGroup_hi_lo_3512 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3513;
  assign dataGroup_hi_lo_3513 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3514;
  assign dataGroup_hi_lo_3514 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3515;
  assign dataGroup_hi_lo_3515 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3516;
  assign dataGroup_hi_lo_3516 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3517;
  assign dataGroup_hi_lo_3517 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3518;
  assign dataGroup_hi_lo_3518 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3519;
  assign dataGroup_hi_lo_3519 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3520;
  assign dataGroup_hi_lo_3520 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3521;
  assign dataGroup_hi_lo_3521 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3522;
  assign dataGroup_hi_lo_3522 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3523;
  assign dataGroup_hi_lo_3523 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3524;
  assign dataGroup_hi_lo_3524 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3525;
  assign dataGroup_hi_lo_3525 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3526;
  assign dataGroup_hi_lo_3526 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3527;
  assign dataGroup_hi_lo_3527 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3528;
  assign dataGroup_hi_lo_3528 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3529;
  assign dataGroup_hi_lo_3529 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3530;
  assign dataGroup_hi_lo_3530 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3531;
  assign dataGroup_hi_lo_3531 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3532;
  assign dataGroup_hi_lo_3532 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3533;
  assign dataGroup_hi_lo_3533 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3534;
  assign dataGroup_hi_lo_3534 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3535;
  assign dataGroup_hi_lo_3535 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3536;
  assign dataGroup_hi_lo_3536 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3537;
  assign dataGroup_hi_lo_3537 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3538;
  assign dataGroup_hi_lo_3538 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3539;
  assign dataGroup_hi_lo_3539 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3540;
  assign dataGroup_hi_lo_3540 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3541;
  assign dataGroup_hi_lo_3541 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3542;
  assign dataGroup_hi_lo_3542 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3543;
  assign dataGroup_hi_lo_3543 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3544;
  assign dataGroup_hi_lo_3544 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3545;
  assign dataGroup_hi_lo_3545 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3546;
  assign dataGroup_hi_lo_3546 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3547;
  assign dataGroup_hi_lo_3547 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3548;
  assign dataGroup_hi_lo_3548 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3549;
  assign dataGroup_hi_lo_3549 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3550;
  assign dataGroup_hi_lo_3550 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3551;
  assign dataGroup_hi_lo_3551 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3552;
  assign dataGroup_hi_lo_3552 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3553;
  assign dataGroup_hi_lo_3553 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3554;
  assign dataGroup_hi_lo_3554 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3555;
  assign dataGroup_hi_lo_3555 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3556;
  assign dataGroup_hi_lo_3556 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3557;
  assign dataGroup_hi_lo_3557 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3558;
  assign dataGroup_hi_lo_3558 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3559;
  assign dataGroup_hi_lo_3559 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3560;
  assign dataGroup_hi_lo_3560 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3561;
  assign dataGroup_hi_lo_3561 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3562;
  assign dataGroup_hi_lo_3562 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3563;
  assign dataGroup_hi_lo_3563 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3564;
  assign dataGroup_hi_lo_3564 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3565;
  assign dataGroup_hi_lo_3565 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3566;
  assign dataGroup_hi_lo_3566 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3567;
  assign dataGroup_hi_lo_3567 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3568;
  assign dataGroup_hi_lo_3568 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3569;
  assign dataGroup_hi_lo_3569 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3570;
  assign dataGroup_hi_lo_3570 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3571;
  assign dataGroup_hi_lo_3571 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3572;
  assign dataGroup_hi_lo_3572 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3573;
  assign dataGroup_hi_lo_3573 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3574;
  assign dataGroup_hi_lo_3574 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3575;
  assign dataGroup_hi_lo_3575 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3576;
  assign dataGroup_hi_lo_3576 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3577;
  assign dataGroup_hi_lo_3577 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3578;
  assign dataGroup_hi_lo_3578 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3579;
  assign dataGroup_hi_lo_3579 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3580;
  assign dataGroup_hi_lo_3580 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3581;
  assign dataGroup_hi_lo_3581 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3582;
  assign dataGroup_hi_lo_3582 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3583;
  assign dataGroup_hi_lo_3583 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3584;
  assign dataGroup_hi_lo_3584 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3585;
  assign dataGroup_hi_lo_3585 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3586;
  assign dataGroup_hi_lo_3586 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3587;
  assign dataGroup_hi_lo_3587 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3588;
  assign dataGroup_hi_lo_3588 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3589;
  assign dataGroup_hi_lo_3589 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3590;
  assign dataGroup_hi_lo_3590 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3591;
  assign dataGroup_hi_lo_3591 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3592;
  assign dataGroup_hi_lo_3592 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3593;
  assign dataGroup_hi_lo_3593 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3594;
  assign dataGroup_hi_lo_3594 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3595;
  assign dataGroup_hi_lo_3595 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3596;
  assign dataGroup_hi_lo_3596 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3597;
  assign dataGroup_hi_lo_3597 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3598;
  assign dataGroup_hi_lo_3598 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3599;
  assign dataGroup_hi_lo_3599 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3600;
  assign dataGroup_hi_lo_3600 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3601;
  assign dataGroup_hi_lo_3601 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3602;
  assign dataGroup_hi_lo_3602 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3603;
  assign dataGroup_hi_lo_3603 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3604;
  assign dataGroup_hi_lo_3604 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3605;
  assign dataGroup_hi_lo_3605 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3606;
  assign dataGroup_hi_lo_3606 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3607;
  assign dataGroup_hi_lo_3607 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3608;
  assign dataGroup_hi_lo_3608 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3609;
  assign dataGroup_hi_lo_3609 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3610;
  assign dataGroup_hi_lo_3610 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3611;
  assign dataGroup_hi_lo_3611 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3612;
  assign dataGroup_hi_lo_3612 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3613;
  assign dataGroup_hi_lo_3613 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3614;
  assign dataGroup_hi_lo_3614 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3615;
  assign dataGroup_hi_lo_3615 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3616;
  assign dataGroup_hi_lo_3616 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3617;
  assign dataGroup_hi_lo_3617 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3618;
  assign dataGroup_hi_lo_3618 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3619;
  assign dataGroup_hi_lo_3619 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3620;
  assign dataGroup_hi_lo_3620 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3621;
  assign dataGroup_hi_lo_3621 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3622;
  assign dataGroup_hi_lo_3622 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3623;
  assign dataGroup_hi_lo_3623 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3624;
  assign dataGroup_hi_lo_3624 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3625;
  assign dataGroup_hi_lo_3625 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3626;
  assign dataGroup_hi_lo_3626 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3627;
  assign dataGroup_hi_lo_3627 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3628;
  assign dataGroup_hi_lo_3628 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3629;
  assign dataGroup_hi_lo_3629 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3630;
  assign dataGroup_hi_lo_3630 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3631;
  assign dataGroup_hi_lo_3631 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3632;
  assign dataGroup_hi_lo_3632 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3633;
  assign dataGroup_hi_lo_3633 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3634;
  assign dataGroup_hi_lo_3634 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3635;
  assign dataGroup_hi_lo_3635 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3636;
  assign dataGroup_hi_lo_3636 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3637;
  assign dataGroup_hi_lo_3637 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3638;
  assign dataGroup_hi_lo_3638 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3639;
  assign dataGroup_hi_lo_3639 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3640;
  assign dataGroup_hi_lo_3640 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3641;
  assign dataGroup_hi_lo_3641 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3642;
  assign dataGroup_hi_lo_3642 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3643;
  assign dataGroup_hi_lo_3643 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3644;
  assign dataGroup_hi_lo_3644 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3645;
  assign dataGroup_hi_lo_3645 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3646;
  assign dataGroup_hi_lo_3646 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3647;
  assign dataGroup_hi_lo_3647 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3648;
  assign dataGroup_hi_lo_3648 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3649;
  assign dataGroup_hi_lo_3649 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3650;
  assign dataGroup_hi_lo_3650 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3651;
  assign dataGroup_hi_lo_3651 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3652;
  assign dataGroup_hi_lo_3652 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3653;
  assign dataGroup_hi_lo_3653 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3654;
  assign dataGroup_hi_lo_3654 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3655;
  assign dataGroup_hi_lo_3655 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3656;
  assign dataGroup_hi_lo_3656 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3657;
  assign dataGroup_hi_lo_3657 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3658;
  assign dataGroup_hi_lo_3658 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3659;
  assign dataGroup_hi_lo_3659 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3660;
  assign dataGroup_hi_lo_3660 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3661;
  assign dataGroup_hi_lo_3661 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3662;
  assign dataGroup_hi_lo_3662 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3663;
  assign dataGroup_hi_lo_3663 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3664;
  assign dataGroup_hi_lo_3664 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3665;
  assign dataGroup_hi_lo_3665 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3666;
  assign dataGroup_hi_lo_3666 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3667;
  assign dataGroup_hi_lo_3667 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3668;
  assign dataGroup_hi_lo_3668 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3669;
  assign dataGroup_hi_lo_3669 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3670;
  assign dataGroup_hi_lo_3670 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3671;
  assign dataGroup_hi_lo_3671 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3672;
  assign dataGroup_hi_lo_3672 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3673;
  assign dataGroup_hi_lo_3673 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3674;
  assign dataGroup_hi_lo_3674 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3675;
  assign dataGroup_hi_lo_3675 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3676;
  assign dataGroup_hi_lo_3676 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3677;
  assign dataGroup_hi_lo_3677 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3678;
  assign dataGroup_hi_lo_3678 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3679;
  assign dataGroup_hi_lo_3679 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3680;
  assign dataGroup_hi_lo_3680 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3681;
  assign dataGroup_hi_lo_3681 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3682;
  assign dataGroup_hi_lo_3682 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3683;
  assign dataGroup_hi_lo_3683 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3684;
  assign dataGroup_hi_lo_3684 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3685;
  assign dataGroup_hi_lo_3685 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3686;
  assign dataGroup_hi_lo_3686 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3687;
  assign dataGroup_hi_lo_3687 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3688;
  assign dataGroup_hi_lo_3688 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3689;
  assign dataGroup_hi_lo_3689 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3690;
  assign dataGroup_hi_lo_3690 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3691;
  assign dataGroup_hi_lo_3691 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3692;
  assign dataGroup_hi_lo_3692 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3693;
  assign dataGroup_hi_lo_3693 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3694;
  assign dataGroup_hi_lo_3694 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3695;
  assign dataGroup_hi_lo_3695 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3696;
  assign dataGroup_hi_lo_3696 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3697;
  assign dataGroup_hi_lo_3697 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3698;
  assign dataGroup_hi_lo_3698 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3699;
  assign dataGroup_hi_lo_3699 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3700;
  assign dataGroup_hi_lo_3700 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3701;
  assign dataGroup_hi_lo_3701 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3702;
  assign dataGroup_hi_lo_3702 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3703;
  assign dataGroup_hi_lo_3703 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3704;
  assign dataGroup_hi_lo_3704 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3705;
  assign dataGroup_hi_lo_3705 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3706;
  assign dataGroup_hi_lo_3706 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3707;
  assign dataGroup_hi_lo_3707 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3708;
  assign dataGroup_hi_lo_3708 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3709;
  assign dataGroup_hi_lo_3709 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3710;
  assign dataGroup_hi_lo_3710 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3711;
  assign dataGroup_hi_lo_3711 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3712;
  assign dataGroup_hi_lo_3712 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3713;
  assign dataGroup_hi_lo_3713 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3714;
  assign dataGroup_hi_lo_3714 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3715;
  assign dataGroup_hi_lo_3715 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3716;
  assign dataGroup_hi_lo_3716 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3717;
  assign dataGroup_hi_lo_3717 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3718;
  assign dataGroup_hi_lo_3718 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3719;
  assign dataGroup_hi_lo_3719 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3720;
  assign dataGroup_hi_lo_3720 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3721;
  assign dataGroup_hi_lo_3721 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3722;
  assign dataGroup_hi_lo_3722 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3723;
  assign dataGroup_hi_lo_3723 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3724;
  assign dataGroup_hi_lo_3724 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3725;
  assign dataGroup_hi_lo_3725 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3726;
  assign dataGroup_hi_lo_3726 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3727;
  assign dataGroup_hi_lo_3727 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3728;
  assign dataGroup_hi_lo_3728 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3729;
  assign dataGroup_hi_lo_3729 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3730;
  assign dataGroup_hi_lo_3730 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3731;
  assign dataGroup_hi_lo_3731 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3732;
  assign dataGroup_hi_lo_3732 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3733;
  assign dataGroup_hi_lo_3733 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3734;
  assign dataGroup_hi_lo_3734 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3735;
  assign dataGroup_hi_lo_3735 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3736;
  assign dataGroup_hi_lo_3736 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3737;
  assign dataGroup_hi_lo_3737 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3738;
  assign dataGroup_hi_lo_3738 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3739;
  assign dataGroup_hi_lo_3739 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3740;
  assign dataGroup_hi_lo_3740 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3741;
  assign dataGroup_hi_lo_3741 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3742;
  assign dataGroup_hi_lo_3742 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3743;
  assign dataGroup_hi_lo_3743 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3744;
  assign dataGroup_hi_lo_3744 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3745;
  assign dataGroup_hi_lo_3745 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3746;
  assign dataGroup_hi_lo_3746 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3747;
  assign dataGroup_hi_lo_3747 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3748;
  assign dataGroup_hi_lo_3748 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3749;
  assign dataGroup_hi_lo_3749 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3750;
  assign dataGroup_hi_lo_3750 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3751;
  assign dataGroup_hi_lo_3751 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3752;
  assign dataGroup_hi_lo_3752 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3753;
  assign dataGroup_hi_lo_3753 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3754;
  assign dataGroup_hi_lo_3754 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3755;
  assign dataGroup_hi_lo_3755 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3756;
  assign dataGroup_hi_lo_3756 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3757;
  assign dataGroup_hi_lo_3757 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3758;
  assign dataGroup_hi_lo_3758 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3759;
  assign dataGroup_hi_lo_3759 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3760;
  assign dataGroup_hi_lo_3760 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3761;
  assign dataGroup_hi_lo_3761 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3762;
  assign dataGroup_hi_lo_3762 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3763;
  assign dataGroup_hi_lo_3763 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3764;
  assign dataGroup_hi_lo_3764 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3765;
  assign dataGroup_hi_lo_3765 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3766;
  assign dataGroup_hi_lo_3766 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3767;
  assign dataGroup_hi_lo_3767 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3768;
  assign dataGroup_hi_lo_3768 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3769;
  assign dataGroup_hi_lo_3769 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3770;
  assign dataGroup_hi_lo_3770 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3771;
  assign dataGroup_hi_lo_3771 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3772;
  assign dataGroup_hi_lo_3772 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3773;
  assign dataGroup_hi_lo_3773 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3774;
  assign dataGroup_hi_lo_3774 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3775;
  assign dataGroup_hi_lo_3775 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3776;
  assign dataGroup_hi_lo_3776 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3777;
  assign dataGroup_hi_lo_3777 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3778;
  assign dataGroup_hi_lo_3778 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3779;
  assign dataGroup_hi_lo_3779 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3780;
  assign dataGroup_hi_lo_3780 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3781;
  assign dataGroup_hi_lo_3781 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3782;
  assign dataGroup_hi_lo_3782 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3783;
  assign dataGroup_hi_lo_3783 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3784;
  assign dataGroup_hi_lo_3784 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3785;
  assign dataGroup_hi_lo_3785 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3786;
  assign dataGroup_hi_lo_3786 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3787;
  assign dataGroup_hi_lo_3787 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3788;
  assign dataGroup_hi_lo_3788 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3789;
  assign dataGroup_hi_lo_3789 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3790;
  assign dataGroup_hi_lo_3790 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3791;
  assign dataGroup_hi_lo_3791 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3792;
  assign dataGroup_hi_lo_3792 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3793;
  assign dataGroup_hi_lo_3793 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3794;
  assign dataGroup_hi_lo_3794 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3795;
  assign dataGroup_hi_lo_3795 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3796;
  assign dataGroup_hi_lo_3796 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3797;
  assign dataGroup_hi_lo_3797 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3798;
  assign dataGroup_hi_lo_3798 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3799;
  assign dataGroup_hi_lo_3799 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3800;
  assign dataGroup_hi_lo_3800 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3801;
  assign dataGroup_hi_lo_3801 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3802;
  assign dataGroup_hi_lo_3802 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3803;
  assign dataGroup_hi_lo_3803 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3804;
  assign dataGroup_hi_lo_3804 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3805;
  assign dataGroup_hi_lo_3805 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3806;
  assign dataGroup_hi_lo_3806 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3807;
  assign dataGroup_hi_lo_3807 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3808;
  assign dataGroup_hi_lo_3808 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3809;
  assign dataGroup_hi_lo_3809 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3810;
  assign dataGroup_hi_lo_3810 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3811;
  assign dataGroup_hi_lo_3811 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3812;
  assign dataGroup_hi_lo_3812 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3813;
  assign dataGroup_hi_lo_3813 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3814;
  assign dataGroup_hi_lo_3814 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3815;
  assign dataGroup_hi_lo_3815 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3816;
  assign dataGroup_hi_lo_3816 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3817;
  assign dataGroup_hi_lo_3817 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3818;
  assign dataGroup_hi_lo_3818 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3819;
  assign dataGroup_hi_lo_3819 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3820;
  assign dataGroup_hi_lo_3820 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3821;
  assign dataGroup_hi_lo_3821 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3822;
  assign dataGroup_hi_lo_3822 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3823;
  assign dataGroup_hi_lo_3823 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3824;
  assign dataGroup_hi_lo_3824 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3825;
  assign dataGroup_hi_lo_3825 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3826;
  assign dataGroup_hi_lo_3826 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3827;
  assign dataGroup_hi_lo_3827 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3828;
  assign dataGroup_hi_lo_3828 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3829;
  assign dataGroup_hi_lo_3829 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3830;
  assign dataGroup_hi_lo_3830 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3831;
  assign dataGroup_hi_lo_3831 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3832;
  assign dataGroup_hi_lo_3832 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3833;
  assign dataGroup_hi_lo_3833 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3834;
  assign dataGroup_hi_lo_3834 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3835;
  assign dataGroup_hi_lo_3835 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3836;
  assign dataGroup_hi_lo_3836 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3837;
  assign dataGroup_hi_lo_3837 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3838;
  assign dataGroup_hi_lo_3838 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3839;
  assign dataGroup_hi_lo_3839 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3840;
  assign dataGroup_hi_lo_3840 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3841;
  assign dataGroup_hi_lo_3841 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3842;
  assign dataGroup_hi_lo_3842 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3843;
  assign dataGroup_hi_lo_3843 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3844;
  assign dataGroup_hi_lo_3844 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3845;
  assign dataGroup_hi_lo_3845 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3846;
  assign dataGroup_hi_lo_3846 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3847;
  assign dataGroup_hi_lo_3847 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3848;
  assign dataGroup_hi_lo_3848 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3849;
  assign dataGroup_hi_lo_3849 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3850;
  assign dataGroup_hi_lo_3850 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3851;
  assign dataGroup_hi_lo_3851 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3852;
  assign dataGroup_hi_lo_3852 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3853;
  assign dataGroup_hi_lo_3853 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3854;
  assign dataGroup_hi_lo_3854 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3855;
  assign dataGroup_hi_lo_3855 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3856;
  assign dataGroup_hi_lo_3856 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3857;
  assign dataGroup_hi_lo_3857 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3858;
  assign dataGroup_hi_lo_3858 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3859;
  assign dataGroup_hi_lo_3859 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3860;
  assign dataGroup_hi_lo_3860 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3861;
  assign dataGroup_hi_lo_3861 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3862;
  assign dataGroup_hi_lo_3862 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3863;
  assign dataGroup_hi_lo_3863 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3864;
  assign dataGroup_hi_lo_3864 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3865;
  assign dataGroup_hi_lo_3865 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3866;
  assign dataGroup_hi_lo_3866 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3867;
  assign dataGroup_hi_lo_3867 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3868;
  assign dataGroup_hi_lo_3868 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3869;
  assign dataGroup_hi_lo_3869 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3870;
  assign dataGroup_hi_lo_3870 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3871;
  assign dataGroup_hi_lo_3871 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3872;
  assign dataGroup_hi_lo_3872 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3873;
  assign dataGroup_hi_lo_3873 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3874;
  assign dataGroup_hi_lo_3874 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3875;
  assign dataGroup_hi_lo_3875 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3876;
  assign dataGroup_hi_lo_3876 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3877;
  assign dataGroup_hi_lo_3877 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3878;
  assign dataGroup_hi_lo_3878 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3879;
  assign dataGroup_hi_lo_3879 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3880;
  assign dataGroup_hi_lo_3880 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3881;
  assign dataGroup_hi_lo_3881 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3882;
  assign dataGroup_hi_lo_3882 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3883;
  assign dataGroup_hi_lo_3883 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3884;
  assign dataGroup_hi_lo_3884 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3885;
  assign dataGroup_hi_lo_3885 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3886;
  assign dataGroup_hi_lo_3886 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3887;
  assign dataGroup_hi_lo_3887 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3888;
  assign dataGroup_hi_lo_3888 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3889;
  assign dataGroup_hi_lo_3889 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3890;
  assign dataGroup_hi_lo_3890 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3891;
  assign dataGroup_hi_lo_3891 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3892;
  assign dataGroup_hi_lo_3892 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3893;
  assign dataGroup_hi_lo_3893 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3894;
  assign dataGroup_hi_lo_3894 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3895;
  assign dataGroup_hi_lo_3895 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3896;
  assign dataGroup_hi_lo_3896 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3897;
  assign dataGroup_hi_lo_3897 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3898;
  assign dataGroup_hi_lo_3898 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3899;
  assign dataGroup_hi_lo_3899 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3900;
  assign dataGroup_hi_lo_3900 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3901;
  assign dataGroup_hi_lo_3901 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3902;
  assign dataGroup_hi_lo_3902 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3903;
  assign dataGroup_hi_lo_3903 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3904;
  assign dataGroup_hi_lo_3904 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3905;
  assign dataGroup_hi_lo_3905 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3906;
  assign dataGroup_hi_lo_3906 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3907;
  assign dataGroup_hi_lo_3907 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3908;
  assign dataGroup_hi_lo_3908 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3909;
  assign dataGroup_hi_lo_3909 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3910;
  assign dataGroup_hi_lo_3910 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3911;
  assign dataGroup_hi_lo_3911 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3912;
  assign dataGroup_hi_lo_3912 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3913;
  assign dataGroup_hi_lo_3913 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3914;
  assign dataGroup_hi_lo_3914 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3915;
  assign dataGroup_hi_lo_3915 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3916;
  assign dataGroup_hi_lo_3916 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3917;
  assign dataGroup_hi_lo_3917 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3918;
  assign dataGroup_hi_lo_3918 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3919;
  assign dataGroup_hi_lo_3919 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3920;
  assign dataGroup_hi_lo_3920 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3921;
  assign dataGroup_hi_lo_3921 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3922;
  assign dataGroup_hi_lo_3922 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3923;
  assign dataGroup_hi_lo_3923 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3924;
  assign dataGroup_hi_lo_3924 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3925;
  assign dataGroup_hi_lo_3925 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3926;
  assign dataGroup_hi_lo_3926 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3927;
  assign dataGroup_hi_lo_3927 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3928;
  assign dataGroup_hi_lo_3928 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3929;
  assign dataGroup_hi_lo_3929 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3930;
  assign dataGroup_hi_lo_3930 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3931;
  assign dataGroup_hi_lo_3931 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3932;
  assign dataGroup_hi_lo_3932 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3933;
  assign dataGroup_hi_lo_3933 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3934;
  assign dataGroup_hi_lo_3934 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3935;
  assign dataGroup_hi_lo_3935 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3936;
  assign dataGroup_hi_lo_3936 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3937;
  assign dataGroup_hi_lo_3937 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3938;
  assign dataGroup_hi_lo_3938 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3939;
  assign dataGroup_hi_lo_3939 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3940;
  assign dataGroup_hi_lo_3940 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3941;
  assign dataGroup_hi_lo_3941 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3942;
  assign dataGroup_hi_lo_3942 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3943;
  assign dataGroup_hi_lo_3943 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3944;
  assign dataGroup_hi_lo_3944 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3945;
  assign dataGroup_hi_lo_3945 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3946;
  assign dataGroup_hi_lo_3946 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3947;
  assign dataGroup_hi_lo_3947 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3948;
  assign dataGroup_hi_lo_3948 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3949;
  assign dataGroup_hi_lo_3949 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3950;
  assign dataGroup_hi_lo_3950 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3951;
  assign dataGroup_hi_lo_3951 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3952;
  assign dataGroup_hi_lo_3952 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3953;
  assign dataGroup_hi_lo_3953 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3954;
  assign dataGroup_hi_lo_3954 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3955;
  assign dataGroup_hi_lo_3955 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3956;
  assign dataGroup_hi_lo_3956 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3957;
  assign dataGroup_hi_lo_3957 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3958;
  assign dataGroup_hi_lo_3958 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3959;
  assign dataGroup_hi_lo_3959 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3960;
  assign dataGroup_hi_lo_3960 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3961;
  assign dataGroup_hi_lo_3961 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3962;
  assign dataGroup_hi_lo_3962 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3963;
  assign dataGroup_hi_lo_3963 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3964;
  assign dataGroup_hi_lo_3964 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3965;
  assign dataGroup_hi_lo_3965 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3966;
  assign dataGroup_hi_lo_3966 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3967;
  assign dataGroup_hi_lo_3967 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3968;
  assign dataGroup_hi_lo_3968 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3969;
  assign dataGroup_hi_lo_3969 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3970;
  assign dataGroup_hi_lo_3970 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3971;
  assign dataGroup_hi_lo_3971 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3972;
  assign dataGroup_hi_lo_3972 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3973;
  assign dataGroup_hi_lo_3973 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3974;
  assign dataGroup_hi_lo_3974 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3975;
  assign dataGroup_hi_lo_3975 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3976;
  assign dataGroup_hi_lo_3976 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3977;
  assign dataGroup_hi_lo_3977 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3978;
  assign dataGroup_hi_lo_3978 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3979;
  assign dataGroup_hi_lo_3979 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3980;
  assign dataGroup_hi_lo_3980 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3981;
  assign dataGroup_hi_lo_3981 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3982;
  assign dataGroup_hi_lo_3982 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3983;
  assign dataGroup_hi_lo_3983 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3984;
  assign dataGroup_hi_lo_3984 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3985;
  assign dataGroup_hi_lo_3985 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3986;
  assign dataGroup_hi_lo_3986 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3987;
  assign dataGroup_hi_lo_3987 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3988;
  assign dataGroup_hi_lo_3988 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3989;
  assign dataGroup_hi_lo_3989 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3990;
  assign dataGroup_hi_lo_3990 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3991;
  assign dataGroup_hi_lo_3991 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3992;
  assign dataGroup_hi_lo_3992 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3993;
  assign dataGroup_hi_lo_3993 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3994;
  assign dataGroup_hi_lo_3994 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3995;
  assign dataGroup_hi_lo_3995 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3996;
  assign dataGroup_hi_lo_3996 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3997;
  assign dataGroup_hi_lo_3997 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3998;
  assign dataGroup_hi_lo_3998 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_3999;
  assign dataGroup_hi_lo_3999 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4000;
  assign dataGroup_hi_lo_4000 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4001;
  assign dataGroup_hi_lo_4001 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4002;
  assign dataGroup_hi_lo_4002 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4003;
  assign dataGroup_hi_lo_4003 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4004;
  assign dataGroup_hi_lo_4004 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4005;
  assign dataGroup_hi_lo_4005 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4006;
  assign dataGroup_hi_lo_4006 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4007;
  assign dataGroup_hi_lo_4007 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4008;
  assign dataGroup_hi_lo_4008 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4009;
  assign dataGroup_hi_lo_4009 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4010;
  assign dataGroup_hi_lo_4010 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4011;
  assign dataGroup_hi_lo_4011 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4012;
  assign dataGroup_hi_lo_4012 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4013;
  assign dataGroup_hi_lo_4013 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4014;
  assign dataGroup_hi_lo_4014 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4015;
  assign dataGroup_hi_lo_4015 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4016;
  assign dataGroup_hi_lo_4016 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4017;
  assign dataGroup_hi_lo_4017 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4018;
  assign dataGroup_hi_lo_4018 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4019;
  assign dataGroup_hi_lo_4019 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4020;
  assign dataGroup_hi_lo_4020 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4021;
  assign dataGroup_hi_lo_4021 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4022;
  assign dataGroup_hi_lo_4022 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4023;
  assign dataGroup_hi_lo_4023 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4024;
  assign dataGroup_hi_lo_4024 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4025;
  assign dataGroup_hi_lo_4025 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4026;
  assign dataGroup_hi_lo_4026 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4027;
  assign dataGroup_hi_lo_4027 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4028;
  assign dataGroup_hi_lo_4028 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4029;
  assign dataGroup_hi_lo_4029 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4030;
  assign dataGroup_hi_lo_4030 = _GEN_7;
  wire [1023:0] dataGroup_hi_lo_4031;
  assign dataGroup_hi_lo_4031 = _GEN_7;
  wire [1023:0] _GEN_8 = {dataSelect_7, dataSelect_6};
  wire [1023:0] dataGroup_hi_hi;
  assign dataGroup_hi_hi = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1;
  assign dataGroup_hi_hi_1 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2;
  assign dataGroup_hi_hi_2 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3;
  assign dataGroup_hi_hi_3 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4;
  assign dataGroup_hi_hi_4 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_5;
  assign dataGroup_hi_hi_5 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_6;
  assign dataGroup_hi_hi_6 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_7;
  assign dataGroup_hi_hi_7 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_8;
  assign dataGroup_hi_hi_8 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_9;
  assign dataGroup_hi_hi_9 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_10;
  assign dataGroup_hi_hi_10 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_11;
  assign dataGroup_hi_hi_11 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_12;
  assign dataGroup_hi_hi_12 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_13;
  assign dataGroup_hi_hi_13 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_14;
  assign dataGroup_hi_hi_14 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_15;
  assign dataGroup_hi_hi_15 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_16;
  assign dataGroup_hi_hi_16 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_17;
  assign dataGroup_hi_hi_17 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_18;
  assign dataGroup_hi_hi_18 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_19;
  assign dataGroup_hi_hi_19 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_20;
  assign dataGroup_hi_hi_20 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_21;
  assign dataGroup_hi_hi_21 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_22;
  assign dataGroup_hi_hi_22 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_23;
  assign dataGroup_hi_hi_23 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_24;
  assign dataGroup_hi_hi_24 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_25;
  assign dataGroup_hi_hi_25 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_26;
  assign dataGroup_hi_hi_26 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_27;
  assign dataGroup_hi_hi_27 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_28;
  assign dataGroup_hi_hi_28 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_29;
  assign dataGroup_hi_hi_29 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_30;
  assign dataGroup_hi_hi_30 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_31;
  assign dataGroup_hi_hi_31 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_32;
  assign dataGroup_hi_hi_32 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_33;
  assign dataGroup_hi_hi_33 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_34;
  assign dataGroup_hi_hi_34 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_35;
  assign dataGroup_hi_hi_35 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_36;
  assign dataGroup_hi_hi_36 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_37;
  assign dataGroup_hi_hi_37 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_38;
  assign dataGroup_hi_hi_38 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_39;
  assign dataGroup_hi_hi_39 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_40;
  assign dataGroup_hi_hi_40 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_41;
  assign dataGroup_hi_hi_41 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_42;
  assign dataGroup_hi_hi_42 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_43;
  assign dataGroup_hi_hi_43 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_44;
  assign dataGroup_hi_hi_44 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_45;
  assign dataGroup_hi_hi_45 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_46;
  assign dataGroup_hi_hi_46 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_47;
  assign dataGroup_hi_hi_47 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_48;
  assign dataGroup_hi_hi_48 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_49;
  assign dataGroup_hi_hi_49 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_50;
  assign dataGroup_hi_hi_50 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_51;
  assign dataGroup_hi_hi_51 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_52;
  assign dataGroup_hi_hi_52 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_53;
  assign dataGroup_hi_hi_53 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_54;
  assign dataGroup_hi_hi_54 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_55;
  assign dataGroup_hi_hi_55 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_56;
  assign dataGroup_hi_hi_56 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_57;
  assign dataGroup_hi_hi_57 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_58;
  assign dataGroup_hi_hi_58 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_59;
  assign dataGroup_hi_hi_59 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_60;
  assign dataGroup_hi_hi_60 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_61;
  assign dataGroup_hi_hi_61 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_62;
  assign dataGroup_hi_hi_62 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_63;
  assign dataGroup_hi_hi_63 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_64;
  assign dataGroup_hi_hi_64 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_65;
  assign dataGroup_hi_hi_65 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_66;
  assign dataGroup_hi_hi_66 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_67;
  assign dataGroup_hi_hi_67 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_68;
  assign dataGroup_hi_hi_68 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_69;
  assign dataGroup_hi_hi_69 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_70;
  assign dataGroup_hi_hi_70 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_71;
  assign dataGroup_hi_hi_71 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_72;
  assign dataGroup_hi_hi_72 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_73;
  assign dataGroup_hi_hi_73 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_74;
  assign dataGroup_hi_hi_74 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_75;
  assign dataGroup_hi_hi_75 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_76;
  assign dataGroup_hi_hi_76 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_77;
  assign dataGroup_hi_hi_77 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_78;
  assign dataGroup_hi_hi_78 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_79;
  assign dataGroup_hi_hi_79 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_80;
  assign dataGroup_hi_hi_80 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_81;
  assign dataGroup_hi_hi_81 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_82;
  assign dataGroup_hi_hi_82 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_83;
  assign dataGroup_hi_hi_83 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_84;
  assign dataGroup_hi_hi_84 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_85;
  assign dataGroup_hi_hi_85 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_86;
  assign dataGroup_hi_hi_86 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_87;
  assign dataGroup_hi_hi_87 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_88;
  assign dataGroup_hi_hi_88 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_89;
  assign dataGroup_hi_hi_89 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_90;
  assign dataGroup_hi_hi_90 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_91;
  assign dataGroup_hi_hi_91 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_92;
  assign dataGroup_hi_hi_92 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_93;
  assign dataGroup_hi_hi_93 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_94;
  assign dataGroup_hi_hi_94 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_95;
  assign dataGroup_hi_hi_95 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_96;
  assign dataGroup_hi_hi_96 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_97;
  assign dataGroup_hi_hi_97 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_98;
  assign dataGroup_hi_hi_98 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_99;
  assign dataGroup_hi_hi_99 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_100;
  assign dataGroup_hi_hi_100 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_101;
  assign dataGroup_hi_hi_101 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_102;
  assign dataGroup_hi_hi_102 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_103;
  assign dataGroup_hi_hi_103 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_104;
  assign dataGroup_hi_hi_104 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_105;
  assign dataGroup_hi_hi_105 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_106;
  assign dataGroup_hi_hi_106 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_107;
  assign dataGroup_hi_hi_107 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_108;
  assign dataGroup_hi_hi_108 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_109;
  assign dataGroup_hi_hi_109 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_110;
  assign dataGroup_hi_hi_110 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_111;
  assign dataGroup_hi_hi_111 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_112;
  assign dataGroup_hi_hi_112 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_113;
  assign dataGroup_hi_hi_113 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_114;
  assign dataGroup_hi_hi_114 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_115;
  assign dataGroup_hi_hi_115 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_116;
  assign dataGroup_hi_hi_116 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_117;
  assign dataGroup_hi_hi_117 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_118;
  assign dataGroup_hi_hi_118 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_119;
  assign dataGroup_hi_hi_119 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_120;
  assign dataGroup_hi_hi_120 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_121;
  assign dataGroup_hi_hi_121 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_122;
  assign dataGroup_hi_hi_122 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_123;
  assign dataGroup_hi_hi_123 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_124;
  assign dataGroup_hi_hi_124 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_125;
  assign dataGroup_hi_hi_125 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_126;
  assign dataGroup_hi_hi_126 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_127;
  assign dataGroup_hi_hi_127 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_128;
  assign dataGroup_hi_hi_128 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_129;
  assign dataGroup_hi_hi_129 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_130;
  assign dataGroup_hi_hi_130 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_131;
  assign dataGroup_hi_hi_131 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_132;
  assign dataGroup_hi_hi_132 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_133;
  assign dataGroup_hi_hi_133 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_134;
  assign dataGroup_hi_hi_134 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_135;
  assign dataGroup_hi_hi_135 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_136;
  assign dataGroup_hi_hi_136 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_137;
  assign dataGroup_hi_hi_137 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_138;
  assign dataGroup_hi_hi_138 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_139;
  assign dataGroup_hi_hi_139 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_140;
  assign dataGroup_hi_hi_140 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_141;
  assign dataGroup_hi_hi_141 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_142;
  assign dataGroup_hi_hi_142 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_143;
  assign dataGroup_hi_hi_143 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_144;
  assign dataGroup_hi_hi_144 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_145;
  assign dataGroup_hi_hi_145 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_146;
  assign dataGroup_hi_hi_146 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_147;
  assign dataGroup_hi_hi_147 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_148;
  assign dataGroup_hi_hi_148 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_149;
  assign dataGroup_hi_hi_149 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_150;
  assign dataGroup_hi_hi_150 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_151;
  assign dataGroup_hi_hi_151 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_152;
  assign dataGroup_hi_hi_152 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_153;
  assign dataGroup_hi_hi_153 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_154;
  assign dataGroup_hi_hi_154 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_155;
  assign dataGroup_hi_hi_155 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_156;
  assign dataGroup_hi_hi_156 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_157;
  assign dataGroup_hi_hi_157 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_158;
  assign dataGroup_hi_hi_158 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_159;
  assign dataGroup_hi_hi_159 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_160;
  assign dataGroup_hi_hi_160 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_161;
  assign dataGroup_hi_hi_161 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_162;
  assign dataGroup_hi_hi_162 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_163;
  assign dataGroup_hi_hi_163 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_164;
  assign dataGroup_hi_hi_164 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_165;
  assign dataGroup_hi_hi_165 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_166;
  assign dataGroup_hi_hi_166 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_167;
  assign dataGroup_hi_hi_167 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_168;
  assign dataGroup_hi_hi_168 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_169;
  assign dataGroup_hi_hi_169 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_170;
  assign dataGroup_hi_hi_170 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_171;
  assign dataGroup_hi_hi_171 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_172;
  assign dataGroup_hi_hi_172 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_173;
  assign dataGroup_hi_hi_173 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_174;
  assign dataGroup_hi_hi_174 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_175;
  assign dataGroup_hi_hi_175 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_176;
  assign dataGroup_hi_hi_176 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_177;
  assign dataGroup_hi_hi_177 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_178;
  assign dataGroup_hi_hi_178 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_179;
  assign dataGroup_hi_hi_179 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_180;
  assign dataGroup_hi_hi_180 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_181;
  assign dataGroup_hi_hi_181 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_182;
  assign dataGroup_hi_hi_182 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_183;
  assign dataGroup_hi_hi_183 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_184;
  assign dataGroup_hi_hi_184 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_185;
  assign dataGroup_hi_hi_185 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_186;
  assign dataGroup_hi_hi_186 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_187;
  assign dataGroup_hi_hi_187 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_188;
  assign dataGroup_hi_hi_188 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_189;
  assign dataGroup_hi_hi_189 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_190;
  assign dataGroup_hi_hi_190 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_191;
  assign dataGroup_hi_hi_191 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_192;
  assign dataGroup_hi_hi_192 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_193;
  assign dataGroup_hi_hi_193 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_194;
  assign dataGroup_hi_hi_194 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_195;
  assign dataGroup_hi_hi_195 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_196;
  assign dataGroup_hi_hi_196 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_197;
  assign dataGroup_hi_hi_197 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_198;
  assign dataGroup_hi_hi_198 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_199;
  assign dataGroup_hi_hi_199 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_200;
  assign dataGroup_hi_hi_200 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_201;
  assign dataGroup_hi_hi_201 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_202;
  assign dataGroup_hi_hi_202 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_203;
  assign dataGroup_hi_hi_203 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_204;
  assign dataGroup_hi_hi_204 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_205;
  assign dataGroup_hi_hi_205 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_206;
  assign dataGroup_hi_hi_206 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_207;
  assign dataGroup_hi_hi_207 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_208;
  assign dataGroup_hi_hi_208 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_209;
  assign dataGroup_hi_hi_209 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_210;
  assign dataGroup_hi_hi_210 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_211;
  assign dataGroup_hi_hi_211 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_212;
  assign dataGroup_hi_hi_212 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_213;
  assign dataGroup_hi_hi_213 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_214;
  assign dataGroup_hi_hi_214 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_215;
  assign dataGroup_hi_hi_215 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_216;
  assign dataGroup_hi_hi_216 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_217;
  assign dataGroup_hi_hi_217 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_218;
  assign dataGroup_hi_hi_218 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_219;
  assign dataGroup_hi_hi_219 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_220;
  assign dataGroup_hi_hi_220 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_221;
  assign dataGroup_hi_hi_221 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_222;
  assign dataGroup_hi_hi_222 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_223;
  assign dataGroup_hi_hi_223 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_224;
  assign dataGroup_hi_hi_224 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_225;
  assign dataGroup_hi_hi_225 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_226;
  assign dataGroup_hi_hi_226 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_227;
  assign dataGroup_hi_hi_227 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_228;
  assign dataGroup_hi_hi_228 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_229;
  assign dataGroup_hi_hi_229 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_230;
  assign dataGroup_hi_hi_230 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_231;
  assign dataGroup_hi_hi_231 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_232;
  assign dataGroup_hi_hi_232 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_233;
  assign dataGroup_hi_hi_233 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_234;
  assign dataGroup_hi_hi_234 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_235;
  assign dataGroup_hi_hi_235 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_236;
  assign dataGroup_hi_hi_236 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_237;
  assign dataGroup_hi_hi_237 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_238;
  assign dataGroup_hi_hi_238 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_239;
  assign dataGroup_hi_hi_239 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_240;
  assign dataGroup_hi_hi_240 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_241;
  assign dataGroup_hi_hi_241 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_242;
  assign dataGroup_hi_hi_242 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_243;
  assign dataGroup_hi_hi_243 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_244;
  assign dataGroup_hi_hi_244 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_245;
  assign dataGroup_hi_hi_245 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_246;
  assign dataGroup_hi_hi_246 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_247;
  assign dataGroup_hi_hi_247 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_248;
  assign dataGroup_hi_hi_248 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_249;
  assign dataGroup_hi_hi_249 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_250;
  assign dataGroup_hi_hi_250 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_251;
  assign dataGroup_hi_hi_251 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_252;
  assign dataGroup_hi_hi_252 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_253;
  assign dataGroup_hi_hi_253 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_254;
  assign dataGroup_hi_hi_254 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_255;
  assign dataGroup_hi_hi_255 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_256;
  assign dataGroup_hi_hi_256 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_257;
  assign dataGroup_hi_hi_257 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_258;
  assign dataGroup_hi_hi_258 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_259;
  assign dataGroup_hi_hi_259 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_260;
  assign dataGroup_hi_hi_260 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_261;
  assign dataGroup_hi_hi_261 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_262;
  assign dataGroup_hi_hi_262 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_263;
  assign dataGroup_hi_hi_263 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_264;
  assign dataGroup_hi_hi_264 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_265;
  assign dataGroup_hi_hi_265 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_266;
  assign dataGroup_hi_hi_266 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_267;
  assign dataGroup_hi_hi_267 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_268;
  assign dataGroup_hi_hi_268 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_269;
  assign dataGroup_hi_hi_269 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_270;
  assign dataGroup_hi_hi_270 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_271;
  assign dataGroup_hi_hi_271 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_272;
  assign dataGroup_hi_hi_272 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_273;
  assign dataGroup_hi_hi_273 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_274;
  assign dataGroup_hi_hi_274 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_275;
  assign dataGroup_hi_hi_275 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_276;
  assign dataGroup_hi_hi_276 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_277;
  assign dataGroup_hi_hi_277 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_278;
  assign dataGroup_hi_hi_278 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_279;
  assign dataGroup_hi_hi_279 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_280;
  assign dataGroup_hi_hi_280 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_281;
  assign dataGroup_hi_hi_281 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_282;
  assign dataGroup_hi_hi_282 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_283;
  assign dataGroup_hi_hi_283 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_284;
  assign dataGroup_hi_hi_284 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_285;
  assign dataGroup_hi_hi_285 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_286;
  assign dataGroup_hi_hi_286 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_287;
  assign dataGroup_hi_hi_287 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_288;
  assign dataGroup_hi_hi_288 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_289;
  assign dataGroup_hi_hi_289 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_290;
  assign dataGroup_hi_hi_290 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_291;
  assign dataGroup_hi_hi_291 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_292;
  assign dataGroup_hi_hi_292 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_293;
  assign dataGroup_hi_hi_293 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_294;
  assign dataGroup_hi_hi_294 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_295;
  assign dataGroup_hi_hi_295 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_296;
  assign dataGroup_hi_hi_296 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_297;
  assign dataGroup_hi_hi_297 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_298;
  assign dataGroup_hi_hi_298 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_299;
  assign dataGroup_hi_hi_299 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_300;
  assign dataGroup_hi_hi_300 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_301;
  assign dataGroup_hi_hi_301 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_302;
  assign dataGroup_hi_hi_302 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_303;
  assign dataGroup_hi_hi_303 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_304;
  assign dataGroup_hi_hi_304 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_305;
  assign dataGroup_hi_hi_305 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_306;
  assign dataGroup_hi_hi_306 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_307;
  assign dataGroup_hi_hi_307 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_308;
  assign dataGroup_hi_hi_308 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_309;
  assign dataGroup_hi_hi_309 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_310;
  assign dataGroup_hi_hi_310 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_311;
  assign dataGroup_hi_hi_311 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_312;
  assign dataGroup_hi_hi_312 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_313;
  assign dataGroup_hi_hi_313 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_314;
  assign dataGroup_hi_hi_314 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_315;
  assign dataGroup_hi_hi_315 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_316;
  assign dataGroup_hi_hi_316 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_317;
  assign dataGroup_hi_hi_317 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_318;
  assign dataGroup_hi_hi_318 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_319;
  assign dataGroup_hi_hi_319 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_320;
  assign dataGroup_hi_hi_320 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_321;
  assign dataGroup_hi_hi_321 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_322;
  assign dataGroup_hi_hi_322 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_323;
  assign dataGroup_hi_hi_323 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_324;
  assign dataGroup_hi_hi_324 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_325;
  assign dataGroup_hi_hi_325 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_326;
  assign dataGroup_hi_hi_326 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_327;
  assign dataGroup_hi_hi_327 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_328;
  assign dataGroup_hi_hi_328 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_329;
  assign dataGroup_hi_hi_329 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_330;
  assign dataGroup_hi_hi_330 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_331;
  assign dataGroup_hi_hi_331 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_332;
  assign dataGroup_hi_hi_332 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_333;
  assign dataGroup_hi_hi_333 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_334;
  assign dataGroup_hi_hi_334 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_335;
  assign dataGroup_hi_hi_335 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_336;
  assign dataGroup_hi_hi_336 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_337;
  assign dataGroup_hi_hi_337 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_338;
  assign dataGroup_hi_hi_338 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_339;
  assign dataGroup_hi_hi_339 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_340;
  assign dataGroup_hi_hi_340 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_341;
  assign dataGroup_hi_hi_341 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_342;
  assign dataGroup_hi_hi_342 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_343;
  assign dataGroup_hi_hi_343 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_344;
  assign dataGroup_hi_hi_344 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_345;
  assign dataGroup_hi_hi_345 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_346;
  assign dataGroup_hi_hi_346 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_347;
  assign dataGroup_hi_hi_347 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_348;
  assign dataGroup_hi_hi_348 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_349;
  assign dataGroup_hi_hi_349 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_350;
  assign dataGroup_hi_hi_350 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_351;
  assign dataGroup_hi_hi_351 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_352;
  assign dataGroup_hi_hi_352 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_353;
  assign dataGroup_hi_hi_353 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_354;
  assign dataGroup_hi_hi_354 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_355;
  assign dataGroup_hi_hi_355 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_356;
  assign dataGroup_hi_hi_356 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_357;
  assign dataGroup_hi_hi_357 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_358;
  assign dataGroup_hi_hi_358 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_359;
  assign dataGroup_hi_hi_359 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_360;
  assign dataGroup_hi_hi_360 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_361;
  assign dataGroup_hi_hi_361 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_362;
  assign dataGroup_hi_hi_362 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_363;
  assign dataGroup_hi_hi_363 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_364;
  assign dataGroup_hi_hi_364 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_365;
  assign dataGroup_hi_hi_365 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_366;
  assign dataGroup_hi_hi_366 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_367;
  assign dataGroup_hi_hi_367 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_368;
  assign dataGroup_hi_hi_368 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_369;
  assign dataGroup_hi_hi_369 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_370;
  assign dataGroup_hi_hi_370 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_371;
  assign dataGroup_hi_hi_371 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_372;
  assign dataGroup_hi_hi_372 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_373;
  assign dataGroup_hi_hi_373 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_374;
  assign dataGroup_hi_hi_374 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_375;
  assign dataGroup_hi_hi_375 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_376;
  assign dataGroup_hi_hi_376 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_377;
  assign dataGroup_hi_hi_377 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_378;
  assign dataGroup_hi_hi_378 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_379;
  assign dataGroup_hi_hi_379 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_380;
  assign dataGroup_hi_hi_380 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_381;
  assign dataGroup_hi_hi_381 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_382;
  assign dataGroup_hi_hi_382 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_383;
  assign dataGroup_hi_hi_383 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_384;
  assign dataGroup_hi_hi_384 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_385;
  assign dataGroup_hi_hi_385 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_386;
  assign dataGroup_hi_hi_386 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_387;
  assign dataGroup_hi_hi_387 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_388;
  assign dataGroup_hi_hi_388 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_389;
  assign dataGroup_hi_hi_389 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_390;
  assign dataGroup_hi_hi_390 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_391;
  assign dataGroup_hi_hi_391 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_392;
  assign dataGroup_hi_hi_392 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_393;
  assign dataGroup_hi_hi_393 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_394;
  assign dataGroup_hi_hi_394 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_395;
  assign dataGroup_hi_hi_395 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_396;
  assign dataGroup_hi_hi_396 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_397;
  assign dataGroup_hi_hi_397 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_398;
  assign dataGroup_hi_hi_398 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_399;
  assign dataGroup_hi_hi_399 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_400;
  assign dataGroup_hi_hi_400 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_401;
  assign dataGroup_hi_hi_401 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_402;
  assign dataGroup_hi_hi_402 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_403;
  assign dataGroup_hi_hi_403 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_404;
  assign dataGroup_hi_hi_404 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_405;
  assign dataGroup_hi_hi_405 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_406;
  assign dataGroup_hi_hi_406 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_407;
  assign dataGroup_hi_hi_407 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_408;
  assign dataGroup_hi_hi_408 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_409;
  assign dataGroup_hi_hi_409 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_410;
  assign dataGroup_hi_hi_410 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_411;
  assign dataGroup_hi_hi_411 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_412;
  assign dataGroup_hi_hi_412 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_413;
  assign dataGroup_hi_hi_413 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_414;
  assign dataGroup_hi_hi_414 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_415;
  assign dataGroup_hi_hi_415 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_416;
  assign dataGroup_hi_hi_416 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_417;
  assign dataGroup_hi_hi_417 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_418;
  assign dataGroup_hi_hi_418 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_419;
  assign dataGroup_hi_hi_419 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_420;
  assign dataGroup_hi_hi_420 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_421;
  assign dataGroup_hi_hi_421 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_422;
  assign dataGroup_hi_hi_422 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_423;
  assign dataGroup_hi_hi_423 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_424;
  assign dataGroup_hi_hi_424 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_425;
  assign dataGroup_hi_hi_425 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_426;
  assign dataGroup_hi_hi_426 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_427;
  assign dataGroup_hi_hi_427 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_428;
  assign dataGroup_hi_hi_428 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_429;
  assign dataGroup_hi_hi_429 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_430;
  assign dataGroup_hi_hi_430 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_431;
  assign dataGroup_hi_hi_431 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_432;
  assign dataGroup_hi_hi_432 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_433;
  assign dataGroup_hi_hi_433 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_434;
  assign dataGroup_hi_hi_434 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_435;
  assign dataGroup_hi_hi_435 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_436;
  assign dataGroup_hi_hi_436 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_437;
  assign dataGroup_hi_hi_437 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_438;
  assign dataGroup_hi_hi_438 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_439;
  assign dataGroup_hi_hi_439 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_440;
  assign dataGroup_hi_hi_440 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_441;
  assign dataGroup_hi_hi_441 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_442;
  assign dataGroup_hi_hi_442 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_443;
  assign dataGroup_hi_hi_443 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_444;
  assign dataGroup_hi_hi_444 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_445;
  assign dataGroup_hi_hi_445 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_446;
  assign dataGroup_hi_hi_446 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_447;
  assign dataGroup_hi_hi_447 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_448;
  assign dataGroup_hi_hi_448 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_449;
  assign dataGroup_hi_hi_449 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_450;
  assign dataGroup_hi_hi_450 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_451;
  assign dataGroup_hi_hi_451 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_452;
  assign dataGroup_hi_hi_452 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_453;
  assign dataGroup_hi_hi_453 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_454;
  assign dataGroup_hi_hi_454 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_455;
  assign dataGroup_hi_hi_455 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_456;
  assign dataGroup_hi_hi_456 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_457;
  assign dataGroup_hi_hi_457 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_458;
  assign dataGroup_hi_hi_458 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_459;
  assign dataGroup_hi_hi_459 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_460;
  assign dataGroup_hi_hi_460 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_461;
  assign dataGroup_hi_hi_461 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_462;
  assign dataGroup_hi_hi_462 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_463;
  assign dataGroup_hi_hi_463 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_464;
  assign dataGroup_hi_hi_464 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_465;
  assign dataGroup_hi_hi_465 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_466;
  assign dataGroup_hi_hi_466 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_467;
  assign dataGroup_hi_hi_467 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_468;
  assign dataGroup_hi_hi_468 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_469;
  assign dataGroup_hi_hi_469 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_470;
  assign dataGroup_hi_hi_470 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_471;
  assign dataGroup_hi_hi_471 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_472;
  assign dataGroup_hi_hi_472 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_473;
  assign dataGroup_hi_hi_473 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_474;
  assign dataGroup_hi_hi_474 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_475;
  assign dataGroup_hi_hi_475 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_476;
  assign dataGroup_hi_hi_476 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_477;
  assign dataGroup_hi_hi_477 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_478;
  assign dataGroup_hi_hi_478 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_479;
  assign dataGroup_hi_hi_479 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_480;
  assign dataGroup_hi_hi_480 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_481;
  assign dataGroup_hi_hi_481 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_482;
  assign dataGroup_hi_hi_482 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_483;
  assign dataGroup_hi_hi_483 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_484;
  assign dataGroup_hi_hi_484 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_485;
  assign dataGroup_hi_hi_485 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_486;
  assign dataGroup_hi_hi_486 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_487;
  assign dataGroup_hi_hi_487 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_488;
  assign dataGroup_hi_hi_488 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_489;
  assign dataGroup_hi_hi_489 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_490;
  assign dataGroup_hi_hi_490 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_491;
  assign dataGroup_hi_hi_491 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_492;
  assign dataGroup_hi_hi_492 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_493;
  assign dataGroup_hi_hi_493 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_494;
  assign dataGroup_hi_hi_494 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_495;
  assign dataGroup_hi_hi_495 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_496;
  assign dataGroup_hi_hi_496 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_497;
  assign dataGroup_hi_hi_497 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_498;
  assign dataGroup_hi_hi_498 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_499;
  assign dataGroup_hi_hi_499 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_500;
  assign dataGroup_hi_hi_500 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_501;
  assign dataGroup_hi_hi_501 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_502;
  assign dataGroup_hi_hi_502 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_503;
  assign dataGroup_hi_hi_503 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_504;
  assign dataGroup_hi_hi_504 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_505;
  assign dataGroup_hi_hi_505 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_506;
  assign dataGroup_hi_hi_506 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_507;
  assign dataGroup_hi_hi_507 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_508;
  assign dataGroup_hi_hi_508 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_509;
  assign dataGroup_hi_hi_509 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_510;
  assign dataGroup_hi_hi_510 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_511;
  assign dataGroup_hi_hi_511 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_512;
  assign dataGroup_hi_hi_512 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_513;
  assign dataGroup_hi_hi_513 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_514;
  assign dataGroup_hi_hi_514 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_515;
  assign dataGroup_hi_hi_515 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_516;
  assign dataGroup_hi_hi_516 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_517;
  assign dataGroup_hi_hi_517 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_518;
  assign dataGroup_hi_hi_518 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_519;
  assign dataGroup_hi_hi_519 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_520;
  assign dataGroup_hi_hi_520 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_521;
  assign dataGroup_hi_hi_521 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_522;
  assign dataGroup_hi_hi_522 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_523;
  assign dataGroup_hi_hi_523 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_524;
  assign dataGroup_hi_hi_524 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_525;
  assign dataGroup_hi_hi_525 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_526;
  assign dataGroup_hi_hi_526 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_527;
  assign dataGroup_hi_hi_527 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_528;
  assign dataGroup_hi_hi_528 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_529;
  assign dataGroup_hi_hi_529 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_530;
  assign dataGroup_hi_hi_530 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_531;
  assign dataGroup_hi_hi_531 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_532;
  assign dataGroup_hi_hi_532 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_533;
  assign dataGroup_hi_hi_533 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_534;
  assign dataGroup_hi_hi_534 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_535;
  assign dataGroup_hi_hi_535 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_536;
  assign dataGroup_hi_hi_536 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_537;
  assign dataGroup_hi_hi_537 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_538;
  assign dataGroup_hi_hi_538 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_539;
  assign dataGroup_hi_hi_539 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_540;
  assign dataGroup_hi_hi_540 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_541;
  assign dataGroup_hi_hi_541 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_542;
  assign dataGroup_hi_hi_542 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_543;
  assign dataGroup_hi_hi_543 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_544;
  assign dataGroup_hi_hi_544 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_545;
  assign dataGroup_hi_hi_545 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_546;
  assign dataGroup_hi_hi_546 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_547;
  assign dataGroup_hi_hi_547 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_548;
  assign dataGroup_hi_hi_548 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_549;
  assign dataGroup_hi_hi_549 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_550;
  assign dataGroup_hi_hi_550 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_551;
  assign dataGroup_hi_hi_551 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_552;
  assign dataGroup_hi_hi_552 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_553;
  assign dataGroup_hi_hi_553 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_554;
  assign dataGroup_hi_hi_554 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_555;
  assign dataGroup_hi_hi_555 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_556;
  assign dataGroup_hi_hi_556 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_557;
  assign dataGroup_hi_hi_557 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_558;
  assign dataGroup_hi_hi_558 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_559;
  assign dataGroup_hi_hi_559 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_560;
  assign dataGroup_hi_hi_560 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_561;
  assign dataGroup_hi_hi_561 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_562;
  assign dataGroup_hi_hi_562 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_563;
  assign dataGroup_hi_hi_563 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_564;
  assign dataGroup_hi_hi_564 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_565;
  assign dataGroup_hi_hi_565 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_566;
  assign dataGroup_hi_hi_566 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_567;
  assign dataGroup_hi_hi_567 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_568;
  assign dataGroup_hi_hi_568 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_569;
  assign dataGroup_hi_hi_569 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_570;
  assign dataGroup_hi_hi_570 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_571;
  assign dataGroup_hi_hi_571 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_572;
  assign dataGroup_hi_hi_572 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_573;
  assign dataGroup_hi_hi_573 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_574;
  assign dataGroup_hi_hi_574 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_575;
  assign dataGroup_hi_hi_575 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_576;
  assign dataGroup_hi_hi_576 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_577;
  assign dataGroup_hi_hi_577 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_578;
  assign dataGroup_hi_hi_578 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_579;
  assign dataGroup_hi_hi_579 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_580;
  assign dataGroup_hi_hi_580 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_581;
  assign dataGroup_hi_hi_581 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_582;
  assign dataGroup_hi_hi_582 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_583;
  assign dataGroup_hi_hi_583 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_584;
  assign dataGroup_hi_hi_584 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_585;
  assign dataGroup_hi_hi_585 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_586;
  assign dataGroup_hi_hi_586 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_587;
  assign dataGroup_hi_hi_587 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_588;
  assign dataGroup_hi_hi_588 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_589;
  assign dataGroup_hi_hi_589 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_590;
  assign dataGroup_hi_hi_590 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_591;
  assign dataGroup_hi_hi_591 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_592;
  assign dataGroup_hi_hi_592 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_593;
  assign dataGroup_hi_hi_593 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_594;
  assign dataGroup_hi_hi_594 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_595;
  assign dataGroup_hi_hi_595 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_596;
  assign dataGroup_hi_hi_596 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_597;
  assign dataGroup_hi_hi_597 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_598;
  assign dataGroup_hi_hi_598 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_599;
  assign dataGroup_hi_hi_599 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_600;
  assign dataGroup_hi_hi_600 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_601;
  assign dataGroup_hi_hi_601 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_602;
  assign dataGroup_hi_hi_602 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_603;
  assign dataGroup_hi_hi_603 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_604;
  assign dataGroup_hi_hi_604 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_605;
  assign dataGroup_hi_hi_605 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_606;
  assign dataGroup_hi_hi_606 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_607;
  assign dataGroup_hi_hi_607 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_608;
  assign dataGroup_hi_hi_608 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_609;
  assign dataGroup_hi_hi_609 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_610;
  assign dataGroup_hi_hi_610 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_611;
  assign dataGroup_hi_hi_611 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_612;
  assign dataGroup_hi_hi_612 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_613;
  assign dataGroup_hi_hi_613 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_614;
  assign dataGroup_hi_hi_614 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_615;
  assign dataGroup_hi_hi_615 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_616;
  assign dataGroup_hi_hi_616 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_617;
  assign dataGroup_hi_hi_617 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_618;
  assign dataGroup_hi_hi_618 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_619;
  assign dataGroup_hi_hi_619 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_620;
  assign dataGroup_hi_hi_620 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_621;
  assign dataGroup_hi_hi_621 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_622;
  assign dataGroup_hi_hi_622 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_623;
  assign dataGroup_hi_hi_623 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_624;
  assign dataGroup_hi_hi_624 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_625;
  assign dataGroup_hi_hi_625 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_626;
  assign dataGroup_hi_hi_626 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_627;
  assign dataGroup_hi_hi_627 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_628;
  assign dataGroup_hi_hi_628 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_629;
  assign dataGroup_hi_hi_629 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_630;
  assign dataGroup_hi_hi_630 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_631;
  assign dataGroup_hi_hi_631 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_632;
  assign dataGroup_hi_hi_632 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_633;
  assign dataGroup_hi_hi_633 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_634;
  assign dataGroup_hi_hi_634 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_635;
  assign dataGroup_hi_hi_635 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_636;
  assign dataGroup_hi_hi_636 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_637;
  assign dataGroup_hi_hi_637 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_638;
  assign dataGroup_hi_hi_638 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_639;
  assign dataGroup_hi_hi_639 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_640;
  assign dataGroup_hi_hi_640 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_641;
  assign dataGroup_hi_hi_641 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_642;
  assign dataGroup_hi_hi_642 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_643;
  assign dataGroup_hi_hi_643 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_644;
  assign dataGroup_hi_hi_644 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_645;
  assign dataGroup_hi_hi_645 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_646;
  assign dataGroup_hi_hi_646 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_647;
  assign dataGroup_hi_hi_647 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_648;
  assign dataGroup_hi_hi_648 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_649;
  assign dataGroup_hi_hi_649 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_650;
  assign dataGroup_hi_hi_650 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_651;
  assign dataGroup_hi_hi_651 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_652;
  assign dataGroup_hi_hi_652 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_653;
  assign dataGroup_hi_hi_653 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_654;
  assign dataGroup_hi_hi_654 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_655;
  assign dataGroup_hi_hi_655 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_656;
  assign dataGroup_hi_hi_656 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_657;
  assign dataGroup_hi_hi_657 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_658;
  assign dataGroup_hi_hi_658 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_659;
  assign dataGroup_hi_hi_659 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_660;
  assign dataGroup_hi_hi_660 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_661;
  assign dataGroup_hi_hi_661 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_662;
  assign dataGroup_hi_hi_662 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_663;
  assign dataGroup_hi_hi_663 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_664;
  assign dataGroup_hi_hi_664 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_665;
  assign dataGroup_hi_hi_665 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_666;
  assign dataGroup_hi_hi_666 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_667;
  assign dataGroup_hi_hi_667 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_668;
  assign dataGroup_hi_hi_668 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_669;
  assign dataGroup_hi_hi_669 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_670;
  assign dataGroup_hi_hi_670 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_671;
  assign dataGroup_hi_hi_671 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_672;
  assign dataGroup_hi_hi_672 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_673;
  assign dataGroup_hi_hi_673 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_674;
  assign dataGroup_hi_hi_674 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_675;
  assign dataGroup_hi_hi_675 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_676;
  assign dataGroup_hi_hi_676 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_677;
  assign dataGroup_hi_hi_677 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_678;
  assign dataGroup_hi_hi_678 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_679;
  assign dataGroup_hi_hi_679 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_680;
  assign dataGroup_hi_hi_680 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_681;
  assign dataGroup_hi_hi_681 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_682;
  assign dataGroup_hi_hi_682 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_683;
  assign dataGroup_hi_hi_683 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_684;
  assign dataGroup_hi_hi_684 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_685;
  assign dataGroup_hi_hi_685 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_686;
  assign dataGroup_hi_hi_686 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_687;
  assign dataGroup_hi_hi_687 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_688;
  assign dataGroup_hi_hi_688 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_689;
  assign dataGroup_hi_hi_689 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_690;
  assign dataGroup_hi_hi_690 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_691;
  assign dataGroup_hi_hi_691 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_692;
  assign dataGroup_hi_hi_692 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_693;
  assign dataGroup_hi_hi_693 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_694;
  assign dataGroup_hi_hi_694 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_695;
  assign dataGroup_hi_hi_695 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_696;
  assign dataGroup_hi_hi_696 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_697;
  assign dataGroup_hi_hi_697 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_698;
  assign dataGroup_hi_hi_698 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_699;
  assign dataGroup_hi_hi_699 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_700;
  assign dataGroup_hi_hi_700 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_701;
  assign dataGroup_hi_hi_701 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_702;
  assign dataGroup_hi_hi_702 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_703;
  assign dataGroup_hi_hi_703 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_704;
  assign dataGroup_hi_hi_704 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_705;
  assign dataGroup_hi_hi_705 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_706;
  assign dataGroup_hi_hi_706 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_707;
  assign dataGroup_hi_hi_707 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_708;
  assign dataGroup_hi_hi_708 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_709;
  assign dataGroup_hi_hi_709 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_710;
  assign dataGroup_hi_hi_710 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_711;
  assign dataGroup_hi_hi_711 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_712;
  assign dataGroup_hi_hi_712 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_713;
  assign dataGroup_hi_hi_713 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_714;
  assign dataGroup_hi_hi_714 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_715;
  assign dataGroup_hi_hi_715 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_716;
  assign dataGroup_hi_hi_716 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_717;
  assign dataGroup_hi_hi_717 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_718;
  assign dataGroup_hi_hi_718 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_719;
  assign dataGroup_hi_hi_719 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_720;
  assign dataGroup_hi_hi_720 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_721;
  assign dataGroup_hi_hi_721 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_722;
  assign dataGroup_hi_hi_722 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_723;
  assign dataGroup_hi_hi_723 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_724;
  assign dataGroup_hi_hi_724 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_725;
  assign dataGroup_hi_hi_725 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_726;
  assign dataGroup_hi_hi_726 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_727;
  assign dataGroup_hi_hi_727 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_728;
  assign dataGroup_hi_hi_728 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_729;
  assign dataGroup_hi_hi_729 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_730;
  assign dataGroup_hi_hi_730 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_731;
  assign dataGroup_hi_hi_731 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_732;
  assign dataGroup_hi_hi_732 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_733;
  assign dataGroup_hi_hi_733 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_734;
  assign dataGroup_hi_hi_734 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_735;
  assign dataGroup_hi_hi_735 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_736;
  assign dataGroup_hi_hi_736 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_737;
  assign dataGroup_hi_hi_737 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_738;
  assign dataGroup_hi_hi_738 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_739;
  assign dataGroup_hi_hi_739 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_740;
  assign dataGroup_hi_hi_740 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_741;
  assign dataGroup_hi_hi_741 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_742;
  assign dataGroup_hi_hi_742 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_743;
  assign dataGroup_hi_hi_743 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_744;
  assign dataGroup_hi_hi_744 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_745;
  assign dataGroup_hi_hi_745 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_746;
  assign dataGroup_hi_hi_746 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_747;
  assign dataGroup_hi_hi_747 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_748;
  assign dataGroup_hi_hi_748 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_749;
  assign dataGroup_hi_hi_749 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_750;
  assign dataGroup_hi_hi_750 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_751;
  assign dataGroup_hi_hi_751 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_752;
  assign dataGroup_hi_hi_752 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_753;
  assign dataGroup_hi_hi_753 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_754;
  assign dataGroup_hi_hi_754 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_755;
  assign dataGroup_hi_hi_755 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_756;
  assign dataGroup_hi_hi_756 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_757;
  assign dataGroup_hi_hi_757 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_758;
  assign dataGroup_hi_hi_758 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_759;
  assign dataGroup_hi_hi_759 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_760;
  assign dataGroup_hi_hi_760 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_761;
  assign dataGroup_hi_hi_761 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_762;
  assign dataGroup_hi_hi_762 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_763;
  assign dataGroup_hi_hi_763 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_764;
  assign dataGroup_hi_hi_764 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_765;
  assign dataGroup_hi_hi_765 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_766;
  assign dataGroup_hi_hi_766 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_767;
  assign dataGroup_hi_hi_767 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_768;
  assign dataGroup_hi_hi_768 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_769;
  assign dataGroup_hi_hi_769 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_770;
  assign dataGroup_hi_hi_770 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_771;
  assign dataGroup_hi_hi_771 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_772;
  assign dataGroup_hi_hi_772 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_773;
  assign dataGroup_hi_hi_773 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_774;
  assign dataGroup_hi_hi_774 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_775;
  assign dataGroup_hi_hi_775 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_776;
  assign dataGroup_hi_hi_776 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_777;
  assign dataGroup_hi_hi_777 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_778;
  assign dataGroup_hi_hi_778 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_779;
  assign dataGroup_hi_hi_779 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_780;
  assign dataGroup_hi_hi_780 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_781;
  assign dataGroup_hi_hi_781 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_782;
  assign dataGroup_hi_hi_782 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_783;
  assign dataGroup_hi_hi_783 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_784;
  assign dataGroup_hi_hi_784 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_785;
  assign dataGroup_hi_hi_785 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_786;
  assign dataGroup_hi_hi_786 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_787;
  assign dataGroup_hi_hi_787 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_788;
  assign dataGroup_hi_hi_788 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_789;
  assign dataGroup_hi_hi_789 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_790;
  assign dataGroup_hi_hi_790 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_791;
  assign dataGroup_hi_hi_791 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_792;
  assign dataGroup_hi_hi_792 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_793;
  assign dataGroup_hi_hi_793 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_794;
  assign dataGroup_hi_hi_794 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_795;
  assign dataGroup_hi_hi_795 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_796;
  assign dataGroup_hi_hi_796 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_797;
  assign dataGroup_hi_hi_797 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_798;
  assign dataGroup_hi_hi_798 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_799;
  assign dataGroup_hi_hi_799 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_800;
  assign dataGroup_hi_hi_800 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_801;
  assign dataGroup_hi_hi_801 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_802;
  assign dataGroup_hi_hi_802 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_803;
  assign dataGroup_hi_hi_803 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_804;
  assign dataGroup_hi_hi_804 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_805;
  assign dataGroup_hi_hi_805 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_806;
  assign dataGroup_hi_hi_806 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_807;
  assign dataGroup_hi_hi_807 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_808;
  assign dataGroup_hi_hi_808 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_809;
  assign dataGroup_hi_hi_809 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_810;
  assign dataGroup_hi_hi_810 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_811;
  assign dataGroup_hi_hi_811 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_812;
  assign dataGroup_hi_hi_812 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_813;
  assign dataGroup_hi_hi_813 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_814;
  assign dataGroup_hi_hi_814 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_815;
  assign dataGroup_hi_hi_815 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_816;
  assign dataGroup_hi_hi_816 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_817;
  assign dataGroup_hi_hi_817 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_818;
  assign dataGroup_hi_hi_818 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_819;
  assign dataGroup_hi_hi_819 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_820;
  assign dataGroup_hi_hi_820 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_821;
  assign dataGroup_hi_hi_821 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_822;
  assign dataGroup_hi_hi_822 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_823;
  assign dataGroup_hi_hi_823 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_824;
  assign dataGroup_hi_hi_824 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_825;
  assign dataGroup_hi_hi_825 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_826;
  assign dataGroup_hi_hi_826 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_827;
  assign dataGroup_hi_hi_827 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_828;
  assign dataGroup_hi_hi_828 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_829;
  assign dataGroup_hi_hi_829 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_830;
  assign dataGroup_hi_hi_830 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_831;
  assign dataGroup_hi_hi_831 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_832;
  assign dataGroup_hi_hi_832 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_833;
  assign dataGroup_hi_hi_833 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_834;
  assign dataGroup_hi_hi_834 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_835;
  assign dataGroup_hi_hi_835 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_836;
  assign dataGroup_hi_hi_836 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_837;
  assign dataGroup_hi_hi_837 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_838;
  assign dataGroup_hi_hi_838 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_839;
  assign dataGroup_hi_hi_839 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_840;
  assign dataGroup_hi_hi_840 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_841;
  assign dataGroup_hi_hi_841 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_842;
  assign dataGroup_hi_hi_842 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_843;
  assign dataGroup_hi_hi_843 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_844;
  assign dataGroup_hi_hi_844 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_845;
  assign dataGroup_hi_hi_845 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_846;
  assign dataGroup_hi_hi_846 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_847;
  assign dataGroup_hi_hi_847 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_848;
  assign dataGroup_hi_hi_848 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_849;
  assign dataGroup_hi_hi_849 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_850;
  assign dataGroup_hi_hi_850 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_851;
  assign dataGroup_hi_hi_851 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_852;
  assign dataGroup_hi_hi_852 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_853;
  assign dataGroup_hi_hi_853 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_854;
  assign dataGroup_hi_hi_854 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_855;
  assign dataGroup_hi_hi_855 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_856;
  assign dataGroup_hi_hi_856 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_857;
  assign dataGroup_hi_hi_857 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_858;
  assign dataGroup_hi_hi_858 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_859;
  assign dataGroup_hi_hi_859 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_860;
  assign dataGroup_hi_hi_860 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_861;
  assign dataGroup_hi_hi_861 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_862;
  assign dataGroup_hi_hi_862 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_863;
  assign dataGroup_hi_hi_863 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_864;
  assign dataGroup_hi_hi_864 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_865;
  assign dataGroup_hi_hi_865 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_866;
  assign dataGroup_hi_hi_866 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_867;
  assign dataGroup_hi_hi_867 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_868;
  assign dataGroup_hi_hi_868 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_869;
  assign dataGroup_hi_hi_869 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_870;
  assign dataGroup_hi_hi_870 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_871;
  assign dataGroup_hi_hi_871 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_872;
  assign dataGroup_hi_hi_872 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_873;
  assign dataGroup_hi_hi_873 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_874;
  assign dataGroup_hi_hi_874 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_875;
  assign dataGroup_hi_hi_875 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_876;
  assign dataGroup_hi_hi_876 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_877;
  assign dataGroup_hi_hi_877 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_878;
  assign dataGroup_hi_hi_878 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_879;
  assign dataGroup_hi_hi_879 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_880;
  assign dataGroup_hi_hi_880 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_881;
  assign dataGroup_hi_hi_881 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_882;
  assign dataGroup_hi_hi_882 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_883;
  assign dataGroup_hi_hi_883 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_884;
  assign dataGroup_hi_hi_884 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_885;
  assign dataGroup_hi_hi_885 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_886;
  assign dataGroup_hi_hi_886 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_887;
  assign dataGroup_hi_hi_887 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_888;
  assign dataGroup_hi_hi_888 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_889;
  assign dataGroup_hi_hi_889 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_890;
  assign dataGroup_hi_hi_890 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_891;
  assign dataGroup_hi_hi_891 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_892;
  assign dataGroup_hi_hi_892 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_893;
  assign dataGroup_hi_hi_893 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_894;
  assign dataGroup_hi_hi_894 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_895;
  assign dataGroup_hi_hi_895 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_896;
  assign dataGroup_hi_hi_896 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_897;
  assign dataGroup_hi_hi_897 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_898;
  assign dataGroup_hi_hi_898 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_899;
  assign dataGroup_hi_hi_899 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_900;
  assign dataGroup_hi_hi_900 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_901;
  assign dataGroup_hi_hi_901 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_902;
  assign dataGroup_hi_hi_902 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_903;
  assign dataGroup_hi_hi_903 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_904;
  assign dataGroup_hi_hi_904 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_905;
  assign dataGroup_hi_hi_905 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_906;
  assign dataGroup_hi_hi_906 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_907;
  assign dataGroup_hi_hi_907 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_908;
  assign dataGroup_hi_hi_908 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_909;
  assign dataGroup_hi_hi_909 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_910;
  assign dataGroup_hi_hi_910 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_911;
  assign dataGroup_hi_hi_911 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_912;
  assign dataGroup_hi_hi_912 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_913;
  assign dataGroup_hi_hi_913 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_914;
  assign dataGroup_hi_hi_914 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_915;
  assign dataGroup_hi_hi_915 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_916;
  assign dataGroup_hi_hi_916 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_917;
  assign dataGroup_hi_hi_917 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_918;
  assign dataGroup_hi_hi_918 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_919;
  assign dataGroup_hi_hi_919 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_920;
  assign dataGroup_hi_hi_920 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_921;
  assign dataGroup_hi_hi_921 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_922;
  assign dataGroup_hi_hi_922 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_923;
  assign dataGroup_hi_hi_923 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_924;
  assign dataGroup_hi_hi_924 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_925;
  assign dataGroup_hi_hi_925 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_926;
  assign dataGroup_hi_hi_926 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_927;
  assign dataGroup_hi_hi_927 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_928;
  assign dataGroup_hi_hi_928 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_929;
  assign dataGroup_hi_hi_929 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_930;
  assign dataGroup_hi_hi_930 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_931;
  assign dataGroup_hi_hi_931 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_932;
  assign dataGroup_hi_hi_932 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_933;
  assign dataGroup_hi_hi_933 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_934;
  assign dataGroup_hi_hi_934 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_935;
  assign dataGroup_hi_hi_935 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_936;
  assign dataGroup_hi_hi_936 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_937;
  assign dataGroup_hi_hi_937 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_938;
  assign dataGroup_hi_hi_938 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_939;
  assign dataGroup_hi_hi_939 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_940;
  assign dataGroup_hi_hi_940 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_941;
  assign dataGroup_hi_hi_941 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_942;
  assign dataGroup_hi_hi_942 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_943;
  assign dataGroup_hi_hi_943 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_944;
  assign dataGroup_hi_hi_944 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_945;
  assign dataGroup_hi_hi_945 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_946;
  assign dataGroup_hi_hi_946 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_947;
  assign dataGroup_hi_hi_947 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_948;
  assign dataGroup_hi_hi_948 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_949;
  assign dataGroup_hi_hi_949 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_950;
  assign dataGroup_hi_hi_950 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_951;
  assign dataGroup_hi_hi_951 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_952;
  assign dataGroup_hi_hi_952 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_953;
  assign dataGroup_hi_hi_953 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_954;
  assign dataGroup_hi_hi_954 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_955;
  assign dataGroup_hi_hi_955 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_956;
  assign dataGroup_hi_hi_956 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_957;
  assign dataGroup_hi_hi_957 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_958;
  assign dataGroup_hi_hi_958 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_959;
  assign dataGroup_hi_hi_959 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_960;
  assign dataGroup_hi_hi_960 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_961;
  assign dataGroup_hi_hi_961 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_962;
  assign dataGroup_hi_hi_962 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_963;
  assign dataGroup_hi_hi_963 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_964;
  assign dataGroup_hi_hi_964 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_965;
  assign dataGroup_hi_hi_965 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_966;
  assign dataGroup_hi_hi_966 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_967;
  assign dataGroup_hi_hi_967 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_968;
  assign dataGroup_hi_hi_968 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_969;
  assign dataGroup_hi_hi_969 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_970;
  assign dataGroup_hi_hi_970 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_971;
  assign dataGroup_hi_hi_971 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_972;
  assign dataGroup_hi_hi_972 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_973;
  assign dataGroup_hi_hi_973 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_974;
  assign dataGroup_hi_hi_974 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_975;
  assign dataGroup_hi_hi_975 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_976;
  assign dataGroup_hi_hi_976 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_977;
  assign dataGroup_hi_hi_977 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_978;
  assign dataGroup_hi_hi_978 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_979;
  assign dataGroup_hi_hi_979 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_980;
  assign dataGroup_hi_hi_980 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_981;
  assign dataGroup_hi_hi_981 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_982;
  assign dataGroup_hi_hi_982 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_983;
  assign dataGroup_hi_hi_983 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_984;
  assign dataGroup_hi_hi_984 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_985;
  assign dataGroup_hi_hi_985 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_986;
  assign dataGroup_hi_hi_986 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_987;
  assign dataGroup_hi_hi_987 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_988;
  assign dataGroup_hi_hi_988 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_989;
  assign dataGroup_hi_hi_989 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_990;
  assign dataGroup_hi_hi_990 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_991;
  assign dataGroup_hi_hi_991 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_992;
  assign dataGroup_hi_hi_992 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_993;
  assign dataGroup_hi_hi_993 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_994;
  assign dataGroup_hi_hi_994 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_995;
  assign dataGroup_hi_hi_995 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_996;
  assign dataGroup_hi_hi_996 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_997;
  assign dataGroup_hi_hi_997 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_998;
  assign dataGroup_hi_hi_998 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_999;
  assign dataGroup_hi_hi_999 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1000;
  assign dataGroup_hi_hi_1000 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1001;
  assign dataGroup_hi_hi_1001 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1002;
  assign dataGroup_hi_hi_1002 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1003;
  assign dataGroup_hi_hi_1003 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1004;
  assign dataGroup_hi_hi_1004 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1005;
  assign dataGroup_hi_hi_1005 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1006;
  assign dataGroup_hi_hi_1006 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1007;
  assign dataGroup_hi_hi_1007 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1008;
  assign dataGroup_hi_hi_1008 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1009;
  assign dataGroup_hi_hi_1009 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1010;
  assign dataGroup_hi_hi_1010 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1011;
  assign dataGroup_hi_hi_1011 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1012;
  assign dataGroup_hi_hi_1012 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1013;
  assign dataGroup_hi_hi_1013 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1014;
  assign dataGroup_hi_hi_1014 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1015;
  assign dataGroup_hi_hi_1015 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1016;
  assign dataGroup_hi_hi_1016 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1017;
  assign dataGroup_hi_hi_1017 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1018;
  assign dataGroup_hi_hi_1018 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1019;
  assign dataGroup_hi_hi_1019 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1020;
  assign dataGroup_hi_hi_1020 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1021;
  assign dataGroup_hi_hi_1021 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1022;
  assign dataGroup_hi_hi_1022 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1023;
  assign dataGroup_hi_hi_1023 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1024;
  assign dataGroup_hi_hi_1024 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1025;
  assign dataGroup_hi_hi_1025 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1026;
  assign dataGroup_hi_hi_1026 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1027;
  assign dataGroup_hi_hi_1027 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1028;
  assign dataGroup_hi_hi_1028 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1029;
  assign dataGroup_hi_hi_1029 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1030;
  assign dataGroup_hi_hi_1030 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1031;
  assign dataGroup_hi_hi_1031 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1032;
  assign dataGroup_hi_hi_1032 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1033;
  assign dataGroup_hi_hi_1033 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1034;
  assign dataGroup_hi_hi_1034 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1035;
  assign dataGroup_hi_hi_1035 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1036;
  assign dataGroup_hi_hi_1036 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1037;
  assign dataGroup_hi_hi_1037 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1038;
  assign dataGroup_hi_hi_1038 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1039;
  assign dataGroup_hi_hi_1039 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1040;
  assign dataGroup_hi_hi_1040 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1041;
  assign dataGroup_hi_hi_1041 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1042;
  assign dataGroup_hi_hi_1042 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1043;
  assign dataGroup_hi_hi_1043 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1044;
  assign dataGroup_hi_hi_1044 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1045;
  assign dataGroup_hi_hi_1045 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1046;
  assign dataGroup_hi_hi_1046 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1047;
  assign dataGroup_hi_hi_1047 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1048;
  assign dataGroup_hi_hi_1048 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1049;
  assign dataGroup_hi_hi_1049 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1050;
  assign dataGroup_hi_hi_1050 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1051;
  assign dataGroup_hi_hi_1051 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1052;
  assign dataGroup_hi_hi_1052 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1053;
  assign dataGroup_hi_hi_1053 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1054;
  assign dataGroup_hi_hi_1054 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1055;
  assign dataGroup_hi_hi_1055 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1056;
  assign dataGroup_hi_hi_1056 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1057;
  assign dataGroup_hi_hi_1057 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1058;
  assign dataGroup_hi_hi_1058 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1059;
  assign dataGroup_hi_hi_1059 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1060;
  assign dataGroup_hi_hi_1060 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1061;
  assign dataGroup_hi_hi_1061 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1062;
  assign dataGroup_hi_hi_1062 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1063;
  assign dataGroup_hi_hi_1063 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1064;
  assign dataGroup_hi_hi_1064 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1065;
  assign dataGroup_hi_hi_1065 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1066;
  assign dataGroup_hi_hi_1066 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1067;
  assign dataGroup_hi_hi_1067 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1068;
  assign dataGroup_hi_hi_1068 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1069;
  assign dataGroup_hi_hi_1069 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1070;
  assign dataGroup_hi_hi_1070 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1071;
  assign dataGroup_hi_hi_1071 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1072;
  assign dataGroup_hi_hi_1072 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1073;
  assign dataGroup_hi_hi_1073 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1074;
  assign dataGroup_hi_hi_1074 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1075;
  assign dataGroup_hi_hi_1075 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1076;
  assign dataGroup_hi_hi_1076 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1077;
  assign dataGroup_hi_hi_1077 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1078;
  assign dataGroup_hi_hi_1078 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1079;
  assign dataGroup_hi_hi_1079 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1080;
  assign dataGroup_hi_hi_1080 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1081;
  assign dataGroup_hi_hi_1081 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1082;
  assign dataGroup_hi_hi_1082 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1083;
  assign dataGroup_hi_hi_1083 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1084;
  assign dataGroup_hi_hi_1084 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1085;
  assign dataGroup_hi_hi_1085 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1086;
  assign dataGroup_hi_hi_1086 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1087;
  assign dataGroup_hi_hi_1087 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1088;
  assign dataGroup_hi_hi_1088 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1089;
  assign dataGroup_hi_hi_1089 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1090;
  assign dataGroup_hi_hi_1090 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1091;
  assign dataGroup_hi_hi_1091 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1092;
  assign dataGroup_hi_hi_1092 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1093;
  assign dataGroup_hi_hi_1093 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1094;
  assign dataGroup_hi_hi_1094 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1095;
  assign dataGroup_hi_hi_1095 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1096;
  assign dataGroup_hi_hi_1096 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1097;
  assign dataGroup_hi_hi_1097 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1098;
  assign dataGroup_hi_hi_1098 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1099;
  assign dataGroup_hi_hi_1099 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1100;
  assign dataGroup_hi_hi_1100 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1101;
  assign dataGroup_hi_hi_1101 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1102;
  assign dataGroup_hi_hi_1102 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1103;
  assign dataGroup_hi_hi_1103 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1104;
  assign dataGroup_hi_hi_1104 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1105;
  assign dataGroup_hi_hi_1105 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1106;
  assign dataGroup_hi_hi_1106 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1107;
  assign dataGroup_hi_hi_1107 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1108;
  assign dataGroup_hi_hi_1108 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1109;
  assign dataGroup_hi_hi_1109 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1110;
  assign dataGroup_hi_hi_1110 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1111;
  assign dataGroup_hi_hi_1111 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1112;
  assign dataGroup_hi_hi_1112 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1113;
  assign dataGroup_hi_hi_1113 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1114;
  assign dataGroup_hi_hi_1114 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1115;
  assign dataGroup_hi_hi_1115 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1116;
  assign dataGroup_hi_hi_1116 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1117;
  assign dataGroup_hi_hi_1117 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1118;
  assign dataGroup_hi_hi_1118 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1119;
  assign dataGroup_hi_hi_1119 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1120;
  assign dataGroup_hi_hi_1120 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1121;
  assign dataGroup_hi_hi_1121 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1122;
  assign dataGroup_hi_hi_1122 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1123;
  assign dataGroup_hi_hi_1123 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1124;
  assign dataGroup_hi_hi_1124 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1125;
  assign dataGroup_hi_hi_1125 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1126;
  assign dataGroup_hi_hi_1126 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1127;
  assign dataGroup_hi_hi_1127 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1128;
  assign dataGroup_hi_hi_1128 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1129;
  assign dataGroup_hi_hi_1129 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1130;
  assign dataGroup_hi_hi_1130 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1131;
  assign dataGroup_hi_hi_1131 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1132;
  assign dataGroup_hi_hi_1132 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1133;
  assign dataGroup_hi_hi_1133 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1134;
  assign dataGroup_hi_hi_1134 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1135;
  assign dataGroup_hi_hi_1135 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1136;
  assign dataGroup_hi_hi_1136 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1137;
  assign dataGroup_hi_hi_1137 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1138;
  assign dataGroup_hi_hi_1138 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1139;
  assign dataGroup_hi_hi_1139 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1140;
  assign dataGroup_hi_hi_1140 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1141;
  assign dataGroup_hi_hi_1141 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1142;
  assign dataGroup_hi_hi_1142 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1143;
  assign dataGroup_hi_hi_1143 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1144;
  assign dataGroup_hi_hi_1144 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1145;
  assign dataGroup_hi_hi_1145 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1146;
  assign dataGroup_hi_hi_1146 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1147;
  assign dataGroup_hi_hi_1147 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1148;
  assign dataGroup_hi_hi_1148 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1149;
  assign dataGroup_hi_hi_1149 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1150;
  assign dataGroup_hi_hi_1150 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1151;
  assign dataGroup_hi_hi_1151 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1152;
  assign dataGroup_hi_hi_1152 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1153;
  assign dataGroup_hi_hi_1153 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1154;
  assign dataGroup_hi_hi_1154 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1155;
  assign dataGroup_hi_hi_1155 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1156;
  assign dataGroup_hi_hi_1156 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1157;
  assign dataGroup_hi_hi_1157 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1158;
  assign dataGroup_hi_hi_1158 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1159;
  assign dataGroup_hi_hi_1159 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1160;
  assign dataGroup_hi_hi_1160 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1161;
  assign dataGroup_hi_hi_1161 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1162;
  assign dataGroup_hi_hi_1162 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1163;
  assign dataGroup_hi_hi_1163 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1164;
  assign dataGroup_hi_hi_1164 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1165;
  assign dataGroup_hi_hi_1165 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1166;
  assign dataGroup_hi_hi_1166 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1167;
  assign dataGroup_hi_hi_1167 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1168;
  assign dataGroup_hi_hi_1168 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1169;
  assign dataGroup_hi_hi_1169 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1170;
  assign dataGroup_hi_hi_1170 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1171;
  assign dataGroup_hi_hi_1171 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1172;
  assign dataGroup_hi_hi_1172 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1173;
  assign dataGroup_hi_hi_1173 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1174;
  assign dataGroup_hi_hi_1174 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1175;
  assign dataGroup_hi_hi_1175 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1176;
  assign dataGroup_hi_hi_1176 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1177;
  assign dataGroup_hi_hi_1177 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1178;
  assign dataGroup_hi_hi_1178 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1179;
  assign dataGroup_hi_hi_1179 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1180;
  assign dataGroup_hi_hi_1180 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1181;
  assign dataGroup_hi_hi_1181 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1182;
  assign dataGroup_hi_hi_1182 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1183;
  assign dataGroup_hi_hi_1183 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1184;
  assign dataGroup_hi_hi_1184 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1185;
  assign dataGroup_hi_hi_1185 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1186;
  assign dataGroup_hi_hi_1186 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1187;
  assign dataGroup_hi_hi_1187 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1188;
  assign dataGroup_hi_hi_1188 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1189;
  assign dataGroup_hi_hi_1189 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1190;
  assign dataGroup_hi_hi_1190 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1191;
  assign dataGroup_hi_hi_1191 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1192;
  assign dataGroup_hi_hi_1192 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1193;
  assign dataGroup_hi_hi_1193 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1194;
  assign dataGroup_hi_hi_1194 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1195;
  assign dataGroup_hi_hi_1195 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1196;
  assign dataGroup_hi_hi_1196 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1197;
  assign dataGroup_hi_hi_1197 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1198;
  assign dataGroup_hi_hi_1198 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1199;
  assign dataGroup_hi_hi_1199 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1200;
  assign dataGroup_hi_hi_1200 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1201;
  assign dataGroup_hi_hi_1201 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1202;
  assign dataGroup_hi_hi_1202 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1203;
  assign dataGroup_hi_hi_1203 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1204;
  assign dataGroup_hi_hi_1204 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1205;
  assign dataGroup_hi_hi_1205 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1206;
  assign dataGroup_hi_hi_1206 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1207;
  assign dataGroup_hi_hi_1207 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1208;
  assign dataGroup_hi_hi_1208 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1209;
  assign dataGroup_hi_hi_1209 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1210;
  assign dataGroup_hi_hi_1210 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1211;
  assign dataGroup_hi_hi_1211 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1212;
  assign dataGroup_hi_hi_1212 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1213;
  assign dataGroup_hi_hi_1213 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1214;
  assign dataGroup_hi_hi_1214 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1215;
  assign dataGroup_hi_hi_1215 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1216;
  assign dataGroup_hi_hi_1216 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1217;
  assign dataGroup_hi_hi_1217 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1218;
  assign dataGroup_hi_hi_1218 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1219;
  assign dataGroup_hi_hi_1219 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1220;
  assign dataGroup_hi_hi_1220 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1221;
  assign dataGroup_hi_hi_1221 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1222;
  assign dataGroup_hi_hi_1222 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1223;
  assign dataGroup_hi_hi_1223 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1224;
  assign dataGroup_hi_hi_1224 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1225;
  assign dataGroup_hi_hi_1225 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1226;
  assign dataGroup_hi_hi_1226 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1227;
  assign dataGroup_hi_hi_1227 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1228;
  assign dataGroup_hi_hi_1228 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1229;
  assign dataGroup_hi_hi_1229 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1230;
  assign dataGroup_hi_hi_1230 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1231;
  assign dataGroup_hi_hi_1231 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1232;
  assign dataGroup_hi_hi_1232 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1233;
  assign dataGroup_hi_hi_1233 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1234;
  assign dataGroup_hi_hi_1234 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1235;
  assign dataGroup_hi_hi_1235 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1236;
  assign dataGroup_hi_hi_1236 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1237;
  assign dataGroup_hi_hi_1237 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1238;
  assign dataGroup_hi_hi_1238 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1239;
  assign dataGroup_hi_hi_1239 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1240;
  assign dataGroup_hi_hi_1240 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1241;
  assign dataGroup_hi_hi_1241 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1242;
  assign dataGroup_hi_hi_1242 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1243;
  assign dataGroup_hi_hi_1243 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1244;
  assign dataGroup_hi_hi_1244 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1245;
  assign dataGroup_hi_hi_1245 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1246;
  assign dataGroup_hi_hi_1246 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1247;
  assign dataGroup_hi_hi_1247 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1248;
  assign dataGroup_hi_hi_1248 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1249;
  assign dataGroup_hi_hi_1249 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1250;
  assign dataGroup_hi_hi_1250 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1251;
  assign dataGroup_hi_hi_1251 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1252;
  assign dataGroup_hi_hi_1252 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1253;
  assign dataGroup_hi_hi_1253 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1254;
  assign dataGroup_hi_hi_1254 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1255;
  assign dataGroup_hi_hi_1255 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1256;
  assign dataGroup_hi_hi_1256 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1257;
  assign dataGroup_hi_hi_1257 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1258;
  assign dataGroup_hi_hi_1258 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1259;
  assign dataGroup_hi_hi_1259 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1260;
  assign dataGroup_hi_hi_1260 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1261;
  assign dataGroup_hi_hi_1261 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1262;
  assign dataGroup_hi_hi_1262 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1263;
  assign dataGroup_hi_hi_1263 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1264;
  assign dataGroup_hi_hi_1264 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1265;
  assign dataGroup_hi_hi_1265 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1266;
  assign dataGroup_hi_hi_1266 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1267;
  assign dataGroup_hi_hi_1267 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1268;
  assign dataGroup_hi_hi_1268 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1269;
  assign dataGroup_hi_hi_1269 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1270;
  assign dataGroup_hi_hi_1270 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1271;
  assign dataGroup_hi_hi_1271 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1272;
  assign dataGroup_hi_hi_1272 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1273;
  assign dataGroup_hi_hi_1273 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1274;
  assign dataGroup_hi_hi_1274 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1275;
  assign dataGroup_hi_hi_1275 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1276;
  assign dataGroup_hi_hi_1276 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1277;
  assign dataGroup_hi_hi_1277 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1278;
  assign dataGroup_hi_hi_1278 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1279;
  assign dataGroup_hi_hi_1279 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1280;
  assign dataGroup_hi_hi_1280 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1281;
  assign dataGroup_hi_hi_1281 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1282;
  assign dataGroup_hi_hi_1282 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1283;
  assign dataGroup_hi_hi_1283 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1284;
  assign dataGroup_hi_hi_1284 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1285;
  assign dataGroup_hi_hi_1285 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1286;
  assign dataGroup_hi_hi_1286 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1287;
  assign dataGroup_hi_hi_1287 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1288;
  assign dataGroup_hi_hi_1288 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1289;
  assign dataGroup_hi_hi_1289 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1290;
  assign dataGroup_hi_hi_1290 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1291;
  assign dataGroup_hi_hi_1291 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1292;
  assign dataGroup_hi_hi_1292 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1293;
  assign dataGroup_hi_hi_1293 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1294;
  assign dataGroup_hi_hi_1294 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1295;
  assign dataGroup_hi_hi_1295 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1296;
  assign dataGroup_hi_hi_1296 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1297;
  assign dataGroup_hi_hi_1297 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1298;
  assign dataGroup_hi_hi_1298 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1299;
  assign dataGroup_hi_hi_1299 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1300;
  assign dataGroup_hi_hi_1300 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1301;
  assign dataGroup_hi_hi_1301 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1302;
  assign dataGroup_hi_hi_1302 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1303;
  assign dataGroup_hi_hi_1303 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1304;
  assign dataGroup_hi_hi_1304 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1305;
  assign dataGroup_hi_hi_1305 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1306;
  assign dataGroup_hi_hi_1306 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1307;
  assign dataGroup_hi_hi_1307 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1308;
  assign dataGroup_hi_hi_1308 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1309;
  assign dataGroup_hi_hi_1309 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1310;
  assign dataGroup_hi_hi_1310 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1311;
  assign dataGroup_hi_hi_1311 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1312;
  assign dataGroup_hi_hi_1312 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1313;
  assign dataGroup_hi_hi_1313 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1314;
  assign dataGroup_hi_hi_1314 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1315;
  assign dataGroup_hi_hi_1315 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1316;
  assign dataGroup_hi_hi_1316 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1317;
  assign dataGroup_hi_hi_1317 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1318;
  assign dataGroup_hi_hi_1318 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1319;
  assign dataGroup_hi_hi_1319 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1320;
  assign dataGroup_hi_hi_1320 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1321;
  assign dataGroup_hi_hi_1321 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1322;
  assign dataGroup_hi_hi_1322 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1323;
  assign dataGroup_hi_hi_1323 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1324;
  assign dataGroup_hi_hi_1324 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1325;
  assign dataGroup_hi_hi_1325 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1326;
  assign dataGroup_hi_hi_1326 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1327;
  assign dataGroup_hi_hi_1327 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1328;
  assign dataGroup_hi_hi_1328 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1329;
  assign dataGroup_hi_hi_1329 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1330;
  assign dataGroup_hi_hi_1330 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1331;
  assign dataGroup_hi_hi_1331 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1332;
  assign dataGroup_hi_hi_1332 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1333;
  assign dataGroup_hi_hi_1333 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1334;
  assign dataGroup_hi_hi_1334 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1335;
  assign dataGroup_hi_hi_1335 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1336;
  assign dataGroup_hi_hi_1336 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1337;
  assign dataGroup_hi_hi_1337 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1338;
  assign dataGroup_hi_hi_1338 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1339;
  assign dataGroup_hi_hi_1339 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1340;
  assign dataGroup_hi_hi_1340 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1341;
  assign dataGroup_hi_hi_1341 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1342;
  assign dataGroup_hi_hi_1342 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1343;
  assign dataGroup_hi_hi_1343 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1344;
  assign dataGroup_hi_hi_1344 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1345;
  assign dataGroup_hi_hi_1345 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1346;
  assign dataGroup_hi_hi_1346 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1347;
  assign dataGroup_hi_hi_1347 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1348;
  assign dataGroup_hi_hi_1348 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1349;
  assign dataGroup_hi_hi_1349 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1350;
  assign dataGroup_hi_hi_1350 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1351;
  assign dataGroup_hi_hi_1351 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1352;
  assign dataGroup_hi_hi_1352 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1353;
  assign dataGroup_hi_hi_1353 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1354;
  assign dataGroup_hi_hi_1354 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1355;
  assign dataGroup_hi_hi_1355 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1356;
  assign dataGroup_hi_hi_1356 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1357;
  assign dataGroup_hi_hi_1357 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1358;
  assign dataGroup_hi_hi_1358 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1359;
  assign dataGroup_hi_hi_1359 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1360;
  assign dataGroup_hi_hi_1360 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1361;
  assign dataGroup_hi_hi_1361 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1362;
  assign dataGroup_hi_hi_1362 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1363;
  assign dataGroup_hi_hi_1363 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1364;
  assign dataGroup_hi_hi_1364 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1365;
  assign dataGroup_hi_hi_1365 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1366;
  assign dataGroup_hi_hi_1366 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1367;
  assign dataGroup_hi_hi_1367 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1368;
  assign dataGroup_hi_hi_1368 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1369;
  assign dataGroup_hi_hi_1369 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1370;
  assign dataGroup_hi_hi_1370 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1371;
  assign dataGroup_hi_hi_1371 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1372;
  assign dataGroup_hi_hi_1372 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1373;
  assign dataGroup_hi_hi_1373 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1374;
  assign dataGroup_hi_hi_1374 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1375;
  assign dataGroup_hi_hi_1375 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1376;
  assign dataGroup_hi_hi_1376 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1377;
  assign dataGroup_hi_hi_1377 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1378;
  assign dataGroup_hi_hi_1378 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1379;
  assign dataGroup_hi_hi_1379 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1380;
  assign dataGroup_hi_hi_1380 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1381;
  assign dataGroup_hi_hi_1381 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1382;
  assign dataGroup_hi_hi_1382 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1383;
  assign dataGroup_hi_hi_1383 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1384;
  assign dataGroup_hi_hi_1384 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1385;
  assign dataGroup_hi_hi_1385 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1386;
  assign dataGroup_hi_hi_1386 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1387;
  assign dataGroup_hi_hi_1387 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1388;
  assign dataGroup_hi_hi_1388 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1389;
  assign dataGroup_hi_hi_1389 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1390;
  assign dataGroup_hi_hi_1390 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1391;
  assign dataGroup_hi_hi_1391 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1392;
  assign dataGroup_hi_hi_1392 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1393;
  assign dataGroup_hi_hi_1393 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1394;
  assign dataGroup_hi_hi_1394 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1395;
  assign dataGroup_hi_hi_1395 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1396;
  assign dataGroup_hi_hi_1396 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1397;
  assign dataGroup_hi_hi_1397 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1398;
  assign dataGroup_hi_hi_1398 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1399;
  assign dataGroup_hi_hi_1399 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1400;
  assign dataGroup_hi_hi_1400 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1401;
  assign dataGroup_hi_hi_1401 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1402;
  assign dataGroup_hi_hi_1402 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1403;
  assign dataGroup_hi_hi_1403 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1404;
  assign dataGroup_hi_hi_1404 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1405;
  assign dataGroup_hi_hi_1405 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1406;
  assign dataGroup_hi_hi_1406 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1407;
  assign dataGroup_hi_hi_1407 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1408;
  assign dataGroup_hi_hi_1408 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1409;
  assign dataGroup_hi_hi_1409 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1410;
  assign dataGroup_hi_hi_1410 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1411;
  assign dataGroup_hi_hi_1411 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1412;
  assign dataGroup_hi_hi_1412 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1413;
  assign dataGroup_hi_hi_1413 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1414;
  assign dataGroup_hi_hi_1414 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1415;
  assign dataGroup_hi_hi_1415 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1416;
  assign dataGroup_hi_hi_1416 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1417;
  assign dataGroup_hi_hi_1417 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1418;
  assign dataGroup_hi_hi_1418 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1419;
  assign dataGroup_hi_hi_1419 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1420;
  assign dataGroup_hi_hi_1420 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1421;
  assign dataGroup_hi_hi_1421 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1422;
  assign dataGroup_hi_hi_1422 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1423;
  assign dataGroup_hi_hi_1423 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1424;
  assign dataGroup_hi_hi_1424 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1425;
  assign dataGroup_hi_hi_1425 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1426;
  assign dataGroup_hi_hi_1426 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1427;
  assign dataGroup_hi_hi_1427 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1428;
  assign dataGroup_hi_hi_1428 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1429;
  assign dataGroup_hi_hi_1429 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1430;
  assign dataGroup_hi_hi_1430 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1431;
  assign dataGroup_hi_hi_1431 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1432;
  assign dataGroup_hi_hi_1432 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1433;
  assign dataGroup_hi_hi_1433 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1434;
  assign dataGroup_hi_hi_1434 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1435;
  assign dataGroup_hi_hi_1435 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1436;
  assign dataGroup_hi_hi_1436 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1437;
  assign dataGroup_hi_hi_1437 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1438;
  assign dataGroup_hi_hi_1438 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1439;
  assign dataGroup_hi_hi_1439 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1440;
  assign dataGroup_hi_hi_1440 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1441;
  assign dataGroup_hi_hi_1441 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1442;
  assign dataGroup_hi_hi_1442 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1443;
  assign dataGroup_hi_hi_1443 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1444;
  assign dataGroup_hi_hi_1444 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1445;
  assign dataGroup_hi_hi_1445 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1446;
  assign dataGroup_hi_hi_1446 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1447;
  assign dataGroup_hi_hi_1447 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1448;
  assign dataGroup_hi_hi_1448 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1449;
  assign dataGroup_hi_hi_1449 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1450;
  assign dataGroup_hi_hi_1450 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1451;
  assign dataGroup_hi_hi_1451 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1452;
  assign dataGroup_hi_hi_1452 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1453;
  assign dataGroup_hi_hi_1453 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1454;
  assign dataGroup_hi_hi_1454 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1455;
  assign dataGroup_hi_hi_1455 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1456;
  assign dataGroup_hi_hi_1456 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1457;
  assign dataGroup_hi_hi_1457 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1458;
  assign dataGroup_hi_hi_1458 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1459;
  assign dataGroup_hi_hi_1459 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1460;
  assign dataGroup_hi_hi_1460 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1461;
  assign dataGroup_hi_hi_1461 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1462;
  assign dataGroup_hi_hi_1462 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1463;
  assign dataGroup_hi_hi_1463 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1464;
  assign dataGroup_hi_hi_1464 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1465;
  assign dataGroup_hi_hi_1465 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1466;
  assign dataGroup_hi_hi_1466 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1467;
  assign dataGroup_hi_hi_1467 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1468;
  assign dataGroup_hi_hi_1468 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1469;
  assign dataGroup_hi_hi_1469 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1470;
  assign dataGroup_hi_hi_1470 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1471;
  assign dataGroup_hi_hi_1471 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1472;
  assign dataGroup_hi_hi_1472 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1473;
  assign dataGroup_hi_hi_1473 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1474;
  assign dataGroup_hi_hi_1474 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1475;
  assign dataGroup_hi_hi_1475 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1476;
  assign dataGroup_hi_hi_1476 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1477;
  assign dataGroup_hi_hi_1477 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1478;
  assign dataGroup_hi_hi_1478 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1479;
  assign dataGroup_hi_hi_1479 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1480;
  assign dataGroup_hi_hi_1480 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1481;
  assign dataGroup_hi_hi_1481 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1482;
  assign dataGroup_hi_hi_1482 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1483;
  assign dataGroup_hi_hi_1483 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1484;
  assign dataGroup_hi_hi_1484 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1485;
  assign dataGroup_hi_hi_1485 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1486;
  assign dataGroup_hi_hi_1486 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1487;
  assign dataGroup_hi_hi_1487 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1488;
  assign dataGroup_hi_hi_1488 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1489;
  assign dataGroup_hi_hi_1489 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1490;
  assign dataGroup_hi_hi_1490 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1491;
  assign dataGroup_hi_hi_1491 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1492;
  assign dataGroup_hi_hi_1492 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1493;
  assign dataGroup_hi_hi_1493 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1494;
  assign dataGroup_hi_hi_1494 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1495;
  assign dataGroup_hi_hi_1495 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1496;
  assign dataGroup_hi_hi_1496 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1497;
  assign dataGroup_hi_hi_1497 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1498;
  assign dataGroup_hi_hi_1498 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1499;
  assign dataGroup_hi_hi_1499 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1500;
  assign dataGroup_hi_hi_1500 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1501;
  assign dataGroup_hi_hi_1501 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1502;
  assign dataGroup_hi_hi_1502 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1503;
  assign dataGroup_hi_hi_1503 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1504;
  assign dataGroup_hi_hi_1504 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1505;
  assign dataGroup_hi_hi_1505 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1506;
  assign dataGroup_hi_hi_1506 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1507;
  assign dataGroup_hi_hi_1507 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1508;
  assign dataGroup_hi_hi_1508 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1509;
  assign dataGroup_hi_hi_1509 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1510;
  assign dataGroup_hi_hi_1510 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1511;
  assign dataGroup_hi_hi_1511 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1512;
  assign dataGroup_hi_hi_1512 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1513;
  assign dataGroup_hi_hi_1513 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1514;
  assign dataGroup_hi_hi_1514 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1515;
  assign dataGroup_hi_hi_1515 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1516;
  assign dataGroup_hi_hi_1516 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1517;
  assign dataGroup_hi_hi_1517 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1518;
  assign dataGroup_hi_hi_1518 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1519;
  assign dataGroup_hi_hi_1519 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1520;
  assign dataGroup_hi_hi_1520 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1521;
  assign dataGroup_hi_hi_1521 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1522;
  assign dataGroup_hi_hi_1522 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1523;
  assign dataGroup_hi_hi_1523 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1524;
  assign dataGroup_hi_hi_1524 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1525;
  assign dataGroup_hi_hi_1525 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1526;
  assign dataGroup_hi_hi_1526 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1527;
  assign dataGroup_hi_hi_1527 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1528;
  assign dataGroup_hi_hi_1528 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1529;
  assign dataGroup_hi_hi_1529 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1530;
  assign dataGroup_hi_hi_1530 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1531;
  assign dataGroup_hi_hi_1531 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1532;
  assign dataGroup_hi_hi_1532 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1533;
  assign dataGroup_hi_hi_1533 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1534;
  assign dataGroup_hi_hi_1534 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1535;
  assign dataGroup_hi_hi_1535 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1536;
  assign dataGroup_hi_hi_1536 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1537;
  assign dataGroup_hi_hi_1537 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1538;
  assign dataGroup_hi_hi_1538 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1539;
  assign dataGroup_hi_hi_1539 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1540;
  assign dataGroup_hi_hi_1540 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1541;
  assign dataGroup_hi_hi_1541 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1542;
  assign dataGroup_hi_hi_1542 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1543;
  assign dataGroup_hi_hi_1543 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1544;
  assign dataGroup_hi_hi_1544 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1545;
  assign dataGroup_hi_hi_1545 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1546;
  assign dataGroup_hi_hi_1546 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1547;
  assign dataGroup_hi_hi_1547 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1548;
  assign dataGroup_hi_hi_1548 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1549;
  assign dataGroup_hi_hi_1549 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1550;
  assign dataGroup_hi_hi_1550 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1551;
  assign dataGroup_hi_hi_1551 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1552;
  assign dataGroup_hi_hi_1552 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1553;
  assign dataGroup_hi_hi_1553 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1554;
  assign dataGroup_hi_hi_1554 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1555;
  assign dataGroup_hi_hi_1555 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1556;
  assign dataGroup_hi_hi_1556 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1557;
  assign dataGroup_hi_hi_1557 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1558;
  assign dataGroup_hi_hi_1558 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1559;
  assign dataGroup_hi_hi_1559 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1560;
  assign dataGroup_hi_hi_1560 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1561;
  assign dataGroup_hi_hi_1561 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1562;
  assign dataGroup_hi_hi_1562 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1563;
  assign dataGroup_hi_hi_1563 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1564;
  assign dataGroup_hi_hi_1564 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1565;
  assign dataGroup_hi_hi_1565 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1566;
  assign dataGroup_hi_hi_1566 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1567;
  assign dataGroup_hi_hi_1567 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1568;
  assign dataGroup_hi_hi_1568 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1569;
  assign dataGroup_hi_hi_1569 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1570;
  assign dataGroup_hi_hi_1570 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1571;
  assign dataGroup_hi_hi_1571 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1572;
  assign dataGroup_hi_hi_1572 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1573;
  assign dataGroup_hi_hi_1573 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1574;
  assign dataGroup_hi_hi_1574 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1575;
  assign dataGroup_hi_hi_1575 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1576;
  assign dataGroup_hi_hi_1576 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1577;
  assign dataGroup_hi_hi_1577 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1578;
  assign dataGroup_hi_hi_1578 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1579;
  assign dataGroup_hi_hi_1579 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1580;
  assign dataGroup_hi_hi_1580 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1581;
  assign dataGroup_hi_hi_1581 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1582;
  assign dataGroup_hi_hi_1582 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1583;
  assign dataGroup_hi_hi_1583 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1584;
  assign dataGroup_hi_hi_1584 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1585;
  assign dataGroup_hi_hi_1585 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1586;
  assign dataGroup_hi_hi_1586 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1587;
  assign dataGroup_hi_hi_1587 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1588;
  assign dataGroup_hi_hi_1588 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1589;
  assign dataGroup_hi_hi_1589 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1590;
  assign dataGroup_hi_hi_1590 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1591;
  assign dataGroup_hi_hi_1591 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1592;
  assign dataGroup_hi_hi_1592 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1593;
  assign dataGroup_hi_hi_1593 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1594;
  assign dataGroup_hi_hi_1594 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1595;
  assign dataGroup_hi_hi_1595 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1596;
  assign dataGroup_hi_hi_1596 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1597;
  assign dataGroup_hi_hi_1597 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1598;
  assign dataGroup_hi_hi_1598 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1599;
  assign dataGroup_hi_hi_1599 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1600;
  assign dataGroup_hi_hi_1600 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1601;
  assign dataGroup_hi_hi_1601 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1602;
  assign dataGroup_hi_hi_1602 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1603;
  assign dataGroup_hi_hi_1603 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1604;
  assign dataGroup_hi_hi_1604 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1605;
  assign dataGroup_hi_hi_1605 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1606;
  assign dataGroup_hi_hi_1606 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1607;
  assign dataGroup_hi_hi_1607 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1608;
  assign dataGroup_hi_hi_1608 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1609;
  assign dataGroup_hi_hi_1609 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1610;
  assign dataGroup_hi_hi_1610 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1611;
  assign dataGroup_hi_hi_1611 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1612;
  assign dataGroup_hi_hi_1612 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1613;
  assign dataGroup_hi_hi_1613 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1614;
  assign dataGroup_hi_hi_1614 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1615;
  assign dataGroup_hi_hi_1615 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1616;
  assign dataGroup_hi_hi_1616 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1617;
  assign dataGroup_hi_hi_1617 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1618;
  assign dataGroup_hi_hi_1618 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1619;
  assign dataGroup_hi_hi_1619 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1620;
  assign dataGroup_hi_hi_1620 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1621;
  assign dataGroup_hi_hi_1621 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1622;
  assign dataGroup_hi_hi_1622 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1623;
  assign dataGroup_hi_hi_1623 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1624;
  assign dataGroup_hi_hi_1624 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1625;
  assign dataGroup_hi_hi_1625 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1626;
  assign dataGroup_hi_hi_1626 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1627;
  assign dataGroup_hi_hi_1627 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1628;
  assign dataGroup_hi_hi_1628 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1629;
  assign dataGroup_hi_hi_1629 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1630;
  assign dataGroup_hi_hi_1630 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1631;
  assign dataGroup_hi_hi_1631 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1632;
  assign dataGroup_hi_hi_1632 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1633;
  assign dataGroup_hi_hi_1633 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1634;
  assign dataGroup_hi_hi_1634 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1635;
  assign dataGroup_hi_hi_1635 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1636;
  assign dataGroup_hi_hi_1636 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1637;
  assign dataGroup_hi_hi_1637 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1638;
  assign dataGroup_hi_hi_1638 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1639;
  assign dataGroup_hi_hi_1639 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1640;
  assign dataGroup_hi_hi_1640 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1641;
  assign dataGroup_hi_hi_1641 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1642;
  assign dataGroup_hi_hi_1642 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1643;
  assign dataGroup_hi_hi_1643 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1644;
  assign dataGroup_hi_hi_1644 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1645;
  assign dataGroup_hi_hi_1645 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1646;
  assign dataGroup_hi_hi_1646 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1647;
  assign dataGroup_hi_hi_1647 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1648;
  assign dataGroup_hi_hi_1648 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1649;
  assign dataGroup_hi_hi_1649 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1650;
  assign dataGroup_hi_hi_1650 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1651;
  assign dataGroup_hi_hi_1651 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1652;
  assign dataGroup_hi_hi_1652 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1653;
  assign dataGroup_hi_hi_1653 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1654;
  assign dataGroup_hi_hi_1654 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1655;
  assign dataGroup_hi_hi_1655 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1656;
  assign dataGroup_hi_hi_1656 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1657;
  assign dataGroup_hi_hi_1657 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1658;
  assign dataGroup_hi_hi_1658 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1659;
  assign dataGroup_hi_hi_1659 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1660;
  assign dataGroup_hi_hi_1660 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1661;
  assign dataGroup_hi_hi_1661 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1662;
  assign dataGroup_hi_hi_1662 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1663;
  assign dataGroup_hi_hi_1663 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1664;
  assign dataGroup_hi_hi_1664 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1665;
  assign dataGroup_hi_hi_1665 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1666;
  assign dataGroup_hi_hi_1666 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1667;
  assign dataGroup_hi_hi_1667 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1668;
  assign dataGroup_hi_hi_1668 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1669;
  assign dataGroup_hi_hi_1669 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1670;
  assign dataGroup_hi_hi_1670 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1671;
  assign dataGroup_hi_hi_1671 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1672;
  assign dataGroup_hi_hi_1672 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1673;
  assign dataGroup_hi_hi_1673 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1674;
  assign dataGroup_hi_hi_1674 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1675;
  assign dataGroup_hi_hi_1675 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1676;
  assign dataGroup_hi_hi_1676 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1677;
  assign dataGroup_hi_hi_1677 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1678;
  assign dataGroup_hi_hi_1678 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1679;
  assign dataGroup_hi_hi_1679 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1680;
  assign dataGroup_hi_hi_1680 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1681;
  assign dataGroup_hi_hi_1681 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1682;
  assign dataGroup_hi_hi_1682 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1683;
  assign dataGroup_hi_hi_1683 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1684;
  assign dataGroup_hi_hi_1684 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1685;
  assign dataGroup_hi_hi_1685 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1686;
  assign dataGroup_hi_hi_1686 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1687;
  assign dataGroup_hi_hi_1687 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1688;
  assign dataGroup_hi_hi_1688 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1689;
  assign dataGroup_hi_hi_1689 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1690;
  assign dataGroup_hi_hi_1690 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1691;
  assign dataGroup_hi_hi_1691 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1692;
  assign dataGroup_hi_hi_1692 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1693;
  assign dataGroup_hi_hi_1693 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1694;
  assign dataGroup_hi_hi_1694 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1695;
  assign dataGroup_hi_hi_1695 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1696;
  assign dataGroup_hi_hi_1696 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1697;
  assign dataGroup_hi_hi_1697 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1698;
  assign dataGroup_hi_hi_1698 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1699;
  assign dataGroup_hi_hi_1699 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1700;
  assign dataGroup_hi_hi_1700 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1701;
  assign dataGroup_hi_hi_1701 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1702;
  assign dataGroup_hi_hi_1702 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1703;
  assign dataGroup_hi_hi_1703 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1704;
  assign dataGroup_hi_hi_1704 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1705;
  assign dataGroup_hi_hi_1705 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1706;
  assign dataGroup_hi_hi_1706 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1707;
  assign dataGroup_hi_hi_1707 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1708;
  assign dataGroup_hi_hi_1708 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1709;
  assign dataGroup_hi_hi_1709 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1710;
  assign dataGroup_hi_hi_1710 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1711;
  assign dataGroup_hi_hi_1711 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1712;
  assign dataGroup_hi_hi_1712 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1713;
  assign dataGroup_hi_hi_1713 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1714;
  assign dataGroup_hi_hi_1714 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1715;
  assign dataGroup_hi_hi_1715 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1716;
  assign dataGroup_hi_hi_1716 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1717;
  assign dataGroup_hi_hi_1717 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1718;
  assign dataGroup_hi_hi_1718 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1719;
  assign dataGroup_hi_hi_1719 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1720;
  assign dataGroup_hi_hi_1720 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1721;
  assign dataGroup_hi_hi_1721 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1722;
  assign dataGroup_hi_hi_1722 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1723;
  assign dataGroup_hi_hi_1723 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1724;
  assign dataGroup_hi_hi_1724 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1725;
  assign dataGroup_hi_hi_1725 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1726;
  assign dataGroup_hi_hi_1726 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1727;
  assign dataGroup_hi_hi_1727 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1728;
  assign dataGroup_hi_hi_1728 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1729;
  assign dataGroup_hi_hi_1729 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1730;
  assign dataGroup_hi_hi_1730 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1731;
  assign dataGroup_hi_hi_1731 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1732;
  assign dataGroup_hi_hi_1732 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1733;
  assign dataGroup_hi_hi_1733 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1734;
  assign dataGroup_hi_hi_1734 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1735;
  assign dataGroup_hi_hi_1735 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1736;
  assign dataGroup_hi_hi_1736 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1737;
  assign dataGroup_hi_hi_1737 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1738;
  assign dataGroup_hi_hi_1738 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1739;
  assign dataGroup_hi_hi_1739 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1740;
  assign dataGroup_hi_hi_1740 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1741;
  assign dataGroup_hi_hi_1741 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1742;
  assign dataGroup_hi_hi_1742 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1743;
  assign dataGroup_hi_hi_1743 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1744;
  assign dataGroup_hi_hi_1744 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1745;
  assign dataGroup_hi_hi_1745 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1746;
  assign dataGroup_hi_hi_1746 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1747;
  assign dataGroup_hi_hi_1747 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1748;
  assign dataGroup_hi_hi_1748 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1749;
  assign dataGroup_hi_hi_1749 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1750;
  assign dataGroup_hi_hi_1750 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1751;
  assign dataGroup_hi_hi_1751 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1752;
  assign dataGroup_hi_hi_1752 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1753;
  assign dataGroup_hi_hi_1753 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1754;
  assign dataGroup_hi_hi_1754 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1755;
  assign dataGroup_hi_hi_1755 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1756;
  assign dataGroup_hi_hi_1756 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1757;
  assign dataGroup_hi_hi_1757 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1758;
  assign dataGroup_hi_hi_1758 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1759;
  assign dataGroup_hi_hi_1759 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1760;
  assign dataGroup_hi_hi_1760 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1761;
  assign dataGroup_hi_hi_1761 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1762;
  assign dataGroup_hi_hi_1762 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1763;
  assign dataGroup_hi_hi_1763 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1764;
  assign dataGroup_hi_hi_1764 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1765;
  assign dataGroup_hi_hi_1765 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1766;
  assign dataGroup_hi_hi_1766 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1767;
  assign dataGroup_hi_hi_1767 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1768;
  assign dataGroup_hi_hi_1768 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1769;
  assign dataGroup_hi_hi_1769 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1770;
  assign dataGroup_hi_hi_1770 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1771;
  assign dataGroup_hi_hi_1771 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1772;
  assign dataGroup_hi_hi_1772 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1773;
  assign dataGroup_hi_hi_1773 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1774;
  assign dataGroup_hi_hi_1774 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1775;
  assign dataGroup_hi_hi_1775 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1776;
  assign dataGroup_hi_hi_1776 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1777;
  assign dataGroup_hi_hi_1777 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1778;
  assign dataGroup_hi_hi_1778 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1779;
  assign dataGroup_hi_hi_1779 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1780;
  assign dataGroup_hi_hi_1780 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1781;
  assign dataGroup_hi_hi_1781 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1782;
  assign dataGroup_hi_hi_1782 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1783;
  assign dataGroup_hi_hi_1783 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1784;
  assign dataGroup_hi_hi_1784 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1785;
  assign dataGroup_hi_hi_1785 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1786;
  assign dataGroup_hi_hi_1786 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1787;
  assign dataGroup_hi_hi_1787 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1788;
  assign dataGroup_hi_hi_1788 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1789;
  assign dataGroup_hi_hi_1789 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1790;
  assign dataGroup_hi_hi_1790 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1791;
  assign dataGroup_hi_hi_1791 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1792;
  assign dataGroup_hi_hi_1792 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1793;
  assign dataGroup_hi_hi_1793 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1794;
  assign dataGroup_hi_hi_1794 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1795;
  assign dataGroup_hi_hi_1795 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1796;
  assign dataGroup_hi_hi_1796 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1797;
  assign dataGroup_hi_hi_1797 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1798;
  assign dataGroup_hi_hi_1798 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1799;
  assign dataGroup_hi_hi_1799 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1800;
  assign dataGroup_hi_hi_1800 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1801;
  assign dataGroup_hi_hi_1801 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1802;
  assign dataGroup_hi_hi_1802 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1803;
  assign dataGroup_hi_hi_1803 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1804;
  assign dataGroup_hi_hi_1804 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1805;
  assign dataGroup_hi_hi_1805 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1806;
  assign dataGroup_hi_hi_1806 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1807;
  assign dataGroup_hi_hi_1807 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1808;
  assign dataGroup_hi_hi_1808 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1809;
  assign dataGroup_hi_hi_1809 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1810;
  assign dataGroup_hi_hi_1810 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1811;
  assign dataGroup_hi_hi_1811 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1812;
  assign dataGroup_hi_hi_1812 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1813;
  assign dataGroup_hi_hi_1813 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1814;
  assign dataGroup_hi_hi_1814 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1815;
  assign dataGroup_hi_hi_1815 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1816;
  assign dataGroup_hi_hi_1816 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1817;
  assign dataGroup_hi_hi_1817 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1818;
  assign dataGroup_hi_hi_1818 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1819;
  assign dataGroup_hi_hi_1819 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1820;
  assign dataGroup_hi_hi_1820 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1821;
  assign dataGroup_hi_hi_1821 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1822;
  assign dataGroup_hi_hi_1822 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1823;
  assign dataGroup_hi_hi_1823 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1824;
  assign dataGroup_hi_hi_1824 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1825;
  assign dataGroup_hi_hi_1825 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1826;
  assign dataGroup_hi_hi_1826 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1827;
  assign dataGroup_hi_hi_1827 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1828;
  assign dataGroup_hi_hi_1828 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1829;
  assign dataGroup_hi_hi_1829 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1830;
  assign dataGroup_hi_hi_1830 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1831;
  assign dataGroup_hi_hi_1831 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1832;
  assign dataGroup_hi_hi_1832 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1833;
  assign dataGroup_hi_hi_1833 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1834;
  assign dataGroup_hi_hi_1834 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1835;
  assign dataGroup_hi_hi_1835 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1836;
  assign dataGroup_hi_hi_1836 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1837;
  assign dataGroup_hi_hi_1837 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1838;
  assign dataGroup_hi_hi_1838 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1839;
  assign dataGroup_hi_hi_1839 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1840;
  assign dataGroup_hi_hi_1840 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1841;
  assign dataGroup_hi_hi_1841 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1842;
  assign dataGroup_hi_hi_1842 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1843;
  assign dataGroup_hi_hi_1843 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1844;
  assign dataGroup_hi_hi_1844 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1845;
  assign dataGroup_hi_hi_1845 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1846;
  assign dataGroup_hi_hi_1846 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1847;
  assign dataGroup_hi_hi_1847 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1848;
  assign dataGroup_hi_hi_1848 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1849;
  assign dataGroup_hi_hi_1849 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1850;
  assign dataGroup_hi_hi_1850 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1851;
  assign dataGroup_hi_hi_1851 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1852;
  assign dataGroup_hi_hi_1852 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1853;
  assign dataGroup_hi_hi_1853 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1854;
  assign dataGroup_hi_hi_1854 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1855;
  assign dataGroup_hi_hi_1855 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1856;
  assign dataGroup_hi_hi_1856 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1857;
  assign dataGroup_hi_hi_1857 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1858;
  assign dataGroup_hi_hi_1858 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1859;
  assign dataGroup_hi_hi_1859 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1860;
  assign dataGroup_hi_hi_1860 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1861;
  assign dataGroup_hi_hi_1861 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1862;
  assign dataGroup_hi_hi_1862 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1863;
  assign dataGroup_hi_hi_1863 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1864;
  assign dataGroup_hi_hi_1864 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1865;
  assign dataGroup_hi_hi_1865 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1866;
  assign dataGroup_hi_hi_1866 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1867;
  assign dataGroup_hi_hi_1867 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1868;
  assign dataGroup_hi_hi_1868 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1869;
  assign dataGroup_hi_hi_1869 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1870;
  assign dataGroup_hi_hi_1870 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1871;
  assign dataGroup_hi_hi_1871 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1872;
  assign dataGroup_hi_hi_1872 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1873;
  assign dataGroup_hi_hi_1873 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1874;
  assign dataGroup_hi_hi_1874 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1875;
  assign dataGroup_hi_hi_1875 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1876;
  assign dataGroup_hi_hi_1876 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1877;
  assign dataGroup_hi_hi_1877 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1878;
  assign dataGroup_hi_hi_1878 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1879;
  assign dataGroup_hi_hi_1879 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1880;
  assign dataGroup_hi_hi_1880 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1881;
  assign dataGroup_hi_hi_1881 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1882;
  assign dataGroup_hi_hi_1882 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1883;
  assign dataGroup_hi_hi_1883 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1884;
  assign dataGroup_hi_hi_1884 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1885;
  assign dataGroup_hi_hi_1885 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1886;
  assign dataGroup_hi_hi_1886 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1887;
  assign dataGroup_hi_hi_1887 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1888;
  assign dataGroup_hi_hi_1888 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1889;
  assign dataGroup_hi_hi_1889 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1890;
  assign dataGroup_hi_hi_1890 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1891;
  assign dataGroup_hi_hi_1891 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1892;
  assign dataGroup_hi_hi_1892 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1893;
  assign dataGroup_hi_hi_1893 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1894;
  assign dataGroup_hi_hi_1894 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1895;
  assign dataGroup_hi_hi_1895 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1896;
  assign dataGroup_hi_hi_1896 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1897;
  assign dataGroup_hi_hi_1897 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1898;
  assign dataGroup_hi_hi_1898 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1899;
  assign dataGroup_hi_hi_1899 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1900;
  assign dataGroup_hi_hi_1900 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1901;
  assign dataGroup_hi_hi_1901 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1902;
  assign dataGroup_hi_hi_1902 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1903;
  assign dataGroup_hi_hi_1903 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1904;
  assign dataGroup_hi_hi_1904 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1905;
  assign dataGroup_hi_hi_1905 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1906;
  assign dataGroup_hi_hi_1906 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1907;
  assign dataGroup_hi_hi_1907 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1908;
  assign dataGroup_hi_hi_1908 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1909;
  assign dataGroup_hi_hi_1909 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1910;
  assign dataGroup_hi_hi_1910 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1911;
  assign dataGroup_hi_hi_1911 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1912;
  assign dataGroup_hi_hi_1912 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1913;
  assign dataGroup_hi_hi_1913 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1914;
  assign dataGroup_hi_hi_1914 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1915;
  assign dataGroup_hi_hi_1915 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1916;
  assign dataGroup_hi_hi_1916 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1917;
  assign dataGroup_hi_hi_1917 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1918;
  assign dataGroup_hi_hi_1918 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1919;
  assign dataGroup_hi_hi_1919 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1920;
  assign dataGroup_hi_hi_1920 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1921;
  assign dataGroup_hi_hi_1921 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1922;
  assign dataGroup_hi_hi_1922 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1923;
  assign dataGroup_hi_hi_1923 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1924;
  assign dataGroup_hi_hi_1924 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1925;
  assign dataGroup_hi_hi_1925 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1926;
  assign dataGroup_hi_hi_1926 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1927;
  assign dataGroup_hi_hi_1927 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1928;
  assign dataGroup_hi_hi_1928 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1929;
  assign dataGroup_hi_hi_1929 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1930;
  assign dataGroup_hi_hi_1930 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1931;
  assign dataGroup_hi_hi_1931 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1932;
  assign dataGroup_hi_hi_1932 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1933;
  assign dataGroup_hi_hi_1933 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1934;
  assign dataGroup_hi_hi_1934 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1935;
  assign dataGroup_hi_hi_1935 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1936;
  assign dataGroup_hi_hi_1936 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1937;
  assign dataGroup_hi_hi_1937 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1938;
  assign dataGroup_hi_hi_1938 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1939;
  assign dataGroup_hi_hi_1939 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1940;
  assign dataGroup_hi_hi_1940 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1941;
  assign dataGroup_hi_hi_1941 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1942;
  assign dataGroup_hi_hi_1942 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1943;
  assign dataGroup_hi_hi_1943 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1944;
  assign dataGroup_hi_hi_1944 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1945;
  assign dataGroup_hi_hi_1945 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1946;
  assign dataGroup_hi_hi_1946 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1947;
  assign dataGroup_hi_hi_1947 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1948;
  assign dataGroup_hi_hi_1948 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1949;
  assign dataGroup_hi_hi_1949 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1950;
  assign dataGroup_hi_hi_1950 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1951;
  assign dataGroup_hi_hi_1951 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1952;
  assign dataGroup_hi_hi_1952 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1953;
  assign dataGroup_hi_hi_1953 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1954;
  assign dataGroup_hi_hi_1954 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1955;
  assign dataGroup_hi_hi_1955 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1956;
  assign dataGroup_hi_hi_1956 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1957;
  assign dataGroup_hi_hi_1957 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1958;
  assign dataGroup_hi_hi_1958 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1959;
  assign dataGroup_hi_hi_1959 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1960;
  assign dataGroup_hi_hi_1960 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1961;
  assign dataGroup_hi_hi_1961 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1962;
  assign dataGroup_hi_hi_1962 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1963;
  assign dataGroup_hi_hi_1963 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1964;
  assign dataGroup_hi_hi_1964 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1965;
  assign dataGroup_hi_hi_1965 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1966;
  assign dataGroup_hi_hi_1966 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1967;
  assign dataGroup_hi_hi_1967 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1968;
  assign dataGroup_hi_hi_1968 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1969;
  assign dataGroup_hi_hi_1969 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1970;
  assign dataGroup_hi_hi_1970 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1971;
  assign dataGroup_hi_hi_1971 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1972;
  assign dataGroup_hi_hi_1972 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1973;
  assign dataGroup_hi_hi_1973 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1974;
  assign dataGroup_hi_hi_1974 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1975;
  assign dataGroup_hi_hi_1975 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1976;
  assign dataGroup_hi_hi_1976 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1977;
  assign dataGroup_hi_hi_1977 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1978;
  assign dataGroup_hi_hi_1978 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1979;
  assign dataGroup_hi_hi_1979 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1980;
  assign dataGroup_hi_hi_1980 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1981;
  assign dataGroup_hi_hi_1981 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1982;
  assign dataGroup_hi_hi_1982 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1983;
  assign dataGroup_hi_hi_1983 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1984;
  assign dataGroup_hi_hi_1984 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1985;
  assign dataGroup_hi_hi_1985 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1986;
  assign dataGroup_hi_hi_1986 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1987;
  assign dataGroup_hi_hi_1987 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1988;
  assign dataGroup_hi_hi_1988 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1989;
  assign dataGroup_hi_hi_1989 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1990;
  assign dataGroup_hi_hi_1990 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1991;
  assign dataGroup_hi_hi_1991 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1992;
  assign dataGroup_hi_hi_1992 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1993;
  assign dataGroup_hi_hi_1993 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1994;
  assign dataGroup_hi_hi_1994 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1995;
  assign dataGroup_hi_hi_1995 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1996;
  assign dataGroup_hi_hi_1996 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1997;
  assign dataGroup_hi_hi_1997 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1998;
  assign dataGroup_hi_hi_1998 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_1999;
  assign dataGroup_hi_hi_1999 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2000;
  assign dataGroup_hi_hi_2000 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2001;
  assign dataGroup_hi_hi_2001 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2002;
  assign dataGroup_hi_hi_2002 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2003;
  assign dataGroup_hi_hi_2003 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2004;
  assign dataGroup_hi_hi_2004 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2005;
  assign dataGroup_hi_hi_2005 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2006;
  assign dataGroup_hi_hi_2006 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2007;
  assign dataGroup_hi_hi_2007 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2008;
  assign dataGroup_hi_hi_2008 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2009;
  assign dataGroup_hi_hi_2009 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2010;
  assign dataGroup_hi_hi_2010 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2011;
  assign dataGroup_hi_hi_2011 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2012;
  assign dataGroup_hi_hi_2012 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2013;
  assign dataGroup_hi_hi_2013 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2014;
  assign dataGroup_hi_hi_2014 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2015;
  assign dataGroup_hi_hi_2015 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2016;
  assign dataGroup_hi_hi_2016 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2017;
  assign dataGroup_hi_hi_2017 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2018;
  assign dataGroup_hi_hi_2018 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2019;
  assign dataGroup_hi_hi_2019 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2020;
  assign dataGroup_hi_hi_2020 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2021;
  assign dataGroup_hi_hi_2021 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2022;
  assign dataGroup_hi_hi_2022 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2023;
  assign dataGroup_hi_hi_2023 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2024;
  assign dataGroup_hi_hi_2024 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2025;
  assign dataGroup_hi_hi_2025 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2026;
  assign dataGroup_hi_hi_2026 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2027;
  assign dataGroup_hi_hi_2027 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2028;
  assign dataGroup_hi_hi_2028 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2029;
  assign dataGroup_hi_hi_2029 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2030;
  assign dataGroup_hi_hi_2030 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2031;
  assign dataGroup_hi_hi_2031 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2032;
  assign dataGroup_hi_hi_2032 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2033;
  assign dataGroup_hi_hi_2033 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2034;
  assign dataGroup_hi_hi_2034 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2035;
  assign dataGroup_hi_hi_2035 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2036;
  assign dataGroup_hi_hi_2036 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2037;
  assign dataGroup_hi_hi_2037 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2038;
  assign dataGroup_hi_hi_2038 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2039;
  assign dataGroup_hi_hi_2039 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2040;
  assign dataGroup_hi_hi_2040 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2041;
  assign dataGroup_hi_hi_2041 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2042;
  assign dataGroup_hi_hi_2042 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2043;
  assign dataGroup_hi_hi_2043 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2044;
  assign dataGroup_hi_hi_2044 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2045;
  assign dataGroup_hi_hi_2045 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2046;
  assign dataGroup_hi_hi_2046 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2047;
  assign dataGroup_hi_hi_2047 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2048;
  assign dataGroup_hi_hi_2048 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2049;
  assign dataGroup_hi_hi_2049 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2050;
  assign dataGroup_hi_hi_2050 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2051;
  assign dataGroup_hi_hi_2051 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2052;
  assign dataGroup_hi_hi_2052 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2053;
  assign dataGroup_hi_hi_2053 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2054;
  assign dataGroup_hi_hi_2054 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2055;
  assign dataGroup_hi_hi_2055 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2056;
  assign dataGroup_hi_hi_2056 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2057;
  assign dataGroup_hi_hi_2057 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2058;
  assign dataGroup_hi_hi_2058 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2059;
  assign dataGroup_hi_hi_2059 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2060;
  assign dataGroup_hi_hi_2060 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2061;
  assign dataGroup_hi_hi_2061 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2062;
  assign dataGroup_hi_hi_2062 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2063;
  assign dataGroup_hi_hi_2063 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2064;
  assign dataGroup_hi_hi_2064 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2065;
  assign dataGroup_hi_hi_2065 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2066;
  assign dataGroup_hi_hi_2066 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2067;
  assign dataGroup_hi_hi_2067 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2068;
  assign dataGroup_hi_hi_2068 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2069;
  assign dataGroup_hi_hi_2069 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2070;
  assign dataGroup_hi_hi_2070 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2071;
  assign dataGroup_hi_hi_2071 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2072;
  assign dataGroup_hi_hi_2072 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2073;
  assign dataGroup_hi_hi_2073 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2074;
  assign dataGroup_hi_hi_2074 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2075;
  assign dataGroup_hi_hi_2075 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2076;
  assign dataGroup_hi_hi_2076 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2077;
  assign dataGroup_hi_hi_2077 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2078;
  assign dataGroup_hi_hi_2078 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2079;
  assign dataGroup_hi_hi_2079 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2080;
  assign dataGroup_hi_hi_2080 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2081;
  assign dataGroup_hi_hi_2081 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2082;
  assign dataGroup_hi_hi_2082 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2083;
  assign dataGroup_hi_hi_2083 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2084;
  assign dataGroup_hi_hi_2084 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2085;
  assign dataGroup_hi_hi_2085 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2086;
  assign dataGroup_hi_hi_2086 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2087;
  assign dataGroup_hi_hi_2087 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2088;
  assign dataGroup_hi_hi_2088 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2089;
  assign dataGroup_hi_hi_2089 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2090;
  assign dataGroup_hi_hi_2090 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2091;
  assign dataGroup_hi_hi_2091 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2092;
  assign dataGroup_hi_hi_2092 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2093;
  assign dataGroup_hi_hi_2093 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2094;
  assign dataGroup_hi_hi_2094 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2095;
  assign dataGroup_hi_hi_2095 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2096;
  assign dataGroup_hi_hi_2096 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2097;
  assign dataGroup_hi_hi_2097 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2098;
  assign dataGroup_hi_hi_2098 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2099;
  assign dataGroup_hi_hi_2099 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2100;
  assign dataGroup_hi_hi_2100 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2101;
  assign dataGroup_hi_hi_2101 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2102;
  assign dataGroup_hi_hi_2102 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2103;
  assign dataGroup_hi_hi_2103 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2104;
  assign dataGroup_hi_hi_2104 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2105;
  assign dataGroup_hi_hi_2105 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2106;
  assign dataGroup_hi_hi_2106 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2107;
  assign dataGroup_hi_hi_2107 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2108;
  assign dataGroup_hi_hi_2108 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2109;
  assign dataGroup_hi_hi_2109 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2110;
  assign dataGroup_hi_hi_2110 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2111;
  assign dataGroup_hi_hi_2111 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2112;
  assign dataGroup_hi_hi_2112 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2113;
  assign dataGroup_hi_hi_2113 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2114;
  assign dataGroup_hi_hi_2114 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2115;
  assign dataGroup_hi_hi_2115 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2116;
  assign dataGroup_hi_hi_2116 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2117;
  assign dataGroup_hi_hi_2117 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2118;
  assign dataGroup_hi_hi_2118 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2119;
  assign dataGroup_hi_hi_2119 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2120;
  assign dataGroup_hi_hi_2120 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2121;
  assign dataGroup_hi_hi_2121 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2122;
  assign dataGroup_hi_hi_2122 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2123;
  assign dataGroup_hi_hi_2123 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2124;
  assign dataGroup_hi_hi_2124 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2125;
  assign dataGroup_hi_hi_2125 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2126;
  assign dataGroup_hi_hi_2126 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2127;
  assign dataGroup_hi_hi_2127 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2128;
  assign dataGroup_hi_hi_2128 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2129;
  assign dataGroup_hi_hi_2129 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2130;
  assign dataGroup_hi_hi_2130 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2131;
  assign dataGroup_hi_hi_2131 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2132;
  assign dataGroup_hi_hi_2132 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2133;
  assign dataGroup_hi_hi_2133 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2134;
  assign dataGroup_hi_hi_2134 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2135;
  assign dataGroup_hi_hi_2135 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2136;
  assign dataGroup_hi_hi_2136 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2137;
  assign dataGroup_hi_hi_2137 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2138;
  assign dataGroup_hi_hi_2138 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2139;
  assign dataGroup_hi_hi_2139 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2140;
  assign dataGroup_hi_hi_2140 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2141;
  assign dataGroup_hi_hi_2141 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2142;
  assign dataGroup_hi_hi_2142 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2143;
  assign dataGroup_hi_hi_2143 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2144;
  assign dataGroup_hi_hi_2144 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2145;
  assign dataGroup_hi_hi_2145 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2146;
  assign dataGroup_hi_hi_2146 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2147;
  assign dataGroup_hi_hi_2147 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2148;
  assign dataGroup_hi_hi_2148 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2149;
  assign dataGroup_hi_hi_2149 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2150;
  assign dataGroup_hi_hi_2150 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2151;
  assign dataGroup_hi_hi_2151 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2152;
  assign dataGroup_hi_hi_2152 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2153;
  assign dataGroup_hi_hi_2153 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2154;
  assign dataGroup_hi_hi_2154 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2155;
  assign dataGroup_hi_hi_2155 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2156;
  assign dataGroup_hi_hi_2156 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2157;
  assign dataGroup_hi_hi_2157 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2158;
  assign dataGroup_hi_hi_2158 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2159;
  assign dataGroup_hi_hi_2159 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2160;
  assign dataGroup_hi_hi_2160 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2161;
  assign dataGroup_hi_hi_2161 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2162;
  assign dataGroup_hi_hi_2162 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2163;
  assign dataGroup_hi_hi_2163 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2164;
  assign dataGroup_hi_hi_2164 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2165;
  assign dataGroup_hi_hi_2165 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2166;
  assign dataGroup_hi_hi_2166 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2167;
  assign dataGroup_hi_hi_2167 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2168;
  assign dataGroup_hi_hi_2168 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2169;
  assign dataGroup_hi_hi_2169 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2170;
  assign dataGroup_hi_hi_2170 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2171;
  assign dataGroup_hi_hi_2171 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2172;
  assign dataGroup_hi_hi_2172 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2173;
  assign dataGroup_hi_hi_2173 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2174;
  assign dataGroup_hi_hi_2174 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2175;
  assign dataGroup_hi_hi_2175 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2176;
  assign dataGroup_hi_hi_2176 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2177;
  assign dataGroup_hi_hi_2177 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2178;
  assign dataGroup_hi_hi_2178 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2179;
  assign dataGroup_hi_hi_2179 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2180;
  assign dataGroup_hi_hi_2180 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2181;
  assign dataGroup_hi_hi_2181 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2182;
  assign dataGroup_hi_hi_2182 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2183;
  assign dataGroup_hi_hi_2183 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2184;
  assign dataGroup_hi_hi_2184 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2185;
  assign dataGroup_hi_hi_2185 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2186;
  assign dataGroup_hi_hi_2186 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2187;
  assign dataGroup_hi_hi_2187 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2188;
  assign dataGroup_hi_hi_2188 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2189;
  assign dataGroup_hi_hi_2189 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2190;
  assign dataGroup_hi_hi_2190 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2191;
  assign dataGroup_hi_hi_2191 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2192;
  assign dataGroup_hi_hi_2192 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2193;
  assign dataGroup_hi_hi_2193 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2194;
  assign dataGroup_hi_hi_2194 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2195;
  assign dataGroup_hi_hi_2195 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2196;
  assign dataGroup_hi_hi_2196 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2197;
  assign dataGroup_hi_hi_2197 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2198;
  assign dataGroup_hi_hi_2198 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2199;
  assign dataGroup_hi_hi_2199 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2200;
  assign dataGroup_hi_hi_2200 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2201;
  assign dataGroup_hi_hi_2201 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2202;
  assign dataGroup_hi_hi_2202 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2203;
  assign dataGroup_hi_hi_2203 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2204;
  assign dataGroup_hi_hi_2204 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2205;
  assign dataGroup_hi_hi_2205 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2206;
  assign dataGroup_hi_hi_2206 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2207;
  assign dataGroup_hi_hi_2207 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2208;
  assign dataGroup_hi_hi_2208 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2209;
  assign dataGroup_hi_hi_2209 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2210;
  assign dataGroup_hi_hi_2210 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2211;
  assign dataGroup_hi_hi_2211 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2212;
  assign dataGroup_hi_hi_2212 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2213;
  assign dataGroup_hi_hi_2213 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2214;
  assign dataGroup_hi_hi_2214 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2215;
  assign dataGroup_hi_hi_2215 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2216;
  assign dataGroup_hi_hi_2216 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2217;
  assign dataGroup_hi_hi_2217 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2218;
  assign dataGroup_hi_hi_2218 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2219;
  assign dataGroup_hi_hi_2219 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2220;
  assign dataGroup_hi_hi_2220 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2221;
  assign dataGroup_hi_hi_2221 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2222;
  assign dataGroup_hi_hi_2222 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2223;
  assign dataGroup_hi_hi_2223 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2224;
  assign dataGroup_hi_hi_2224 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2225;
  assign dataGroup_hi_hi_2225 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2226;
  assign dataGroup_hi_hi_2226 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2227;
  assign dataGroup_hi_hi_2227 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2228;
  assign dataGroup_hi_hi_2228 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2229;
  assign dataGroup_hi_hi_2229 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2230;
  assign dataGroup_hi_hi_2230 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2231;
  assign dataGroup_hi_hi_2231 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2232;
  assign dataGroup_hi_hi_2232 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2233;
  assign dataGroup_hi_hi_2233 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2234;
  assign dataGroup_hi_hi_2234 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2235;
  assign dataGroup_hi_hi_2235 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2236;
  assign dataGroup_hi_hi_2236 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2237;
  assign dataGroup_hi_hi_2237 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2238;
  assign dataGroup_hi_hi_2238 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2239;
  assign dataGroup_hi_hi_2239 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2240;
  assign dataGroup_hi_hi_2240 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2241;
  assign dataGroup_hi_hi_2241 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2242;
  assign dataGroup_hi_hi_2242 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2243;
  assign dataGroup_hi_hi_2243 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2244;
  assign dataGroup_hi_hi_2244 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2245;
  assign dataGroup_hi_hi_2245 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2246;
  assign dataGroup_hi_hi_2246 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2247;
  assign dataGroup_hi_hi_2247 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2248;
  assign dataGroup_hi_hi_2248 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2249;
  assign dataGroup_hi_hi_2249 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2250;
  assign dataGroup_hi_hi_2250 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2251;
  assign dataGroup_hi_hi_2251 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2252;
  assign dataGroup_hi_hi_2252 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2253;
  assign dataGroup_hi_hi_2253 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2254;
  assign dataGroup_hi_hi_2254 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2255;
  assign dataGroup_hi_hi_2255 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2256;
  assign dataGroup_hi_hi_2256 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2257;
  assign dataGroup_hi_hi_2257 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2258;
  assign dataGroup_hi_hi_2258 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2259;
  assign dataGroup_hi_hi_2259 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2260;
  assign dataGroup_hi_hi_2260 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2261;
  assign dataGroup_hi_hi_2261 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2262;
  assign dataGroup_hi_hi_2262 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2263;
  assign dataGroup_hi_hi_2263 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2264;
  assign dataGroup_hi_hi_2264 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2265;
  assign dataGroup_hi_hi_2265 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2266;
  assign dataGroup_hi_hi_2266 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2267;
  assign dataGroup_hi_hi_2267 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2268;
  assign dataGroup_hi_hi_2268 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2269;
  assign dataGroup_hi_hi_2269 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2270;
  assign dataGroup_hi_hi_2270 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2271;
  assign dataGroup_hi_hi_2271 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2272;
  assign dataGroup_hi_hi_2272 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2273;
  assign dataGroup_hi_hi_2273 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2274;
  assign dataGroup_hi_hi_2274 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2275;
  assign dataGroup_hi_hi_2275 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2276;
  assign dataGroup_hi_hi_2276 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2277;
  assign dataGroup_hi_hi_2277 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2278;
  assign dataGroup_hi_hi_2278 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2279;
  assign dataGroup_hi_hi_2279 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2280;
  assign dataGroup_hi_hi_2280 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2281;
  assign dataGroup_hi_hi_2281 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2282;
  assign dataGroup_hi_hi_2282 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2283;
  assign dataGroup_hi_hi_2283 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2284;
  assign dataGroup_hi_hi_2284 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2285;
  assign dataGroup_hi_hi_2285 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2286;
  assign dataGroup_hi_hi_2286 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2287;
  assign dataGroup_hi_hi_2287 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2288;
  assign dataGroup_hi_hi_2288 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2289;
  assign dataGroup_hi_hi_2289 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2290;
  assign dataGroup_hi_hi_2290 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2291;
  assign dataGroup_hi_hi_2291 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2292;
  assign dataGroup_hi_hi_2292 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2293;
  assign dataGroup_hi_hi_2293 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2294;
  assign dataGroup_hi_hi_2294 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2295;
  assign dataGroup_hi_hi_2295 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2296;
  assign dataGroup_hi_hi_2296 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2297;
  assign dataGroup_hi_hi_2297 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2298;
  assign dataGroup_hi_hi_2298 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2299;
  assign dataGroup_hi_hi_2299 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2300;
  assign dataGroup_hi_hi_2300 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2301;
  assign dataGroup_hi_hi_2301 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2302;
  assign dataGroup_hi_hi_2302 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2303;
  assign dataGroup_hi_hi_2303 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2304;
  assign dataGroup_hi_hi_2304 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2305;
  assign dataGroup_hi_hi_2305 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2306;
  assign dataGroup_hi_hi_2306 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2307;
  assign dataGroup_hi_hi_2307 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2308;
  assign dataGroup_hi_hi_2308 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2309;
  assign dataGroup_hi_hi_2309 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2310;
  assign dataGroup_hi_hi_2310 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2311;
  assign dataGroup_hi_hi_2311 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2312;
  assign dataGroup_hi_hi_2312 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2313;
  assign dataGroup_hi_hi_2313 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2314;
  assign dataGroup_hi_hi_2314 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2315;
  assign dataGroup_hi_hi_2315 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2316;
  assign dataGroup_hi_hi_2316 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2317;
  assign dataGroup_hi_hi_2317 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2318;
  assign dataGroup_hi_hi_2318 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2319;
  assign dataGroup_hi_hi_2319 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2320;
  assign dataGroup_hi_hi_2320 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2321;
  assign dataGroup_hi_hi_2321 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2322;
  assign dataGroup_hi_hi_2322 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2323;
  assign dataGroup_hi_hi_2323 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2324;
  assign dataGroup_hi_hi_2324 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2325;
  assign dataGroup_hi_hi_2325 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2326;
  assign dataGroup_hi_hi_2326 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2327;
  assign dataGroup_hi_hi_2327 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2328;
  assign dataGroup_hi_hi_2328 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2329;
  assign dataGroup_hi_hi_2329 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2330;
  assign dataGroup_hi_hi_2330 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2331;
  assign dataGroup_hi_hi_2331 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2332;
  assign dataGroup_hi_hi_2332 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2333;
  assign dataGroup_hi_hi_2333 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2334;
  assign dataGroup_hi_hi_2334 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2335;
  assign dataGroup_hi_hi_2335 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2336;
  assign dataGroup_hi_hi_2336 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2337;
  assign dataGroup_hi_hi_2337 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2338;
  assign dataGroup_hi_hi_2338 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2339;
  assign dataGroup_hi_hi_2339 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2340;
  assign dataGroup_hi_hi_2340 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2341;
  assign dataGroup_hi_hi_2341 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2342;
  assign dataGroup_hi_hi_2342 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2343;
  assign dataGroup_hi_hi_2343 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2344;
  assign dataGroup_hi_hi_2344 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2345;
  assign dataGroup_hi_hi_2345 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2346;
  assign dataGroup_hi_hi_2346 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2347;
  assign dataGroup_hi_hi_2347 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2348;
  assign dataGroup_hi_hi_2348 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2349;
  assign dataGroup_hi_hi_2349 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2350;
  assign dataGroup_hi_hi_2350 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2351;
  assign dataGroup_hi_hi_2351 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2352;
  assign dataGroup_hi_hi_2352 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2353;
  assign dataGroup_hi_hi_2353 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2354;
  assign dataGroup_hi_hi_2354 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2355;
  assign dataGroup_hi_hi_2355 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2356;
  assign dataGroup_hi_hi_2356 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2357;
  assign dataGroup_hi_hi_2357 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2358;
  assign dataGroup_hi_hi_2358 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2359;
  assign dataGroup_hi_hi_2359 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2360;
  assign dataGroup_hi_hi_2360 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2361;
  assign dataGroup_hi_hi_2361 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2362;
  assign dataGroup_hi_hi_2362 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2363;
  assign dataGroup_hi_hi_2363 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2364;
  assign dataGroup_hi_hi_2364 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2365;
  assign dataGroup_hi_hi_2365 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2366;
  assign dataGroup_hi_hi_2366 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2367;
  assign dataGroup_hi_hi_2367 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2368;
  assign dataGroup_hi_hi_2368 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2369;
  assign dataGroup_hi_hi_2369 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2370;
  assign dataGroup_hi_hi_2370 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2371;
  assign dataGroup_hi_hi_2371 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2372;
  assign dataGroup_hi_hi_2372 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2373;
  assign dataGroup_hi_hi_2373 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2374;
  assign dataGroup_hi_hi_2374 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2375;
  assign dataGroup_hi_hi_2375 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2376;
  assign dataGroup_hi_hi_2376 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2377;
  assign dataGroup_hi_hi_2377 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2378;
  assign dataGroup_hi_hi_2378 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2379;
  assign dataGroup_hi_hi_2379 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2380;
  assign dataGroup_hi_hi_2380 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2381;
  assign dataGroup_hi_hi_2381 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2382;
  assign dataGroup_hi_hi_2382 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2383;
  assign dataGroup_hi_hi_2383 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2384;
  assign dataGroup_hi_hi_2384 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2385;
  assign dataGroup_hi_hi_2385 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2386;
  assign dataGroup_hi_hi_2386 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2387;
  assign dataGroup_hi_hi_2387 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2388;
  assign dataGroup_hi_hi_2388 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2389;
  assign dataGroup_hi_hi_2389 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2390;
  assign dataGroup_hi_hi_2390 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2391;
  assign dataGroup_hi_hi_2391 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2392;
  assign dataGroup_hi_hi_2392 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2393;
  assign dataGroup_hi_hi_2393 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2394;
  assign dataGroup_hi_hi_2394 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2395;
  assign dataGroup_hi_hi_2395 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2396;
  assign dataGroup_hi_hi_2396 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2397;
  assign dataGroup_hi_hi_2397 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2398;
  assign dataGroup_hi_hi_2398 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2399;
  assign dataGroup_hi_hi_2399 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2400;
  assign dataGroup_hi_hi_2400 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2401;
  assign dataGroup_hi_hi_2401 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2402;
  assign dataGroup_hi_hi_2402 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2403;
  assign dataGroup_hi_hi_2403 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2404;
  assign dataGroup_hi_hi_2404 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2405;
  assign dataGroup_hi_hi_2405 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2406;
  assign dataGroup_hi_hi_2406 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2407;
  assign dataGroup_hi_hi_2407 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2408;
  assign dataGroup_hi_hi_2408 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2409;
  assign dataGroup_hi_hi_2409 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2410;
  assign dataGroup_hi_hi_2410 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2411;
  assign dataGroup_hi_hi_2411 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2412;
  assign dataGroup_hi_hi_2412 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2413;
  assign dataGroup_hi_hi_2413 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2414;
  assign dataGroup_hi_hi_2414 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2415;
  assign dataGroup_hi_hi_2415 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2416;
  assign dataGroup_hi_hi_2416 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2417;
  assign dataGroup_hi_hi_2417 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2418;
  assign dataGroup_hi_hi_2418 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2419;
  assign dataGroup_hi_hi_2419 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2420;
  assign dataGroup_hi_hi_2420 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2421;
  assign dataGroup_hi_hi_2421 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2422;
  assign dataGroup_hi_hi_2422 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2423;
  assign dataGroup_hi_hi_2423 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2424;
  assign dataGroup_hi_hi_2424 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2425;
  assign dataGroup_hi_hi_2425 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2426;
  assign dataGroup_hi_hi_2426 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2427;
  assign dataGroup_hi_hi_2427 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2428;
  assign dataGroup_hi_hi_2428 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2429;
  assign dataGroup_hi_hi_2429 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2430;
  assign dataGroup_hi_hi_2430 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2431;
  assign dataGroup_hi_hi_2431 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2432;
  assign dataGroup_hi_hi_2432 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2433;
  assign dataGroup_hi_hi_2433 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2434;
  assign dataGroup_hi_hi_2434 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2435;
  assign dataGroup_hi_hi_2435 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2436;
  assign dataGroup_hi_hi_2436 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2437;
  assign dataGroup_hi_hi_2437 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2438;
  assign dataGroup_hi_hi_2438 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2439;
  assign dataGroup_hi_hi_2439 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2440;
  assign dataGroup_hi_hi_2440 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2441;
  assign dataGroup_hi_hi_2441 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2442;
  assign dataGroup_hi_hi_2442 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2443;
  assign dataGroup_hi_hi_2443 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2444;
  assign dataGroup_hi_hi_2444 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2445;
  assign dataGroup_hi_hi_2445 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2446;
  assign dataGroup_hi_hi_2446 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2447;
  assign dataGroup_hi_hi_2447 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2448;
  assign dataGroup_hi_hi_2448 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2449;
  assign dataGroup_hi_hi_2449 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2450;
  assign dataGroup_hi_hi_2450 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2451;
  assign dataGroup_hi_hi_2451 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2452;
  assign dataGroup_hi_hi_2452 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2453;
  assign dataGroup_hi_hi_2453 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2454;
  assign dataGroup_hi_hi_2454 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2455;
  assign dataGroup_hi_hi_2455 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2456;
  assign dataGroup_hi_hi_2456 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2457;
  assign dataGroup_hi_hi_2457 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2458;
  assign dataGroup_hi_hi_2458 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2459;
  assign dataGroup_hi_hi_2459 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2460;
  assign dataGroup_hi_hi_2460 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2461;
  assign dataGroup_hi_hi_2461 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2462;
  assign dataGroup_hi_hi_2462 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2463;
  assign dataGroup_hi_hi_2463 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2464;
  assign dataGroup_hi_hi_2464 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2465;
  assign dataGroup_hi_hi_2465 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2466;
  assign dataGroup_hi_hi_2466 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2467;
  assign dataGroup_hi_hi_2467 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2468;
  assign dataGroup_hi_hi_2468 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2469;
  assign dataGroup_hi_hi_2469 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2470;
  assign dataGroup_hi_hi_2470 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2471;
  assign dataGroup_hi_hi_2471 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2472;
  assign dataGroup_hi_hi_2472 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2473;
  assign dataGroup_hi_hi_2473 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2474;
  assign dataGroup_hi_hi_2474 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2475;
  assign dataGroup_hi_hi_2475 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2476;
  assign dataGroup_hi_hi_2476 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2477;
  assign dataGroup_hi_hi_2477 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2478;
  assign dataGroup_hi_hi_2478 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2479;
  assign dataGroup_hi_hi_2479 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2480;
  assign dataGroup_hi_hi_2480 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2481;
  assign dataGroup_hi_hi_2481 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2482;
  assign dataGroup_hi_hi_2482 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2483;
  assign dataGroup_hi_hi_2483 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2484;
  assign dataGroup_hi_hi_2484 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2485;
  assign dataGroup_hi_hi_2485 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2486;
  assign dataGroup_hi_hi_2486 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2487;
  assign dataGroup_hi_hi_2487 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2488;
  assign dataGroup_hi_hi_2488 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2489;
  assign dataGroup_hi_hi_2489 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2490;
  assign dataGroup_hi_hi_2490 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2491;
  assign dataGroup_hi_hi_2491 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2492;
  assign dataGroup_hi_hi_2492 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2493;
  assign dataGroup_hi_hi_2493 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2494;
  assign dataGroup_hi_hi_2494 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2495;
  assign dataGroup_hi_hi_2495 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2496;
  assign dataGroup_hi_hi_2496 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2497;
  assign dataGroup_hi_hi_2497 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2498;
  assign dataGroup_hi_hi_2498 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2499;
  assign dataGroup_hi_hi_2499 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2500;
  assign dataGroup_hi_hi_2500 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2501;
  assign dataGroup_hi_hi_2501 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2502;
  assign dataGroup_hi_hi_2502 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2503;
  assign dataGroup_hi_hi_2503 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2504;
  assign dataGroup_hi_hi_2504 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2505;
  assign dataGroup_hi_hi_2505 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2506;
  assign dataGroup_hi_hi_2506 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2507;
  assign dataGroup_hi_hi_2507 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2508;
  assign dataGroup_hi_hi_2508 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2509;
  assign dataGroup_hi_hi_2509 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2510;
  assign dataGroup_hi_hi_2510 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2511;
  assign dataGroup_hi_hi_2511 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2512;
  assign dataGroup_hi_hi_2512 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2513;
  assign dataGroup_hi_hi_2513 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2514;
  assign dataGroup_hi_hi_2514 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2515;
  assign dataGroup_hi_hi_2515 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2516;
  assign dataGroup_hi_hi_2516 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2517;
  assign dataGroup_hi_hi_2517 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2518;
  assign dataGroup_hi_hi_2518 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2519;
  assign dataGroup_hi_hi_2519 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2520;
  assign dataGroup_hi_hi_2520 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2521;
  assign dataGroup_hi_hi_2521 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2522;
  assign dataGroup_hi_hi_2522 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2523;
  assign dataGroup_hi_hi_2523 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2524;
  assign dataGroup_hi_hi_2524 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2525;
  assign dataGroup_hi_hi_2525 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2526;
  assign dataGroup_hi_hi_2526 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2527;
  assign dataGroup_hi_hi_2527 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2528;
  assign dataGroup_hi_hi_2528 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2529;
  assign dataGroup_hi_hi_2529 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2530;
  assign dataGroup_hi_hi_2530 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2531;
  assign dataGroup_hi_hi_2531 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2532;
  assign dataGroup_hi_hi_2532 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2533;
  assign dataGroup_hi_hi_2533 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2534;
  assign dataGroup_hi_hi_2534 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2535;
  assign dataGroup_hi_hi_2535 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2536;
  assign dataGroup_hi_hi_2536 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2537;
  assign dataGroup_hi_hi_2537 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2538;
  assign dataGroup_hi_hi_2538 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2539;
  assign dataGroup_hi_hi_2539 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2540;
  assign dataGroup_hi_hi_2540 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2541;
  assign dataGroup_hi_hi_2541 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2542;
  assign dataGroup_hi_hi_2542 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2543;
  assign dataGroup_hi_hi_2543 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2544;
  assign dataGroup_hi_hi_2544 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2545;
  assign dataGroup_hi_hi_2545 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2546;
  assign dataGroup_hi_hi_2546 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2547;
  assign dataGroup_hi_hi_2547 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2548;
  assign dataGroup_hi_hi_2548 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2549;
  assign dataGroup_hi_hi_2549 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2550;
  assign dataGroup_hi_hi_2550 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2551;
  assign dataGroup_hi_hi_2551 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2552;
  assign dataGroup_hi_hi_2552 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2553;
  assign dataGroup_hi_hi_2553 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2554;
  assign dataGroup_hi_hi_2554 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2555;
  assign dataGroup_hi_hi_2555 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2556;
  assign dataGroup_hi_hi_2556 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2557;
  assign dataGroup_hi_hi_2557 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2558;
  assign dataGroup_hi_hi_2558 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2559;
  assign dataGroup_hi_hi_2559 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2560;
  assign dataGroup_hi_hi_2560 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2561;
  assign dataGroup_hi_hi_2561 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2562;
  assign dataGroup_hi_hi_2562 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2563;
  assign dataGroup_hi_hi_2563 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2564;
  assign dataGroup_hi_hi_2564 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2565;
  assign dataGroup_hi_hi_2565 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2566;
  assign dataGroup_hi_hi_2566 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2567;
  assign dataGroup_hi_hi_2567 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2568;
  assign dataGroup_hi_hi_2568 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2569;
  assign dataGroup_hi_hi_2569 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2570;
  assign dataGroup_hi_hi_2570 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2571;
  assign dataGroup_hi_hi_2571 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2572;
  assign dataGroup_hi_hi_2572 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2573;
  assign dataGroup_hi_hi_2573 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2574;
  assign dataGroup_hi_hi_2574 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2575;
  assign dataGroup_hi_hi_2575 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2576;
  assign dataGroup_hi_hi_2576 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2577;
  assign dataGroup_hi_hi_2577 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2578;
  assign dataGroup_hi_hi_2578 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2579;
  assign dataGroup_hi_hi_2579 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2580;
  assign dataGroup_hi_hi_2580 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2581;
  assign dataGroup_hi_hi_2581 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2582;
  assign dataGroup_hi_hi_2582 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2583;
  assign dataGroup_hi_hi_2583 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2584;
  assign dataGroup_hi_hi_2584 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2585;
  assign dataGroup_hi_hi_2585 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2586;
  assign dataGroup_hi_hi_2586 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2587;
  assign dataGroup_hi_hi_2587 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2588;
  assign dataGroup_hi_hi_2588 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2589;
  assign dataGroup_hi_hi_2589 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2590;
  assign dataGroup_hi_hi_2590 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2591;
  assign dataGroup_hi_hi_2591 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2592;
  assign dataGroup_hi_hi_2592 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2593;
  assign dataGroup_hi_hi_2593 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2594;
  assign dataGroup_hi_hi_2594 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2595;
  assign dataGroup_hi_hi_2595 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2596;
  assign dataGroup_hi_hi_2596 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2597;
  assign dataGroup_hi_hi_2597 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2598;
  assign dataGroup_hi_hi_2598 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2599;
  assign dataGroup_hi_hi_2599 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2600;
  assign dataGroup_hi_hi_2600 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2601;
  assign dataGroup_hi_hi_2601 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2602;
  assign dataGroup_hi_hi_2602 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2603;
  assign dataGroup_hi_hi_2603 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2604;
  assign dataGroup_hi_hi_2604 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2605;
  assign dataGroup_hi_hi_2605 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2606;
  assign dataGroup_hi_hi_2606 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2607;
  assign dataGroup_hi_hi_2607 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2608;
  assign dataGroup_hi_hi_2608 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2609;
  assign dataGroup_hi_hi_2609 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2610;
  assign dataGroup_hi_hi_2610 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2611;
  assign dataGroup_hi_hi_2611 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2612;
  assign dataGroup_hi_hi_2612 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2613;
  assign dataGroup_hi_hi_2613 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2614;
  assign dataGroup_hi_hi_2614 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2615;
  assign dataGroup_hi_hi_2615 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2616;
  assign dataGroup_hi_hi_2616 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2617;
  assign dataGroup_hi_hi_2617 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2618;
  assign dataGroup_hi_hi_2618 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2619;
  assign dataGroup_hi_hi_2619 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2620;
  assign dataGroup_hi_hi_2620 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2621;
  assign dataGroup_hi_hi_2621 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2622;
  assign dataGroup_hi_hi_2622 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2623;
  assign dataGroup_hi_hi_2623 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2624;
  assign dataGroup_hi_hi_2624 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2625;
  assign dataGroup_hi_hi_2625 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2626;
  assign dataGroup_hi_hi_2626 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2627;
  assign dataGroup_hi_hi_2627 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2628;
  assign dataGroup_hi_hi_2628 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2629;
  assign dataGroup_hi_hi_2629 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2630;
  assign dataGroup_hi_hi_2630 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2631;
  assign dataGroup_hi_hi_2631 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2632;
  assign dataGroup_hi_hi_2632 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2633;
  assign dataGroup_hi_hi_2633 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2634;
  assign dataGroup_hi_hi_2634 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2635;
  assign dataGroup_hi_hi_2635 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2636;
  assign dataGroup_hi_hi_2636 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2637;
  assign dataGroup_hi_hi_2637 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2638;
  assign dataGroup_hi_hi_2638 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2639;
  assign dataGroup_hi_hi_2639 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2640;
  assign dataGroup_hi_hi_2640 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2641;
  assign dataGroup_hi_hi_2641 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2642;
  assign dataGroup_hi_hi_2642 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2643;
  assign dataGroup_hi_hi_2643 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2644;
  assign dataGroup_hi_hi_2644 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2645;
  assign dataGroup_hi_hi_2645 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2646;
  assign dataGroup_hi_hi_2646 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2647;
  assign dataGroup_hi_hi_2647 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2648;
  assign dataGroup_hi_hi_2648 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2649;
  assign dataGroup_hi_hi_2649 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2650;
  assign dataGroup_hi_hi_2650 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2651;
  assign dataGroup_hi_hi_2651 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2652;
  assign dataGroup_hi_hi_2652 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2653;
  assign dataGroup_hi_hi_2653 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2654;
  assign dataGroup_hi_hi_2654 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2655;
  assign dataGroup_hi_hi_2655 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2656;
  assign dataGroup_hi_hi_2656 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2657;
  assign dataGroup_hi_hi_2657 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2658;
  assign dataGroup_hi_hi_2658 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2659;
  assign dataGroup_hi_hi_2659 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2660;
  assign dataGroup_hi_hi_2660 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2661;
  assign dataGroup_hi_hi_2661 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2662;
  assign dataGroup_hi_hi_2662 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2663;
  assign dataGroup_hi_hi_2663 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2664;
  assign dataGroup_hi_hi_2664 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2665;
  assign dataGroup_hi_hi_2665 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2666;
  assign dataGroup_hi_hi_2666 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2667;
  assign dataGroup_hi_hi_2667 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2668;
  assign dataGroup_hi_hi_2668 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2669;
  assign dataGroup_hi_hi_2669 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2670;
  assign dataGroup_hi_hi_2670 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2671;
  assign dataGroup_hi_hi_2671 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2672;
  assign dataGroup_hi_hi_2672 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2673;
  assign dataGroup_hi_hi_2673 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2674;
  assign dataGroup_hi_hi_2674 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2675;
  assign dataGroup_hi_hi_2675 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2676;
  assign dataGroup_hi_hi_2676 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2677;
  assign dataGroup_hi_hi_2677 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2678;
  assign dataGroup_hi_hi_2678 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2679;
  assign dataGroup_hi_hi_2679 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2680;
  assign dataGroup_hi_hi_2680 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2681;
  assign dataGroup_hi_hi_2681 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2682;
  assign dataGroup_hi_hi_2682 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2683;
  assign dataGroup_hi_hi_2683 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2684;
  assign dataGroup_hi_hi_2684 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2685;
  assign dataGroup_hi_hi_2685 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2686;
  assign dataGroup_hi_hi_2686 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2687;
  assign dataGroup_hi_hi_2687 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2688;
  assign dataGroup_hi_hi_2688 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2689;
  assign dataGroup_hi_hi_2689 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2690;
  assign dataGroup_hi_hi_2690 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2691;
  assign dataGroup_hi_hi_2691 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2692;
  assign dataGroup_hi_hi_2692 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2693;
  assign dataGroup_hi_hi_2693 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2694;
  assign dataGroup_hi_hi_2694 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2695;
  assign dataGroup_hi_hi_2695 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2696;
  assign dataGroup_hi_hi_2696 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2697;
  assign dataGroup_hi_hi_2697 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2698;
  assign dataGroup_hi_hi_2698 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2699;
  assign dataGroup_hi_hi_2699 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2700;
  assign dataGroup_hi_hi_2700 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2701;
  assign dataGroup_hi_hi_2701 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2702;
  assign dataGroup_hi_hi_2702 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2703;
  assign dataGroup_hi_hi_2703 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2704;
  assign dataGroup_hi_hi_2704 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2705;
  assign dataGroup_hi_hi_2705 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2706;
  assign dataGroup_hi_hi_2706 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2707;
  assign dataGroup_hi_hi_2707 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2708;
  assign dataGroup_hi_hi_2708 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2709;
  assign dataGroup_hi_hi_2709 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2710;
  assign dataGroup_hi_hi_2710 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2711;
  assign dataGroup_hi_hi_2711 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2712;
  assign dataGroup_hi_hi_2712 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2713;
  assign dataGroup_hi_hi_2713 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2714;
  assign dataGroup_hi_hi_2714 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2715;
  assign dataGroup_hi_hi_2715 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2716;
  assign dataGroup_hi_hi_2716 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2717;
  assign dataGroup_hi_hi_2717 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2718;
  assign dataGroup_hi_hi_2718 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2719;
  assign dataGroup_hi_hi_2719 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2720;
  assign dataGroup_hi_hi_2720 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2721;
  assign dataGroup_hi_hi_2721 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2722;
  assign dataGroup_hi_hi_2722 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2723;
  assign dataGroup_hi_hi_2723 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2724;
  assign dataGroup_hi_hi_2724 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2725;
  assign dataGroup_hi_hi_2725 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2726;
  assign dataGroup_hi_hi_2726 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2727;
  assign dataGroup_hi_hi_2727 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2728;
  assign dataGroup_hi_hi_2728 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2729;
  assign dataGroup_hi_hi_2729 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2730;
  assign dataGroup_hi_hi_2730 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2731;
  assign dataGroup_hi_hi_2731 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2732;
  assign dataGroup_hi_hi_2732 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2733;
  assign dataGroup_hi_hi_2733 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2734;
  assign dataGroup_hi_hi_2734 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2735;
  assign dataGroup_hi_hi_2735 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2736;
  assign dataGroup_hi_hi_2736 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2737;
  assign dataGroup_hi_hi_2737 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2738;
  assign dataGroup_hi_hi_2738 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2739;
  assign dataGroup_hi_hi_2739 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2740;
  assign dataGroup_hi_hi_2740 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2741;
  assign dataGroup_hi_hi_2741 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2742;
  assign dataGroup_hi_hi_2742 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2743;
  assign dataGroup_hi_hi_2743 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2744;
  assign dataGroup_hi_hi_2744 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2745;
  assign dataGroup_hi_hi_2745 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2746;
  assign dataGroup_hi_hi_2746 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2747;
  assign dataGroup_hi_hi_2747 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2748;
  assign dataGroup_hi_hi_2748 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2749;
  assign dataGroup_hi_hi_2749 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2750;
  assign dataGroup_hi_hi_2750 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2751;
  assign dataGroup_hi_hi_2751 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2752;
  assign dataGroup_hi_hi_2752 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2753;
  assign dataGroup_hi_hi_2753 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2754;
  assign dataGroup_hi_hi_2754 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2755;
  assign dataGroup_hi_hi_2755 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2756;
  assign dataGroup_hi_hi_2756 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2757;
  assign dataGroup_hi_hi_2757 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2758;
  assign dataGroup_hi_hi_2758 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2759;
  assign dataGroup_hi_hi_2759 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2760;
  assign dataGroup_hi_hi_2760 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2761;
  assign dataGroup_hi_hi_2761 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2762;
  assign dataGroup_hi_hi_2762 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2763;
  assign dataGroup_hi_hi_2763 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2764;
  assign dataGroup_hi_hi_2764 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2765;
  assign dataGroup_hi_hi_2765 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2766;
  assign dataGroup_hi_hi_2766 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2767;
  assign dataGroup_hi_hi_2767 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2768;
  assign dataGroup_hi_hi_2768 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2769;
  assign dataGroup_hi_hi_2769 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2770;
  assign dataGroup_hi_hi_2770 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2771;
  assign dataGroup_hi_hi_2771 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2772;
  assign dataGroup_hi_hi_2772 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2773;
  assign dataGroup_hi_hi_2773 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2774;
  assign dataGroup_hi_hi_2774 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2775;
  assign dataGroup_hi_hi_2775 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2776;
  assign dataGroup_hi_hi_2776 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2777;
  assign dataGroup_hi_hi_2777 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2778;
  assign dataGroup_hi_hi_2778 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2779;
  assign dataGroup_hi_hi_2779 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2780;
  assign dataGroup_hi_hi_2780 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2781;
  assign dataGroup_hi_hi_2781 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2782;
  assign dataGroup_hi_hi_2782 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2783;
  assign dataGroup_hi_hi_2783 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2784;
  assign dataGroup_hi_hi_2784 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2785;
  assign dataGroup_hi_hi_2785 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2786;
  assign dataGroup_hi_hi_2786 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2787;
  assign dataGroup_hi_hi_2787 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2788;
  assign dataGroup_hi_hi_2788 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2789;
  assign dataGroup_hi_hi_2789 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2790;
  assign dataGroup_hi_hi_2790 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2791;
  assign dataGroup_hi_hi_2791 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2792;
  assign dataGroup_hi_hi_2792 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2793;
  assign dataGroup_hi_hi_2793 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2794;
  assign dataGroup_hi_hi_2794 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2795;
  assign dataGroup_hi_hi_2795 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2796;
  assign dataGroup_hi_hi_2796 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2797;
  assign dataGroup_hi_hi_2797 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2798;
  assign dataGroup_hi_hi_2798 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2799;
  assign dataGroup_hi_hi_2799 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2800;
  assign dataGroup_hi_hi_2800 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2801;
  assign dataGroup_hi_hi_2801 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2802;
  assign dataGroup_hi_hi_2802 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2803;
  assign dataGroup_hi_hi_2803 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2804;
  assign dataGroup_hi_hi_2804 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2805;
  assign dataGroup_hi_hi_2805 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2806;
  assign dataGroup_hi_hi_2806 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2807;
  assign dataGroup_hi_hi_2807 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2808;
  assign dataGroup_hi_hi_2808 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2809;
  assign dataGroup_hi_hi_2809 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2810;
  assign dataGroup_hi_hi_2810 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2811;
  assign dataGroup_hi_hi_2811 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2812;
  assign dataGroup_hi_hi_2812 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2813;
  assign dataGroup_hi_hi_2813 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2814;
  assign dataGroup_hi_hi_2814 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2815;
  assign dataGroup_hi_hi_2815 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2816;
  assign dataGroup_hi_hi_2816 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2817;
  assign dataGroup_hi_hi_2817 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2818;
  assign dataGroup_hi_hi_2818 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2819;
  assign dataGroup_hi_hi_2819 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2820;
  assign dataGroup_hi_hi_2820 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2821;
  assign dataGroup_hi_hi_2821 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2822;
  assign dataGroup_hi_hi_2822 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2823;
  assign dataGroup_hi_hi_2823 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2824;
  assign dataGroup_hi_hi_2824 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2825;
  assign dataGroup_hi_hi_2825 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2826;
  assign dataGroup_hi_hi_2826 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2827;
  assign dataGroup_hi_hi_2827 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2828;
  assign dataGroup_hi_hi_2828 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2829;
  assign dataGroup_hi_hi_2829 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2830;
  assign dataGroup_hi_hi_2830 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2831;
  assign dataGroup_hi_hi_2831 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2832;
  assign dataGroup_hi_hi_2832 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2833;
  assign dataGroup_hi_hi_2833 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2834;
  assign dataGroup_hi_hi_2834 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2835;
  assign dataGroup_hi_hi_2835 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2836;
  assign dataGroup_hi_hi_2836 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2837;
  assign dataGroup_hi_hi_2837 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2838;
  assign dataGroup_hi_hi_2838 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2839;
  assign dataGroup_hi_hi_2839 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2840;
  assign dataGroup_hi_hi_2840 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2841;
  assign dataGroup_hi_hi_2841 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2842;
  assign dataGroup_hi_hi_2842 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2843;
  assign dataGroup_hi_hi_2843 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2844;
  assign dataGroup_hi_hi_2844 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2845;
  assign dataGroup_hi_hi_2845 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2846;
  assign dataGroup_hi_hi_2846 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2847;
  assign dataGroup_hi_hi_2847 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2848;
  assign dataGroup_hi_hi_2848 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2849;
  assign dataGroup_hi_hi_2849 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2850;
  assign dataGroup_hi_hi_2850 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2851;
  assign dataGroup_hi_hi_2851 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2852;
  assign dataGroup_hi_hi_2852 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2853;
  assign dataGroup_hi_hi_2853 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2854;
  assign dataGroup_hi_hi_2854 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2855;
  assign dataGroup_hi_hi_2855 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2856;
  assign dataGroup_hi_hi_2856 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2857;
  assign dataGroup_hi_hi_2857 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2858;
  assign dataGroup_hi_hi_2858 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2859;
  assign dataGroup_hi_hi_2859 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2860;
  assign dataGroup_hi_hi_2860 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2861;
  assign dataGroup_hi_hi_2861 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2862;
  assign dataGroup_hi_hi_2862 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2863;
  assign dataGroup_hi_hi_2863 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2864;
  assign dataGroup_hi_hi_2864 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2865;
  assign dataGroup_hi_hi_2865 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2866;
  assign dataGroup_hi_hi_2866 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2867;
  assign dataGroup_hi_hi_2867 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2868;
  assign dataGroup_hi_hi_2868 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2869;
  assign dataGroup_hi_hi_2869 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2870;
  assign dataGroup_hi_hi_2870 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2871;
  assign dataGroup_hi_hi_2871 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2872;
  assign dataGroup_hi_hi_2872 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2873;
  assign dataGroup_hi_hi_2873 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2874;
  assign dataGroup_hi_hi_2874 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2875;
  assign dataGroup_hi_hi_2875 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2876;
  assign dataGroup_hi_hi_2876 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2877;
  assign dataGroup_hi_hi_2877 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2878;
  assign dataGroup_hi_hi_2878 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2879;
  assign dataGroup_hi_hi_2879 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2880;
  assign dataGroup_hi_hi_2880 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2881;
  assign dataGroup_hi_hi_2881 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2882;
  assign dataGroup_hi_hi_2882 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2883;
  assign dataGroup_hi_hi_2883 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2884;
  assign dataGroup_hi_hi_2884 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2885;
  assign dataGroup_hi_hi_2885 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2886;
  assign dataGroup_hi_hi_2886 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2887;
  assign dataGroup_hi_hi_2887 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2888;
  assign dataGroup_hi_hi_2888 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2889;
  assign dataGroup_hi_hi_2889 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2890;
  assign dataGroup_hi_hi_2890 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2891;
  assign dataGroup_hi_hi_2891 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2892;
  assign dataGroup_hi_hi_2892 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2893;
  assign dataGroup_hi_hi_2893 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2894;
  assign dataGroup_hi_hi_2894 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2895;
  assign dataGroup_hi_hi_2895 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2896;
  assign dataGroup_hi_hi_2896 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2897;
  assign dataGroup_hi_hi_2897 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2898;
  assign dataGroup_hi_hi_2898 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2899;
  assign dataGroup_hi_hi_2899 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2900;
  assign dataGroup_hi_hi_2900 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2901;
  assign dataGroup_hi_hi_2901 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2902;
  assign dataGroup_hi_hi_2902 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2903;
  assign dataGroup_hi_hi_2903 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2904;
  assign dataGroup_hi_hi_2904 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2905;
  assign dataGroup_hi_hi_2905 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2906;
  assign dataGroup_hi_hi_2906 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2907;
  assign dataGroup_hi_hi_2907 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2908;
  assign dataGroup_hi_hi_2908 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2909;
  assign dataGroup_hi_hi_2909 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2910;
  assign dataGroup_hi_hi_2910 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2911;
  assign dataGroup_hi_hi_2911 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2912;
  assign dataGroup_hi_hi_2912 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2913;
  assign dataGroup_hi_hi_2913 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2914;
  assign dataGroup_hi_hi_2914 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2915;
  assign dataGroup_hi_hi_2915 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2916;
  assign dataGroup_hi_hi_2916 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2917;
  assign dataGroup_hi_hi_2917 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2918;
  assign dataGroup_hi_hi_2918 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2919;
  assign dataGroup_hi_hi_2919 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2920;
  assign dataGroup_hi_hi_2920 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2921;
  assign dataGroup_hi_hi_2921 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2922;
  assign dataGroup_hi_hi_2922 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2923;
  assign dataGroup_hi_hi_2923 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2924;
  assign dataGroup_hi_hi_2924 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2925;
  assign dataGroup_hi_hi_2925 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2926;
  assign dataGroup_hi_hi_2926 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2927;
  assign dataGroup_hi_hi_2927 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2928;
  assign dataGroup_hi_hi_2928 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2929;
  assign dataGroup_hi_hi_2929 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2930;
  assign dataGroup_hi_hi_2930 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2931;
  assign dataGroup_hi_hi_2931 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2932;
  assign dataGroup_hi_hi_2932 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2933;
  assign dataGroup_hi_hi_2933 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2934;
  assign dataGroup_hi_hi_2934 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2935;
  assign dataGroup_hi_hi_2935 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2936;
  assign dataGroup_hi_hi_2936 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2937;
  assign dataGroup_hi_hi_2937 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2938;
  assign dataGroup_hi_hi_2938 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2939;
  assign dataGroup_hi_hi_2939 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2940;
  assign dataGroup_hi_hi_2940 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2941;
  assign dataGroup_hi_hi_2941 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2942;
  assign dataGroup_hi_hi_2942 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2943;
  assign dataGroup_hi_hi_2943 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2944;
  assign dataGroup_hi_hi_2944 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2945;
  assign dataGroup_hi_hi_2945 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2946;
  assign dataGroup_hi_hi_2946 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2947;
  assign dataGroup_hi_hi_2947 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2948;
  assign dataGroup_hi_hi_2948 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2949;
  assign dataGroup_hi_hi_2949 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2950;
  assign dataGroup_hi_hi_2950 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2951;
  assign dataGroup_hi_hi_2951 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2952;
  assign dataGroup_hi_hi_2952 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2953;
  assign dataGroup_hi_hi_2953 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2954;
  assign dataGroup_hi_hi_2954 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2955;
  assign dataGroup_hi_hi_2955 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2956;
  assign dataGroup_hi_hi_2956 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2957;
  assign dataGroup_hi_hi_2957 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2958;
  assign dataGroup_hi_hi_2958 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2959;
  assign dataGroup_hi_hi_2959 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2960;
  assign dataGroup_hi_hi_2960 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2961;
  assign dataGroup_hi_hi_2961 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2962;
  assign dataGroup_hi_hi_2962 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2963;
  assign dataGroup_hi_hi_2963 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2964;
  assign dataGroup_hi_hi_2964 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2965;
  assign dataGroup_hi_hi_2965 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2966;
  assign dataGroup_hi_hi_2966 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2967;
  assign dataGroup_hi_hi_2967 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2968;
  assign dataGroup_hi_hi_2968 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2969;
  assign dataGroup_hi_hi_2969 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2970;
  assign dataGroup_hi_hi_2970 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2971;
  assign dataGroup_hi_hi_2971 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2972;
  assign dataGroup_hi_hi_2972 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2973;
  assign dataGroup_hi_hi_2973 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2974;
  assign dataGroup_hi_hi_2974 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2975;
  assign dataGroup_hi_hi_2975 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2976;
  assign dataGroup_hi_hi_2976 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2977;
  assign dataGroup_hi_hi_2977 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2978;
  assign dataGroup_hi_hi_2978 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2979;
  assign dataGroup_hi_hi_2979 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2980;
  assign dataGroup_hi_hi_2980 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2981;
  assign dataGroup_hi_hi_2981 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2982;
  assign dataGroup_hi_hi_2982 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2983;
  assign dataGroup_hi_hi_2983 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2984;
  assign dataGroup_hi_hi_2984 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2985;
  assign dataGroup_hi_hi_2985 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2986;
  assign dataGroup_hi_hi_2986 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2987;
  assign dataGroup_hi_hi_2987 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2988;
  assign dataGroup_hi_hi_2988 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2989;
  assign dataGroup_hi_hi_2989 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2990;
  assign dataGroup_hi_hi_2990 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2991;
  assign dataGroup_hi_hi_2991 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2992;
  assign dataGroup_hi_hi_2992 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2993;
  assign dataGroup_hi_hi_2993 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2994;
  assign dataGroup_hi_hi_2994 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2995;
  assign dataGroup_hi_hi_2995 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2996;
  assign dataGroup_hi_hi_2996 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2997;
  assign dataGroup_hi_hi_2997 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2998;
  assign dataGroup_hi_hi_2998 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_2999;
  assign dataGroup_hi_hi_2999 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3000;
  assign dataGroup_hi_hi_3000 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3001;
  assign dataGroup_hi_hi_3001 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3002;
  assign dataGroup_hi_hi_3002 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3003;
  assign dataGroup_hi_hi_3003 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3004;
  assign dataGroup_hi_hi_3004 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3005;
  assign dataGroup_hi_hi_3005 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3006;
  assign dataGroup_hi_hi_3006 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3007;
  assign dataGroup_hi_hi_3007 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3008;
  assign dataGroup_hi_hi_3008 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3009;
  assign dataGroup_hi_hi_3009 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3010;
  assign dataGroup_hi_hi_3010 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3011;
  assign dataGroup_hi_hi_3011 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3012;
  assign dataGroup_hi_hi_3012 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3013;
  assign dataGroup_hi_hi_3013 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3014;
  assign dataGroup_hi_hi_3014 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3015;
  assign dataGroup_hi_hi_3015 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3016;
  assign dataGroup_hi_hi_3016 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3017;
  assign dataGroup_hi_hi_3017 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3018;
  assign dataGroup_hi_hi_3018 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3019;
  assign dataGroup_hi_hi_3019 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3020;
  assign dataGroup_hi_hi_3020 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3021;
  assign dataGroup_hi_hi_3021 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3022;
  assign dataGroup_hi_hi_3022 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3023;
  assign dataGroup_hi_hi_3023 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3024;
  assign dataGroup_hi_hi_3024 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3025;
  assign dataGroup_hi_hi_3025 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3026;
  assign dataGroup_hi_hi_3026 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3027;
  assign dataGroup_hi_hi_3027 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3028;
  assign dataGroup_hi_hi_3028 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3029;
  assign dataGroup_hi_hi_3029 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3030;
  assign dataGroup_hi_hi_3030 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3031;
  assign dataGroup_hi_hi_3031 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3032;
  assign dataGroup_hi_hi_3032 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3033;
  assign dataGroup_hi_hi_3033 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3034;
  assign dataGroup_hi_hi_3034 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3035;
  assign dataGroup_hi_hi_3035 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3036;
  assign dataGroup_hi_hi_3036 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3037;
  assign dataGroup_hi_hi_3037 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3038;
  assign dataGroup_hi_hi_3038 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3039;
  assign dataGroup_hi_hi_3039 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3040;
  assign dataGroup_hi_hi_3040 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3041;
  assign dataGroup_hi_hi_3041 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3042;
  assign dataGroup_hi_hi_3042 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3043;
  assign dataGroup_hi_hi_3043 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3044;
  assign dataGroup_hi_hi_3044 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3045;
  assign dataGroup_hi_hi_3045 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3046;
  assign dataGroup_hi_hi_3046 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3047;
  assign dataGroup_hi_hi_3047 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3048;
  assign dataGroup_hi_hi_3048 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3049;
  assign dataGroup_hi_hi_3049 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3050;
  assign dataGroup_hi_hi_3050 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3051;
  assign dataGroup_hi_hi_3051 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3052;
  assign dataGroup_hi_hi_3052 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3053;
  assign dataGroup_hi_hi_3053 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3054;
  assign dataGroup_hi_hi_3054 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3055;
  assign dataGroup_hi_hi_3055 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3056;
  assign dataGroup_hi_hi_3056 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3057;
  assign dataGroup_hi_hi_3057 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3058;
  assign dataGroup_hi_hi_3058 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3059;
  assign dataGroup_hi_hi_3059 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3060;
  assign dataGroup_hi_hi_3060 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3061;
  assign dataGroup_hi_hi_3061 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3062;
  assign dataGroup_hi_hi_3062 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3063;
  assign dataGroup_hi_hi_3063 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3064;
  assign dataGroup_hi_hi_3064 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3065;
  assign dataGroup_hi_hi_3065 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3066;
  assign dataGroup_hi_hi_3066 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3067;
  assign dataGroup_hi_hi_3067 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3068;
  assign dataGroup_hi_hi_3068 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3069;
  assign dataGroup_hi_hi_3069 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3070;
  assign dataGroup_hi_hi_3070 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3071;
  assign dataGroup_hi_hi_3071 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3072;
  assign dataGroup_hi_hi_3072 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3073;
  assign dataGroup_hi_hi_3073 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3074;
  assign dataGroup_hi_hi_3074 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3075;
  assign dataGroup_hi_hi_3075 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3076;
  assign dataGroup_hi_hi_3076 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3077;
  assign dataGroup_hi_hi_3077 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3078;
  assign dataGroup_hi_hi_3078 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3079;
  assign dataGroup_hi_hi_3079 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3080;
  assign dataGroup_hi_hi_3080 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3081;
  assign dataGroup_hi_hi_3081 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3082;
  assign dataGroup_hi_hi_3082 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3083;
  assign dataGroup_hi_hi_3083 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3084;
  assign dataGroup_hi_hi_3084 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3085;
  assign dataGroup_hi_hi_3085 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3086;
  assign dataGroup_hi_hi_3086 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3087;
  assign dataGroup_hi_hi_3087 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3088;
  assign dataGroup_hi_hi_3088 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3089;
  assign dataGroup_hi_hi_3089 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3090;
  assign dataGroup_hi_hi_3090 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3091;
  assign dataGroup_hi_hi_3091 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3092;
  assign dataGroup_hi_hi_3092 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3093;
  assign dataGroup_hi_hi_3093 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3094;
  assign dataGroup_hi_hi_3094 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3095;
  assign dataGroup_hi_hi_3095 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3096;
  assign dataGroup_hi_hi_3096 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3097;
  assign dataGroup_hi_hi_3097 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3098;
  assign dataGroup_hi_hi_3098 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3099;
  assign dataGroup_hi_hi_3099 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3100;
  assign dataGroup_hi_hi_3100 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3101;
  assign dataGroup_hi_hi_3101 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3102;
  assign dataGroup_hi_hi_3102 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3103;
  assign dataGroup_hi_hi_3103 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3104;
  assign dataGroup_hi_hi_3104 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3105;
  assign dataGroup_hi_hi_3105 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3106;
  assign dataGroup_hi_hi_3106 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3107;
  assign dataGroup_hi_hi_3107 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3108;
  assign dataGroup_hi_hi_3108 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3109;
  assign dataGroup_hi_hi_3109 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3110;
  assign dataGroup_hi_hi_3110 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3111;
  assign dataGroup_hi_hi_3111 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3112;
  assign dataGroup_hi_hi_3112 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3113;
  assign dataGroup_hi_hi_3113 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3114;
  assign dataGroup_hi_hi_3114 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3115;
  assign dataGroup_hi_hi_3115 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3116;
  assign dataGroup_hi_hi_3116 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3117;
  assign dataGroup_hi_hi_3117 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3118;
  assign dataGroup_hi_hi_3118 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3119;
  assign dataGroup_hi_hi_3119 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3120;
  assign dataGroup_hi_hi_3120 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3121;
  assign dataGroup_hi_hi_3121 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3122;
  assign dataGroup_hi_hi_3122 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3123;
  assign dataGroup_hi_hi_3123 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3124;
  assign dataGroup_hi_hi_3124 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3125;
  assign dataGroup_hi_hi_3125 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3126;
  assign dataGroup_hi_hi_3126 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3127;
  assign dataGroup_hi_hi_3127 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3128;
  assign dataGroup_hi_hi_3128 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3129;
  assign dataGroup_hi_hi_3129 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3130;
  assign dataGroup_hi_hi_3130 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3131;
  assign dataGroup_hi_hi_3131 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3132;
  assign dataGroup_hi_hi_3132 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3133;
  assign dataGroup_hi_hi_3133 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3134;
  assign dataGroup_hi_hi_3134 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3135;
  assign dataGroup_hi_hi_3135 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3136;
  assign dataGroup_hi_hi_3136 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3137;
  assign dataGroup_hi_hi_3137 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3138;
  assign dataGroup_hi_hi_3138 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3139;
  assign dataGroup_hi_hi_3139 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3140;
  assign dataGroup_hi_hi_3140 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3141;
  assign dataGroup_hi_hi_3141 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3142;
  assign dataGroup_hi_hi_3142 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3143;
  assign dataGroup_hi_hi_3143 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3144;
  assign dataGroup_hi_hi_3144 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3145;
  assign dataGroup_hi_hi_3145 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3146;
  assign dataGroup_hi_hi_3146 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3147;
  assign dataGroup_hi_hi_3147 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3148;
  assign dataGroup_hi_hi_3148 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3149;
  assign dataGroup_hi_hi_3149 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3150;
  assign dataGroup_hi_hi_3150 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3151;
  assign dataGroup_hi_hi_3151 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3152;
  assign dataGroup_hi_hi_3152 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3153;
  assign dataGroup_hi_hi_3153 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3154;
  assign dataGroup_hi_hi_3154 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3155;
  assign dataGroup_hi_hi_3155 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3156;
  assign dataGroup_hi_hi_3156 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3157;
  assign dataGroup_hi_hi_3157 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3158;
  assign dataGroup_hi_hi_3158 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3159;
  assign dataGroup_hi_hi_3159 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3160;
  assign dataGroup_hi_hi_3160 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3161;
  assign dataGroup_hi_hi_3161 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3162;
  assign dataGroup_hi_hi_3162 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3163;
  assign dataGroup_hi_hi_3163 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3164;
  assign dataGroup_hi_hi_3164 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3165;
  assign dataGroup_hi_hi_3165 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3166;
  assign dataGroup_hi_hi_3166 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3167;
  assign dataGroup_hi_hi_3167 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3168;
  assign dataGroup_hi_hi_3168 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3169;
  assign dataGroup_hi_hi_3169 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3170;
  assign dataGroup_hi_hi_3170 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3171;
  assign dataGroup_hi_hi_3171 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3172;
  assign dataGroup_hi_hi_3172 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3173;
  assign dataGroup_hi_hi_3173 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3174;
  assign dataGroup_hi_hi_3174 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3175;
  assign dataGroup_hi_hi_3175 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3176;
  assign dataGroup_hi_hi_3176 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3177;
  assign dataGroup_hi_hi_3177 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3178;
  assign dataGroup_hi_hi_3178 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3179;
  assign dataGroup_hi_hi_3179 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3180;
  assign dataGroup_hi_hi_3180 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3181;
  assign dataGroup_hi_hi_3181 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3182;
  assign dataGroup_hi_hi_3182 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3183;
  assign dataGroup_hi_hi_3183 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3184;
  assign dataGroup_hi_hi_3184 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3185;
  assign dataGroup_hi_hi_3185 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3186;
  assign dataGroup_hi_hi_3186 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3187;
  assign dataGroup_hi_hi_3187 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3188;
  assign dataGroup_hi_hi_3188 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3189;
  assign dataGroup_hi_hi_3189 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3190;
  assign dataGroup_hi_hi_3190 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3191;
  assign dataGroup_hi_hi_3191 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3192;
  assign dataGroup_hi_hi_3192 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3193;
  assign dataGroup_hi_hi_3193 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3194;
  assign dataGroup_hi_hi_3194 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3195;
  assign dataGroup_hi_hi_3195 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3196;
  assign dataGroup_hi_hi_3196 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3197;
  assign dataGroup_hi_hi_3197 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3198;
  assign dataGroup_hi_hi_3198 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3199;
  assign dataGroup_hi_hi_3199 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3200;
  assign dataGroup_hi_hi_3200 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3201;
  assign dataGroup_hi_hi_3201 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3202;
  assign dataGroup_hi_hi_3202 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3203;
  assign dataGroup_hi_hi_3203 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3204;
  assign dataGroup_hi_hi_3204 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3205;
  assign dataGroup_hi_hi_3205 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3206;
  assign dataGroup_hi_hi_3206 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3207;
  assign dataGroup_hi_hi_3207 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3208;
  assign dataGroup_hi_hi_3208 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3209;
  assign dataGroup_hi_hi_3209 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3210;
  assign dataGroup_hi_hi_3210 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3211;
  assign dataGroup_hi_hi_3211 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3212;
  assign dataGroup_hi_hi_3212 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3213;
  assign dataGroup_hi_hi_3213 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3214;
  assign dataGroup_hi_hi_3214 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3215;
  assign dataGroup_hi_hi_3215 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3216;
  assign dataGroup_hi_hi_3216 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3217;
  assign dataGroup_hi_hi_3217 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3218;
  assign dataGroup_hi_hi_3218 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3219;
  assign dataGroup_hi_hi_3219 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3220;
  assign dataGroup_hi_hi_3220 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3221;
  assign dataGroup_hi_hi_3221 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3222;
  assign dataGroup_hi_hi_3222 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3223;
  assign dataGroup_hi_hi_3223 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3224;
  assign dataGroup_hi_hi_3224 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3225;
  assign dataGroup_hi_hi_3225 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3226;
  assign dataGroup_hi_hi_3226 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3227;
  assign dataGroup_hi_hi_3227 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3228;
  assign dataGroup_hi_hi_3228 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3229;
  assign dataGroup_hi_hi_3229 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3230;
  assign dataGroup_hi_hi_3230 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3231;
  assign dataGroup_hi_hi_3231 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3232;
  assign dataGroup_hi_hi_3232 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3233;
  assign dataGroup_hi_hi_3233 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3234;
  assign dataGroup_hi_hi_3234 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3235;
  assign dataGroup_hi_hi_3235 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3236;
  assign dataGroup_hi_hi_3236 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3237;
  assign dataGroup_hi_hi_3237 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3238;
  assign dataGroup_hi_hi_3238 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3239;
  assign dataGroup_hi_hi_3239 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3240;
  assign dataGroup_hi_hi_3240 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3241;
  assign dataGroup_hi_hi_3241 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3242;
  assign dataGroup_hi_hi_3242 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3243;
  assign dataGroup_hi_hi_3243 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3244;
  assign dataGroup_hi_hi_3244 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3245;
  assign dataGroup_hi_hi_3245 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3246;
  assign dataGroup_hi_hi_3246 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3247;
  assign dataGroup_hi_hi_3247 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3248;
  assign dataGroup_hi_hi_3248 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3249;
  assign dataGroup_hi_hi_3249 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3250;
  assign dataGroup_hi_hi_3250 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3251;
  assign dataGroup_hi_hi_3251 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3252;
  assign dataGroup_hi_hi_3252 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3253;
  assign dataGroup_hi_hi_3253 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3254;
  assign dataGroup_hi_hi_3254 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3255;
  assign dataGroup_hi_hi_3255 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3256;
  assign dataGroup_hi_hi_3256 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3257;
  assign dataGroup_hi_hi_3257 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3258;
  assign dataGroup_hi_hi_3258 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3259;
  assign dataGroup_hi_hi_3259 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3260;
  assign dataGroup_hi_hi_3260 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3261;
  assign dataGroup_hi_hi_3261 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3262;
  assign dataGroup_hi_hi_3262 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3263;
  assign dataGroup_hi_hi_3263 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3264;
  assign dataGroup_hi_hi_3264 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3265;
  assign dataGroup_hi_hi_3265 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3266;
  assign dataGroup_hi_hi_3266 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3267;
  assign dataGroup_hi_hi_3267 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3268;
  assign dataGroup_hi_hi_3268 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3269;
  assign dataGroup_hi_hi_3269 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3270;
  assign dataGroup_hi_hi_3270 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3271;
  assign dataGroup_hi_hi_3271 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3272;
  assign dataGroup_hi_hi_3272 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3273;
  assign dataGroup_hi_hi_3273 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3274;
  assign dataGroup_hi_hi_3274 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3275;
  assign dataGroup_hi_hi_3275 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3276;
  assign dataGroup_hi_hi_3276 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3277;
  assign dataGroup_hi_hi_3277 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3278;
  assign dataGroup_hi_hi_3278 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3279;
  assign dataGroup_hi_hi_3279 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3280;
  assign dataGroup_hi_hi_3280 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3281;
  assign dataGroup_hi_hi_3281 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3282;
  assign dataGroup_hi_hi_3282 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3283;
  assign dataGroup_hi_hi_3283 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3284;
  assign dataGroup_hi_hi_3284 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3285;
  assign dataGroup_hi_hi_3285 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3286;
  assign dataGroup_hi_hi_3286 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3287;
  assign dataGroup_hi_hi_3287 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3288;
  assign dataGroup_hi_hi_3288 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3289;
  assign dataGroup_hi_hi_3289 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3290;
  assign dataGroup_hi_hi_3290 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3291;
  assign dataGroup_hi_hi_3291 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3292;
  assign dataGroup_hi_hi_3292 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3293;
  assign dataGroup_hi_hi_3293 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3294;
  assign dataGroup_hi_hi_3294 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3295;
  assign dataGroup_hi_hi_3295 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3296;
  assign dataGroup_hi_hi_3296 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3297;
  assign dataGroup_hi_hi_3297 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3298;
  assign dataGroup_hi_hi_3298 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3299;
  assign dataGroup_hi_hi_3299 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3300;
  assign dataGroup_hi_hi_3300 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3301;
  assign dataGroup_hi_hi_3301 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3302;
  assign dataGroup_hi_hi_3302 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3303;
  assign dataGroup_hi_hi_3303 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3304;
  assign dataGroup_hi_hi_3304 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3305;
  assign dataGroup_hi_hi_3305 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3306;
  assign dataGroup_hi_hi_3306 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3307;
  assign dataGroup_hi_hi_3307 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3308;
  assign dataGroup_hi_hi_3308 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3309;
  assign dataGroup_hi_hi_3309 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3310;
  assign dataGroup_hi_hi_3310 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3311;
  assign dataGroup_hi_hi_3311 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3312;
  assign dataGroup_hi_hi_3312 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3313;
  assign dataGroup_hi_hi_3313 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3314;
  assign dataGroup_hi_hi_3314 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3315;
  assign dataGroup_hi_hi_3315 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3316;
  assign dataGroup_hi_hi_3316 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3317;
  assign dataGroup_hi_hi_3317 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3318;
  assign dataGroup_hi_hi_3318 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3319;
  assign dataGroup_hi_hi_3319 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3320;
  assign dataGroup_hi_hi_3320 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3321;
  assign dataGroup_hi_hi_3321 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3322;
  assign dataGroup_hi_hi_3322 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3323;
  assign dataGroup_hi_hi_3323 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3324;
  assign dataGroup_hi_hi_3324 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3325;
  assign dataGroup_hi_hi_3325 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3326;
  assign dataGroup_hi_hi_3326 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3327;
  assign dataGroup_hi_hi_3327 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3328;
  assign dataGroup_hi_hi_3328 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3329;
  assign dataGroup_hi_hi_3329 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3330;
  assign dataGroup_hi_hi_3330 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3331;
  assign dataGroup_hi_hi_3331 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3332;
  assign dataGroup_hi_hi_3332 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3333;
  assign dataGroup_hi_hi_3333 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3334;
  assign dataGroup_hi_hi_3334 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3335;
  assign dataGroup_hi_hi_3335 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3336;
  assign dataGroup_hi_hi_3336 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3337;
  assign dataGroup_hi_hi_3337 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3338;
  assign dataGroup_hi_hi_3338 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3339;
  assign dataGroup_hi_hi_3339 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3340;
  assign dataGroup_hi_hi_3340 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3341;
  assign dataGroup_hi_hi_3341 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3342;
  assign dataGroup_hi_hi_3342 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3343;
  assign dataGroup_hi_hi_3343 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3344;
  assign dataGroup_hi_hi_3344 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3345;
  assign dataGroup_hi_hi_3345 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3346;
  assign dataGroup_hi_hi_3346 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3347;
  assign dataGroup_hi_hi_3347 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3348;
  assign dataGroup_hi_hi_3348 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3349;
  assign dataGroup_hi_hi_3349 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3350;
  assign dataGroup_hi_hi_3350 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3351;
  assign dataGroup_hi_hi_3351 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3352;
  assign dataGroup_hi_hi_3352 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3353;
  assign dataGroup_hi_hi_3353 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3354;
  assign dataGroup_hi_hi_3354 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3355;
  assign dataGroup_hi_hi_3355 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3356;
  assign dataGroup_hi_hi_3356 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3357;
  assign dataGroup_hi_hi_3357 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3358;
  assign dataGroup_hi_hi_3358 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3359;
  assign dataGroup_hi_hi_3359 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3360;
  assign dataGroup_hi_hi_3360 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3361;
  assign dataGroup_hi_hi_3361 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3362;
  assign dataGroup_hi_hi_3362 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3363;
  assign dataGroup_hi_hi_3363 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3364;
  assign dataGroup_hi_hi_3364 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3365;
  assign dataGroup_hi_hi_3365 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3366;
  assign dataGroup_hi_hi_3366 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3367;
  assign dataGroup_hi_hi_3367 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3368;
  assign dataGroup_hi_hi_3368 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3369;
  assign dataGroup_hi_hi_3369 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3370;
  assign dataGroup_hi_hi_3370 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3371;
  assign dataGroup_hi_hi_3371 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3372;
  assign dataGroup_hi_hi_3372 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3373;
  assign dataGroup_hi_hi_3373 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3374;
  assign dataGroup_hi_hi_3374 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3375;
  assign dataGroup_hi_hi_3375 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3376;
  assign dataGroup_hi_hi_3376 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3377;
  assign dataGroup_hi_hi_3377 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3378;
  assign dataGroup_hi_hi_3378 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3379;
  assign dataGroup_hi_hi_3379 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3380;
  assign dataGroup_hi_hi_3380 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3381;
  assign dataGroup_hi_hi_3381 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3382;
  assign dataGroup_hi_hi_3382 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3383;
  assign dataGroup_hi_hi_3383 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3384;
  assign dataGroup_hi_hi_3384 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3385;
  assign dataGroup_hi_hi_3385 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3386;
  assign dataGroup_hi_hi_3386 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3387;
  assign dataGroup_hi_hi_3387 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3388;
  assign dataGroup_hi_hi_3388 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3389;
  assign dataGroup_hi_hi_3389 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3390;
  assign dataGroup_hi_hi_3390 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3391;
  assign dataGroup_hi_hi_3391 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3392;
  assign dataGroup_hi_hi_3392 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3393;
  assign dataGroup_hi_hi_3393 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3394;
  assign dataGroup_hi_hi_3394 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3395;
  assign dataGroup_hi_hi_3395 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3396;
  assign dataGroup_hi_hi_3396 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3397;
  assign dataGroup_hi_hi_3397 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3398;
  assign dataGroup_hi_hi_3398 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3399;
  assign dataGroup_hi_hi_3399 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3400;
  assign dataGroup_hi_hi_3400 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3401;
  assign dataGroup_hi_hi_3401 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3402;
  assign dataGroup_hi_hi_3402 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3403;
  assign dataGroup_hi_hi_3403 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3404;
  assign dataGroup_hi_hi_3404 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3405;
  assign dataGroup_hi_hi_3405 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3406;
  assign dataGroup_hi_hi_3406 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3407;
  assign dataGroup_hi_hi_3407 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3408;
  assign dataGroup_hi_hi_3408 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3409;
  assign dataGroup_hi_hi_3409 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3410;
  assign dataGroup_hi_hi_3410 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3411;
  assign dataGroup_hi_hi_3411 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3412;
  assign dataGroup_hi_hi_3412 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3413;
  assign dataGroup_hi_hi_3413 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3414;
  assign dataGroup_hi_hi_3414 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3415;
  assign dataGroup_hi_hi_3415 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3416;
  assign dataGroup_hi_hi_3416 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3417;
  assign dataGroup_hi_hi_3417 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3418;
  assign dataGroup_hi_hi_3418 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3419;
  assign dataGroup_hi_hi_3419 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3420;
  assign dataGroup_hi_hi_3420 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3421;
  assign dataGroup_hi_hi_3421 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3422;
  assign dataGroup_hi_hi_3422 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3423;
  assign dataGroup_hi_hi_3423 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3424;
  assign dataGroup_hi_hi_3424 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3425;
  assign dataGroup_hi_hi_3425 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3426;
  assign dataGroup_hi_hi_3426 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3427;
  assign dataGroup_hi_hi_3427 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3428;
  assign dataGroup_hi_hi_3428 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3429;
  assign dataGroup_hi_hi_3429 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3430;
  assign dataGroup_hi_hi_3430 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3431;
  assign dataGroup_hi_hi_3431 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3432;
  assign dataGroup_hi_hi_3432 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3433;
  assign dataGroup_hi_hi_3433 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3434;
  assign dataGroup_hi_hi_3434 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3435;
  assign dataGroup_hi_hi_3435 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3436;
  assign dataGroup_hi_hi_3436 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3437;
  assign dataGroup_hi_hi_3437 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3438;
  assign dataGroup_hi_hi_3438 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3439;
  assign dataGroup_hi_hi_3439 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3440;
  assign dataGroup_hi_hi_3440 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3441;
  assign dataGroup_hi_hi_3441 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3442;
  assign dataGroup_hi_hi_3442 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3443;
  assign dataGroup_hi_hi_3443 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3444;
  assign dataGroup_hi_hi_3444 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3445;
  assign dataGroup_hi_hi_3445 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3446;
  assign dataGroup_hi_hi_3446 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3447;
  assign dataGroup_hi_hi_3447 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3448;
  assign dataGroup_hi_hi_3448 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3449;
  assign dataGroup_hi_hi_3449 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3450;
  assign dataGroup_hi_hi_3450 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3451;
  assign dataGroup_hi_hi_3451 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3452;
  assign dataGroup_hi_hi_3452 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3453;
  assign dataGroup_hi_hi_3453 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3454;
  assign dataGroup_hi_hi_3454 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3455;
  assign dataGroup_hi_hi_3455 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3456;
  assign dataGroup_hi_hi_3456 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3457;
  assign dataGroup_hi_hi_3457 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3458;
  assign dataGroup_hi_hi_3458 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3459;
  assign dataGroup_hi_hi_3459 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3460;
  assign dataGroup_hi_hi_3460 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3461;
  assign dataGroup_hi_hi_3461 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3462;
  assign dataGroup_hi_hi_3462 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3463;
  assign dataGroup_hi_hi_3463 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3464;
  assign dataGroup_hi_hi_3464 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3465;
  assign dataGroup_hi_hi_3465 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3466;
  assign dataGroup_hi_hi_3466 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3467;
  assign dataGroup_hi_hi_3467 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3468;
  assign dataGroup_hi_hi_3468 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3469;
  assign dataGroup_hi_hi_3469 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3470;
  assign dataGroup_hi_hi_3470 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3471;
  assign dataGroup_hi_hi_3471 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3472;
  assign dataGroup_hi_hi_3472 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3473;
  assign dataGroup_hi_hi_3473 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3474;
  assign dataGroup_hi_hi_3474 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3475;
  assign dataGroup_hi_hi_3475 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3476;
  assign dataGroup_hi_hi_3476 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3477;
  assign dataGroup_hi_hi_3477 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3478;
  assign dataGroup_hi_hi_3478 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3479;
  assign dataGroup_hi_hi_3479 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3480;
  assign dataGroup_hi_hi_3480 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3481;
  assign dataGroup_hi_hi_3481 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3482;
  assign dataGroup_hi_hi_3482 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3483;
  assign dataGroup_hi_hi_3483 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3484;
  assign dataGroup_hi_hi_3484 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3485;
  assign dataGroup_hi_hi_3485 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3486;
  assign dataGroup_hi_hi_3486 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3487;
  assign dataGroup_hi_hi_3487 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3488;
  assign dataGroup_hi_hi_3488 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3489;
  assign dataGroup_hi_hi_3489 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3490;
  assign dataGroup_hi_hi_3490 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3491;
  assign dataGroup_hi_hi_3491 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3492;
  assign dataGroup_hi_hi_3492 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3493;
  assign dataGroup_hi_hi_3493 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3494;
  assign dataGroup_hi_hi_3494 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3495;
  assign dataGroup_hi_hi_3495 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3496;
  assign dataGroup_hi_hi_3496 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3497;
  assign dataGroup_hi_hi_3497 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3498;
  assign dataGroup_hi_hi_3498 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3499;
  assign dataGroup_hi_hi_3499 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3500;
  assign dataGroup_hi_hi_3500 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3501;
  assign dataGroup_hi_hi_3501 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3502;
  assign dataGroup_hi_hi_3502 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3503;
  assign dataGroup_hi_hi_3503 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3504;
  assign dataGroup_hi_hi_3504 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3505;
  assign dataGroup_hi_hi_3505 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3506;
  assign dataGroup_hi_hi_3506 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3507;
  assign dataGroup_hi_hi_3507 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3508;
  assign dataGroup_hi_hi_3508 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3509;
  assign dataGroup_hi_hi_3509 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3510;
  assign dataGroup_hi_hi_3510 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3511;
  assign dataGroup_hi_hi_3511 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3512;
  assign dataGroup_hi_hi_3512 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3513;
  assign dataGroup_hi_hi_3513 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3514;
  assign dataGroup_hi_hi_3514 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3515;
  assign dataGroup_hi_hi_3515 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3516;
  assign dataGroup_hi_hi_3516 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3517;
  assign dataGroup_hi_hi_3517 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3518;
  assign dataGroup_hi_hi_3518 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3519;
  assign dataGroup_hi_hi_3519 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3520;
  assign dataGroup_hi_hi_3520 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3521;
  assign dataGroup_hi_hi_3521 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3522;
  assign dataGroup_hi_hi_3522 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3523;
  assign dataGroup_hi_hi_3523 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3524;
  assign dataGroup_hi_hi_3524 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3525;
  assign dataGroup_hi_hi_3525 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3526;
  assign dataGroup_hi_hi_3526 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3527;
  assign dataGroup_hi_hi_3527 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3528;
  assign dataGroup_hi_hi_3528 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3529;
  assign dataGroup_hi_hi_3529 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3530;
  assign dataGroup_hi_hi_3530 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3531;
  assign dataGroup_hi_hi_3531 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3532;
  assign dataGroup_hi_hi_3532 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3533;
  assign dataGroup_hi_hi_3533 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3534;
  assign dataGroup_hi_hi_3534 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3535;
  assign dataGroup_hi_hi_3535 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3536;
  assign dataGroup_hi_hi_3536 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3537;
  assign dataGroup_hi_hi_3537 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3538;
  assign dataGroup_hi_hi_3538 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3539;
  assign dataGroup_hi_hi_3539 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3540;
  assign dataGroup_hi_hi_3540 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3541;
  assign dataGroup_hi_hi_3541 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3542;
  assign dataGroup_hi_hi_3542 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3543;
  assign dataGroup_hi_hi_3543 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3544;
  assign dataGroup_hi_hi_3544 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3545;
  assign dataGroup_hi_hi_3545 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3546;
  assign dataGroup_hi_hi_3546 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3547;
  assign dataGroup_hi_hi_3547 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3548;
  assign dataGroup_hi_hi_3548 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3549;
  assign dataGroup_hi_hi_3549 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3550;
  assign dataGroup_hi_hi_3550 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3551;
  assign dataGroup_hi_hi_3551 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3552;
  assign dataGroup_hi_hi_3552 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3553;
  assign dataGroup_hi_hi_3553 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3554;
  assign dataGroup_hi_hi_3554 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3555;
  assign dataGroup_hi_hi_3555 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3556;
  assign dataGroup_hi_hi_3556 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3557;
  assign dataGroup_hi_hi_3557 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3558;
  assign dataGroup_hi_hi_3558 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3559;
  assign dataGroup_hi_hi_3559 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3560;
  assign dataGroup_hi_hi_3560 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3561;
  assign dataGroup_hi_hi_3561 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3562;
  assign dataGroup_hi_hi_3562 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3563;
  assign dataGroup_hi_hi_3563 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3564;
  assign dataGroup_hi_hi_3564 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3565;
  assign dataGroup_hi_hi_3565 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3566;
  assign dataGroup_hi_hi_3566 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3567;
  assign dataGroup_hi_hi_3567 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3568;
  assign dataGroup_hi_hi_3568 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3569;
  assign dataGroup_hi_hi_3569 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3570;
  assign dataGroup_hi_hi_3570 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3571;
  assign dataGroup_hi_hi_3571 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3572;
  assign dataGroup_hi_hi_3572 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3573;
  assign dataGroup_hi_hi_3573 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3574;
  assign dataGroup_hi_hi_3574 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3575;
  assign dataGroup_hi_hi_3575 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3576;
  assign dataGroup_hi_hi_3576 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3577;
  assign dataGroup_hi_hi_3577 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3578;
  assign dataGroup_hi_hi_3578 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3579;
  assign dataGroup_hi_hi_3579 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3580;
  assign dataGroup_hi_hi_3580 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3581;
  assign dataGroup_hi_hi_3581 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3582;
  assign dataGroup_hi_hi_3582 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3583;
  assign dataGroup_hi_hi_3583 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3584;
  assign dataGroup_hi_hi_3584 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3585;
  assign dataGroup_hi_hi_3585 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3586;
  assign dataGroup_hi_hi_3586 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3587;
  assign dataGroup_hi_hi_3587 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3588;
  assign dataGroup_hi_hi_3588 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3589;
  assign dataGroup_hi_hi_3589 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3590;
  assign dataGroup_hi_hi_3590 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3591;
  assign dataGroup_hi_hi_3591 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3592;
  assign dataGroup_hi_hi_3592 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3593;
  assign dataGroup_hi_hi_3593 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3594;
  assign dataGroup_hi_hi_3594 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3595;
  assign dataGroup_hi_hi_3595 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3596;
  assign dataGroup_hi_hi_3596 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3597;
  assign dataGroup_hi_hi_3597 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3598;
  assign dataGroup_hi_hi_3598 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3599;
  assign dataGroup_hi_hi_3599 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3600;
  assign dataGroup_hi_hi_3600 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3601;
  assign dataGroup_hi_hi_3601 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3602;
  assign dataGroup_hi_hi_3602 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3603;
  assign dataGroup_hi_hi_3603 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3604;
  assign dataGroup_hi_hi_3604 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3605;
  assign dataGroup_hi_hi_3605 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3606;
  assign dataGroup_hi_hi_3606 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3607;
  assign dataGroup_hi_hi_3607 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3608;
  assign dataGroup_hi_hi_3608 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3609;
  assign dataGroup_hi_hi_3609 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3610;
  assign dataGroup_hi_hi_3610 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3611;
  assign dataGroup_hi_hi_3611 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3612;
  assign dataGroup_hi_hi_3612 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3613;
  assign dataGroup_hi_hi_3613 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3614;
  assign dataGroup_hi_hi_3614 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3615;
  assign dataGroup_hi_hi_3615 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3616;
  assign dataGroup_hi_hi_3616 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3617;
  assign dataGroup_hi_hi_3617 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3618;
  assign dataGroup_hi_hi_3618 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3619;
  assign dataGroup_hi_hi_3619 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3620;
  assign dataGroup_hi_hi_3620 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3621;
  assign dataGroup_hi_hi_3621 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3622;
  assign dataGroup_hi_hi_3622 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3623;
  assign dataGroup_hi_hi_3623 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3624;
  assign dataGroup_hi_hi_3624 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3625;
  assign dataGroup_hi_hi_3625 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3626;
  assign dataGroup_hi_hi_3626 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3627;
  assign dataGroup_hi_hi_3627 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3628;
  assign dataGroup_hi_hi_3628 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3629;
  assign dataGroup_hi_hi_3629 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3630;
  assign dataGroup_hi_hi_3630 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3631;
  assign dataGroup_hi_hi_3631 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3632;
  assign dataGroup_hi_hi_3632 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3633;
  assign dataGroup_hi_hi_3633 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3634;
  assign dataGroup_hi_hi_3634 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3635;
  assign dataGroup_hi_hi_3635 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3636;
  assign dataGroup_hi_hi_3636 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3637;
  assign dataGroup_hi_hi_3637 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3638;
  assign dataGroup_hi_hi_3638 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3639;
  assign dataGroup_hi_hi_3639 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3640;
  assign dataGroup_hi_hi_3640 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3641;
  assign dataGroup_hi_hi_3641 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3642;
  assign dataGroup_hi_hi_3642 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3643;
  assign dataGroup_hi_hi_3643 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3644;
  assign dataGroup_hi_hi_3644 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3645;
  assign dataGroup_hi_hi_3645 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3646;
  assign dataGroup_hi_hi_3646 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3647;
  assign dataGroup_hi_hi_3647 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3648;
  assign dataGroup_hi_hi_3648 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3649;
  assign dataGroup_hi_hi_3649 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3650;
  assign dataGroup_hi_hi_3650 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3651;
  assign dataGroup_hi_hi_3651 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3652;
  assign dataGroup_hi_hi_3652 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3653;
  assign dataGroup_hi_hi_3653 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3654;
  assign dataGroup_hi_hi_3654 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3655;
  assign dataGroup_hi_hi_3655 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3656;
  assign dataGroup_hi_hi_3656 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3657;
  assign dataGroup_hi_hi_3657 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3658;
  assign dataGroup_hi_hi_3658 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3659;
  assign dataGroup_hi_hi_3659 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3660;
  assign dataGroup_hi_hi_3660 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3661;
  assign dataGroup_hi_hi_3661 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3662;
  assign dataGroup_hi_hi_3662 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3663;
  assign dataGroup_hi_hi_3663 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3664;
  assign dataGroup_hi_hi_3664 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3665;
  assign dataGroup_hi_hi_3665 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3666;
  assign dataGroup_hi_hi_3666 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3667;
  assign dataGroup_hi_hi_3667 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3668;
  assign dataGroup_hi_hi_3668 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3669;
  assign dataGroup_hi_hi_3669 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3670;
  assign dataGroup_hi_hi_3670 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3671;
  assign dataGroup_hi_hi_3671 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3672;
  assign dataGroup_hi_hi_3672 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3673;
  assign dataGroup_hi_hi_3673 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3674;
  assign dataGroup_hi_hi_3674 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3675;
  assign dataGroup_hi_hi_3675 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3676;
  assign dataGroup_hi_hi_3676 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3677;
  assign dataGroup_hi_hi_3677 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3678;
  assign dataGroup_hi_hi_3678 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3679;
  assign dataGroup_hi_hi_3679 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3680;
  assign dataGroup_hi_hi_3680 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3681;
  assign dataGroup_hi_hi_3681 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3682;
  assign dataGroup_hi_hi_3682 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3683;
  assign dataGroup_hi_hi_3683 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3684;
  assign dataGroup_hi_hi_3684 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3685;
  assign dataGroup_hi_hi_3685 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3686;
  assign dataGroup_hi_hi_3686 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3687;
  assign dataGroup_hi_hi_3687 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3688;
  assign dataGroup_hi_hi_3688 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3689;
  assign dataGroup_hi_hi_3689 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3690;
  assign dataGroup_hi_hi_3690 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3691;
  assign dataGroup_hi_hi_3691 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3692;
  assign dataGroup_hi_hi_3692 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3693;
  assign dataGroup_hi_hi_3693 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3694;
  assign dataGroup_hi_hi_3694 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3695;
  assign dataGroup_hi_hi_3695 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3696;
  assign dataGroup_hi_hi_3696 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3697;
  assign dataGroup_hi_hi_3697 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3698;
  assign dataGroup_hi_hi_3698 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3699;
  assign dataGroup_hi_hi_3699 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3700;
  assign dataGroup_hi_hi_3700 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3701;
  assign dataGroup_hi_hi_3701 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3702;
  assign dataGroup_hi_hi_3702 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3703;
  assign dataGroup_hi_hi_3703 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3704;
  assign dataGroup_hi_hi_3704 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3705;
  assign dataGroup_hi_hi_3705 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3706;
  assign dataGroup_hi_hi_3706 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3707;
  assign dataGroup_hi_hi_3707 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3708;
  assign dataGroup_hi_hi_3708 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3709;
  assign dataGroup_hi_hi_3709 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3710;
  assign dataGroup_hi_hi_3710 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3711;
  assign dataGroup_hi_hi_3711 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3712;
  assign dataGroup_hi_hi_3712 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3713;
  assign dataGroup_hi_hi_3713 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3714;
  assign dataGroup_hi_hi_3714 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3715;
  assign dataGroup_hi_hi_3715 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3716;
  assign dataGroup_hi_hi_3716 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3717;
  assign dataGroup_hi_hi_3717 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3718;
  assign dataGroup_hi_hi_3718 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3719;
  assign dataGroup_hi_hi_3719 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3720;
  assign dataGroup_hi_hi_3720 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3721;
  assign dataGroup_hi_hi_3721 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3722;
  assign dataGroup_hi_hi_3722 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3723;
  assign dataGroup_hi_hi_3723 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3724;
  assign dataGroup_hi_hi_3724 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3725;
  assign dataGroup_hi_hi_3725 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3726;
  assign dataGroup_hi_hi_3726 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3727;
  assign dataGroup_hi_hi_3727 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3728;
  assign dataGroup_hi_hi_3728 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3729;
  assign dataGroup_hi_hi_3729 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3730;
  assign dataGroup_hi_hi_3730 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3731;
  assign dataGroup_hi_hi_3731 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3732;
  assign dataGroup_hi_hi_3732 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3733;
  assign dataGroup_hi_hi_3733 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3734;
  assign dataGroup_hi_hi_3734 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3735;
  assign dataGroup_hi_hi_3735 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3736;
  assign dataGroup_hi_hi_3736 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3737;
  assign dataGroup_hi_hi_3737 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3738;
  assign dataGroup_hi_hi_3738 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3739;
  assign dataGroup_hi_hi_3739 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3740;
  assign dataGroup_hi_hi_3740 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3741;
  assign dataGroup_hi_hi_3741 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3742;
  assign dataGroup_hi_hi_3742 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3743;
  assign dataGroup_hi_hi_3743 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3744;
  assign dataGroup_hi_hi_3744 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3745;
  assign dataGroup_hi_hi_3745 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3746;
  assign dataGroup_hi_hi_3746 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3747;
  assign dataGroup_hi_hi_3747 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3748;
  assign dataGroup_hi_hi_3748 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3749;
  assign dataGroup_hi_hi_3749 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3750;
  assign dataGroup_hi_hi_3750 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3751;
  assign dataGroup_hi_hi_3751 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3752;
  assign dataGroup_hi_hi_3752 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3753;
  assign dataGroup_hi_hi_3753 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3754;
  assign dataGroup_hi_hi_3754 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3755;
  assign dataGroup_hi_hi_3755 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3756;
  assign dataGroup_hi_hi_3756 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3757;
  assign dataGroup_hi_hi_3757 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3758;
  assign dataGroup_hi_hi_3758 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3759;
  assign dataGroup_hi_hi_3759 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3760;
  assign dataGroup_hi_hi_3760 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3761;
  assign dataGroup_hi_hi_3761 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3762;
  assign dataGroup_hi_hi_3762 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3763;
  assign dataGroup_hi_hi_3763 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3764;
  assign dataGroup_hi_hi_3764 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3765;
  assign dataGroup_hi_hi_3765 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3766;
  assign dataGroup_hi_hi_3766 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3767;
  assign dataGroup_hi_hi_3767 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3768;
  assign dataGroup_hi_hi_3768 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3769;
  assign dataGroup_hi_hi_3769 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3770;
  assign dataGroup_hi_hi_3770 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3771;
  assign dataGroup_hi_hi_3771 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3772;
  assign dataGroup_hi_hi_3772 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3773;
  assign dataGroup_hi_hi_3773 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3774;
  assign dataGroup_hi_hi_3774 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3775;
  assign dataGroup_hi_hi_3775 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3776;
  assign dataGroup_hi_hi_3776 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3777;
  assign dataGroup_hi_hi_3777 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3778;
  assign dataGroup_hi_hi_3778 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3779;
  assign dataGroup_hi_hi_3779 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3780;
  assign dataGroup_hi_hi_3780 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3781;
  assign dataGroup_hi_hi_3781 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3782;
  assign dataGroup_hi_hi_3782 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3783;
  assign dataGroup_hi_hi_3783 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3784;
  assign dataGroup_hi_hi_3784 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3785;
  assign dataGroup_hi_hi_3785 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3786;
  assign dataGroup_hi_hi_3786 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3787;
  assign dataGroup_hi_hi_3787 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3788;
  assign dataGroup_hi_hi_3788 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3789;
  assign dataGroup_hi_hi_3789 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3790;
  assign dataGroup_hi_hi_3790 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3791;
  assign dataGroup_hi_hi_3791 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3792;
  assign dataGroup_hi_hi_3792 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3793;
  assign dataGroup_hi_hi_3793 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3794;
  assign dataGroup_hi_hi_3794 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3795;
  assign dataGroup_hi_hi_3795 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3796;
  assign dataGroup_hi_hi_3796 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3797;
  assign dataGroup_hi_hi_3797 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3798;
  assign dataGroup_hi_hi_3798 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3799;
  assign dataGroup_hi_hi_3799 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3800;
  assign dataGroup_hi_hi_3800 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3801;
  assign dataGroup_hi_hi_3801 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3802;
  assign dataGroup_hi_hi_3802 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3803;
  assign dataGroup_hi_hi_3803 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3804;
  assign dataGroup_hi_hi_3804 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3805;
  assign dataGroup_hi_hi_3805 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3806;
  assign dataGroup_hi_hi_3806 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3807;
  assign dataGroup_hi_hi_3807 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3808;
  assign dataGroup_hi_hi_3808 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3809;
  assign dataGroup_hi_hi_3809 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3810;
  assign dataGroup_hi_hi_3810 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3811;
  assign dataGroup_hi_hi_3811 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3812;
  assign dataGroup_hi_hi_3812 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3813;
  assign dataGroup_hi_hi_3813 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3814;
  assign dataGroup_hi_hi_3814 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3815;
  assign dataGroup_hi_hi_3815 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3816;
  assign dataGroup_hi_hi_3816 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3817;
  assign dataGroup_hi_hi_3817 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3818;
  assign dataGroup_hi_hi_3818 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3819;
  assign dataGroup_hi_hi_3819 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3820;
  assign dataGroup_hi_hi_3820 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3821;
  assign dataGroup_hi_hi_3821 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3822;
  assign dataGroup_hi_hi_3822 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3823;
  assign dataGroup_hi_hi_3823 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3824;
  assign dataGroup_hi_hi_3824 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3825;
  assign dataGroup_hi_hi_3825 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3826;
  assign dataGroup_hi_hi_3826 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3827;
  assign dataGroup_hi_hi_3827 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3828;
  assign dataGroup_hi_hi_3828 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3829;
  assign dataGroup_hi_hi_3829 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3830;
  assign dataGroup_hi_hi_3830 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3831;
  assign dataGroup_hi_hi_3831 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3832;
  assign dataGroup_hi_hi_3832 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3833;
  assign dataGroup_hi_hi_3833 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3834;
  assign dataGroup_hi_hi_3834 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3835;
  assign dataGroup_hi_hi_3835 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3836;
  assign dataGroup_hi_hi_3836 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3837;
  assign dataGroup_hi_hi_3837 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3838;
  assign dataGroup_hi_hi_3838 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3839;
  assign dataGroup_hi_hi_3839 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3840;
  assign dataGroup_hi_hi_3840 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3841;
  assign dataGroup_hi_hi_3841 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3842;
  assign dataGroup_hi_hi_3842 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3843;
  assign dataGroup_hi_hi_3843 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3844;
  assign dataGroup_hi_hi_3844 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3845;
  assign dataGroup_hi_hi_3845 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3846;
  assign dataGroup_hi_hi_3846 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3847;
  assign dataGroup_hi_hi_3847 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3848;
  assign dataGroup_hi_hi_3848 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3849;
  assign dataGroup_hi_hi_3849 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3850;
  assign dataGroup_hi_hi_3850 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3851;
  assign dataGroup_hi_hi_3851 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3852;
  assign dataGroup_hi_hi_3852 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3853;
  assign dataGroup_hi_hi_3853 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3854;
  assign dataGroup_hi_hi_3854 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3855;
  assign dataGroup_hi_hi_3855 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3856;
  assign dataGroup_hi_hi_3856 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3857;
  assign dataGroup_hi_hi_3857 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3858;
  assign dataGroup_hi_hi_3858 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3859;
  assign dataGroup_hi_hi_3859 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3860;
  assign dataGroup_hi_hi_3860 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3861;
  assign dataGroup_hi_hi_3861 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3862;
  assign dataGroup_hi_hi_3862 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3863;
  assign dataGroup_hi_hi_3863 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3864;
  assign dataGroup_hi_hi_3864 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3865;
  assign dataGroup_hi_hi_3865 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3866;
  assign dataGroup_hi_hi_3866 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3867;
  assign dataGroup_hi_hi_3867 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3868;
  assign dataGroup_hi_hi_3868 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3869;
  assign dataGroup_hi_hi_3869 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3870;
  assign dataGroup_hi_hi_3870 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3871;
  assign dataGroup_hi_hi_3871 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3872;
  assign dataGroup_hi_hi_3872 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3873;
  assign dataGroup_hi_hi_3873 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3874;
  assign dataGroup_hi_hi_3874 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3875;
  assign dataGroup_hi_hi_3875 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3876;
  assign dataGroup_hi_hi_3876 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3877;
  assign dataGroup_hi_hi_3877 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3878;
  assign dataGroup_hi_hi_3878 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3879;
  assign dataGroup_hi_hi_3879 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3880;
  assign dataGroup_hi_hi_3880 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3881;
  assign dataGroup_hi_hi_3881 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3882;
  assign dataGroup_hi_hi_3882 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3883;
  assign dataGroup_hi_hi_3883 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3884;
  assign dataGroup_hi_hi_3884 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3885;
  assign dataGroup_hi_hi_3885 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3886;
  assign dataGroup_hi_hi_3886 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3887;
  assign dataGroup_hi_hi_3887 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3888;
  assign dataGroup_hi_hi_3888 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3889;
  assign dataGroup_hi_hi_3889 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3890;
  assign dataGroup_hi_hi_3890 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3891;
  assign dataGroup_hi_hi_3891 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3892;
  assign dataGroup_hi_hi_3892 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3893;
  assign dataGroup_hi_hi_3893 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3894;
  assign dataGroup_hi_hi_3894 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3895;
  assign dataGroup_hi_hi_3895 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3896;
  assign dataGroup_hi_hi_3896 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3897;
  assign dataGroup_hi_hi_3897 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3898;
  assign dataGroup_hi_hi_3898 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3899;
  assign dataGroup_hi_hi_3899 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3900;
  assign dataGroup_hi_hi_3900 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3901;
  assign dataGroup_hi_hi_3901 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3902;
  assign dataGroup_hi_hi_3902 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3903;
  assign dataGroup_hi_hi_3903 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3904;
  assign dataGroup_hi_hi_3904 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3905;
  assign dataGroup_hi_hi_3905 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3906;
  assign dataGroup_hi_hi_3906 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3907;
  assign dataGroup_hi_hi_3907 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3908;
  assign dataGroup_hi_hi_3908 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3909;
  assign dataGroup_hi_hi_3909 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3910;
  assign dataGroup_hi_hi_3910 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3911;
  assign dataGroup_hi_hi_3911 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3912;
  assign dataGroup_hi_hi_3912 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3913;
  assign dataGroup_hi_hi_3913 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3914;
  assign dataGroup_hi_hi_3914 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3915;
  assign dataGroup_hi_hi_3915 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3916;
  assign dataGroup_hi_hi_3916 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3917;
  assign dataGroup_hi_hi_3917 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3918;
  assign dataGroup_hi_hi_3918 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3919;
  assign dataGroup_hi_hi_3919 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3920;
  assign dataGroup_hi_hi_3920 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3921;
  assign dataGroup_hi_hi_3921 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3922;
  assign dataGroup_hi_hi_3922 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3923;
  assign dataGroup_hi_hi_3923 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3924;
  assign dataGroup_hi_hi_3924 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3925;
  assign dataGroup_hi_hi_3925 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3926;
  assign dataGroup_hi_hi_3926 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3927;
  assign dataGroup_hi_hi_3927 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3928;
  assign dataGroup_hi_hi_3928 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3929;
  assign dataGroup_hi_hi_3929 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3930;
  assign dataGroup_hi_hi_3930 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3931;
  assign dataGroup_hi_hi_3931 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3932;
  assign dataGroup_hi_hi_3932 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3933;
  assign dataGroup_hi_hi_3933 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3934;
  assign dataGroup_hi_hi_3934 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3935;
  assign dataGroup_hi_hi_3935 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3936;
  assign dataGroup_hi_hi_3936 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3937;
  assign dataGroup_hi_hi_3937 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3938;
  assign dataGroup_hi_hi_3938 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3939;
  assign dataGroup_hi_hi_3939 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3940;
  assign dataGroup_hi_hi_3940 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3941;
  assign dataGroup_hi_hi_3941 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3942;
  assign dataGroup_hi_hi_3942 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3943;
  assign dataGroup_hi_hi_3943 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3944;
  assign dataGroup_hi_hi_3944 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3945;
  assign dataGroup_hi_hi_3945 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3946;
  assign dataGroup_hi_hi_3946 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3947;
  assign dataGroup_hi_hi_3947 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3948;
  assign dataGroup_hi_hi_3948 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3949;
  assign dataGroup_hi_hi_3949 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3950;
  assign dataGroup_hi_hi_3950 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3951;
  assign dataGroup_hi_hi_3951 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3952;
  assign dataGroup_hi_hi_3952 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3953;
  assign dataGroup_hi_hi_3953 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3954;
  assign dataGroup_hi_hi_3954 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3955;
  assign dataGroup_hi_hi_3955 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3956;
  assign dataGroup_hi_hi_3956 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3957;
  assign dataGroup_hi_hi_3957 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3958;
  assign dataGroup_hi_hi_3958 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3959;
  assign dataGroup_hi_hi_3959 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3960;
  assign dataGroup_hi_hi_3960 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3961;
  assign dataGroup_hi_hi_3961 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3962;
  assign dataGroup_hi_hi_3962 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3963;
  assign dataGroup_hi_hi_3963 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3964;
  assign dataGroup_hi_hi_3964 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3965;
  assign dataGroup_hi_hi_3965 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3966;
  assign dataGroup_hi_hi_3966 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3967;
  assign dataGroup_hi_hi_3967 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3968;
  assign dataGroup_hi_hi_3968 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3969;
  assign dataGroup_hi_hi_3969 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3970;
  assign dataGroup_hi_hi_3970 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3971;
  assign dataGroup_hi_hi_3971 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3972;
  assign dataGroup_hi_hi_3972 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3973;
  assign dataGroup_hi_hi_3973 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3974;
  assign dataGroup_hi_hi_3974 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3975;
  assign dataGroup_hi_hi_3975 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3976;
  assign dataGroup_hi_hi_3976 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3977;
  assign dataGroup_hi_hi_3977 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3978;
  assign dataGroup_hi_hi_3978 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3979;
  assign dataGroup_hi_hi_3979 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3980;
  assign dataGroup_hi_hi_3980 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3981;
  assign dataGroup_hi_hi_3981 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3982;
  assign dataGroup_hi_hi_3982 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3983;
  assign dataGroup_hi_hi_3983 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3984;
  assign dataGroup_hi_hi_3984 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3985;
  assign dataGroup_hi_hi_3985 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3986;
  assign dataGroup_hi_hi_3986 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3987;
  assign dataGroup_hi_hi_3987 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3988;
  assign dataGroup_hi_hi_3988 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3989;
  assign dataGroup_hi_hi_3989 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3990;
  assign dataGroup_hi_hi_3990 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3991;
  assign dataGroup_hi_hi_3991 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3992;
  assign dataGroup_hi_hi_3992 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3993;
  assign dataGroup_hi_hi_3993 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3994;
  assign dataGroup_hi_hi_3994 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3995;
  assign dataGroup_hi_hi_3995 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3996;
  assign dataGroup_hi_hi_3996 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3997;
  assign dataGroup_hi_hi_3997 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3998;
  assign dataGroup_hi_hi_3998 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_3999;
  assign dataGroup_hi_hi_3999 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4000;
  assign dataGroup_hi_hi_4000 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4001;
  assign dataGroup_hi_hi_4001 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4002;
  assign dataGroup_hi_hi_4002 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4003;
  assign dataGroup_hi_hi_4003 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4004;
  assign dataGroup_hi_hi_4004 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4005;
  assign dataGroup_hi_hi_4005 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4006;
  assign dataGroup_hi_hi_4006 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4007;
  assign dataGroup_hi_hi_4007 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4008;
  assign dataGroup_hi_hi_4008 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4009;
  assign dataGroup_hi_hi_4009 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4010;
  assign dataGroup_hi_hi_4010 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4011;
  assign dataGroup_hi_hi_4011 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4012;
  assign dataGroup_hi_hi_4012 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4013;
  assign dataGroup_hi_hi_4013 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4014;
  assign dataGroup_hi_hi_4014 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4015;
  assign dataGroup_hi_hi_4015 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4016;
  assign dataGroup_hi_hi_4016 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4017;
  assign dataGroup_hi_hi_4017 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4018;
  assign dataGroup_hi_hi_4018 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4019;
  assign dataGroup_hi_hi_4019 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4020;
  assign dataGroup_hi_hi_4020 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4021;
  assign dataGroup_hi_hi_4021 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4022;
  assign dataGroup_hi_hi_4022 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4023;
  assign dataGroup_hi_hi_4023 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4024;
  assign dataGroup_hi_hi_4024 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4025;
  assign dataGroup_hi_hi_4025 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4026;
  assign dataGroup_hi_hi_4026 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4027;
  assign dataGroup_hi_hi_4027 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4028;
  assign dataGroup_hi_hi_4028 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4029;
  assign dataGroup_hi_hi_4029 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4030;
  assign dataGroup_hi_hi_4030 = _GEN_8;
  wire [1023:0] dataGroup_hi_hi_4031;
  assign dataGroup_hi_hi_4031 = _GEN_8;
  wire [2047:0] dataGroup_hi = {dataGroup_hi_hi, dataGroup_hi_lo};
  wire [7:0]    dataGroup_0 = dataGroup_lo[7:0];
  wire [2047:0] dataGroup_lo_1 = {dataGroup_lo_hi_1, dataGroup_lo_lo_1};
  wire [2047:0] dataGroup_hi_1 = {dataGroup_hi_hi_1, dataGroup_hi_lo_1};
  wire [7:0]    dataGroup_1 = dataGroup_lo_1[15:8];
  wire [2047:0] dataGroup_lo_2 = {dataGroup_lo_hi_2, dataGroup_lo_lo_2};
  wire [2047:0] dataGroup_hi_2 = {dataGroup_hi_hi_2, dataGroup_hi_lo_2};
  wire [7:0]    dataGroup_2 = dataGroup_lo_2[23:16];
  wire [2047:0] dataGroup_lo_3 = {dataGroup_lo_hi_3, dataGroup_lo_lo_3};
  wire [2047:0] dataGroup_hi_3 = {dataGroup_hi_hi_3, dataGroup_hi_lo_3};
  wire [7:0]    dataGroup_3 = dataGroup_lo_3[31:24];
  wire [2047:0] dataGroup_lo_4 = {dataGroup_lo_hi_4, dataGroup_lo_lo_4};
  wire [2047:0] dataGroup_hi_4 = {dataGroup_hi_hi_4, dataGroup_hi_lo_4};
  wire [7:0]    dataGroup_4 = dataGroup_lo_4[39:32];
  wire [2047:0] dataGroup_lo_5 = {dataGroup_lo_hi_5, dataGroup_lo_lo_5};
  wire [2047:0] dataGroup_hi_5 = {dataGroup_hi_hi_5, dataGroup_hi_lo_5};
  wire [7:0]    dataGroup_5 = dataGroup_lo_5[47:40];
  wire [2047:0] dataGroup_lo_6 = {dataGroup_lo_hi_6, dataGroup_lo_lo_6};
  wire [2047:0] dataGroup_hi_6 = {dataGroup_hi_hi_6, dataGroup_hi_lo_6};
  wire [7:0]    dataGroup_6 = dataGroup_lo_6[55:48];
  wire [2047:0] dataGroup_lo_7 = {dataGroup_lo_hi_7, dataGroup_lo_lo_7};
  wire [2047:0] dataGroup_hi_7 = {dataGroup_hi_hi_7, dataGroup_hi_lo_7};
  wire [7:0]    dataGroup_7 = dataGroup_lo_7[63:56];
  wire [2047:0] dataGroup_lo_8 = {dataGroup_lo_hi_8, dataGroup_lo_lo_8};
  wire [2047:0] dataGroup_hi_8 = {dataGroup_hi_hi_8, dataGroup_hi_lo_8};
  wire [7:0]    dataGroup_8 = dataGroup_lo_8[71:64];
  wire [2047:0] dataGroup_lo_9 = {dataGroup_lo_hi_9, dataGroup_lo_lo_9};
  wire [2047:0] dataGroup_hi_9 = {dataGroup_hi_hi_9, dataGroup_hi_lo_9};
  wire [7:0]    dataGroup_9 = dataGroup_lo_9[79:72];
  wire [2047:0] dataGroup_lo_10 = {dataGroup_lo_hi_10, dataGroup_lo_lo_10};
  wire [2047:0] dataGroup_hi_10 = {dataGroup_hi_hi_10, dataGroup_hi_lo_10};
  wire [7:0]    dataGroup_10 = dataGroup_lo_10[87:80];
  wire [2047:0] dataGroup_lo_11 = {dataGroup_lo_hi_11, dataGroup_lo_lo_11};
  wire [2047:0] dataGroup_hi_11 = {dataGroup_hi_hi_11, dataGroup_hi_lo_11};
  wire [7:0]    dataGroup_11 = dataGroup_lo_11[95:88];
  wire [2047:0] dataGroup_lo_12 = {dataGroup_lo_hi_12, dataGroup_lo_lo_12};
  wire [2047:0] dataGroup_hi_12 = {dataGroup_hi_hi_12, dataGroup_hi_lo_12};
  wire [7:0]    dataGroup_12 = dataGroup_lo_12[103:96];
  wire [2047:0] dataGroup_lo_13 = {dataGroup_lo_hi_13, dataGroup_lo_lo_13};
  wire [2047:0] dataGroup_hi_13 = {dataGroup_hi_hi_13, dataGroup_hi_lo_13};
  wire [7:0]    dataGroup_13 = dataGroup_lo_13[111:104];
  wire [2047:0] dataGroup_lo_14 = {dataGroup_lo_hi_14, dataGroup_lo_lo_14};
  wire [2047:0] dataGroup_hi_14 = {dataGroup_hi_hi_14, dataGroup_hi_lo_14};
  wire [7:0]    dataGroup_14 = dataGroup_lo_14[119:112];
  wire [2047:0] dataGroup_lo_15 = {dataGroup_lo_hi_15, dataGroup_lo_lo_15};
  wire [2047:0] dataGroup_hi_15 = {dataGroup_hi_hi_15, dataGroup_hi_lo_15};
  wire [7:0]    dataGroup_15 = dataGroup_lo_15[127:120];
  wire [2047:0] dataGroup_lo_16 = {dataGroup_lo_hi_16, dataGroup_lo_lo_16};
  wire [2047:0] dataGroup_hi_16 = {dataGroup_hi_hi_16, dataGroup_hi_lo_16};
  wire [7:0]    dataGroup_16 = dataGroup_lo_16[135:128];
  wire [2047:0] dataGroup_lo_17 = {dataGroup_lo_hi_17, dataGroup_lo_lo_17};
  wire [2047:0] dataGroup_hi_17 = {dataGroup_hi_hi_17, dataGroup_hi_lo_17};
  wire [7:0]    dataGroup_17 = dataGroup_lo_17[143:136];
  wire [2047:0] dataGroup_lo_18 = {dataGroup_lo_hi_18, dataGroup_lo_lo_18};
  wire [2047:0] dataGroup_hi_18 = {dataGroup_hi_hi_18, dataGroup_hi_lo_18};
  wire [7:0]    dataGroup_18 = dataGroup_lo_18[151:144];
  wire [2047:0] dataGroup_lo_19 = {dataGroup_lo_hi_19, dataGroup_lo_lo_19};
  wire [2047:0] dataGroup_hi_19 = {dataGroup_hi_hi_19, dataGroup_hi_lo_19};
  wire [7:0]    dataGroup_19 = dataGroup_lo_19[159:152];
  wire [2047:0] dataGroup_lo_20 = {dataGroup_lo_hi_20, dataGroup_lo_lo_20};
  wire [2047:0] dataGroup_hi_20 = {dataGroup_hi_hi_20, dataGroup_hi_lo_20};
  wire [7:0]    dataGroup_20 = dataGroup_lo_20[167:160];
  wire [2047:0] dataGroup_lo_21 = {dataGroup_lo_hi_21, dataGroup_lo_lo_21};
  wire [2047:0] dataGroup_hi_21 = {dataGroup_hi_hi_21, dataGroup_hi_lo_21};
  wire [7:0]    dataGroup_21 = dataGroup_lo_21[175:168];
  wire [2047:0] dataGroup_lo_22 = {dataGroup_lo_hi_22, dataGroup_lo_lo_22};
  wire [2047:0] dataGroup_hi_22 = {dataGroup_hi_hi_22, dataGroup_hi_lo_22};
  wire [7:0]    dataGroup_22 = dataGroup_lo_22[183:176];
  wire [2047:0] dataGroup_lo_23 = {dataGroup_lo_hi_23, dataGroup_lo_lo_23};
  wire [2047:0] dataGroup_hi_23 = {dataGroup_hi_hi_23, dataGroup_hi_lo_23};
  wire [7:0]    dataGroup_23 = dataGroup_lo_23[191:184];
  wire [2047:0] dataGroup_lo_24 = {dataGroup_lo_hi_24, dataGroup_lo_lo_24};
  wire [2047:0] dataGroup_hi_24 = {dataGroup_hi_hi_24, dataGroup_hi_lo_24};
  wire [7:0]    dataGroup_24 = dataGroup_lo_24[199:192];
  wire [2047:0] dataGroup_lo_25 = {dataGroup_lo_hi_25, dataGroup_lo_lo_25};
  wire [2047:0] dataGroup_hi_25 = {dataGroup_hi_hi_25, dataGroup_hi_lo_25};
  wire [7:0]    dataGroup_25 = dataGroup_lo_25[207:200];
  wire [2047:0] dataGroup_lo_26 = {dataGroup_lo_hi_26, dataGroup_lo_lo_26};
  wire [2047:0] dataGroup_hi_26 = {dataGroup_hi_hi_26, dataGroup_hi_lo_26};
  wire [7:0]    dataGroup_26 = dataGroup_lo_26[215:208];
  wire [2047:0] dataGroup_lo_27 = {dataGroup_lo_hi_27, dataGroup_lo_lo_27};
  wire [2047:0] dataGroup_hi_27 = {dataGroup_hi_hi_27, dataGroup_hi_lo_27};
  wire [7:0]    dataGroup_27 = dataGroup_lo_27[223:216];
  wire [2047:0] dataGroup_lo_28 = {dataGroup_lo_hi_28, dataGroup_lo_lo_28};
  wire [2047:0] dataGroup_hi_28 = {dataGroup_hi_hi_28, dataGroup_hi_lo_28};
  wire [7:0]    dataGroup_28 = dataGroup_lo_28[231:224];
  wire [2047:0] dataGroup_lo_29 = {dataGroup_lo_hi_29, dataGroup_lo_lo_29};
  wire [2047:0] dataGroup_hi_29 = {dataGroup_hi_hi_29, dataGroup_hi_lo_29};
  wire [7:0]    dataGroup_29 = dataGroup_lo_29[239:232];
  wire [2047:0] dataGroup_lo_30 = {dataGroup_lo_hi_30, dataGroup_lo_lo_30};
  wire [2047:0] dataGroup_hi_30 = {dataGroup_hi_hi_30, dataGroup_hi_lo_30};
  wire [7:0]    dataGroup_30 = dataGroup_lo_30[247:240];
  wire [2047:0] dataGroup_lo_31 = {dataGroup_lo_hi_31, dataGroup_lo_lo_31};
  wire [2047:0] dataGroup_hi_31 = {dataGroup_hi_hi_31, dataGroup_hi_lo_31};
  wire [7:0]    dataGroup_31 = dataGroup_lo_31[255:248];
  wire [2047:0] dataGroup_lo_32 = {dataGroup_lo_hi_32, dataGroup_lo_lo_32};
  wire [2047:0] dataGroup_hi_32 = {dataGroup_hi_hi_32, dataGroup_hi_lo_32};
  wire [7:0]    dataGroup_32 = dataGroup_lo_32[263:256];
  wire [2047:0] dataGroup_lo_33 = {dataGroup_lo_hi_33, dataGroup_lo_lo_33};
  wire [2047:0] dataGroup_hi_33 = {dataGroup_hi_hi_33, dataGroup_hi_lo_33};
  wire [7:0]    dataGroup_33 = dataGroup_lo_33[271:264];
  wire [2047:0] dataGroup_lo_34 = {dataGroup_lo_hi_34, dataGroup_lo_lo_34};
  wire [2047:0] dataGroup_hi_34 = {dataGroup_hi_hi_34, dataGroup_hi_lo_34};
  wire [7:0]    dataGroup_34 = dataGroup_lo_34[279:272];
  wire [2047:0] dataGroup_lo_35 = {dataGroup_lo_hi_35, dataGroup_lo_lo_35};
  wire [2047:0] dataGroup_hi_35 = {dataGroup_hi_hi_35, dataGroup_hi_lo_35};
  wire [7:0]    dataGroup_35 = dataGroup_lo_35[287:280];
  wire [2047:0] dataGroup_lo_36 = {dataGroup_lo_hi_36, dataGroup_lo_lo_36};
  wire [2047:0] dataGroup_hi_36 = {dataGroup_hi_hi_36, dataGroup_hi_lo_36};
  wire [7:0]    dataGroup_36 = dataGroup_lo_36[295:288];
  wire [2047:0] dataGroup_lo_37 = {dataGroup_lo_hi_37, dataGroup_lo_lo_37};
  wire [2047:0] dataGroup_hi_37 = {dataGroup_hi_hi_37, dataGroup_hi_lo_37};
  wire [7:0]    dataGroup_37 = dataGroup_lo_37[303:296];
  wire [2047:0] dataGroup_lo_38 = {dataGroup_lo_hi_38, dataGroup_lo_lo_38};
  wire [2047:0] dataGroup_hi_38 = {dataGroup_hi_hi_38, dataGroup_hi_lo_38};
  wire [7:0]    dataGroup_38 = dataGroup_lo_38[311:304];
  wire [2047:0] dataGroup_lo_39 = {dataGroup_lo_hi_39, dataGroup_lo_lo_39};
  wire [2047:0] dataGroup_hi_39 = {dataGroup_hi_hi_39, dataGroup_hi_lo_39};
  wire [7:0]    dataGroup_39 = dataGroup_lo_39[319:312];
  wire [2047:0] dataGroup_lo_40 = {dataGroup_lo_hi_40, dataGroup_lo_lo_40};
  wire [2047:0] dataGroup_hi_40 = {dataGroup_hi_hi_40, dataGroup_hi_lo_40};
  wire [7:0]    dataGroup_40 = dataGroup_lo_40[327:320];
  wire [2047:0] dataGroup_lo_41 = {dataGroup_lo_hi_41, dataGroup_lo_lo_41};
  wire [2047:0] dataGroup_hi_41 = {dataGroup_hi_hi_41, dataGroup_hi_lo_41};
  wire [7:0]    dataGroup_41 = dataGroup_lo_41[335:328];
  wire [2047:0] dataGroup_lo_42 = {dataGroup_lo_hi_42, dataGroup_lo_lo_42};
  wire [2047:0] dataGroup_hi_42 = {dataGroup_hi_hi_42, dataGroup_hi_lo_42};
  wire [7:0]    dataGroup_42 = dataGroup_lo_42[343:336];
  wire [2047:0] dataGroup_lo_43 = {dataGroup_lo_hi_43, dataGroup_lo_lo_43};
  wire [2047:0] dataGroup_hi_43 = {dataGroup_hi_hi_43, dataGroup_hi_lo_43};
  wire [7:0]    dataGroup_43 = dataGroup_lo_43[351:344];
  wire [2047:0] dataGroup_lo_44 = {dataGroup_lo_hi_44, dataGroup_lo_lo_44};
  wire [2047:0] dataGroup_hi_44 = {dataGroup_hi_hi_44, dataGroup_hi_lo_44};
  wire [7:0]    dataGroup_44 = dataGroup_lo_44[359:352];
  wire [2047:0] dataGroup_lo_45 = {dataGroup_lo_hi_45, dataGroup_lo_lo_45};
  wire [2047:0] dataGroup_hi_45 = {dataGroup_hi_hi_45, dataGroup_hi_lo_45};
  wire [7:0]    dataGroup_45 = dataGroup_lo_45[367:360];
  wire [2047:0] dataGroup_lo_46 = {dataGroup_lo_hi_46, dataGroup_lo_lo_46};
  wire [2047:0] dataGroup_hi_46 = {dataGroup_hi_hi_46, dataGroup_hi_lo_46};
  wire [7:0]    dataGroup_46 = dataGroup_lo_46[375:368];
  wire [2047:0] dataGroup_lo_47 = {dataGroup_lo_hi_47, dataGroup_lo_lo_47};
  wire [2047:0] dataGroup_hi_47 = {dataGroup_hi_hi_47, dataGroup_hi_lo_47};
  wire [7:0]    dataGroup_47 = dataGroup_lo_47[383:376];
  wire [2047:0] dataGroup_lo_48 = {dataGroup_lo_hi_48, dataGroup_lo_lo_48};
  wire [2047:0] dataGroup_hi_48 = {dataGroup_hi_hi_48, dataGroup_hi_lo_48};
  wire [7:0]    dataGroup_48 = dataGroup_lo_48[391:384];
  wire [2047:0] dataGroup_lo_49 = {dataGroup_lo_hi_49, dataGroup_lo_lo_49};
  wire [2047:0] dataGroup_hi_49 = {dataGroup_hi_hi_49, dataGroup_hi_lo_49};
  wire [7:0]    dataGroup_49 = dataGroup_lo_49[399:392];
  wire [2047:0] dataGroup_lo_50 = {dataGroup_lo_hi_50, dataGroup_lo_lo_50};
  wire [2047:0] dataGroup_hi_50 = {dataGroup_hi_hi_50, dataGroup_hi_lo_50};
  wire [7:0]    dataGroup_50 = dataGroup_lo_50[407:400];
  wire [2047:0] dataGroup_lo_51 = {dataGroup_lo_hi_51, dataGroup_lo_lo_51};
  wire [2047:0] dataGroup_hi_51 = {dataGroup_hi_hi_51, dataGroup_hi_lo_51};
  wire [7:0]    dataGroup_51 = dataGroup_lo_51[415:408];
  wire [2047:0] dataGroup_lo_52 = {dataGroup_lo_hi_52, dataGroup_lo_lo_52};
  wire [2047:0] dataGroup_hi_52 = {dataGroup_hi_hi_52, dataGroup_hi_lo_52};
  wire [7:0]    dataGroup_52 = dataGroup_lo_52[423:416];
  wire [2047:0] dataGroup_lo_53 = {dataGroup_lo_hi_53, dataGroup_lo_lo_53};
  wire [2047:0] dataGroup_hi_53 = {dataGroup_hi_hi_53, dataGroup_hi_lo_53};
  wire [7:0]    dataGroup_53 = dataGroup_lo_53[431:424];
  wire [2047:0] dataGroup_lo_54 = {dataGroup_lo_hi_54, dataGroup_lo_lo_54};
  wire [2047:0] dataGroup_hi_54 = {dataGroup_hi_hi_54, dataGroup_hi_lo_54};
  wire [7:0]    dataGroup_54 = dataGroup_lo_54[439:432];
  wire [2047:0] dataGroup_lo_55 = {dataGroup_lo_hi_55, dataGroup_lo_lo_55};
  wire [2047:0] dataGroup_hi_55 = {dataGroup_hi_hi_55, dataGroup_hi_lo_55};
  wire [7:0]    dataGroup_55 = dataGroup_lo_55[447:440];
  wire [2047:0] dataGroup_lo_56 = {dataGroup_lo_hi_56, dataGroup_lo_lo_56};
  wire [2047:0] dataGroup_hi_56 = {dataGroup_hi_hi_56, dataGroup_hi_lo_56};
  wire [7:0]    dataGroup_56 = dataGroup_lo_56[455:448];
  wire [2047:0] dataGroup_lo_57 = {dataGroup_lo_hi_57, dataGroup_lo_lo_57};
  wire [2047:0] dataGroup_hi_57 = {dataGroup_hi_hi_57, dataGroup_hi_lo_57};
  wire [7:0]    dataGroup_57 = dataGroup_lo_57[463:456];
  wire [2047:0] dataGroup_lo_58 = {dataGroup_lo_hi_58, dataGroup_lo_lo_58};
  wire [2047:0] dataGroup_hi_58 = {dataGroup_hi_hi_58, dataGroup_hi_lo_58};
  wire [7:0]    dataGroup_58 = dataGroup_lo_58[471:464];
  wire [2047:0] dataGroup_lo_59 = {dataGroup_lo_hi_59, dataGroup_lo_lo_59};
  wire [2047:0] dataGroup_hi_59 = {dataGroup_hi_hi_59, dataGroup_hi_lo_59};
  wire [7:0]    dataGroup_59 = dataGroup_lo_59[479:472];
  wire [2047:0] dataGroup_lo_60 = {dataGroup_lo_hi_60, dataGroup_lo_lo_60};
  wire [2047:0] dataGroup_hi_60 = {dataGroup_hi_hi_60, dataGroup_hi_lo_60};
  wire [7:0]    dataGroup_60 = dataGroup_lo_60[487:480];
  wire [2047:0] dataGroup_lo_61 = {dataGroup_lo_hi_61, dataGroup_lo_lo_61};
  wire [2047:0] dataGroup_hi_61 = {dataGroup_hi_hi_61, dataGroup_hi_lo_61};
  wire [7:0]    dataGroup_61 = dataGroup_lo_61[495:488];
  wire [2047:0] dataGroup_lo_62 = {dataGroup_lo_hi_62, dataGroup_lo_lo_62};
  wire [2047:0] dataGroup_hi_62 = {dataGroup_hi_hi_62, dataGroup_hi_lo_62};
  wire [7:0]    dataGroup_62 = dataGroup_lo_62[503:496];
  wire [2047:0] dataGroup_lo_63 = {dataGroup_lo_hi_63, dataGroup_lo_lo_63};
  wire [2047:0] dataGroup_hi_63 = {dataGroup_hi_hi_63, dataGroup_hi_lo_63};
  wire [7:0]    dataGroup_63 = dataGroup_lo_63[511:504];
  wire [15:0]   res_lo_lo_lo_lo_lo = {dataGroup_1, dataGroup_0};
  wire [15:0]   res_lo_lo_lo_lo_hi = {dataGroup_3, dataGroup_2};
  wire [31:0]   res_lo_lo_lo_lo = {res_lo_lo_lo_lo_hi, res_lo_lo_lo_lo_lo};
  wire [15:0]   res_lo_lo_lo_hi_lo = {dataGroup_5, dataGroup_4};
  wire [15:0]   res_lo_lo_lo_hi_hi = {dataGroup_7, dataGroup_6};
  wire [31:0]   res_lo_lo_lo_hi = {res_lo_lo_lo_hi_hi, res_lo_lo_lo_hi_lo};
  wire [63:0]   res_lo_lo_lo = {res_lo_lo_lo_hi, res_lo_lo_lo_lo};
  wire [15:0]   res_lo_lo_hi_lo_lo = {dataGroup_9, dataGroup_8};
  wire [15:0]   res_lo_lo_hi_lo_hi = {dataGroup_11, dataGroup_10};
  wire [31:0]   res_lo_lo_hi_lo = {res_lo_lo_hi_lo_hi, res_lo_lo_hi_lo_lo};
  wire [15:0]   res_lo_lo_hi_hi_lo = {dataGroup_13, dataGroup_12};
  wire [15:0]   res_lo_lo_hi_hi_hi = {dataGroup_15, dataGroup_14};
  wire [31:0]   res_lo_lo_hi_hi = {res_lo_lo_hi_hi_hi, res_lo_lo_hi_hi_lo};
  wire [63:0]   res_lo_lo_hi = {res_lo_lo_hi_hi, res_lo_lo_hi_lo};
  wire [127:0]  res_lo_lo = {res_lo_lo_hi, res_lo_lo_lo};
  wire [15:0]   res_lo_hi_lo_lo_lo = {dataGroup_17, dataGroup_16};
  wire [15:0]   res_lo_hi_lo_lo_hi = {dataGroup_19, dataGroup_18};
  wire [31:0]   res_lo_hi_lo_lo = {res_lo_hi_lo_lo_hi, res_lo_hi_lo_lo_lo};
  wire [15:0]   res_lo_hi_lo_hi_lo = {dataGroup_21, dataGroup_20};
  wire [15:0]   res_lo_hi_lo_hi_hi = {dataGroup_23, dataGroup_22};
  wire [31:0]   res_lo_hi_lo_hi = {res_lo_hi_lo_hi_hi, res_lo_hi_lo_hi_lo};
  wire [63:0]   res_lo_hi_lo = {res_lo_hi_lo_hi, res_lo_hi_lo_lo};
  wire [15:0]   res_lo_hi_hi_lo_lo = {dataGroup_25, dataGroup_24};
  wire [15:0]   res_lo_hi_hi_lo_hi = {dataGroup_27, dataGroup_26};
  wire [31:0]   res_lo_hi_hi_lo = {res_lo_hi_hi_lo_hi, res_lo_hi_hi_lo_lo};
  wire [15:0]   res_lo_hi_hi_hi_lo = {dataGroup_29, dataGroup_28};
  wire [15:0]   res_lo_hi_hi_hi_hi = {dataGroup_31, dataGroup_30};
  wire [31:0]   res_lo_hi_hi_hi = {res_lo_hi_hi_hi_hi, res_lo_hi_hi_hi_lo};
  wire [63:0]   res_lo_hi_hi = {res_lo_hi_hi_hi, res_lo_hi_hi_lo};
  wire [127:0]  res_lo_hi = {res_lo_hi_hi, res_lo_hi_lo};
  wire [255:0]  res_lo = {res_lo_hi, res_lo_lo};
  wire [15:0]   res_hi_lo_lo_lo_lo = {dataGroup_33, dataGroup_32};
  wire [15:0]   res_hi_lo_lo_lo_hi = {dataGroup_35, dataGroup_34};
  wire [31:0]   res_hi_lo_lo_lo = {res_hi_lo_lo_lo_hi, res_hi_lo_lo_lo_lo};
  wire [15:0]   res_hi_lo_lo_hi_lo = {dataGroup_37, dataGroup_36};
  wire [15:0]   res_hi_lo_lo_hi_hi = {dataGroup_39, dataGroup_38};
  wire [31:0]   res_hi_lo_lo_hi = {res_hi_lo_lo_hi_hi, res_hi_lo_lo_hi_lo};
  wire [63:0]   res_hi_lo_lo = {res_hi_lo_lo_hi, res_hi_lo_lo_lo};
  wire [15:0]   res_hi_lo_hi_lo_lo = {dataGroup_41, dataGroup_40};
  wire [15:0]   res_hi_lo_hi_lo_hi = {dataGroup_43, dataGroup_42};
  wire [31:0]   res_hi_lo_hi_lo = {res_hi_lo_hi_lo_hi, res_hi_lo_hi_lo_lo};
  wire [15:0]   res_hi_lo_hi_hi_lo = {dataGroup_45, dataGroup_44};
  wire [15:0]   res_hi_lo_hi_hi_hi = {dataGroup_47, dataGroup_46};
  wire [31:0]   res_hi_lo_hi_hi = {res_hi_lo_hi_hi_hi, res_hi_lo_hi_hi_lo};
  wire [63:0]   res_hi_lo_hi = {res_hi_lo_hi_hi, res_hi_lo_hi_lo};
  wire [127:0]  res_hi_lo = {res_hi_lo_hi, res_hi_lo_lo};
  wire [15:0]   res_hi_hi_lo_lo_lo = {dataGroup_49, dataGroup_48};
  wire [15:0]   res_hi_hi_lo_lo_hi = {dataGroup_51, dataGroup_50};
  wire [31:0]   res_hi_hi_lo_lo = {res_hi_hi_lo_lo_hi, res_hi_hi_lo_lo_lo};
  wire [15:0]   res_hi_hi_lo_hi_lo = {dataGroup_53, dataGroup_52};
  wire [15:0]   res_hi_hi_lo_hi_hi = {dataGroup_55, dataGroup_54};
  wire [31:0]   res_hi_hi_lo_hi = {res_hi_hi_lo_hi_hi, res_hi_hi_lo_hi_lo};
  wire [63:0]   res_hi_hi_lo = {res_hi_hi_lo_hi, res_hi_hi_lo_lo};
  wire [15:0]   res_hi_hi_hi_lo_lo = {dataGroup_57, dataGroup_56};
  wire [15:0]   res_hi_hi_hi_lo_hi = {dataGroup_59, dataGroup_58};
  wire [31:0]   res_hi_hi_hi_lo = {res_hi_hi_hi_lo_hi, res_hi_hi_hi_lo_lo};
  wire [15:0]   res_hi_hi_hi_hi_lo = {dataGroup_61, dataGroup_60};
  wire [15:0]   res_hi_hi_hi_hi_hi = {dataGroup_63, dataGroup_62};
  wire [31:0]   res_hi_hi_hi_hi = {res_hi_hi_hi_hi_hi, res_hi_hi_hi_hi_lo};
  wire [63:0]   res_hi_hi_hi = {res_hi_hi_hi_hi, res_hi_hi_hi_lo};
  wire [127:0]  res_hi_hi = {res_hi_hi_hi, res_hi_hi_lo};
  wire [255:0]  res_hi = {res_hi_hi, res_hi_lo};
  wire [511:0]  res = {res_hi, res_lo};
  wire [1023:0] lo_lo = {512'h0, res};
  wire [2047:0] lo = {1024'h0, lo_lo};
  wire [4095:0] regroupLoadData_0_0 = {2048'h0, lo};
  wire [2047:0] dataGroup_lo_64 = {dataGroup_lo_hi_64, dataGroup_lo_lo_64};
  wire [2047:0] dataGroup_hi_64 = {dataGroup_hi_hi_64, dataGroup_hi_lo_64};
  wire [7:0]    dataGroup_0_1 = dataGroup_lo_64[7:0];
  wire [2047:0] dataGroup_lo_65 = {dataGroup_lo_hi_65, dataGroup_lo_lo_65};
  wire [2047:0] dataGroup_hi_65 = {dataGroup_hi_hi_65, dataGroup_hi_lo_65};
  wire [7:0]    dataGroup_1_1 = dataGroup_lo_65[23:16];
  wire [2047:0] dataGroup_lo_66 = {dataGroup_lo_hi_66, dataGroup_lo_lo_66};
  wire [2047:0] dataGroup_hi_66 = {dataGroup_hi_hi_66, dataGroup_hi_lo_66};
  wire [7:0]    dataGroup_2_1 = dataGroup_lo_66[39:32];
  wire [2047:0] dataGroup_lo_67 = {dataGroup_lo_hi_67, dataGroup_lo_lo_67};
  wire [2047:0] dataGroup_hi_67 = {dataGroup_hi_hi_67, dataGroup_hi_lo_67};
  wire [7:0]    dataGroup_3_1 = dataGroup_lo_67[55:48];
  wire [2047:0] dataGroup_lo_68 = {dataGroup_lo_hi_68, dataGroup_lo_lo_68};
  wire [2047:0] dataGroup_hi_68 = {dataGroup_hi_hi_68, dataGroup_hi_lo_68};
  wire [7:0]    dataGroup_4_1 = dataGroup_lo_68[71:64];
  wire [2047:0] dataGroup_lo_69 = {dataGroup_lo_hi_69, dataGroup_lo_lo_69};
  wire [2047:0] dataGroup_hi_69 = {dataGroup_hi_hi_69, dataGroup_hi_lo_69};
  wire [7:0]    dataGroup_5_1 = dataGroup_lo_69[87:80];
  wire [2047:0] dataGroup_lo_70 = {dataGroup_lo_hi_70, dataGroup_lo_lo_70};
  wire [2047:0] dataGroup_hi_70 = {dataGroup_hi_hi_70, dataGroup_hi_lo_70};
  wire [7:0]    dataGroup_6_1 = dataGroup_lo_70[103:96];
  wire [2047:0] dataGroup_lo_71 = {dataGroup_lo_hi_71, dataGroup_lo_lo_71};
  wire [2047:0] dataGroup_hi_71 = {dataGroup_hi_hi_71, dataGroup_hi_lo_71};
  wire [7:0]    dataGroup_7_1 = dataGroup_lo_71[119:112];
  wire [2047:0] dataGroup_lo_72 = {dataGroup_lo_hi_72, dataGroup_lo_lo_72};
  wire [2047:0] dataGroup_hi_72 = {dataGroup_hi_hi_72, dataGroup_hi_lo_72};
  wire [7:0]    dataGroup_8_1 = dataGroup_lo_72[135:128];
  wire [2047:0] dataGroup_lo_73 = {dataGroup_lo_hi_73, dataGroup_lo_lo_73};
  wire [2047:0] dataGroup_hi_73 = {dataGroup_hi_hi_73, dataGroup_hi_lo_73};
  wire [7:0]    dataGroup_9_1 = dataGroup_lo_73[151:144];
  wire [2047:0] dataGroup_lo_74 = {dataGroup_lo_hi_74, dataGroup_lo_lo_74};
  wire [2047:0] dataGroup_hi_74 = {dataGroup_hi_hi_74, dataGroup_hi_lo_74};
  wire [7:0]    dataGroup_10_1 = dataGroup_lo_74[167:160];
  wire [2047:0] dataGroup_lo_75 = {dataGroup_lo_hi_75, dataGroup_lo_lo_75};
  wire [2047:0] dataGroup_hi_75 = {dataGroup_hi_hi_75, dataGroup_hi_lo_75};
  wire [7:0]    dataGroup_11_1 = dataGroup_lo_75[183:176];
  wire [2047:0] dataGroup_lo_76 = {dataGroup_lo_hi_76, dataGroup_lo_lo_76};
  wire [2047:0] dataGroup_hi_76 = {dataGroup_hi_hi_76, dataGroup_hi_lo_76};
  wire [7:0]    dataGroup_12_1 = dataGroup_lo_76[199:192];
  wire [2047:0] dataGroup_lo_77 = {dataGroup_lo_hi_77, dataGroup_lo_lo_77};
  wire [2047:0] dataGroup_hi_77 = {dataGroup_hi_hi_77, dataGroup_hi_lo_77};
  wire [7:0]    dataGroup_13_1 = dataGroup_lo_77[215:208];
  wire [2047:0] dataGroup_lo_78 = {dataGroup_lo_hi_78, dataGroup_lo_lo_78};
  wire [2047:0] dataGroup_hi_78 = {dataGroup_hi_hi_78, dataGroup_hi_lo_78};
  wire [7:0]    dataGroup_14_1 = dataGroup_lo_78[231:224];
  wire [2047:0] dataGroup_lo_79 = {dataGroup_lo_hi_79, dataGroup_lo_lo_79};
  wire [2047:0] dataGroup_hi_79 = {dataGroup_hi_hi_79, dataGroup_hi_lo_79};
  wire [7:0]    dataGroup_15_1 = dataGroup_lo_79[247:240];
  wire [2047:0] dataGroup_lo_80 = {dataGroup_lo_hi_80, dataGroup_lo_lo_80};
  wire [2047:0] dataGroup_hi_80 = {dataGroup_hi_hi_80, dataGroup_hi_lo_80};
  wire [7:0]    dataGroup_16_1 = dataGroup_lo_80[263:256];
  wire [2047:0] dataGroup_lo_81 = {dataGroup_lo_hi_81, dataGroup_lo_lo_81};
  wire [2047:0] dataGroup_hi_81 = {dataGroup_hi_hi_81, dataGroup_hi_lo_81};
  wire [7:0]    dataGroup_17_1 = dataGroup_lo_81[279:272];
  wire [2047:0] dataGroup_lo_82 = {dataGroup_lo_hi_82, dataGroup_lo_lo_82};
  wire [2047:0] dataGroup_hi_82 = {dataGroup_hi_hi_82, dataGroup_hi_lo_82};
  wire [7:0]    dataGroup_18_1 = dataGroup_lo_82[295:288];
  wire [2047:0] dataGroup_lo_83 = {dataGroup_lo_hi_83, dataGroup_lo_lo_83};
  wire [2047:0] dataGroup_hi_83 = {dataGroup_hi_hi_83, dataGroup_hi_lo_83};
  wire [7:0]    dataGroup_19_1 = dataGroup_lo_83[311:304];
  wire [2047:0] dataGroup_lo_84 = {dataGroup_lo_hi_84, dataGroup_lo_lo_84};
  wire [2047:0] dataGroup_hi_84 = {dataGroup_hi_hi_84, dataGroup_hi_lo_84};
  wire [7:0]    dataGroup_20_1 = dataGroup_lo_84[327:320];
  wire [2047:0] dataGroup_lo_85 = {dataGroup_lo_hi_85, dataGroup_lo_lo_85};
  wire [2047:0] dataGroup_hi_85 = {dataGroup_hi_hi_85, dataGroup_hi_lo_85};
  wire [7:0]    dataGroup_21_1 = dataGroup_lo_85[343:336];
  wire [2047:0] dataGroup_lo_86 = {dataGroup_lo_hi_86, dataGroup_lo_lo_86};
  wire [2047:0] dataGroup_hi_86 = {dataGroup_hi_hi_86, dataGroup_hi_lo_86};
  wire [7:0]    dataGroup_22_1 = dataGroup_lo_86[359:352];
  wire [2047:0] dataGroup_lo_87 = {dataGroup_lo_hi_87, dataGroup_lo_lo_87};
  wire [2047:0] dataGroup_hi_87 = {dataGroup_hi_hi_87, dataGroup_hi_lo_87};
  wire [7:0]    dataGroup_23_1 = dataGroup_lo_87[375:368];
  wire [2047:0] dataGroup_lo_88 = {dataGroup_lo_hi_88, dataGroup_lo_lo_88};
  wire [2047:0] dataGroup_hi_88 = {dataGroup_hi_hi_88, dataGroup_hi_lo_88};
  wire [7:0]    dataGroup_24_1 = dataGroup_lo_88[391:384];
  wire [2047:0] dataGroup_lo_89 = {dataGroup_lo_hi_89, dataGroup_lo_lo_89};
  wire [2047:0] dataGroup_hi_89 = {dataGroup_hi_hi_89, dataGroup_hi_lo_89};
  wire [7:0]    dataGroup_25_1 = dataGroup_lo_89[407:400];
  wire [2047:0] dataGroup_lo_90 = {dataGroup_lo_hi_90, dataGroup_lo_lo_90};
  wire [2047:0] dataGroup_hi_90 = {dataGroup_hi_hi_90, dataGroup_hi_lo_90};
  wire [7:0]    dataGroup_26_1 = dataGroup_lo_90[423:416];
  wire [2047:0] dataGroup_lo_91 = {dataGroup_lo_hi_91, dataGroup_lo_lo_91};
  wire [2047:0] dataGroup_hi_91 = {dataGroup_hi_hi_91, dataGroup_hi_lo_91};
  wire [7:0]    dataGroup_27_1 = dataGroup_lo_91[439:432];
  wire [2047:0] dataGroup_lo_92 = {dataGroup_lo_hi_92, dataGroup_lo_lo_92};
  wire [2047:0] dataGroup_hi_92 = {dataGroup_hi_hi_92, dataGroup_hi_lo_92};
  wire [7:0]    dataGroup_28_1 = dataGroup_lo_92[455:448];
  wire [2047:0] dataGroup_lo_93 = {dataGroup_lo_hi_93, dataGroup_lo_lo_93};
  wire [2047:0] dataGroup_hi_93 = {dataGroup_hi_hi_93, dataGroup_hi_lo_93};
  wire [7:0]    dataGroup_29_1 = dataGroup_lo_93[471:464];
  wire [2047:0] dataGroup_lo_94 = {dataGroup_lo_hi_94, dataGroup_lo_lo_94};
  wire [2047:0] dataGroup_hi_94 = {dataGroup_hi_hi_94, dataGroup_hi_lo_94};
  wire [7:0]    dataGroup_30_1 = dataGroup_lo_94[487:480];
  wire [2047:0] dataGroup_lo_95 = {dataGroup_lo_hi_95, dataGroup_lo_lo_95};
  wire [2047:0] dataGroup_hi_95 = {dataGroup_hi_hi_95, dataGroup_hi_lo_95};
  wire [7:0]    dataGroup_31_1 = dataGroup_lo_95[503:496];
  wire [2047:0] dataGroup_lo_96 = {dataGroup_lo_hi_96, dataGroup_lo_lo_96};
  wire [2047:0] dataGroup_hi_96 = {dataGroup_hi_hi_96, dataGroup_hi_lo_96};
  wire [7:0]    dataGroup_32_1 = dataGroup_lo_96[519:512];
  wire [2047:0] dataGroup_lo_97 = {dataGroup_lo_hi_97, dataGroup_lo_lo_97};
  wire [2047:0] dataGroup_hi_97 = {dataGroup_hi_hi_97, dataGroup_hi_lo_97};
  wire [7:0]    dataGroup_33_1 = dataGroup_lo_97[535:528];
  wire [2047:0] dataGroup_lo_98 = {dataGroup_lo_hi_98, dataGroup_lo_lo_98};
  wire [2047:0] dataGroup_hi_98 = {dataGroup_hi_hi_98, dataGroup_hi_lo_98};
  wire [7:0]    dataGroup_34_1 = dataGroup_lo_98[551:544];
  wire [2047:0] dataGroup_lo_99 = {dataGroup_lo_hi_99, dataGroup_lo_lo_99};
  wire [2047:0] dataGroup_hi_99 = {dataGroup_hi_hi_99, dataGroup_hi_lo_99};
  wire [7:0]    dataGroup_35_1 = dataGroup_lo_99[567:560];
  wire [2047:0] dataGroup_lo_100 = {dataGroup_lo_hi_100, dataGroup_lo_lo_100};
  wire [2047:0] dataGroup_hi_100 = {dataGroup_hi_hi_100, dataGroup_hi_lo_100};
  wire [7:0]    dataGroup_36_1 = dataGroup_lo_100[583:576];
  wire [2047:0] dataGroup_lo_101 = {dataGroup_lo_hi_101, dataGroup_lo_lo_101};
  wire [2047:0] dataGroup_hi_101 = {dataGroup_hi_hi_101, dataGroup_hi_lo_101};
  wire [7:0]    dataGroup_37_1 = dataGroup_lo_101[599:592];
  wire [2047:0] dataGroup_lo_102 = {dataGroup_lo_hi_102, dataGroup_lo_lo_102};
  wire [2047:0] dataGroup_hi_102 = {dataGroup_hi_hi_102, dataGroup_hi_lo_102};
  wire [7:0]    dataGroup_38_1 = dataGroup_lo_102[615:608];
  wire [2047:0] dataGroup_lo_103 = {dataGroup_lo_hi_103, dataGroup_lo_lo_103};
  wire [2047:0] dataGroup_hi_103 = {dataGroup_hi_hi_103, dataGroup_hi_lo_103};
  wire [7:0]    dataGroup_39_1 = dataGroup_lo_103[631:624];
  wire [2047:0] dataGroup_lo_104 = {dataGroup_lo_hi_104, dataGroup_lo_lo_104};
  wire [2047:0] dataGroup_hi_104 = {dataGroup_hi_hi_104, dataGroup_hi_lo_104};
  wire [7:0]    dataGroup_40_1 = dataGroup_lo_104[647:640];
  wire [2047:0] dataGroup_lo_105 = {dataGroup_lo_hi_105, dataGroup_lo_lo_105};
  wire [2047:0] dataGroup_hi_105 = {dataGroup_hi_hi_105, dataGroup_hi_lo_105};
  wire [7:0]    dataGroup_41_1 = dataGroup_lo_105[663:656];
  wire [2047:0] dataGroup_lo_106 = {dataGroup_lo_hi_106, dataGroup_lo_lo_106};
  wire [2047:0] dataGroup_hi_106 = {dataGroup_hi_hi_106, dataGroup_hi_lo_106};
  wire [7:0]    dataGroup_42_1 = dataGroup_lo_106[679:672];
  wire [2047:0] dataGroup_lo_107 = {dataGroup_lo_hi_107, dataGroup_lo_lo_107};
  wire [2047:0] dataGroup_hi_107 = {dataGroup_hi_hi_107, dataGroup_hi_lo_107};
  wire [7:0]    dataGroup_43_1 = dataGroup_lo_107[695:688];
  wire [2047:0] dataGroup_lo_108 = {dataGroup_lo_hi_108, dataGroup_lo_lo_108};
  wire [2047:0] dataGroup_hi_108 = {dataGroup_hi_hi_108, dataGroup_hi_lo_108};
  wire [7:0]    dataGroup_44_1 = dataGroup_lo_108[711:704];
  wire [2047:0] dataGroup_lo_109 = {dataGroup_lo_hi_109, dataGroup_lo_lo_109};
  wire [2047:0] dataGroup_hi_109 = {dataGroup_hi_hi_109, dataGroup_hi_lo_109};
  wire [7:0]    dataGroup_45_1 = dataGroup_lo_109[727:720];
  wire [2047:0] dataGroup_lo_110 = {dataGroup_lo_hi_110, dataGroup_lo_lo_110};
  wire [2047:0] dataGroup_hi_110 = {dataGroup_hi_hi_110, dataGroup_hi_lo_110};
  wire [7:0]    dataGroup_46_1 = dataGroup_lo_110[743:736];
  wire [2047:0] dataGroup_lo_111 = {dataGroup_lo_hi_111, dataGroup_lo_lo_111};
  wire [2047:0] dataGroup_hi_111 = {dataGroup_hi_hi_111, dataGroup_hi_lo_111};
  wire [7:0]    dataGroup_47_1 = dataGroup_lo_111[759:752];
  wire [2047:0] dataGroup_lo_112 = {dataGroup_lo_hi_112, dataGroup_lo_lo_112};
  wire [2047:0] dataGroup_hi_112 = {dataGroup_hi_hi_112, dataGroup_hi_lo_112};
  wire [7:0]    dataGroup_48_1 = dataGroup_lo_112[775:768];
  wire [2047:0] dataGroup_lo_113 = {dataGroup_lo_hi_113, dataGroup_lo_lo_113};
  wire [2047:0] dataGroup_hi_113 = {dataGroup_hi_hi_113, dataGroup_hi_lo_113};
  wire [7:0]    dataGroup_49_1 = dataGroup_lo_113[791:784];
  wire [2047:0] dataGroup_lo_114 = {dataGroup_lo_hi_114, dataGroup_lo_lo_114};
  wire [2047:0] dataGroup_hi_114 = {dataGroup_hi_hi_114, dataGroup_hi_lo_114};
  wire [7:0]    dataGroup_50_1 = dataGroup_lo_114[807:800];
  wire [2047:0] dataGroup_lo_115 = {dataGroup_lo_hi_115, dataGroup_lo_lo_115};
  wire [2047:0] dataGroup_hi_115 = {dataGroup_hi_hi_115, dataGroup_hi_lo_115};
  wire [7:0]    dataGroup_51_1 = dataGroup_lo_115[823:816];
  wire [2047:0] dataGroup_lo_116 = {dataGroup_lo_hi_116, dataGroup_lo_lo_116};
  wire [2047:0] dataGroup_hi_116 = {dataGroup_hi_hi_116, dataGroup_hi_lo_116};
  wire [7:0]    dataGroup_52_1 = dataGroup_lo_116[839:832];
  wire [2047:0] dataGroup_lo_117 = {dataGroup_lo_hi_117, dataGroup_lo_lo_117};
  wire [2047:0] dataGroup_hi_117 = {dataGroup_hi_hi_117, dataGroup_hi_lo_117};
  wire [7:0]    dataGroup_53_1 = dataGroup_lo_117[855:848];
  wire [2047:0] dataGroup_lo_118 = {dataGroup_lo_hi_118, dataGroup_lo_lo_118};
  wire [2047:0] dataGroup_hi_118 = {dataGroup_hi_hi_118, dataGroup_hi_lo_118};
  wire [7:0]    dataGroup_54_1 = dataGroup_lo_118[871:864];
  wire [2047:0] dataGroup_lo_119 = {dataGroup_lo_hi_119, dataGroup_lo_lo_119};
  wire [2047:0] dataGroup_hi_119 = {dataGroup_hi_hi_119, dataGroup_hi_lo_119};
  wire [7:0]    dataGroup_55_1 = dataGroup_lo_119[887:880];
  wire [2047:0] dataGroup_lo_120 = {dataGroup_lo_hi_120, dataGroup_lo_lo_120};
  wire [2047:0] dataGroup_hi_120 = {dataGroup_hi_hi_120, dataGroup_hi_lo_120};
  wire [7:0]    dataGroup_56_1 = dataGroup_lo_120[903:896];
  wire [2047:0] dataGroup_lo_121 = {dataGroup_lo_hi_121, dataGroup_lo_lo_121};
  wire [2047:0] dataGroup_hi_121 = {dataGroup_hi_hi_121, dataGroup_hi_lo_121};
  wire [7:0]    dataGroup_57_1 = dataGroup_lo_121[919:912];
  wire [2047:0] dataGroup_lo_122 = {dataGroup_lo_hi_122, dataGroup_lo_lo_122};
  wire [2047:0] dataGroup_hi_122 = {dataGroup_hi_hi_122, dataGroup_hi_lo_122};
  wire [7:0]    dataGroup_58_1 = dataGroup_lo_122[935:928];
  wire [2047:0] dataGroup_lo_123 = {dataGroup_lo_hi_123, dataGroup_lo_lo_123};
  wire [2047:0] dataGroup_hi_123 = {dataGroup_hi_hi_123, dataGroup_hi_lo_123};
  wire [7:0]    dataGroup_59_1 = dataGroup_lo_123[951:944];
  wire [2047:0] dataGroup_lo_124 = {dataGroup_lo_hi_124, dataGroup_lo_lo_124};
  wire [2047:0] dataGroup_hi_124 = {dataGroup_hi_hi_124, dataGroup_hi_lo_124};
  wire [7:0]    dataGroup_60_1 = dataGroup_lo_124[967:960];
  wire [2047:0] dataGroup_lo_125 = {dataGroup_lo_hi_125, dataGroup_lo_lo_125};
  wire [2047:0] dataGroup_hi_125 = {dataGroup_hi_hi_125, dataGroup_hi_lo_125};
  wire [7:0]    dataGroup_61_1 = dataGroup_lo_125[983:976];
  wire [2047:0] dataGroup_lo_126 = {dataGroup_lo_hi_126, dataGroup_lo_lo_126};
  wire [2047:0] dataGroup_hi_126 = {dataGroup_hi_hi_126, dataGroup_hi_lo_126};
  wire [7:0]    dataGroup_62_1 = dataGroup_lo_126[999:992];
  wire [2047:0] dataGroup_lo_127 = {dataGroup_lo_hi_127, dataGroup_lo_lo_127};
  wire [2047:0] dataGroup_hi_127 = {dataGroup_hi_hi_127, dataGroup_hi_lo_127};
  wire [7:0]    dataGroup_63_1 = dataGroup_lo_127[1015:1008];
  wire [15:0]   res_lo_lo_lo_lo_lo_1 = {dataGroup_1_1, dataGroup_0_1};
  wire [15:0]   res_lo_lo_lo_lo_hi_1 = {dataGroup_3_1, dataGroup_2_1};
  wire [31:0]   res_lo_lo_lo_lo_1 = {res_lo_lo_lo_lo_hi_1, res_lo_lo_lo_lo_lo_1};
  wire [15:0]   res_lo_lo_lo_hi_lo_1 = {dataGroup_5_1, dataGroup_4_1};
  wire [15:0]   res_lo_lo_lo_hi_hi_1 = {dataGroup_7_1, dataGroup_6_1};
  wire [31:0]   res_lo_lo_lo_hi_1 = {res_lo_lo_lo_hi_hi_1, res_lo_lo_lo_hi_lo_1};
  wire [63:0]   res_lo_lo_lo_1 = {res_lo_lo_lo_hi_1, res_lo_lo_lo_lo_1};
  wire [15:0]   res_lo_lo_hi_lo_lo_1 = {dataGroup_9_1, dataGroup_8_1};
  wire [15:0]   res_lo_lo_hi_lo_hi_1 = {dataGroup_11_1, dataGroup_10_1};
  wire [31:0]   res_lo_lo_hi_lo_1 = {res_lo_lo_hi_lo_hi_1, res_lo_lo_hi_lo_lo_1};
  wire [15:0]   res_lo_lo_hi_hi_lo_1 = {dataGroup_13_1, dataGroup_12_1};
  wire [15:0]   res_lo_lo_hi_hi_hi_1 = {dataGroup_15_1, dataGroup_14_1};
  wire [31:0]   res_lo_lo_hi_hi_1 = {res_lo_lo_hi_hi_hi_1, res_lo_lo_hi_hi_lo_1};
  wire [63:0]   res_lo_lo_hi_1 = {res_lo_lo_hi_hi_1, res_lo_lo_hi_lo_1};
  wire [127:0]  res_lo_lo_1 = {res_lo_lo_hi_1, res_lo_lo_lo_1};
  wire [15:0]   res_lo_hi_lo_lo_lo_1 = {dataGroup_17_1, dataGroup_16_1};
  wire [15:0]   res_lo_hi_lo_lo_hi_1 = {dataGroup_19_1, dataGroup_18_1};
  wire [31:0]   res_lo_hi_lo_lo_1 = {res_lo_hi_lo_lo_hi_1, res_lo_hi_lo_lo_lo_1};
  wire [15:0]   res_lo_hi_lo_hi_lo_1 = {dataGroup_21_1, dataGroup_20_1};
  wire [15:0]   res_lo_hi_lo_hi_hi_1 = {dataGroup_23_1, dataGroup_22_1};
  wire [31:0]   res_lo_hi_lo_hi_1 = {res_lo_hi_lo_hi_hi_1, res_lo_hi_lo_hi_lo_1};
  wire [63:0]   res_lo_hi_lo_1 = {res_lo_hi_lo_hi_1, res_lo_hi_lo_lo_1};
  wire [15:0]   res_lo_hi_hi_lo_lo_1 = {dataGroup_25_1, dataGroup_24_1};
  wire [15:0]   res_lo_hi_hi_lo_hi_1 = {dataGroup_27_1, dataGroup_26_1};
  wire [31:0]   res_lo_hi_hi_lo_1 = {res_lo_hi_hi_lo_hi_1, res_lo_hi_hi_lo_lo_1};
  wire [15:0]   res_lo_hi_hi_hi_lo_1 = {dataGroup_29_1, dataGroup_28_1};
  wire [15:0]   res_lo_hi_hi_hi_hi_1 = {dataGroup_31_1, dataGroup_30_1};
  wire [31:0]   res_lo_hi_hi_hi_1 = {res_lo_hi_hi_hi_hi_1, res_lo_hi_hi_hi_lo_1};
  wire [63:0]   res_lo_hi_hi_1 = {res_lo_hi_hi_hi_1, res_lo_hi_hi_lo_1};
  wire [127:0]  res_lo_hi_1 = {res_lo_hi_hi_1, res_lo_hi_lo_1};
  wire [255:0]  res_lo_1 = {res_lo_hi_1, res_lo_lo_1};
  wire [15:0]   res_hi_lo_lo_lo_lo_1 = {dataGroup_33_1, dataGroup_32_1};
  wire [15:0]   res_hi_lo_lo_lo_hi_1 = {dataGroup_35_1, dataGroup_34_1};
  wire [31:0]   res_hi_lo_lo_lo_1 = {res_hi_lo_lo_lo_hi_1, res_hi_lo_lo_lo_lo_1};
  wire [15:0]   res_hi_lo_lo_hi_lo_1 = {dataGroup_37_1, dataGroup_36_1};
  wire [15:0]   res_hi_lo_lo_hi_hi_1 = {dataGroup_39_1, dataGroup_38_1};
  wire [31:0]   res_hi_lo_lo_hi_1 = {res_hi_lo_lo_hi_hi_1, res_hi_lo_lo_hi_lo_1};
  wire [63:0]   res_hi_lo_lo_1 = {res_hi_lo_lo_hi_1, res_hi_lo_lo_lo_1};
  wire [15:0]   res_hi_lo_hi_lo_lo_1 = {dataGroup_41_1, dataGroup_40_1};
  wire [15:0]   res_hi_lo_hi_lo_hi_1 = {dataGroup_43_1, dataGroup_42_1};
  wire [31:0]   res_hi_lo_hi_lo_1 = {res_hi_lo_hi_lo_hi_1, res_hi_lo_hi_lo_lo_1};
  wire [15:0]   res_hi_lo_hi_hi_lo_1 = {dataGroup_45_1, dataGroup_44_1};
  wire [15:0]   res_hi_lo_hi_hi_hi_1 = {dataGroup_47_1, dataGroup_46_1};
  wire [31:0]   res_hi_lo_hi_hi_1 = {res_hi_lo_hi_hi_hi_1, res_hi_lo_hi_hi_lo_1};
  wire [63:0]   res_hi_lo_hi_1 = {res_hi_lo_hi_hi_1, res_hi_lo_hi_lo_1};
  wire [127:0]  res_hi_lo_1 = {res_hi_lo_hi_1, res_hi_lo_lo_1};
  wire [15:0]   res_hi_hi_lo_lo_lo_1 = {dataGroup_49_1, dataGroup_48_1};
  wire [15:0]   res_hi_hi_lo_lo_hi_1 = {dataGroup_51_1, dataGroup_50_1};
  wire [31:0]   res_hi_hi_lo_lo_1 = {res_hi_hi_lo_lo_hi_1, res_hi_hi_lo_lo_lo_1};
  wire [15:0]   res_hi_hi_lo_hi_lo_1 = {dataGroup_53_1, dataGroup_52_1};
  wire [15:0]   res_hi_hi_lo_hi_hi_1 = {dataGroup_55_1, dataGroup_54_1};
  wire [31:0]   res_hi_hi_lo_hi_1 = {res_hi_hi_lo_hi_hi_1, res_hi_hi_lo_hi_lo_1};
  wire [63:0]   res_hi_hi_lo_1 = {res_hi_hi_lo_hi_1, res_hi_hi_lo_lo_1};
  wire [15:0]   res_hi_hi_hi_lo_lo_1 = {dataGroup_57_1, dataGroup_56_1};
  wire [15:0]   res_hi_hi_hi_lo_hi_1 = {dataGroup_59_1, dataGroup_58_1};
  wire [31:0]   res_hi_hi_hi_lo_1 = {res_hi_hi_hi_lo_hi_1, res_hi_hi_hi_lo_lo_1};
  wire [15:0]   res_hi_hi_hi_hi_lo_1 = {dataGroup_61_1, dataGroup_60_1};
  wire [15:0]   res_hi_hi_hi_hi_hi_1 = {dataGroup_63_1, dataGroup_62_1};
  wire [31:0]   res_hi_hi_hi_hi_1 = {res_hi_hi_hi_hi_hi_1, res_hi_hi_hi_hi_lo_1};
  wire [63:0]   res_hi_hi_hi_1 = {res_hi_hi_hi_hi_1, res_hi_hi_hi_lo_1};
  wire [127:0]  res_hi_hi_1 = {res_hi_hi_hi_1, res_hi_hi_lo_1};
  wire [255:0]  res_hi_1 = {res_hi_hi_1, res_hi_lo_1};
  wire [511:0]  res_8 = {res_hi_1, res_lo_1};
  wire [2047:0] dataGroup_lo_128 = {dataGroup_lo_hi_128, dataGroup_lo_lo_128};
  wire [2047:0] dataGroup_hi_128 = {dataGroup_hi_hi_128, dataGroup_hi_lo_128};
  wire [7:0]    dataGroup_0_2 = dataGroup_lo_128[15:8];
  wire [2047:0] dataGroup_lo_129 = {dataGroup_lo_hi_129, dataGroup_lo_lo_129};
  wire [2047:0] dataGroup_hi_129 = {dataGroup_hi_hi_129, dataGroup_hi_lo_129};
  wire [7:0]    dataGroup_1_2 = dataGroup_lo_129[31:24];
  wire [2047:0] dataGroup_lo_130 = {dataGroup_lo_hi_130, dataGroup_lo_lo_130};
  wire [2047:0] dataGroup_hi_130 = {dataGroup_hi_hi_130, dataGroup_hi_lo_130};
  wire [7:0]    dataGroup_2_2 = dataGroup_lo_130[47:40];
  wire [2047:0] dataGroup_lo_131 = {dataGroup_lo_hi_131, dataGroup_lo_lo_131};
  wire [2047:0] dataGroup_hi_131 = {dataGroup_hi_hi_131, dataGroup_hi_lo_131};
  wire [7:0]    dataGroup_3_2 = dataGroup_lo_131[63:56];
  wire [2047:0] dataGroup_lo_132 = {dataGroup_lo_hi_132, dataGroup_lo_lo_132};
  wire [2047:0] dataGroup_hi_132 = {dataGroup_hi_hi_132, dataGroup_hi_lo_132};
  wire [7:0]    dataGroup_4_2 = dataGroup_lo_132[79:72];
  wire [2047:0] dataGroup_lo_133 = {dataGroup_lo_hi_133, dataGroup_lo_lo_133};
  wire [2047:0] dataGroup_hi_133 = {dataGroup_hi_hi_133, dataGroup_hi_lo_133};
  wire [7:0]    dataGroup_5_2 = dataGroup_lo_133[95:88];
  wire [2047:0] dataGroup_lo_134 = {dataGroup_lo_hi_134, dataGroup_lo_lo_134};
  wire [2047:0] dataGroup_hi_134 = {dataGroup_hi_hi_134, dataGroup_hi_lo_134};
  wire [7:0]    dataGroup_6_2 = dataGroup_lo_134[111:104];
  wire [2047:0] dataGroup_lo_135 = {dataGroup_lo_hi_135, dataGroup_lo_lo_135};
  wire [2047:0] dataGroup_hi_135 = {dataGroup_hi_hi_135, dataGroup_hi_lo_135};
  wire [7:0]    dataGroup_7_2 = dataGroup_lo_135[127:120];
  wire [2047:0] dataGroup_lo_136 = {dataGroup_lo_hi_136, dataGroup_lo_lo_136};
  wire [2047:0] dataGroup_hi_136 = {dataGroup_hi_hi_136, dataGroup_hi_lo_136};
  wire [7:0]    dataGroup_8_2 = dataGroup_lo_136[143:136];
  wire [2047:0] dataGroup_lo_137 = {dataGroup_lo_hi_137, dataGroup_lo_lo_137};
  wire [2047:0] dataGroup_hi_137 = {dataGroup_hi_hi_137, dataGroup_hi_lo_137};
  wire [7:0]    dataGroup_9_2 = dataGroup_lo_137[159:152];
  wire [2047:0] dataGroup_lo_138 = {dataGroup_lo_hi_138, dataGroup_lo_lo_138};
  wire [2047:0] dataGroup_hi_138 = {dataGroup_hi_hi_138, dataGroup_hi_lo_138};
  wire [7:0]    dataGroup_10_2 = dataGroup_lo_138[175:168];
  wire [2047:0] dataGroup_lo_139 = {dataGroup_lo_hi_139, dataGroup_lo_lo_139};
  wire [2047:0] dataGroup_hi_139 = {dataGroup_hi_hi_139, dataGroup_hi_lo_139};
  wire [7:0]    dataGroup_11_2 = dataGroup_lo_139[191:184];
  wire [2047:0] dataGroup_lo_140 = {dataGroup_lo_hi_140, dataGroup_lo_lo_140};
  wire [2047:0] dataGroup_hi_140 = {dataGroup_hi_hi_140, dataGroup_hi_lo_140};
  wire [7:0]    dataGroup_12_2 = dataGroup_lo_140[207:200];
  wire [2047:0] dataGroup_lo_141 = {dataGroup_lo_hi_141, dataGroup_lo_lo_141};
  wire [2047:0] dataGroup_hi_141 = {dataGroup_hi_hi_141, dataGroup_hi_lo_141};
  wire [7:0]    dataGroup_13_2 = dataGroup_lo_141[223:216];
  wire [2047:0] dataGroup_lo_142 = {dataGroup_lo_hi_142, dataGroup_lo_lo_142};
  wire [2047:0] dataGroup_hi_142 = {dataGroup_hi_hi_142, dataGroup_hi_lo_142};
  wire [7:0]    dataGroup_14_2 = dataGroup_lo_142[239:232];
  wire [2047:0] dataGroup_lo_143 = {dataGroup_lo_hi_143, dataGroup_lo_lo_143};
  wire [2047:0] dataGroup_hi_143 = {dataGroup_hi_hi_143, dataGroup_hi_lo_143};
  wire [7:0]    dataGroup_15_2 = dataGroup_lo_143[255:248];
  wire [2047:0] dataGroup_lo_144 = {dataGroup_lo_hi_144, dataGroup_lo_lo_144};
  wire [2047:0] dataGroup_hi_144 = {dataGroup_hi_hi_144, dataGroup_hi_lo_144};
  wire [7:0]    dataGroup_16_2 = dataGroup_lo_144[271:264];
  wire [2047:0] dataGroup_lo_145 = {dataGroup_lo_hi_145, dataGroup_lo_lo_145};
  wire [2047:0] dataGroup_hi_145 = {dataGroup_hi_hi_145, dataGroup_hi_lo_145};
  wire [7:0]    dataGroup_17_2 = dataGroup_lo_145[287:280];
  wire [2047:0] dataGroup_lo_146 = {dataGroup_lo_hi_146, dataGroup_lo_lo_146};
  wire [2047:0] dataGroup_hi_146 = {dataGroup_hi_hi_146, dataGroup_hi_lo_146};
  wire [7:0]    dataGroup_18_2 = dataGroup_lo_146[303:296];
  wire [2047:0] dataGroup_lo_147 = {dataGroup_lo_hi_147, dataGroup_lo_lo_147};
  wire [2047:0] dataGroup_hi_147 = {dataGroup_hi_hi_147, dataGroup_hi_lo_147};
  wire [7:0]    dataGroup_19_2 = dataGroup_lo_147[319:312];
  wire [2047:0] dataGroup_lo_148 = {dataGroup_lo_hi_148, dataGroup_lo_lo_148};
  wire [2047:0] dataGroup_hi_148 = {dataGroup_hi_hi_148, dataGroup_hi_lo_148};
  wire [7:0]    dataGroup_20_2 = dataGroup_lo_148[335:328];
  wire [2047:0] dataGroup_lo_149 = {dataGroup_lo_hi_149, dataGroup_lo_lo_149};
  wire [2047:0] dataGroup_hi_149 = {dataGroup_hi_hi_149, dataGroup_hi_lo_149};
  wire [7:0]    dataGroup_21_2 = dataGroup_lo_149[351:344];
  wire [2047:0] dataGroup_lo_150 = {dataGroup_lo_hi_150, dataGroup_lo_lo_150};
  wire [2047:0] dataGroup_hi_150 = {dataGroup_hi_hi_150, dataGroup_hi_lo_150};
  wire [7:0]    dataGroup_22_2 = dataGroup_lo_150[367:360];
  wire [2047:0] dataGroup_lo_151 = {dataGroup_lo_hi_151, dataGroup_lo_lo_151};
  wire [2047:0] dataGroup_hi_151 = {dataGroup_hi_hi_151, dataGroup_hi_lo_151};
  wire [7:0]    dataGroup_23_2 = dataGroup_lo_151[383:376];
  wire [2047:0] dataGroup_lo_152 = {dataGroup_lo_hi_152, dataGroup_lo_lo_152};
  wire [2047:0] dataGroup_hi_152 = {dataGroup_hi_hi_152, dataGroup_hi_lo_152};
  wire [7:0]    dataGroup_24_2 = dataGroup_lo_152[399:392];
  wire [2047:0] dataGroup_lo_153 = {dataGroup_lo_hi_153, dataGroup_lo_lo_153};
  wire [2047:0] dataGroup_hi_153 = {dataGroup_hi_hi_153, dataGroup_hi_lo_153};
  wire [7:0]    dataGroup_25_2 = dataGroup_lo_153[415:408];
  wire [2047:0] dataGroup_lo_154 = {dataGroup_lo_hi_154, dataGroup_lo_lo_154};
  wire [2047:0] dataGroup_hi_154 = {dataGroup_hi_hi_154, dataGroup_hi_lo_154};
  wire [7:0]    dataGroup_26_2 = dataGroup_lo_154[431:424];
  wire [2047:0] dataGroup_lo_155 = {dataGroup_lo_hi_155, dataGroup_lo_lo_155};
  wire [2047:0] dataGroup_hi_155 = {dataGroup_hi_hi_155, dataGroup_hi_lo_155};
  wire [7:0]    dataGroup_27_2 = dataGroup_lo_155[447:440];
  wire [2047:0] dataGroup_lo_156 = {dataGroup_lo_hi_156, dataGroup_lo_lo_156};
  wire [2047:0] dataGroup_hi_156 = {dataGroup_hi_hi_156, dataGroup_hi_lo_156};
  wire [7:0]    dataGroup_28_2 = dataGroup_lo_156[463:456];
  wire [2047:0] dataGroup_lo_157 = {dataGroup_lo_hi_157, dataGroup_lo_lo_157};
  wire [2047:0] dataGroup_hi_157 = {dataGroup_hi_hi_157, dataGroup_hi_lo_157};
  wire [7:0]    dataGroup_29_2 = dataGroup_lo_157[479:472];
  wire [2047:0] dataGroup_lo_158 = {dataGroup_lo_hi_158, dataGroup_lo_lo_158};
  wire [2047:0] dataGroup_hi_158 = {dataGroup_hi_hi_158, dataGroup_hi_lo_158};
  wire [7:0]    dataGroup_30_2 = dataGroup_lo_158[495:488];
  wire [2047:0] dataGroup_lo_159 = {dataGroup_lo_hi_159, dataGroup_lo_lo_159};
  wire [2047:0] dataGroup_hi_159 = {dataGroup_hi_hi_159, dataGroup_hi_lo_159};
  wire [7:0]    dataGroup_31_2 = dataGroup_lo_159[511:504];
  wire [2047:0] dataGroup_lo_160 = {dataGroup_lo_hi_160, dataGroup_lo_lo_160};
  wire [2047:0] dataGroup_hi_160 = {dataGroup_hi_hi_160, dataGroup_hi_lo_160};
  wire [7:0]    dataGroup_32_2 = dataGroup_lo_160[527:520];
  wire [2047:0] dataGroup_lo_161 = {dataGroup_lo_hi_161, dataGroup_lo_lo_161};
  wire [2047:0] dataGroup_hi_161 = {dataGroup_hi_hi_161, dataGroup_hi_lo_161};
  wire [7:0]    dataGroup_33_2 = dataGroup_lo_161[543:536];
  wire [2047:0] dataGroup_lo_162 = {dataGroup_lo_hi_162, dataGroup_lo_lo_162};
  wire [2047:0] dataGroup_hi_162 = {dataGroup_hi_hi_162, dataGroup_hi_lo_162};
  wire [7:0]    dataGroup_34_2 = dataGroup_lo_162[559:552];
  wire [2047:0] dataGroup_lo_163 = {dataGroup_lo_hi_163, dataGroup_lo_lo_163};
  wire [2047:0] dataGroup_hi_163 = {dataGroup_hi_hi_163, dataGroup_hi_lo_163};
  wire [7:0]    dataGroup_35_2 = dataGroup_lo_163[575:568];
  wire [2047:0] dataGroup_lo_164 = {dataGroup_lo_hi_164, dataGroup_lo_lo_164};
  wire [2047:0] dataGroup_hi_164 = {dataGroup_hi_hi_164, dataGroup_hi_lo_164};
  wire [7:0]    dataGroup_36_2 = dataGroup_lo_164[591:584];
  wire [2047:0] dataGroup_lo_165 = {dataGroup_lo_hi_165, dataGroup_lo_lo_165};
  wire [2047:0] dataGroup_hi_165 = {dataGroup_hi_hi_165, dataGroup_hi_lo_165};
  wire [7:0]    dataGroup_37_2 = dataGroup_lo_165[607:600];
  wire [2047:0] dataGroup_lo_166 = {dataGroup_lo_hi_166, dataGroup_lo_lo_166};
  wire [2047:0] dataGroup_hi_166 = {dataGroup_hi_hi_166, dataGroup_hi_lo_166};
  wire [7:0]    dataGroup_38_2 = dataGroup_lo_166[623:616];
  wire [2047:0] dataGroup_lo_167 = {dataGroup_lo_hi_167, dataGroup_lo_lo_167};
  wire [2047:0] dataGroup_hi_167 = {dataGroup_hi_hi_167, dataGroup_hi_lo_167};
  wire [7:0]    dataGroup_39_2 = dataGroup_lo_167[639:632];
  wire [2047:0] dataGroup_lo_168 = {dataGroup_lo_hi_168, dataGroup_lo_lo_168};
  wire [2047:0] dataGroup_hi_168 = {dataGroup_hi_hi_168, dataGroup_hi_lo_168};
  wire [7:0]    dataGroup_40_2 = dataGroup_lo_168[655:648];
  wire [2047:0] dataGroup_lo_169 = {dataGroup_lo_hi_169, dataGroup_lo_lo_169};
  wire [2047:0] dataGroup_hi_169 = {dataGroup_hi_hi_169, dataGroup_hi_lo_169};
  wire [7:0]    dataGroup_41_2 = dataGroup_lo_169[671:664];
  wire [2047:0] dataGroup_lo_170 = {dataGroup_lo_hi_170, dataGroup_lo_lo_170};
  wire [2047:0] dataGroup_hi_170 = {dataGroup_hi_hi_170, dataGroup_hi_lo_170};
  wire [7:0]    dataGroup_42_2 = dataGroup_lo_170[687:680];
  wire [2047:0] dataGroup_lo_171 = {dataGroup_lo_hi_171, dataGroup_lo_lo_171};
  wire [2047:0] dataGroup_hi_171 = {dataGroup_hi_hi_171, dataGroup_hi_lo_171};
  wire [7:0]    dataGroup_43_2 = dataGroup_lo_171[703:696];
  wire [2047:0] dataGroup_lo_172 = {dataGroup_lo_hi_172, dataGroup_lo_lo_172};
  wire [2047:0] dataGroup_hi_172 = {dataGroup_hi_hi_172, dataGroup_hi_lo_172};
  wire [7:0]    dataGroup_44_2 = dataGroup_lo_172[719:712];
  wire [2047:0] dataGroup_lo_173 = {dataGroup_lo_hi_173, dataGroup_lo_lo_173};
  wire [2047:0] dataGroup_hi_173 = {dataGroup_hi_hi_173, dataGroup_hi_lo_173};
  wire [7:0]    dataGroup_45_2 = dataGroup_lo_173[735:728];
  wire [2047:0] dataGroup_lo_174 = {dataGroup_lo_hi_174, dataGroup_lo_lo_174};
  wire [2047:0] dataGroup_hi_174 = {dataGroup_hi_hi_174, dataGroup_hi_lo_174};
  wire [7:0]    dataGroup_46_2 = dataGroup_lo_174[751:744];
  wire [2047:0] dataGroup_lo_175 = {dataGroup_lo_hi_175, dataGroup_lo_lo_175};
  wire [2047:0] dataGroup_hi_175 = {dataGroup_hi_hi_175, dataGroup_hi_lo_175};
  wire [7:0]    dataGroup_47_2 = dataGroup_lo_175[767:760];
  wire [2047:0] dataGroup_lo_176 = {dataGroup_lo_hi_176, dataGroup_lo_lo_176};
  wire [2047:0] dataGroup_hi_176 = {dataGroup_hi_hi_176, dataGroup_hi_lo_176};
  wire [7:0]    dataGroup_48_2 = dataGroup_lo_176[783:776];
  wire [2047:0] dataGroup_lo_177 = {dataGroup_lo_hi_177, dataGroup_lo_lo_177};
  wire [2047:0] dataGroup_hi_177 = {dataGroup_hi_hi_177, dataGroup_hi_lo_177};
  wire [7:0]    dataGroup_49_2 = dataGroup_lo_177[799:792];
  wire [2047:0] dataGroup_lo_178 = {dataGroup_lo_hi_178, dataGroup_lo_lo_178};
  wire [2047:0] dataGroup_hi_178 = {dataGroup_hi_hi_178, dataGroup_hi_lo_178};
  wire [7:0]    dataGroup_50_2 = dataGroup_lo_178[815:808];
  wire [2047:0] dataGroup_lo_179 = {dataGroup_lo_hi_179, dataGroup_lo_lo_179};
  wire [2047:0] dataGroup_hi_179 = {dataGroup_hi_hi_179, dataGroup_hi_lo_179};
  wire [7:0]    dataGroup_51_2 = dataGroup_lo_179[831:824];
  wire [2047:0] dataGroup_lo_180 = {dataGroup_lo_hi_180, dataGroup_lo_lo_180};
  wire [2047:0] dataGroup_hi_180 = {dataGroup_hi_hi_180, dataGroup_hi_lo_180};
  wire [7:0]    dataGroup_52_2 = dataGroup_lo_180[847:840];
  wire [2047:0] dataGroup_lo_181 = {dataGroup_lo_hi_181, dataGroup_lo_lo_181};
  wire [2047:0] dataGroup_hi_181 = {dataGroup_hi_hi_181, dataGroup_hi_lo_181};
  wire [7:0]    dataGroup_53_2 = dataGroup_lo_181[863:856];
  wire [2047:0] dataGroup_lo_182 = {dataGroup_lo_hi_182, dataGroup_lo_lo_182};
  wire [2047:0] dataGroup_hi_182 = {dataGroup_hi_hi_182, dataGroup_hi_lo_182};
  wire [7:0]    dataGroup_54_2 = dataGroup_lo_182[879:872];
  wire [2047:0] dataGroup_lo_183 = {dataGroup_lo_hi_183, dataGroup_lo_lo_183};
  wire [2047:0] dataGroup_hi_183 = {dataGroup_hi_hi_183, dataGroup_hi_lo_183};
  wire [7:0]    dataGroup_55_2 = dataGroup_lo_183[895:888];
  wire [2047:0] dataGroup_lo_184 = {dataGroup_lo_hi_184, dataGroup_lo_lo_184};
  wire [2047:0] dataGroup_hi_184 = {dataGroup_hi_hi_184, dataGroup_hi_lo_184};
  wire [7:0]    dataGroup_56_2 = dataGroup_lo_184[911:904];
  wire [2047:0] dataGroup_lo_185 = {dataGroup_lo_hi_185, dataGroup_lo_lo_185};
  wire [2047:0] dataGroup_hi_185 = {dataGroup_hi_hi_185, dataGroup_hi_lo_185};
  wire [7:0]    dataGroup_57_2 = dataGroup_lo_185[927:920];
  wire [2047:0] dataGroup_lo_186 = {dataGroup_lo_hi_186, dataGroup_lo_lo_186};
  wire [2047:0] dataGroup_hi_186 = {dataGroup_hi_hi_186, dataGroup_hi_lo_186};
  wire [7:0]    dataGroup_58_2 = dataGroup_lo_186[943:936];
  wire [2047:0] dataGroup_lo_187 = {dataGroup_lo_hi_187, dataGroup_lo_lo_187};
  wire [2047:0] dataGroup_hi_187 = {dataGroup_hi_hi_187, dataGroup_hi_lo_187};
  wire [7:0]    dataGroup_59_2 = dataGroup_lo_187[959:952];
  wire [2047:0] dataGroup_lo_188 = {dataGroup_lo_hi_188, dataGroup_lo_lo_188};
  wire [2047:0] dataGroup_hi_188 = {dataGroup_hi_hi_188, dataGroup_hi_lo_188};
  wire [7:0]    dataGroup_60_2 = dataGroup_lo_188[975:968];
  wire [2047:0] dataGroup_lo_189 = {dataGroup_lo_hi_189, dataGroup_lo_lo_189};
  wire [2047:0] dataGroup_hi_189 = {dataGroup_hi_hi_189, dataGroup_hi_lo_189};
  wire [7:0]    dataGroup_61_2 = dataGroup_lo_189[991:984];
  wire [2047:0] dataGroup_lo_190 = {dataGroup_lo_hi_190, dataGroup_lo_lo_190};
  wire [2047:0] dataGroup_hi_190 = {dataGroup_hi_hi_190, dataGroup_hi_lo_190};
  wire [7:0]    dataGroup_62_2 = dataGroup_lo_190[1007:1000];
  wire [2047:0] dataGroup_lo_191 = {dataGroup_lo_hi_191, dataGroup_lo_lo_191};
  wire [2047:0] dataGroup_hi_191 = {dataGroup_hi_hi_191, dataGroup_hi_lo_191};
  wire [7:0]    dataGroup_63_2 = dataGroup_lo_191[1023:1016];
  wire [15:0]   res_lo_lo_lo_lo_lo_2 = {dataGroup_1_2, dataGroup_0_2};
  wire [15:0]   res_lo_lo_lo_lo_hi_2 = {dataGroup_3_2, dataGroup_2_2};
  wire [31:0]   res_lo_lo_lo_lo_2 = {res_lo_lo_lo_lo_hi_2, res_lo_lo_lo_lo_lo_2};
  wire [15:0]   res_lo_lo_lo_hi_lo_2 = {dataGroup_5_2, dataGroup_4_2};
  wire [15:0]   res_lo_lo_lo_hi_hi_2 = {dataGroup_7_2, dataGroup_6_2};
  wire [31:0]   res_lo_lo_lo_hi_2 = {res_lo_lo_lo_hi_hi_2, res_lo_lo_lo_hi_lo_2};
  wire [63:0]   res_lo_lo_lo_2 = {res_lo_lo_lo_hi_2, res_lo_lo_lo_lo_2};
  wire [15:0]   res_lo_lo_hi_lo_lo_2 = {dataGroup_9_2, dataGroup_8_2};
  wire [15:0]   res_lo_lo_hi_lo_hi_2 = {dataGroup_11_2, dataGroup_10_2};
  wire [31:0]   res_lo_lo_hi_lo_2 = {res_lo_lo_hi_lo_hi_2, res_lo_lo_hi_lo_lo_2};
  wire [15:0]   res_lo_lo_hi_hi_lo_2 = {dataGroup_13_2, dataGroup_12_2};
  wire [15:0]   res_lo_lo_hi_hi_hi_2 = {dataGroup_15_2, dataGroup_14_2};
  wire [31:0]   res_lo_lo_hi_hi_2 = {res_lo_lo_hi_hi_hi_2, res_lo_lo_hi_hi_lo_2};
  wire [63:0]   res_lo_lo_hi_2 = {res_lo_lo_hi_hi_2, res_lo_lo_hi_lo_2};
  wire [127:0]  res_lo_lo_2 = {res_lo_lo_hi_2, res_lo_lo_lo_2};
  wire [15:0]   res_lo_hi_lo_lo_lo_2 = {dataGroup_17_2, dataGroup_16_2};
  wire [15:0]   res_lo_hi_lo_lo_hi_2 = {dataGroup_19_2, dataGroup_18_2};
  wire [31:0]   res_lo_hi_lo_lo_2 = {res_lo_hi_lo_lo_hi_2, res_lo_hi_lo_lo_lo_2};
  wire [15:0]   res_lo_hi_lo_hi_lo_2 = {dataGroup_21_2, dataGroup_20_2};
  wire [15:0]   res_lo_hi_lo_hi_hi_2 = {dataGroup_23_2, dataGroup_22_2};
  wire [31:0]   res_lo_hi_lo_hi_2 = {res_lo_hi_lo_hi_hi_2, res_lo_hi_lo_hi_lo_2};
  wire [63:0]   res_lo_hi_lo_2 = {res_lo_hi_lo_hi_2, res_lo_hi_lo_lo_2};
  wire [15:0]   res_lo_hi_hi_lo_lo_2 = {dataGroup_25_2, dataGroup_24_2};
  wire [15:0]   res_lo_hi_hi_lo_hi_2 = {dataGroup_27_2, dataGroup_26_2};
  wire [31:0]   res_lo_hi_hi_lo_2 = {res_lo_hi_hi_lo_hi_2, res_lo_hi_hi_lo_lo_2};
  wire [15:0]   res_lo_hi_hi_hi_lo_2 = {dataGroup_29_2, dataGroup_28_2};
  wire [15:0]   res_lo_hi_hi_hi_hi_2 = {dataGroup_31_2, dataGroup_30_2};
  wire [31:0]   res_lo_hi_hi_hi_2 = {res_lo_hi_hi_hi_hi_2, res_lo_hi_hi_hi_lo_2};
  wire [63:0]   res_lo_hi_hi_2 = {res_lo_hi_hi_hi_2, res_lo_hi_hi_lo_2};
  wire [127:0]  res_lo_hi_2 = {res_lo_hi_hi_2, res_lo_hi_lo_2};
  wire [255:0]  res_lo_2 = {res_lo_hi_2, res_lo_lo_2};
  wire [15:0]   res_hi_lo_lo_lo_lo_2 = {dataGroup_33_2, dataGroup_32_2};
  wire [15:0]   res_hi_lo_lo_lo_hi_2 = {dataGroup_35_2, dataGroup_34_2};
  wire [31:0]   res_hi_lo_lo_lo_2 = {res_hi_lo_lo_lo_hi_2, res_hi_lo_lo_lo_lo_2};
  wire [15:0]   res_hi_lo_lo_hi_lo_2 = {dataGroup_37_2, dataGroup_36_2};
  wire [15:0]   res_hi_lo_lo_hi_hi_2 = {dataGroup_39_2, dataGroup_38_2};
  wire [31:0]   res_hi_lo_lo_hi_2 = {res_hi_lo_lo_hi_hi_2, res_hi_lo_lo_hi_lo_2};
  wire [63:0]   res_hi_lo_lo_2 = {res_hi_lo_lo_hi_2, res_hi_lo_lo_lo_2};
  wire [15:0]   res_hi_lo_hi_lo_lo_2 = {dataGroup_41_2, dataGroup_40_2};
  wire [15:0]   res_hi_lo_hi_lo_hi_2 = {dataGroup_43_2, dataGroup_42_2};
  wire [31:0]   res_hi_lo_hi_lo_2 = {res_hi_lo_hi_lo_hi_2, res_hi_lo_hi_lo_lo_2};
  wire [15:0]   res_hi_lo_hi_hi_lo_2 = {dataGroup_45_2, dataGroup_44_2};
  wire [15:0]   res_hi_lo_hi_hi_hi_2 = {dataGroup_47_2, dataGroup_46_2};
  wire [31:0]   res_hi_lo_hi_hi_2 = {res_hi_lo_hi_hi_hi_2, res_hi_lo_hi_hi_lo_2};
  wire [63:0]   res_hi_lo_hi_2 = {res_hi_lo_hi_hi_2, res_hi_lo_hi_lo_2};
  wire [127:0]  res_hi_lo_2 = {res_hi_lo_hi_2, res_hi_lo_lo_2};
  wire [15:0]   res_hi_hi_lo_lo_lo_2 = {dataGroup_49_2, dataGroup_48_2};
  wire [15:0]   res_hi_hi_lo_lo_hi_2 = {dataGroup_51_2, dataGroup_50_2};
  wire [31:0]   res_hi_hi_lo_lo_2 = {res_hi_hi_lo_lo_hi_2, res_hi_hi_lo_lo_lo_2};
  wire [15:0]   res_hi_hi_lo_hi_lo_2 = {dataGroup_53_2, dataGroup_52_2};
  wire [15:0]   res_hi_hi_lo_hi_hi_2 = {dataGroup_55_2, dataGroup_54_2};
  wire [31:0]   res_hi_hi_lo_hi_2 = {res_hi_hi_lo_hi_hi_2, res_hi_hi_lo_hi_lo_2};
  wire [63:0]   res_hi_hi_lo_2 = {res_hi_hi_lo_hi_2, res_hi_hi_lo_lo_2};
  wire [15:0]   res_hi_hi_hi_lo_lo_2 = {dataGroup_57_2, dataGroup_56_2};
  wire [15:0]   res_hi_hi_hi_lo_hi_2 = {dataGroup_59_2, dataGroup_58_2};
  wire [31:0]   res_hi_hi_hi_lo_2 = {res_hi_hi_hi_lo_hi_2, res_hi_hi_hi_lo_lo_2};
  wire [15:0]   res_hi_hi_hi_hi_lo_2 = {dataGroup_61_2, dataGroup_60_2};
  wire [15:0]   res_hi_hi_hi_hi_hi_2 = {dataGroup_63_2, dataGroup_62_2};
  wire [31:0]   res_hi_hi_hi_hi_2 = {res_hi_hi_hi_hi_hi_2, res_hi_hi_hi_hi_lo_2};
  wire [63:0]   res_hi_hi_hi_2 = {res_hi_hi_hi_hi_2, res_hi_hi_hi_lo_2};
  wire [127:0]  res_hi_hi_2 = {res_hi_hi_hi_2, res_hi_hi_lo_2};
  wire [255:0]  res_hi_2 = {res_hi_hi_2, res_hi_lo_2};
  wire [511:0]  res_9 = {res_hi_2, res_lo_2};
  wire [1023:0] lo_lo_1 = {res_9, res_8};
  wire [2047:0] lo_1 = {1024'h0, lo_lo_1};
  wire [4095:0] regroupLoadData_0_1 = {2048'h0, lo_1};
  wire [2047:0] dataGroup_lo_192 = {dataGroup_lo_hi_192, dataGroup_lo_lo_192};
  wire [2047:0] dataGroup_hi_192 = {dataGroup_hi_hi_192, dataGroup_hi_lo_192};
  wire [7:0]    dataGroup_0_3 = dataGroup_lo_192[7:0];
  wire [2047:0] dataGroup_lo_193 = {dataGroup_lo_hi_193, dataGroup_lo_lo_193};
  wire [2047:0] dataGroup_hi_193 = {dataGroup_hi_hi_193, dataGroup_hi_lo_193};
  wire [7:0]    dataGroup_1_3 = dataGroup_lo_193[31:24];
  wire [2047:0] dataGroup_lo_194 = {dataGroup_lo_hi_194, dataGroup_lo_lo_194};
  wire [2047:0] dataGroup_hi_194 = {dataGroup_hi_hi_194, dataGroup_hi_lo_194};
  wire [7:0]    dataGroup_2_3 = dataGroup_lo_194[55:48];
  wire [2047:0] dataGroup_lo_195 = {dataGroup_lo_hi_195, dataGroup_lo_lo_195};
  wire [2047:0] dataGroup_hi_195 = {dataGroup_hi_hi_195, dataGroup_hi_lo_195};
  wire [7:0]    dataGroup_3_3 = dataGroup_lo_195[79:72];
  wire [2047:0] dataGroup_lo_196 = {dataGroup_lo_hi_196, dataGroup_lo_lo_196};
  wire [2047:0] dataGroup_hi_196 = {dataGroup_hi_hi_196, dataGroup_hi_lo_196};
  wire [7:0]    dataGroup_4_3 = dataGroup_lo_196[103:96];
  wire [2047:0] dataGroup_lo_197 = {dataGroup_lo_hi_197, dataGroup_lo_lo_197};
  wire [2047:0] dataGroup_hi_197 = {dataGroup_hi_hi_197, dataGroup_hi_lo_197};
  wire [7:0]    dataGroup_5_3 = dataGroup_lo_197[127:120];
  wire [2047:0] dataGroup_lo_198 = {dataGroup_lo_hi_198, dataGroup_lo_lo_198};
  wire [2047:0] dataGroup_hi_198 = {dataGroup_hi_hi_198, dataGroup_hi_lo_198};
  wire [7:0]    dataGroup_6_3 = dataGroup_lo_198[151:144];
  wire [2047:0] dataGroup_lo_199 = {dataGroup_lo_hi_199, dataGroup_lo_lo_199};
  wire [2047:0] dataGroup_hi_199 = {dataGroup_hi_hi_199, dataGroup_hi_lo_199};
  wire [7:0]    dataGroup_7_3 = dataGroup_lo_199[175:168];
  wire [2047:0] dataGroup_lo_200 = {dataGroup_lo_hi_200, dataGroup_lo_lo_200};
  wire [2047:0] dataGroup_hi_200 = {dataGroup_hi_hi_200, dataGroup_hi_lo_200};
  wire [7:0]    dataGroup_8_3 = dataGroup_lo_200[199:192];
  wire [2047:0] dataGroup_lo_201 = {dataGroup_lo_hi_201, dataGroup_lo_lo_201};
  wire [2047:0] dataGroup_hi_201 = {dataGroup_hi_hi_201, dataGroup_hi_lo_201};
  wire [7:0]    dataGroup_9_3 = dataGroup_lo_201[223:216];
  wire [2047:0] dataGroup_lo_202 = {dataGroup_lo_hi_202, dataGroup_lo_lo_202};
  wire [2047:0] dataGroup_hi_202 = {dataGroup_hi_hi_202, dataGroup_hi_lo_202};
  wire [7:0]    dataGroup_10_3 = dataGroup_lo_202[247:240];
  wire [2047:0] dataGroup_lo_203 = {dataGroup_lo_hi_203, dataGroup_lo_lo_203};
  wire [2047:0] dataGroup_hi_203 = {dataGroup_hi_hi_203, dataGroup_hi_lo_203};
  wire [7:0]    dataGroup_11_3 = dataGroup_lo_203[271:264];
  wire [2047:0] dataGroup_lo_204 = {dataGroup_lo_hi_204, dataGroup_lo_lo_204};
  wire [2047:0] dataGroup_hi_204 = {dataGroup_hi_hi_204, dataGroup_hi_lo_204};
  wire [7:0]    dataGroup_12_3 = dataGroup_lo_204[295:288];
  wire [2047:0] dataGroup_lo_205 = {dataGroup_lo_hi_205, dataGroup_lo_lo_205};
  wire [2047:0] dataGroup_hi_205 = {dataGroup_hi_hi_205, dataGroup_hi_lo_205};
  wire [7:0]    dataGroup_13_3 = dataGroup_lo_205[319:312];
  wire [2047:0] dataGroup_lo_206 = {dataGroup_lo_hi_206, dataGroup_lo_lo_206};
  wire [2047:0] dataGroup_hi_206 = {dataGroup_hi_hi_206, dataGroup_hi_lo_206};
  wire [7:0]    dataGroup_14_3 = dataGroup_lo_206[343:336];
  wire [2047:0] dataGroup_lo_207 = {dataGroup_lo_hi_207, dataGroup_lo_lo_207};
  wire [2047:0] dataGroup_hi_207 = {dataGroup_hi_hi_207, dataGroup_hi_lo_207};
  wire [7:0]    dataGroup_15_3 = dataGroup_lo_207[367:360];
  wire [2047:0] dataGroup_lo_208 = {dataGroup_lo_hi_208, dataGroup_lo_lo_208};
  wire [2047:0] dataGroup_hi_208 = {dataGroup_hi_hi_208, dataGroup_hi_lo_208};
  wire [7:0]    dataGroup_16_3 = dataGroup_lo_208[391:384];
  wire [2047:0] dataGroup_lo_209 = {dataGroup_lo_hi_209, dataGroup_lo_lo_209};
  wire [2047:0] dataGroup_hi_209 = {dataGroup_hi_hi_209, dataGroup_hi_lo_209};
  wire [7:0]    dataGroup_17_3 = dataGroup_lo_209[415:408];
  wire [2047:0] dataGroup_lo_210 = {dataGroup_lo_hi_210, dataGroup_lo_lo_210};
  wire [2047:0] dataGroup_hi_210 = {dataGroup_hi_hi_210, dataGroup_hi_lo_210};
  wire [7:0]    dataGroup_18_3 = dataGroup_lo_210[439:432];
  wire [2047:0] dataGroup_lo_211 = {dataGroup_lo_hi_211, dataGroup_lo_lo_211};
  wire [2047:0] dataGroup_hi_211 = {dataGroup_hi_hi_211, dataGroup_hi_lo_211};
  wire [7:0]    dataGroup_19_3 = dataGroup_lo_211[463:456];
  wire [2047:0] dataGroup_lo_212 = {dataGroup_lo_hi_212, dataGroup_lo_lo_212};
  wire [2047:0] dataGroup_hi_212 = {dataGroup_hi_hi_212, dataGroup_hi_lo_212};
  wire [7:0]    dataGroup_20_3 = dataGroup_lo_212[487:480];
  wire [2047:0] dataGroup_lo_213 = {dataGroup_lo_hi_213, dataGroup_lo_lo_213};
  wire [2047:0] dataGroup_hi_213 = {dataGroup_hi_hi_213, dataGroup_hi_lo_213};
  wire [7:0]    dataGroup_21_3 = dataGroup_lo_213[511:504];
  wire [2047:0] dataGroup_lo_214 = {dataGroup_lo_hi_214, dataGroup_lo_lo_214};
  wire [2047:0] dataGroup_hi_214 = {dataGroup_hi_hi_214, dataGroup_hi_lo_214};
  wire [7:0]    dataGroup_22_3 = dataGroup_lo_214[535:528];
  wire [2047:0] dataGroup_lo_215 = {dataGroup_lo_hi_215, dataGroup_lo_lo_215};
  wire [2047:0] dataGroup_hi_215 = {dataGroup_hi_hi_215, dataGroup_hi_lo_215};
  wire [7:0]    dataGroup_23_3 = dataGroup_lo_215[559:552];
  wire [2047:0] dataGroup_lo_216 = {dataGroup_lo_hi_216, dataGroup_lo_lo_216};
  wire [2047:0] dataGroup_hi_216 = {dataGroup_hi_hi_216, dataGroup_hi_lo_216};
  wire [7:0]    dataGroup_24_3 = dataGroup_lo_216[583:576];
  wire [2047:0] dataGroup_lo_217 = {dataGroup_lo_hi_217, dataGroup_lo_lo_217};
  wire [2047:0] dataGroup_hi_217 = {dataGroup_hi_hi_217, dataGroup_hi_lo_217};
  wire [7:0]    dataGroup_25_3 = dataGroup_lo_217[607:600];
  wire [2047:0] dataGroup_lo_218 = {dataGroup_lo_hi_218, dataGroup_lo_lo_218};
  wire [2047:0] dataGroup_hi_218 = {dataGroup_hi_hi_218, dataGroup_hi_lo_218};
  wire [7:0]    dataGroup_26_3 = dataGroup_lo_218[631:624];
  wire [2047:0] dataGroup_lo_219 = {dataGroup_lo_hi_219, dataGroup_lo_lo_219};
  wire [2047:0] dataGroup_hi_219 = {dataGroup_hi_hi_219, dataGroup_hi_lo_219};
  wire [7:0]    dataGroup_27_3 = dataGroup_lo_219[655:648];
  wire [2047:0] dataGroup_lo_220 = {dataGroup_lo_hi_220, dataGroup_lo_lo_220};
  wire [2047:0] dataGroup_hi_220 = {dataGroup_hi_hi_220, dataGroup_hi_lo_220};
  wire [7:0]    dataGroup_28_3 = dataGroup_lo_220[679:672];
  wire [2047:0] dataGroup_lo_221 = {dataGroup_lo_hi_221, dataGroup_lo_lo_221};
  wire [2047:0] dataGroup_hi_221 = {dataGroup_hi_hi_221, dataGroup_hi_lo_221};
  wire [7:0]    dataGroup_29_3 = dataGroup_lo_221[703:696];
  wire [2047:0] dataGroup_lo_222 = {dataGroup_lo_hi_222, dataGroup_lo_lo_222};
  wire [2047:0] dataGroup_hi_222 = {dataGroup_hi_hi_222, dataGroup_hi_lo_222};
  wire [7:0]    dataGroup_30_3 = dataGroup_lo_222[727:720];
  wire [2047:0] dataGroup_lo_223 = {dataGroup_lo_hi_223, dataGroup_lo_lo_223};
  wire [2047:0] dataGroup_hi_223 = {dataGroup_hi_hi_223, dataGroup_hi_lo_223};
  wire [7:0]    dataGroup_31_3 = dataGroup_lo_223[751:744];
  wire [2047:0] dataGroup_lo_224 = {dataGroup_lo_hi_224, dataGroup_lo_lo_224};
  wire [2047:0] dataGroup_hi_224 = {dataGroup_hi_hi_224, dataGroup_hi_lo_224};
  wire [7:0]    dataGroup_32_3 = dataGroup_lo_224[775:768];
  wire [2047:0] dataGroup_lo_225 = {dataGroup_lo_hi_225, dataGroup_lo_lo_225};
  wire [2047:0] dataGroup_hi_225 = {dataGroup_hi_hi_225, dataGroup_hi_lo_225};
  wire [7:0]    dataGroup_33_3 = dataGroup_lo_225[799:792];
  wire [2047:0] dataGroup_lo_226 = {dataGroup_lo_hi_226, dataGroup_lo_lo_226};
  wire [2047:0] dataGroup_hi_226 = {dataGroup_hi_hi_226, dataGroup_hi_lo_226};
  wire [7:0]    dataGroup_34_3 = dataGroup_lo_226[823:816];
  wire [2047:0] dataGroup_lo_227 = {dataGroup_lo_hi_227, dataGroup_lo_lo_227};
  wire [2047:0] dataGroup_hi_227 = {dataGroup_hi_hi_227, dataGroup_hi_lo_227};
  wire [7:0]    dataGroup_35_3 = dataGroup_lo_227[847:840];
  wire [2047:0] dataGroup_lo_228 = {dataGroup_lo_hi_228, dataGroup_lo_lo_228};
  wire [2047:0] dataGroup_hi_228 = {dataGroup_hi_hi_228, dataGroup_hi_lo_228};
  wire [7:0]    dataGroup_36_3 = dataGroup_lo_228[871:864];
  wire [2047:0] dataGroup_lo_229 = {dataGroup_lo_hi_229, dataGroup_lo_lo_229};
  wire [2047:0] dataGroup_hi_229 = {dataGroup_hi_hi_229, dataGroup_hi_lo_229};
  wire [7:0]    dataGroup_37_3 = dataGroup_lo_229[895:888];
  wire [2047:0] dataGroup_lo_230 = {dataGroup_lo_hi_230, dataGroup_lo_lo_230};
  wire [2047:0] dataGroup_hi_230 = {dataGroup_hi_hi_230, dataGroup_hi_lo_230};
  wire [7:0]    dataGroup_38_3 = dataGroup_lo_230[919:912];
  wire [2047:0] dataGroup_lo_231 = {dataGroup_lo_hi_231, dataGroup_lo_lo_231};
  wire [2047:0] dataGroup_hi_231 = {dataGroup_hi_hi_231, dataGroup_hi_lo_231};
  wire [7:0]    dataGroup_39_3 = dataGroup_lo_231[943:936];
  wire [2047:0] dataGroup_lo_232 = {dataGroup_lo_hi_232, dataGroup_lo_lo_232};
  wire [2047:0] dataGroup_hi_232 = {dataGroup_hi_hi_232, dataGroup_hi_lo_232};
  wire [7:0]    dataGroup_40_3 = dataGroup_lo_232[967:960];
  wire [2047:0] dataGroup_lo_233 = {dataGroup_lo_hi_233, dataGroup_lo_lo_233};
  wire [2047:0] dataGroup_hi_233 = {dataGroup_hi_hi_233, dataGroup_hi_lo_233};
  wire [7:0]    dataGroup_41_3 = dataGroup_lo_233[991:984];
  wire [2047:0] dataGroup_lo_234 = {dataGroup_lo_hi_234, dataGroup_lo_lo_234};
  wire [2047:0] dataGroup_hi_234 = {dataGroup_hi_hi_234, dataGroup_hi_lo_234};
  wire [7:0]    dataGroup_42_3 = dataGroup_lo_234[1015:1008];
  wire [2047:0] dataGroup_lo_235 = {dataGroup_lo_hi_235, dataGroup_lo_lo_235};
  wire [2047:0] dataGroup_hi_235 = {dataGroup_hi_hi_235, dataGroup_hi_lo_235};
  wire [7:0]    dataGroup_43_3 = dataGroup_lo_235[1039:1032];
  wire [2047:0] dataGroup_lo_236 = {dataGroup_lo_hi_236, dataGroup_lo_lo_236};
  wire [2047:0] dataGroup_hi_236 = {dataGroup_hi_hi_236, dataGroup_hi_lo_236};
  wire [7:0]    dataGroup_44_3 = dataGroup_lo_236[1063:1056];
  wire [2047:0] dataGroup_lo_237 = {dataGroup_lo_hi_237, dataGroup_lo_lo_237};
  wire [2047:0] dataGroup_hi_237 = {dataGroup_hi_hi_237, dataGroup_hi_lo_237};
  wire [7:0]    dataGroup_45_3 = dataGroup_lo_237[1087:1080];
  wire [2047:0] dataGroup_lo_238 = {dataGroup_lo_hi_238, dataGroup_lo_lo_238};
  wire [2047:0] dataGroup_hi_238 = {dataGroup_hi_hi_238, dataGroup_hi_lo_238};
  wire [7:0]    dataGroup_46_3 = dataGroup_lo_238[1111:1104];
  wire [2047:0] dataGroup_lo_239 = {dataGroup_lo_hi_239, dataGroup_lo_lo_239};
  wire [2047:0] dataGroup_hi_239 = {dataGroup_hi_hi_239, dataGroup_hi_lo_239};
  wire [7:0]    dataGroup_47_3 = dataGroup_lo_239[1135:1128];
  wire [2047:0] dataGroup_lo_240 = {dataGroup_lo_hi_240, dataGroup_lo_lo_240};
  wire [2047:0] dataGroup_hi_240 = {dataGroup_hi_hi_240, dataGroup_hi_lo_240};
  wire [7:0]    dataGroup_48_3 = dataGroup_lo_240[1159:1152];
  wire [2047:0] dataGroup_lo_241 = {dataGroup_lo_hi_241, dataGroup_lo_lo_241};
  wire [2047:0] dataGroup_hi_241 = {dataGroup_hi_hi_241, dataGroup_hi_lo_241};
  wire [7:0]    dataGroup_49_3 = dataGroup_lo_241[1183:1176];
  wire [2047:0] dataGroup_lo_242 = {dataGroup_lo_hi_242, dataGroup_lo_lo_242};
  wire [2047:0] dataGroup_hi_242 = {dataGroup_hi_hi_242, dataGroup_hi_lo_242};
  wire [7:0]    dataGroup_50_3 = dataGroup_lo_242[1207:1200];
  wire [2047:0] dataGroup_lo_243 = {dataGroup_lo_hi_243, dataGroup_lo_lo_243};
  wire [2047:0] dataGroup_hi_243 = {dataGroup_hi_hi_243, dataGroup_hi_lo_243};
  wire [7:0]    dataGroup_51_3 = dataGroup_lo_243[1231:1224];
  wire [2047:0] dataGroup_lo_244 = {dataGroup_lo_hi_244, dataGroup_lo_lo_244};
  wire [2047:0] dataGroup_hi_244 = {dataGroup_hi_hi_244, dataGroup_hi_lo_244};
  wire [7:0]    dataGroup_52_3 = dataGroup_lo_244[1255:1248];
  wire [2047:0] dataGroup_lo_245 = {dataGroup_lo_hi_245, dataGroup_lo_lo_245};
  wire [2047:0] dataGroup_hi_245 = {dataGroup_hi_hi_245, dataGroup_hi_lo_245};
  wire [7:0]    dataGroup_53_3 = dataGroup_lo_245[1279:1272];
  wire [2047:0] dataGroup_lo_246 = {dataGroup_lo_hi_246, dataGroup_lo_lo_246};
  wire [2047:0] dataGroup_hi_246 = {dataGroup_hi_hi_246, dataGroup_hi_lo_246};
  wire [7:0]    dataGroup_54_3 = dataGroup_lo_246[1303:1296];
  wire [2047:0] dataGroup_lo_247 = {dataGroup_lo_hi_247, dataGroup_lo_lo_247};
  wire [2047:0] dataGroup_hi_247 = {dataGroup_hi_hi_247, dataGroup_hi_lo_247};
  wire [7:0]    dataGroup_55_3 = dataGroup_lo_247[1327:1320];
  wire [2047:0] dataGroup_lo_248 = {dataGroup_lo_hi_248, dataGroup_lo_lo_248};
  wire [2047:0] dataGroup_hi_248 = {dataGroup_hi_hi_248, dataGroup_hi_lo_248};
  wire [7:0]    dataGroup_56_3 = dataGroup_lo_248[1351:1344];
  wire [2047:0] dataGroup_lo_249 = {dataGroup_lo_hi_249, dataGroup_lo_lo_249};
  wire [2047:0] dataGroup_hi_249 = {dataGroup_hi_hi_249, dataGroup_hi_lo_249};
  wire [7:0]    dataGroup_57_3 = dataGroup_lo_249[1375:1368];
  wire [2047:0] dataGroup_lo_250 = {dataGroup_lo_hi_250, dataGroup_lo_lo_250};
  wire [2047:0] dataGroup_hi_250 = {dataGroup_hi_hi_250, dataGroup_hi_lo_250};
  wire [7:0]    dataGroup_58_3 = dataGroup_lo_250[1399:1392];
  wire [2047:0] dataGroup_lo_251 = {dataGroup_lo_hi_251, dataGroup_lo_lo_251};
  wire [2047:0] dataGroup_hi_251 = {dataGroup_hi_hi_251, dataGroup_hi_lo_251};
  wire [7:0]    dataGroup_59_3 = dataGroup_lo_251[1423:1416];
  wire [2047:0] dataGroup_lo_252 = {dataGroup_lo_hi_252, dataGroup_lo_lo_252};
  wire [2047:0] dataGroup_hi_252 = {dataGroup_hi_hi_252, dataGroup_hi_lo_252};
  wire [7:0]    dataGroup_60_3 = dataGroup_lo_252[1447:1440];
  wire [2047:0] dataGroup_lo_253 = {dataGroup_lo_hi_253, dataGroup_lo_lo_253};
  wire [2047:0] dataGroup_hi_253 = {dataGroup_hi_hi_253, dataGroup_hi_lo_253};
  wire [7:0]    dataGroup_61_3 = dataGroup_lo_253[1471:1464];
  wire [2047:0] dataGroup_lo_254 = {dataGroup_lo_hi_254, dataGroup_lo_lo_254};
  wire [2047:0] dataGroup_hi_254 = {dataGroup_hi_hi_254, dataGroup_hi_lo_254};
  wire [7:0]    dataGroup_62_3 = dataGroup_lo_254[1495:1488];
  wire [2047:0] dataGroup_lo_255 = {dataGroup_lo_hi_255, dataGroup_lo_lo_255};
  wire [2047:0] dataGroup_hi_255 = {dataGroup_hi_hi_255, dataGroup_hi_lo_255};
  wire [7:0]    dataGroup_63_3 = dataGroup_lo_255[1519:1512];
  wire [15:0]   res_lo_lo_lo_lo_lo_3 = {dataGroup_1_3, dataGroup_0_3};
  wire [15:0]   res_lo_lo_lo_lo_hi_3 = {dataGroup_3_3, dataGroup_2_3};
  wire [31:0]   res_lo_lo_lo_lo_3 = {res_lo_lo_lo_lo_hi_3, res_lo_lo_lo_lo_lo_3};
  wire [15:0]   res_lo_lo_lo_hi_lo_3 = {dataGroup_5_3, dataGroup_4_3};
  wire [15:0]   res_lo_lo_lo_hi_hi_3 = {dataGroup_7_3, dataGroup_6_3};
  wire [31:0]   res_lo_lo_lo_hi_3 = {res_lo_lo_lo_hi_hi_3, res_lo_lo_lo_hi_lo_3};
  wire [63:0]   res_lo_lo_lo_3 = {res_lo_lo_lo_hi_3, res_lo_lo_lo_lo_3};
  wire [15:0]   res_lo_lo_hi_lo_lo_3 = {dataGroup_9_3, dataGroup_8_3};
  wire [15:0]   res_lo_lo_hi_lo_hi_3 = {dataGroup_11_3, dataGroup_10_3};
  wire [31:0]   res_lo_lo_hi_lo_3 = {res_lo_lo_hi_lo_hi_3, res_lo_lo_hi_lo_lo_3};
  wire [15:0]   res_lo_lo_hi_hi_lo_3 = {dataGroup_13_3, dataGroup_12_3};
  wire [15:0]   res_lo_lo_hi_hi_hi_3 = {dataGroup_15_3, dataGroup_14_3};
  wire [31:0]   res_lo_lo_hi_hi_3 = {res_lo_lo_hi_hi_hi_3, res_lo_lo_hi_hi_lo_3};
  wire [63:0]   res_lo_lo_hi_3 = {res_lo_lo_hi_hi_3, res_lo_lo_hi_lo_3};
  wire [127:0]  res_lo_lo_3 = {res_lo_lo_hi_3, res_lo_lo_lo_3};
  wire [15:0]   res_lo_hi_lo_lo_lo_3 = {dataGroup_17_3, dataGroup_16_3};
  wire [15:0]   res_lo_hi_lo_lo_hi_3 = {dataGroup_19_3, dataGroup_18_3};
  wire [31:0]   res_lo_hi_lo_lo_3 = {res_lo_hi_lo_lo_hi_3, res_lo_hi_lo_lo_lo_3};
  wire [15:0]   res_lo_hi_lo_hi_lo_3 = {dataGroup_21_3, dataGroup_20_3};
  wire [15:0]   res_lo_hi_lo_hi_hi_3 = {dataGroup_23_3, dataGroup_22_3};
  wire [31:0]   res_lo_hi_lo_hi_3 = {res_lo_hi_lo_hi_hi_3, res_lo_hi_lo_hi_lo_3};
  wire [63:0]   res_lo_hi_lo_3 = {res_lo_hi_lo_hi_3, res_lo_hi_lo_lo_3};
  wire [15:0]   res_lo_hi_hi_lo_lo_3 = {dataGroup_25_3, dataGroup_24_3};
  wire [15:0]   res_lo_hi_hi_lo_hi_3 = {dataGroup_27_3, dataGroup_26_3};
  wire [31:0]   res_lo_hi_hi_lo_3 = {res_lo_hi_hi_lo_hi_3, res_lo_hi_hi_lo_lo_3};
  wire [15:0]   res_lo_hi_hi_hi_lo_3 = {dataGroup_29_3, dataGroup_28_3};
  wire [15:0]   res_lo_hi_hi_hi_hi_3 = {dataGroup_31_3, dataGroup_30_3};
  wire [31:0]   res_lo_hi_hi_hi_3 = {res_lo_hi_hi_hi_hi_3, res_lo_hi_hi_hi_lo_3};
  wire [63:0]   res_lo_hi_hi_3 = {res_lo_hi_hi_hi_3, res_lo_hi_hi_lo_3};
  wire [127:0]  res_lo_hi_3 = {res_lo_hi_hi_3, res_lo_hi_lo_3};
  wire [255:0]  res_lo_3 = {res_lo_hi_3, res_lo_lo_3};
  wire [15:0]   res_hi_lo_lo_lo_lo_3 = {dataGroup_33_3, dataGroup_32_3};
  wire [15:0]   res_hi_lo_lo_lo_hi_3 = {dataGroup_35_3, dataGroup_34_3};
  wire [31:0]   res_hi_lo_lo_lo_3 = {res_hi_lo_lo_lo_hi_3, res_hi_lo_lo_lo_lo_3};
  wire [15:0]   res_hi_lo_lo_hi_lo_3 = {dataGroup_37_3, dataGroup_36_3};
  wire [15:0]   res_hi_lo_lo_hi_hi_3 = {dataGroup_39_3, dataGroup_38_3};
  wire [31:0]   res_hi_lo_lo_hi_3 = {res_hi_lo_lo_hi_hi_3, res_hi_lo_lo_hi_lo_3};
  wire [63:0]   res_hi_lo_lo_3 = {res_hi_lo_lo_hi_3, res_hi_lo_lo_lo_3};
  wire [15:0]   res_hi_lo_hi_lo_lo_3 = {dataGroup_41_3, dataGroup_40_3};
  wire [15:0]   res_hi_lo_hi_lo_hi_3 = {dataGroup_43_3, dataGroup_42_3};
  wire [31:0]   res_hi_lo_hi_lo_3 = {res_hi_lo_hi_lo_hi_3, res_hi_lo_hi_lo_lo_3};
  wire [15:0]   res_hi_lo_hi_hi_lo_3 = {dataGroup_45_3, dataGroup_44_3};
  wire [15:0]   res_hi_lo_hi_hi_hi_3 = {dataGroup_47_3, dataGroup_46_3};
  wire [31:0]   res_hi_lo_hi_hi_3 = {res_hi_lo_hi_hi_hi_3, res_hi_lo_hi_hi_lo_3};
  wire [63:0]   res_hi_lo_hi_3 = {res_hi_lo_hi_hi_3, res_hi_lo_hi_lo_3};
  wire [127:0]  res_hi_lo_3 = {res_hi_lo_hi_3, res_hi_lo_lo_3};
  wire [15:0]   res_hi_hi_lo_lo_lo_3 = {dataGroup_49_3, dataGroup_48_3};
  wire [15:0]   res_hi_hi_lo_lo_hi_3 = {dataGroup_51_3, dataGroup_50_3};
  wire [31:0]   res_hi_hi_lo_lo_3 = {res_hi_hi_lo_lo_hi_3, res_hi_hi_lo_lo_lo_3};
  wire [15:0]   res_hi_hi_lo_hi_lo_3 = {dataGroup_53_3, dataGroup_52_3};
  wire [15:0]   res_hi_hi_lo_hi_hi_3 = {dataGroup_55_3, dataGroup_54_3};
  wire [31:0]   res_hi_hi_lo_hi_3 = {res_hi_hi_lo_hi_hi_3, res_hi_hi_lo_hi_lo_3};
  wire [63:0]   res_hi_hi_lo_3 = {res_hi_hi_lo_hi_3, res_hi_hi_lo_lo_3};
  wire [15:0]   res_hi_hi_hi_lo_lo_3 = {dataGroup_57_3, dataGroup_56_3};
  wire [15:0]   res_hi_hi_hi_lo_hi_3 = {dataGroup_59_3, dataGroup_58_3};
  wire [31:0]   res_hi_hi_hi_lo_3 = {res_hi_hi_hi_lo_hi_3, res_hi_hi_hi_lo_lo_3};
  wire [15:0]   res_hi_hi_hi_hi_lo_3 = {dataGroup_61_3, dataGroup_60_3};
  wire [15:0]   res_hi_hi_hi_hi_hi_3 = {dataGroup_63_3, dataGroup_62_3};
  wire [31:0]   res_hi_hi_hi_hi_3 = {res_hi_hi_hi_hi_hi_3, res_hi_hi_hi_hi_lo_3};
  wire [63:0]   res_hi_hi_hi_3 = {res_hi_hi_hi_hi_3, res_hi_hi_hi_lo_3};
  wire [127:0]  res_hi_hi_3 = {res_hi_hi_hi_3, res_hi_hi_lo_3};
  wire [255:0]  res_hi_3 = {res_hi_hi_3, res_hi_lo_3};
  wire [511:0]  res_16 = {res_hi_3, res_lo_3};
  wire [2047:0] dataGroup_lo_256 = {dataGroup_lo_hi_256, dataGroup_lo_lo_256};
  wire [2047:0] dataGroup_hi_256 = {dataGroup_hi_hi_256, dataGroup_hi_lo_256};
  wire [7:0]    dataGroup_0_4 = dataGroup_lo_256[15:8];
  wire [2047:0] dataGroup_lo_257 = {dataGroup_lo_hi_257, dataGroup_lo_lo_257};
  wire [2047:0] dataGroup_hi_257 = {dataGroup_hi_hi_257, dataGroup_hi_lo_257};
  wire [7:0]    dataGroup_1_4 = dataGroup_lo_257[39:32];
  wire [2047:0] dataGroup_lo_258 = {dataGroup_lo_hi_258, dataGroup_lo_lo_258};
  wire [2047:0] dataGroup_hi_258 = {dataGroup_hi_hi_258, dataGroup_hi_lo_258};
  wire [7:0]    dataGroup_2_4 = dataGroup_lo_258[63:56];
  wire [2047:0] dataGroup_lo_259 = {dataGroup_lo_hi_259, dataGroup_lo_lo_259};
  wire [2047:0] dataGroup_hi_259 = {dataGroup_hi_hi_259, dataGroup_hi_lo_259};
  wire [7:0]    dataGroup_3_4 = dataGroup_lo_259[87:80];
  wire [2047:0] dataGroup_lo_260 = {dataGroup_lo_hi_260, dataGroup_lo_lo_260};
  wire [2047:0] dataGroup_hi_260 = {dataGroup_hi_hi_260, dataGroup_hi_lo_260};
  wire [7:0]    dataGroup_4_4 = dataGroup_lo_260[111:104];
  wire [2047:0] dataGroup_lo_261 = {dataGroup_lo_hi_261, dataGroup_lo_lo_261};
  wire [2047:0] dataGroup_hi_261 = {dataGroup_hi_hi_261, dataGroup_hi_lo_261};
  wire [7:0]    dataGroup_5_4 = dataGroup_lo_261[135:128];
  wire [2047:0] dataGroup_lo_262 = {dataGroup_lo_hi_262, dataGroup_lo_lo_262};
  wire [2047:0] dataGroup_hi_262 = {dataGroup_hi_hi_262, dataGroup_hi_lo_262};
  wire [7:0]    dataGroup_6_4 = dataGroup_lo_262[159:152];
  wire [2047:0] dataGroup_lo_263 = {dataGroup_lo_hi_263, dataGroup_lo_lo_263};
  wire [2047:0] dataGroup_hi_263 = {dataGroup_hi_hi_263, dataGroup_hi_lo_263};
  wire [7:0]    dataGroup_7_4 = dataGroup_lo_263[183:176];
  wire [2047:0] dataGroup_lo_264 = {dataGroup_lo_hi_264, dataGroup_lo_lo_264};
  wire [2047:0] dataGroup_hi_264 = {dataGroup_hi_hi_264, dataGroup_hi_lo_264};
  wire [7:0]    dataGroup_8_4 = dataGroup_lo_264[207:200];
  wire [2047:0] dataGroup_lo_265 = {dataGroup_lo_hi_265, dataGroup_lo_lo_265};
  wire [2047:0] dataGroup_hi_265 = {dataGroup_hi_hi_265, dataGroup_hi_lo_265};
  wire [7:0]    dataGroup_9_4 = dataGroup_lo_265[231:224];
  wire [2047:0] dataGroup_lo_266 = {dataGroup_lo_hi_266, dataGroup_lo_lo_266};
  wire [2047:0] dataGroup_hi_266 = {dataGroup_hi_hi_266, dataGroup_hi_lo_266};
  wire [7:0]    dataGroup_10_4 = dataGroup_lo_266[255:248];
  wire [2047:0] dataGroup_lo_267 = {dataGroup_lo_hi_267, dataGroup_lo_lo_267};
  wire [2047:0] dataGroup_hi_267 = {dataGroup_hi_hi_267, dataGroup_hi_lo_267};
  wire [7:0]    dataGroup_11_4 = dataGroup_lo_267[279:272];
  wire [2047:0] dataGroup_lo_268 = {dataGroup_lo_hi_268, dataGroup_lo_lo_268};
  wire [2047:0] dataGroup_hi_268 = {dataGroup_hi_hi_268, dataGroup_hi_lo_268};
  wire [7:0]    dataGroup_12_4 = dataGroup_lo_268[303:296];
  wire [2047:0] dataGroup_lo_269 = {dataGroup_lo_hi_269, dataGroup_lo_lo_269};
  wire [2047:0] dataGroup_hi_269 = {dataGroup_hi_hi_269, dataGroup_hi_lo_269};
  wire [7:0]    dataGroup_13_4 = dataGroup_lo_269[327:320];
  wire [2047:0] dataGroup_lo_270 = {dataGroup_lo_hi_270, dataGroup_lo_lo_270};
  wire [2047:0] dataGroup_hi_270 = {dataGroup_hi_hi_270, dataGroup_hi_lo_270};
  wire [7:0]    dataGroup_14_4 = dataGroup_lo_270[351:344];
  wire [2047:0] dataGroup_lo_271 = {dataGroup_lo_hi_271, dataGroup_lo_lo_271};
  wire [2047:0] dataGroup_hi_271 = {dataGroup_hi_hi_271, dataGroup_hi_lo_271};
  wire [7:0]    dataGroup_15_4 = dataGroup_lo_271[375:368];
  wire [2047:0] dataGroup_lo_272 = {dataGroup_lo_hi_272, dataGroup_lo_lo_272};
  wire [2047:0] dataGroup_hi_272 = {dataGroup_hi_hi_272, dataGroup_hi_lo_272};
  wire [7:0]    dataGroup_16_4 = dataGroup_lo_272[399:392];
  wire [2047:0] dataGroup_lo_273 = {dataGroup_lo_hi_273, dataGroup_lo_lo_273};
  wire [2047:0] dataGroup_hi_273 = {dataGroup_hi_hi_273, dataGroup_hi_lo_273};
  wire [7:0]    dataGroup_17_4 = dataGroup_lo_273[423:416];
  wire [2047:0] dataGroup_lo_274 = {dataGroup_lo_hi_274, dataGroup_lo_lo_274};
  wire [2047:0] dataGroup_hi_274 = {dataGroup_hi_hi_274, dataGroup_hi_lo_274};
  wire [7:0]    dataGroup_18_4 = dataGroup_lo_274[447:440];
  wire [2047:0] dataGroup_lo_275 = {dataGroup_lo_hi_275, dataGroup_lo_lo_275};
  wire [2047:0] dataGroup_hi_275 = {dataGroup_hi_hi_275, dataGroup_hi_lo_275};
  wire [7:0]    dataGroup_19_4 = dataGroup_lo_275[471:464];
  wire [2047:0] dataGroup_lo_276 = {dataGroup_lo_hi_276, dataGroup_lo_lo_276};
  wire [2047:0] dataGroup_hi_276 = {dataGroup_hi_hi_276, dataGroup_hi_lo_276};
  wire [7:0]    dataGroup_20_4 = dataGroup_lo_276[495:488];
  wire [2047:0] dataGroup_lo_277 = {dataGroup_lo_hi_277, dataGroup_lo_lo_277};
  wire [2047:0] dataGroup_hi_277 = {dataGroup_hi_hi_277, dataGroup_hi_lo_277};
  wire [7:0]    dataGroup_21_4 = dataGroup_lo_277[519:512];
  wire [2047:0] dataGroup_lo_278 = {dataGroup_lo_hi_278, dataGroup_lo_lo_278};
  wire [2047:0] dataGroup_hi_278 = {dataGroup_hi_hi_278, dataGroup_hi_lo_278};
  wire [7:0]    dataGroup_22_4 = dataGroup_lo_278[543:536];
  wire [2047:0] dataGroup_lo_279 = {dataGroup_lo_hi_279, dataGroup_lo_lo_279};
  wire [2047:0] dataGroup_hi_279 = {dataGroup_hi_hi_279, dataGroup_hi_lo_279};
  wire [7:0]    dataGroup_23_4 = dataGroup_lo_279[567:560];
  wire [2047:0] dataGroup_lo_280 = {dataGroup_lo_hi_280, dataGroup_lo_lo_280};
  wire [2047:0] dataGroup_hi_280 = {dataGroup_hi_hi_280, dataGroup_hi_lo_280};
  wire [7:0]    dataGroup_24_4 = dataGroup_lo_280[591:584];
  wire [2047:0] dataGroup_lo_281 = {dataGroup_lo_hi_281, dataGroup_lo_lo_281};
  wire [2047:0] dataGroup_hi_281 = {dataGroup_hi_hi_281, dataGroup_hi_lo_281};
  wire [7:0]    dataGroup_25_4 = dataGroup_lo_281[615:608];
  wire [2047:0] dataGroup_lo_282 = {dataGroup_lo_hi_282, dataGroup_lo_lo_282};
  wire [2047:0] dataGroup_hi_282 = {dataGroup_hi_hi_282, dataGroup_hi_lo_282};
  wire [7:0]    dataGroup_26_4 = dataGroup_lo_282[639:632];
  wire [2047:0] dataGroup_lo_283 = {dataGroup_lo_hi_283, dataGroup_lo_lo_283};
  wire [2047:0] dataGroup_hi_283 = {dataGroup_hi_hi_283, dataGroup_hi_lo_283};
  wire [7:0]    dataGroup_27_4 = dataGroup_lo_283[663:656];
  wire [2047:0] dataGroup_lo_284 = {dataGroup_lo_hi_284, dataGroup_lo_lo_284};
  wire [2047:0] dataGroup_hi_284 = {dataGroup_hi_hi_284, dataGroup_hi_lo_284};
  wire [7:0]    dataGroup_28_4 = dataGroup_lo_284[687:680];
  wire [2047:0] dataGroup_lo_285 = {dataGroup_lo_hi_285, dataGroup_lo_lo_285};
  wire [2047:0] dataGroup_hi_285 = {dataGroup_hi_hi_285, dataGroup_hi_lo_285};
  wire [7:0]    dataGroup_29_4 = dataGroup_lo_285[711:704];
  wire [2047:0] dataGroup_lo_286 = {dataGroup_lo_hi_286, dataGroup_lo_lo_286};
  wire [2047:0] dataGroup_hi_286 = {dataGroup_hi_hi_286, dataGroup_hi_lo_286};
  wire [7:0]    dataGroup_30_4 = dataGroup_lo_286[735:728];
  wire [2047:0] dataGroup_lo_287 = {dataGroup_lo_hi_287, dataGroup_lo_lo_287};
  wire [2047:0] dataGroup_hi_287 = {dataGroup_hi_hi_287, dataGroup_hi_lo_287};
  wire [7:0]    dataGroup_31_4 = dataGroup_lo_287[759:752];
  wire [2047:0] dataGroup_lo_288 = {dataGroup_lo_hi_288, dataGroup_lo_lo_288};
  wire [2047:0] dataGroup_hi_288 = {dataGroup_hi_hi_288, dataGroup_hi_lo_288};
  wire [7:0]    dataGroup_32_4 = dataGroup_lo_288[783:776];
  wire [2047:0] dataGroup_lo_289 = {dataGroup_lo_hi_289, dataGroup_lo_lo_289};
  wire [2047:0] dataGroup_hi_289 = {dataGroup_hi_hi_289, dataGroup_hi_lo_289};
  wire [7:0]    dataGroup_33_4 = dataGroup_lo_289[807:800];
  wire [2047:0] dataGroup_lo_290 = {dataGroup_lo_hi_290, dataGroup_lo_lo_290};
  wire [2047:0] dataGroup_hi_290 = {dataGroup_hi_hi_290, dataGroup_hi_lo_290};
  wire [7:0]    dataGroup_34_4 = dataGroup_lo_290[831:824];
  wire [2047:0] dataGroup_lo_291 = {dataGroup_lo_hi_291, dataGroup_lo_lo_291};
  wire [2047:0] dataGroup_hi_291 = {dataGroup_hi_hi_291, dataGroup_hi_lo_291};
  wire [7:0]    dataGroup_35_4 = dataGroup_lo_291[855:848];
  wire [2047:0] dataGroup_lo_292 = {dataGroup_lo_hi_292, dataGroup_lo_lo_292};
  wire [2047:0] dataGroup_hi_292 = {dataGroup_hi_hi_292, dataGroup_hi_lo_292};
  wire [7:0]    dataGroup_36_4 = dataGroup_lo_292[879:872];
  wire [2047:0] dataGroup_lo_293 = {dataGroup_lo_hi_293, dataGroup_lo_lo_293};
  wire [2047:0] dataGroup_hi_293 = {dataGroup_hi_hi_293, dataGroup_hi_lo_293};
  wire [7:0]    dataGroup_37_4 = dataGroup_lo_293[903:896];
  wire [2047:0] dataGroup_lo_294 = {dataGroup_lo_hi_294, dataGroup_lo_lo_294};
  wire [2047:0] dataGroup_hi_294 = {dataGroup_hi_hi_294, dataGroup_hi_lo_294};
  wire [7:0]    dataGroup_38_4 = dataGroup_lo_294[927:920];
  wire [2047:0] dataGroup_lo_295 = {dataGroup_lo_hi_295, dataGroup_lo_lo_295};
  wire [2047:0] dataGroup_hi_295 = {dataGroup_hi_hi_295, dataGroup_hi_lo_295};
  wire [7:0]    dataGroup_39_4 = dataGroup_lo_295[951:944];
  wire [2047:0] dataGroup_lo_296 = {dataGroup_lo_hi_296, dataGroup_lo_lo_296};
  wire [2047:0] dataGroup_hi_296 = {dataGroup_hi_hi_296, dataGroup_hi_lo_296};
  wire [7:0]    dataGroup_40_4 = dataGroup_lo_296[975:968];
  wire [2047:0] dataGroup_lo_297 = {dataGroup_lo_hi_297, dataGroup_lo_lo_297};
  wire [2047:0] dataGroup_hi_297 = {dataGroup_hi_hi_297, dataGroup_hi_lo_297};
  wire [7:0]    dataGroup_41_4 = dataGroup_lo_297[999:992];
  wire [2047:0] dataGroup_lo_298 = {dataGroup_lo_hi_298, dataGroup_lo_lo_298};
  wire [2047:0] dataGroup_hi_298 = {dataGroup_hi_hi_298, dataGroup_hi_lo_298};
  wire [7:0]    dataGroup_42_4 = dataGroup_lo_298[1023:1016];
  wire [2047:0] dataGroup_lo_299 = {dataGroup_lo_hi_299, dataGroup_lo_lo_299};
  wire [2047:0] dataGroup_hi_299 = {dataGroup_hi_hi_299, dataGroup_hi_lo_299};
  wire [7:0]    dataGroup_43_4 = dataGroup_lo_299[1047:1040];
  wire [2047:0] dataGroup_lo_300 = {dataGroup_lo_hi_300, dataGroup_lo_lo_300};
  wire [2047:0] dataGroup_hi_300 = {dataGroup_hi_hi_300, dataGroup_hi_lo_300};
  wire [7:0]    dataGroup_44_4 = dataGroup_lo_300[1071:1064];
  wire [2047:0] dataGroup_lo_301 = {dataGroup_lo_hi_301, dataGroup_lo_lo_301};
  wire [2047:0] dataGroup_hi_301 = {dataGroup_hi_hi_301, dataGroup_hi_lo_301};
  wire [7:0]    dataGroup_45_4 = dataGroup_lo_301[1095:1088];
  wire [2047:0] dataGroup_lo_302 = {dataGroup_lo_hi_302, dataGroup_lo_lo_302};
  wire [2047:0] dataGroup_hi_302 = {dataGroup_hi_hi_302, dataGroup_hi_lo_302};
  wire [7:0]    dataGroup_46_4 = dataGroup_lo_302[1119:1112];
  wire [2047:0] dataGroup_lo_303 = {dataGroup_lo_hi_303, dataGroup_lo_lo_303};
  wire [2047:0] dataGroup_hi_303 = {dataGroup_hi_hi_303, dataGroup_hi_lo_303};
  wire [7:0]    dataGroup_47_4 = dataGroup_lo_303[1143:1136];
  wire [2047:0] dataGroup_lo_304 = {dataGroup_lo_hi_304, dataGroup_lo_lo_304};
  wire [2047:0] dataGroup_hi_304 = {dataGroup_hi_hi_304, dataGroup_hi_lo_304};
  wire [7:0]    dataGroup_48_4 = dataGroup_lo_304[1167:1160];
  wire [2047:0] dataGroup_lo_305 = {dataGroup_lo_hi_305, dataGroup_lo_lo_305};
  wire [2047:0] dataGroup_hi_305 = {dataGroup_hi_hi_305, dataGroup_hi_lo_305};
  wire [7:0]    dataGroup_49_4 = dataGroup_lo_305[1191:1184];
  wire [2047:0] dataGroup_lo_306 = {dataGroup_lo_hi_306, dataGroup_lo_lo_306};
  wire [2047:0] dataGroup_hi_306 = {dataGroup_hi_hi_306, dataGroup_hi_lo_306};
  wire [7:0]    dataGroup_50_4 = dataGroup_lo_306[1215:1208];
  wire [2047:0] dataGroup_lo_307 = {dataGroup_lo_hi_307, dataGroup_lo_lo_307};
  wire [2047:0] dataGroup_hi_307 = {dataGroup_hi_hi_307, dataGroup_hi_lo_307};
  wire [7:0]    dataGroup_51_4 = dataGroup_lo_307[1239:1232];
  wire [2047:0] dataGroup_lo_308 = {dataGroup_lo_hi_308, dataGroup_lo_lo_308};
  wire [2047:0] dataGroup_hi_308 = {dataGroup_hi_hi_308, dataGroup_hi_lo_308};
  wire [7:0]    dataGroup_52_4 = dataGroup_lo_308[1263:1256];
  wire [2047:0] dataGroup_lo_309 = {dataGroup_lo_hi_309, dataGroup_lo_lo_309};
  wire [2047:0] dataGroup_hi_309 = {dataGroup_hi_hi_309, dataGroup_hi_lo_309};
  wire [7:0]    dataGroup_53_4 = dataGroup_lo_309[1287:1280];
  wire [2047:0] dataGroup_lo_310 = {dataGroup_lo_hi_310, dataGroup_lo_lo_310};
  wire [2047:0] dataGroup_hi_310 = {dataGroup_hi_hi_310, dataGroup_hi_lo_310};
  wire [7:0]    dataGroup_54_4 = dataGroup_lo_310[1311:1304];
  wire [2047:0] dataGroup_lo_311 = {dataGroup_lo_hi_311, dataGroup_lo_lo_311};
  wire [2047:0] dataGroup_hi_311 = {dataGroup_hi_hi_311, dataGroup_hi_lo_311};
  wire [7:0]    dataGroup_55_4 = dataGroup_lo_311[1335:1328];
  wire [2047:0] dataGroup_lo_312 = {dataGroup_lo_hi_312, dataGroup_lo_lo_312};
  wire [2047:0] dataGroup_hi_312 = {dataGroup_hi_hi_312, dataGroup_hi_lo_312};
  wire [7:0]    dataGroup_56_4 = dataGroup_lo_312[1359:1352];
  wire [2047:0] dataGroup_lo_313 = {dataGroup_lo_hi_313, dataGroup_lo_lo_313};
  wire [2047:0] dataGroup_hi_313 = {dataGroup_hi_hi_313, dataGroup_hi_lo_313};
  wire [7:0]    dataGroup_57_4 = dataGroup_lo_313[1383:1376];
  wire [2047:0] dataGroup_lo_314 = {dataGroup_lo_hi_314, dataGroup_lo_lo_314};
  wire [2047:0] dataGroup_hi_314 = {dataGroup_hi_hi_314, dataGroup_hi_lo_314};
  wire [7:0]    dataGroup_58_4 = dataGroup_lo_314[1407:1400];
  wire [2047:0] dataGroup_lo_315 = {dataGroup_lo_hi_315, dataGroup_lo_lo_315};
  wire [2047:0] dataGroup_hi_315 = {dataGroup_hi_hi_315, dataGroup_hi_lo_315};
  wire [7:0]    dataGroup_59_4 = dataGroup_lo_315[1431:1424];
  wire [2047:0] dataGroup_lo_316 = {dataGroup_lo_hi_316, dataGroup_lo_lo_316};
  wire [2047:0] dataGroup_hi_316 = {dataGroup_hi_hi_316, dataGroup_hi_lo_316};
  wire [7:0]    dataGroup_60_4 = dataGroup_lo_316[1455:1448];
  wire [2047:0] dataGroup_lo_317 = {dataGroup_lo_hi_317, dataGroup_lo_lo_317};
  wire [2047:0] dataGroup_hi_317 = {dataGroup_hi_hi_317, dataGroup_hi_lo_317};
  wire [7:0]    dataGroup_61_4 = dataGroup_lo_317[1479:1472];
  wire [2047:0] dataGroup_lo_318 = {dataGroup_lo_hi_318, dataGroup_lo_lo_318};
  wire [2047:0] dataGroup_hi_318 = {dataGroup_hi_hi_318, dataGroup_hi_lo_318};
  wire [7:0]    dataGroup_62_4 = dataGroup_lo_318[1503:1496];
  wire [2047:0] dataGroup_lo_319 = {dataGroup_lo_hi_319, dataGroup_lo_lo_319};
  wire [2047:0] dataGroup_hi_319 = {dataGroup_hi_hi_319, dataGroup_hi_lo_319};
  wire [7:0]    dataGroup_63_4 = dataGroup_lo_319[1527:1520];
  wire [15:0]   res_lo_lo_lo_lo_lo_4 = {dataGroup_1_4, dataGroup_0_4};
  wire [15:0]   res_lo_lo_lo_lo_hi_4 = {dataGroup_3_4, dataGroup_2_4};
  wire [31:0]   res_lo_lo_lo_lo_4 = {res_lo_lo_lo_lo_hi_4, res_lo_lo_lo_lo_lo_4};
  wire [15:0]   res_lo_lo_lo_hi_lo_4 = {dataGroup_5_4, dataGroup_4_4};
  wire [15:0]   res_lo_lo_lo_hi_hi_4 = {dataGroup_7_4, dataGroup_6_4};
  wire [31:0]   res_lo_lo_lo_hi_4 = {res_lo_lo_lo_hi_hi_4, res_lo_lo_lo_hi_lo_4};
  wire [63:0]   res_lo_lo_lo_4 = {res_lo_lo_lo_hi_4, res_lo_lo_lo_lo_4};
  wire [15:0]   res_lo_lo_hi_lo_lo_4 = {dataGroup_9_4, dataGroup_8_4};
  wire [15:0]   res_lo_lo_hi_lo_hi_4 = {dataGroup_11_4, dataGroup_10_4};
  wire [31:0]   res_lo_lo_hi_lo_4 = {res_lo_lo_hi_lo_hi_4, res_lo_lo_hi_lo_lo_4};
  wire [15:0]   res_lo_lo_hi_hi_lo_4 = {dataGroup_13_4, dataGroup_12_4};
  wire [15:0]   res_lo_lo_hi_hi_hi_4 = {dataGroup_15_4, dataGroup_14_4};
  wire [31:0]   res_lo_lo_hi_hi_4 = {res_lo_lo_hi_hi_hi_4, res_lo_lo_hi_hi_lo_4};
  wire [63:0]   res_lo_lo_hi_4 = {res_lo_lo_hi_hi_4, res_lo_lo_hi_lo_4};
  wire [127:0]  res_lo_lo_4 = {res_lo_lo_hi_4, res_lo_lo_lo_4};
  wire [15:0]   res_lo_hi_lo_lo_lo_4 = {dataGroup_17_4, dataGroup_16_4};
  wire [15:0]   res_lo_hi_lo_lo_hi_4 = {dataGroup_19_4, dataGroup_18_4};
  wire [31:0]   res_lo_hi_lo_lo_4 = {res_lo_hi_lo_lo_hi_4, res_lo_hi_lo_lo_lo_4};
  wire [15:0]   res_lo_hi_lo_hi_lo_4 = {dataGroup_21_4, dataGroup_20_4};
  wire [15:0]   res_lo_hi_lo_hi_hi_4 = {dataGroup_23_4, dataGroup_22_4};
  wire [31:0]   res_lo_hi_lo_hi_4 = {res_lo_hi_lo_hi_hi_4, res_lo_hi_lo_hi_lo_4};
  wire [63:0]   res_lo_hi_lo_4 = {res_lo_hi_lo_hi_4, res_lo_hi_lo_lo_4};
  wire [15:0]   res_lo_hi_hi_lo_lo_4 = {dataGroup_25_4, dataGroup_24_4};
  wire [15:0]   res_lo_hi_hi_lo_hi_4 = {dataGroup_27_4, dataGroup_26_4};
  wire [31:0]   res_lo_hi_hi_lo_4 = {res_lo_hi_hi_lo_hi_4, res_lo_hi_hi_lo_lo_4};
  wire [15:0]   res_lo_hi_hi_hi_lo_4 = {dataGroup_29_4, dataGroup_28_4};
  wire [15:0]   res_lo_hi_hi_hi_hi_4 = {dataGroup_31_4, dataGroup_30_4};
  wire [31:0]   res_lo_hi_hi_hi_4 = {res_lo_hi_hi_hi_hi_4, res_lo_hi_hi_hi_lo_4};
  wire [63:0]   res_lo_hi_hi_4 = {res_lo_hi_hi_hi_4, res_lo_hi_hi_lo_4};
  wire [127:0]  res_lo_hi_4 = {res_lo_hi_hi_4, res_lo_hi_lo_4};
  wire [255:0]  res_lo_4 = {res_lo_hi_4, res_lo_lo_4};
  wire [15:0]   res_hi_lo_lo_lo_lo_4 = {dataGroup_33_4, dataGroup_32_4};
  wire [15:0]   res_hi_lo_lo_lo_hi_4 = {dataGroup_35_4, dataGroup_34_4};
  wire [31:0]   res_hi_lo_lo_lo_4 = {res_hi_lo_lo_lo_hi_4, res_hi_lo_lo_lo_lo_4};
  wire [15:0]   res_hi_lo_lo_hi_lo_4 = {dataGroup_37_4, dataGroup_36_4};
  wire [15:0]   res_hi_lo_lo_hi_hi_4 = {dataGroup_39_4, dataGroup_38_4};
  wire [31:0]   res_hi_lo_lo_hi_4 = {res_hi_lo_lo_hi_hi_4, res_hi_lo_lo_hi_lo_4};
  wire [63:0]   res_hi_lo_lo_4 = {res_hi_lo_lo_hi_4, res_hi_lo_lo_lo_4};
  wire [15:0]   res_hi_lo_hi_lo_lo_4 = {dataGroup_41_4, dataGroup_40_4};
  wire [15:0]   res_hi_lo_hi_lo_hi_4 = {dataGroup_43_4, dataGroup_42_4};
  wire [31:0]   res_hi_lo_hi_lo_4 = {res_hi_lo_hi_lo_hi_4, res_hi_lo_hi_lo_lo_4};
  wire [15:0]   res_hi_lo_hi_hi_lo_4 = {dataGroup_45_4, dataGroup_44_4};
  wire [15:0]   res_hi_lo_hi_hi_hi_4 = {dataGroup_47_4, dataGroup_46_4};
  wire [31:0]   res_hi_lo_hi_hi_4 = {res_hi_lo_hi_hi_hi_4, res_hi_lo_hi_hi_lo_4};
  wire [63:0]   res_hi_lo_hi_4 = {res_hi_lo_hi_hi_4, res_hi_lo_hi_lo_4};
  wire [127:0]  res_hi_lo_4 = {res_hi_lo_hi_4, res_hi_lo_lo_4};
  wire [15:0]   res_hi_hi_lo_lo_lo_4 = {dataGroup_49_4, dataGroup_48_4};
  wire [15:0]   res_hi_hi_lo_lo_hi_4 = {dataGroup_51_4, dataGroup_50_4};
  wire [31:0]   res_hi_hi_lo_lo_4 = {res_hi_hi_lo_lo_hi_4, res_hi_hi_lo_lo_lo_4};
  wire [15:0]   res_hi_hi_lo_hi_lo_4 = {dataGroup_53_4, dataGroup_52_4};
  wire [15:0]   res_hi_hi_lo_hi_hi_4 = {dataGroup_55_4, dataGroup_54_4};
  wire [31:0]   res_hi_hi_lo_hi_4 = {res_hi_hi_lo_hi_hi_4, res_hi_hi_lo_hi_lo_4};
  wire [63:0]   res_hi_hi_lo_4 = {res_hi_hi_lo_hi_4, res_hi_hi_lo_lo_4};
  wire [15:0]   res_hi_hi_hi_lo_lo_4 = {dataGroup_57_4, dataGroup_56_4};
  wire [15:0]   res_hi_hi_hi_lo_hi_4 = {dataGroup_59_4, dataGroup_58_4};
  wire [31:0]   res_hi_hi_hi_lo_4 = {res_hi_hi_hi_lo_hi_4, res_hi_hi_hi_lo_lo_4};
  wire [15:0]   res_hi_hi_hi_hi_lo_4 = {dataGroup_61_4, dataGroup_60_4};
  wire [15:0]   res_hi_hi_hi_hi_hi_4 = {dataGroup_63_4, dataGroup_62_4};
  wire [31:0]   res_hi_hi_hi_hi_4 = {res_hi_hi_hi_hi_hi_4, res_hi_hi_hi_hi_lo_4};
  wire [63:0]   res_hi_hi_hi_4 = {res_hi_hi_hi_hi_4, res_hi_hi_hi_lo_4};
  wire [127:0]  res_hi_hi_4 = {res_hi_hi_hi_4, res_hi_hi_lo_4};
  wire [255:0]  res_hi_4 = {res_hi_hi_4, res_hi_lo_4};
  wire [511:0]  res_17 = {res_hi_4, res_lo_4};
  wire [2047:0] dataGroup_lo_320 = {dataGroup_lo_hi_320, dataGroup_lo_lo_320};
  wire [2047:0] dataGroup_hi_320 = {dataGroup_hi_hi_320, dataGroup_hi_lo_320};
  wire [7:0]    dataGroup_0_5 = dataGroup_lo_320[23:16];
  wire [2047:0] dataGroup_lo_321 = {dataGroup_lo_hi_321, dataGroup_lo_lo_321};
  wire [2047:0] dataGroup_hi_321 = {dataGroup_hi_hi_321, dataGroup_hi_lo_321};
  wire [7:0]    dataGroup_1_5 = dataGroup_lo_321[47:40];
  wire [2047:0] dataGroup_lo_322 = {dataGroup_lo_hi_322, dataGroup_lo_lo_322};
  wire [2047:0] dataGroup_hi_322 = {dataGroup_hi_hi_322, dataGroup_hi_lo_322};
  wire [7:0]    dataGroup_2_5 = dataGroup_lo_322[71:64];
  wire [2047:0] dataGroup_lo_323 = {dataGroup_lo_hi_323, dataGroup_lo_lo_323};
  wire [2047:0] dataGroup_hi_323 = {dataGroup_hi_hi_323, dataGroup_hi_lo_323};
  wire [7:0]    dataGroup_3_5 = dataGroup_lo_323[95:88];
  wire [2047:0] dataGroup_lo_324 = {dataGroup_lo_hi_324, dataGroup_lo_lo_324};
  wire [2047:0] dataGroup_hi_324 = {dataGroup_hi_hi_324, dataGroup_hi_lo_324};
  wire [7:0]    dataGroup_4_5 = dataGroup_lo_324[119:112];
  wire [2047:0] dataGroup_lo_325 = {dataGroup_lo_hi_325, dataGroup_lo_lo_325};
  wire [2047:0] dataGroup_hi_325 = {dataGroup_hi_hi_325, dataGroup_hi_lo_325};
  wire [7:0]    dataGroup_5_5 = dataGroup_lo_325[143:136];
  wire [2047:0] dataGroup_lo_326 = {dataGroup_lo_hi_326, dataGroup_lo_lo_326};
  wire [2047:0] dataGroup_hi_326 = {dataGroup_hi_hi_326, dataGroup_hi_lo_326};
  wire [7:0]    dataGroup_6_5 = dataGroup_lo_326[167:160];
  wire [2047:0] dataGroup_lo_327 = {dataGroup_lo_hi_327, dataGroup_lo_lo_327};
  wire [2047:0] dataGroup_hi_327 = {dataGroup_hi_hi_327, dataGroup_hi_lo_327};
  wire [7:0]    dataGroup_7_5 = dataGroup_lo_327[191:184];
  wire [2047:0] dataGroup_lo_328 = {dataGroup_lo_hi_328, dataGroup_lo_lo_328};
  wire [2047:0] dataGroup_hi_328 = {dataGroup_hi_hi_328, dataGroup_hi_lo_328};
  wire [7:0]    dataGroup_8_5 = dataGroup_lo_328[215:208];
  wire [2047:0] dataGroup_lo_329 = {dataGroup_lo_hi_329, dataGroup_lo_lo_329};
  wire [2047:0] dataGroup_hi_329 = {dataGroup_hi_hi_329, dataGroup_hi_lo_329};
  wire [7:0]    dataGroup_9_5 = dataGroup_lo_329[239:232];
  wire [2047:0] dataGroup_lo_330 = {dataGroup_lo_hi_330, dataGroup_lo_lo_330};
  wire [2047:0] dataGroup_hi_330 = {dataGroup_hi_hi_330, dataGroup_hi_lo_330};
  wire [7:0]    dataGroup_10_5 = dataGroup_lo_330[263:256];
  wire [2047:0] dataGroup_lo_331 = {dataGroup_lo_hi_331, dataGroup_lo_lo_331};
  wire [2047:0] dataGroup_hi_331 = {dataGroup_hi_hi_331, dataGroup_hi_lo_331};
  wire [7:0]    dataGroup_11_5 = dataGroup_lo_331[287:280];
  wire [2047:0] dataGroup_lo_332 = {dataGroup_lo_hi_332, dataGroup_lo_lo_332};
  wire [2047:0] dataGroup_hi_332 = {dataGroup_hi_hi_332, dataGroup_hi_lo_332};
  wire [7:0]    dataGroup_12_5 = dataGroup_lo_332[311:304];
  wire [2047:0] dataGroup_lo_333 = {dataGroup_lo_hi_333, dataGroup_lo_lo_333};
  wire [2047:0] dataGroup_hi_333 = {dataGroup_hi_hi_333, dataGroup_hi_lo_333};
  wire [7:0]    dataGroup_13_5 = dataGroup_lo_333[335:328];
  wire [2047:0] dataGroup_lo_334 = {dataGroup_lo_hi_334, dataGroup_lo_lo_334};
  wire [2047:0] dataGroup_hi_334 = {dataGroup_hi_hi_334, dataGroup_hi_lo_334};
  wire [7:0]    dataGroup_14_5 = dataGroup_lo_334[359:352];
  wire [2047:0] dataGroup_lo_335 = {dataGroup_lo_hi_335, dataGroup_lo_lo_335};
  wire [2047:0] dataGroup_hi_335 = {dataGroup_hi_hi_335, dataGroup_hi_lo_335};
  wire [7:0]    dataGroup_15_5 = dataGroup_lo_335[383:376];
  wire [2047:0] dataGroup_lo_336 = {dataGroup_lo_hi_336, dataGroup_lo_lo_336};
  wire [2047:0] dataGroup_hi_336 = {dataGroup_hi_hi_336, dataGroup_hi_lo_336};
  wire [7:0]    dataGroup_16_5 = dataGroup_lo_336[407:400];
  wire [2047:0] dataGroup_lo_337 = {dataGroup_lo_hi_337, dataGroup_lo_lo_337};
  wire [2047:0] dataGroup_hi_337 = {dataGroup_hi_hi_337, dataGroup_hi_lo_337};
  wire [7:0]    dataGroup_17_5 = dataGroup_lo_337[431:424];
  wire [2047:0] dataGroup_lo_338 = {dataGroup_lo_hi_338, dataGroup_lo_lo_338};
  wire [2047:0] dataGroup_hi_338 = {dataGroup_hi_hi_338, dataGroup_hi_lo_338};
  wire [7:0]    dataGroup_18_5 = dataGroup_lo_338[455:448];
  wire [2047:0] dataGroup_lo_339 = {dataGroup_lo_hi_339, dataGroup_lo_lo_339};
  wire [2047:0] dataGroup_hi_339 = {dataGroup_hi_hi_339, dataGroup_hi_lo_339};
  wire [7:0]    dataGroup_19_5 = dataGroup_lo_339[479:472];
  wire [2047:0] dataGroup_lo_340 = {dataGroup_lo_hi_340, dataGroup_lo_lo_340};
  wire [2047:0] dataGroup_hi_340 = {dataGroup_hi_hi_340, dataGroup_hi_lo_340};
  wire [7:0]    dataGroup_20_5 = dataGroup_lo_340[503:496];
  wire [2047:0] dataGroup_lo_341 = {dataGroup_lo_hi_341, dataGroup_lo_lo_341};
  wire [2047:0] dataGroup_hi_341 = {dataGroup_hi_hi_341, dataGroup_hi_lo_341};
  wire [7:0]    dataGroup_21_5 = dataGroup_lo_341[527:520];
  wire [2047:0] dataGroup_lo_342 = {dataGroup_lo_hi_342, dataGroup_lo_lo_342};
  wire [2047:0] dataGroup_hi_342 = {dataGroup_hi_hi_342, dataGroup_hi_lo_342};
  wire [7:0]    dataGroup_22_5 = dataGroup_lo_342[551:544];
  wire [2047:0] dataGroup_lo_343 = {dataGroup_lo_hi_343, dataGroup_lo_lo_343};
  wire [2047:0] dataGroup_hi_343 = {dataGroup_hi_hi_343, dataGroup_hi_lo_343};
  wire [7:0]    dataGroup_23_5 = dataGroup_lo_343[575:568];
  wire [2047:0] dataGroup_lo_344 = {dataGroup_lo_hi_344, dataGroup_lo_lo_344};
  wire [2047:0] dataGroup_hi_344 = {dataGroup_hi_hi_344, dataGroup_hi_lo_344};
  wire [7:0]    dataGroup_24_5 = dataGroup_lo_344[599:592];
  wire [2047:0] dataGroup_lo_345 = {dataGroup_lo_hi_345, dataGroup_lo_lo_345};
  wire [2047:0] dataGroup_hi_345 = {dataGroup_hi_hi_345, dataGroup_hi_lo_345};
  wire [7:0]    dataGroup_25_5 = dataGroup_lo_345[623:616];
  wire [2047:0] dataGroup_lo_346 = {dataGroup_lo_hi_346, dataGroup_lo_lo_346};
  wire [2047:0] dataGroup_hi_346 = {dataGroup_hi_hi_346, dataGroup_hi_lo_346};
  wire [7:0]    dataGroup_26_5 = dataGroup_lo_346[647:640];
  wire [2047:0] dataGroup_lo_347 = {dataGroup_lo_hi_347, dataGroup_lo_lo_347};
  wire [2047:0] dataGroup_hi_347 = {dataGroup_hi_hi_347, dataGroup_hi_lo_347};
  wire [7:0]    dataGroup_27_5 = dataGroup_lo_347[671:664];
  wire [2047:0] dataGroup_lo_348 = {dataGroup_lo_hi_348, dataGroup_lo_lo_348};
  wire [2047:0] dataGroup_hi_348 = {dataGroup_hi_hi_348, dataGroup_hi_lo_348};
  wire [7:0]    dataGroup_28_5 = dataGroup_lo_348[695:688];
  wire [2047:0] dataGroup_lo_349 = {dataGroup_lo_hi_349, dataGroup_lo_lo_349};
  wire [2047:0] dataGroup_hi_349 = {dataGroup_hi_hi_349, dataGroup_hi_lo_349};
  wire [7:0]    dataGroup_29_5 = dataGroup_lo_349[719:712];
  wire [2047:0] dataGroup_lo_350 = {dataGroup_lo_hi_350, dataGroup_lo_lo_350};
  wire [2047:0] dataGroup_hi_350 = {dataGroup_hi_hi_350, dataGroup_hi_lo_350};
  wire [7:0]    dataGroup_30_5 = dataGroup_lo_350[743:736];
  wire [2047:0] dataGroup_lo_351 = {dataGroup_lo_hi_351, dataGroup_lo_lo_351};
  wire [2047:0] dataGroup_hi_351 = {dataGroup_hi_hi_351, dataGroup_hi_lo_351};
  wire [7:0]    dataGroup_31_5 = dataGroup_lo_351[767:760];
  wire [2047:0] dataGroup_lo_352 = {dataGroup_lo_hi_352, dataGroup_lo_lo_352};
  wire [2047:0] dataGroup_hi_352 = {dataGroup_hi_hi_352, dataGroup_hi_lo_352};
  wire [7:0]    dataGroup_32_5 = dataGroup_lo_352[791:784];
  wire [2047:0] dataGroup_lo_353 = {dataGroup_lo_hi_353, dataGroup_lo_lo_353};
  wire [2047:0] dataGroup_hi_353 = {dataGroup_hi_hi_353, dataGroup_hi_lo_353};
  wire [7:0]    dataGroup_33_5 = dataGroup_lo_353[815:808];
  wire [2047:0] dataGroup_lo_354 = {dataGroup_lo_hi_354, dataGroup_lo_lo_354};
  wire [2047:0] dataGroup_hi_354 = {dataGroup_hi_hi_354, dataGroup_hi_lo_354};
  wire [7:0]    dataGroup_34_5 = dataGroup_lo_354[839:832];
  wire [2047:0] dataGroup_lo_355 = {dataGroup_lo_hi_355, dataGroup_lo_lo_355};
  wire [2047:0] dataGroup_hi_355 = {dataGroup_hi_hi_355, dataGroup_hi_lo_355};
  wire [7:0]    dataGroup_35_5 = dataGroup_lo_355[863:856];
  wire [2047:0] dataGroup_lo_356 = {dataGroup_lo_hi_356, dataGroup_lo_lo_356};
  wire [2047:0] dataGroup_hi_356 = {dataGroup_hi_hi_356, dataGroup_hi_lo_356};
  wire [7:0]    dataGroup_36_5 = dataGroup_lo_356[887:880];
  wire [2047:0] dataGroup_lo_357 = {dataGroup_lo_hi_357, dataGroup_lo_lo_357};
  wire [2047:0] dataGroup_hi_357 = {dataGroup_hi_hi_357, dataGroup_hi_lo_357};
  wire [7:0]    dataGroup_37_5 = dataGroup_lo_357[911:904];
  wire [2047:0] dataGroup_lo_358 = {dataGroup_lo_hi_358, dataGroup_lo_lo_358};
  wire [2047:0] dataGroup_hi_358 = {dataGroup_hi_hi_358, dataGroup_hi_lo_358};
  wire [7:0]    dataGroup_38_5 = dataGroup_lo_358[935:928];
  wire [2047:0] dataGroup_lo_359 = {dataGroup_lo_hi_359, dataGroup_lo_lo_359};
  wire [2047:0] dataGroup_hi_359 = {dataGroup_hi_hi_359, dataGroup_hi_lo_359};
  wire [7:0]    dataGroup_39_5 = dataGroup_lo_359[959:952];
  wire [2047:0] dataGroup_lo_360 = {dataGroup_lo_hi_360, dataGroup_lo_lo_360};
  wire [2047:0] dataGroup_hi_360 = {dataGroup_hi_hi_360, dataGroup_hi_lo_360};
  wire [7:0]    dataGroup_40_5 = dataGroup_lo_360[983:976];
  wire [2047:0] dataGroup_lo_361 = {dataGroup_lo_hi_361, dataGroup_lo_lo_361};
  wire [2047:0] dataGroup_hi_361 = {dataGroup_hi_hi_361, dataGroup_hi_lo_361};
  wire [7:0]    dataGroup_41_5 = dataGroup_lo_361[1007:1000];
  wire [2047:0] dataGroup_lo_362 = {dataGroup_lo_hi_362, dataGroup_lo_lo_362};
  wire [2047:0] dataGroup_hi_362 = {dataGroup_hi_hi_362, dataGroup_hi_lo_362};
  wire [7:0]    dataGroup_42_5 = dataGroup_lo_362[1031:1024];
  wire [2047:0] dataGroup_lo_363 = {dataGroup_lo_hi_363, dataGroup_lo_lo_363};
  wire [2047:0] dataGroup_hi_363 = {dataGroup_hi_hi_363, dataGroup_hi_lo_363};
  wire [7:0]    dataGroup_43_5 = dataGroup_lo_363[1055:1048];
  wire [2047:0] dataGroup_lo_364 = {dataGroup_lo_hi_364, dataGroup_lo_lo_364};
  wire [2047:0] dataGroup_hi_364 = {dataGroup_hi_hi_364, dataGroup_hi_lo_364};
  wire [7:0]    dataGroup_44_5 = dataGroup_lo_364[1079:1072];
  wire [2047:0] dataGroup_lo_365 = {dataGroup_lo_hi_365, dataGroup_lo_lo_365};
  wire [2047:0] dataGroup_hi_365 = {dataGroup_hi_hi_365, dataGroup_hi_lo_365};
  wire [7:0]    dataGroup_45_5 = dataGroup_lo_365[1103:1096];
  wire [2047:0] dataGroup_lo_366 = {dataGroup_lo_hi_366, dataGroup_lo_lo_366};
  wire [2047:0] dataGroup_hi_366 = {dataGroup_hi_hi_366, dataGroup_hi_lo_366};
  wire [7:0]    dataGroup_46_5 = dataGroup_lo_366[1127:1120];
  wire [2047:0] dataGroup_lo_367 = {dataGroup_lo_hi_367, dataGroup_lo_lo_367};
  wire [2047:0] dataGroup_hi_367 = {dataGroup_hi_hi_367, dataGroup_hi_lo_367};
  wire [7:0]    dataGroup_47_5 = dataGroup_lo_367[1151:1144];
  wire [2047:0] dataGroup_lo_368 = {dataGroup_lo_hi_368, dataGroup_lo_lo_368};
  wire [2047:0] dataGroup_hi_368 = {dataGroup_hi_hi_368, dataGroup_hi_lo_368};
  wire [7:0]    dataGroup_48_5 = dataGroup_lo_368[1175:1168];
  wire [2047:0] dataGroup_lo_369 = {dataGroup_lo_hi_369, dataGroup_lo_lo_369};
  wire [2047:0] dataGroup_hi_369 = {dataGroup_hi_hi_369, dataGroup_hi_lo_369};
  wire [7:0]    dataGroup_49_5 = dataGroup_lo_369[1199:1192];
  wire [2047:0] dataGroup_lo_370 = {dataGroup_lo_hi_370, dataGroup_lo_lo_370};
  wire [2047:0] dataGroup_hi_370 = {dataGroup_hi_hi_370, dataGroup_hi_lo_370};
  wire [7:0]    dataGroup_50_5 = dataGroup_lo_370[1223:1216];
  wire [2047:0] dataGroup_lo_371 = {dataGroup_lo_hi_371, dataGroup_lo_lo_371};
  wire [2047:0] dataGroup_hi_371 = {dataGroup_hi_hi_371, dataGroup_hi_lo_371};
  wire [7:0]    dataGroup_51_5 = dataGroup_lo_371[1247:1240];
  wire [2047:0] dataGroup_lo_372 = {dataGroup_lo_hi_372, dataGroup_lo_lo_372};
  wire [2047:0] dataGroup_hi_372 = {dataGroup_hi_hi_372, dataGroup_hi_lo_372};
  wire [7:0]    dataGroup_52_5 = dataGroup_lo_372[1271:1264];
  wire [2047:0] dataGroup_lo_373 = {dataGroup_lo_hi_373, dataGroup_lo_lo_373};
  wire [2047:0] dataGroup_hi_373 = {dataGroup_hi_hi_373, dataGroup_hi_lo_373};
  wire [7:0]    dataGroup_53_5 = dataGroup_lo_373[1295:1288];
  wire [2047:0] dataGroup_lo_374 = {dataGroup_lo_hi_374, dataGroup_lo_lo_374};
  wire [2047:0] dataGroup_hi_374 = {dataGroup_hi_hi_374, dataGroup_hi_lo_374};
  wire [7:0]    dataGroup_54_5 = dataGroup_lo_374[1319:1312];
  wire [2047:0] dataGroup_lo_375 = {dataGroup_lo_hi_375, dataGroup_lo_lo_375};
  wire [2047:0] dataGroup_hi_375 = {dataGroup_hi_hi_375, dataGroup_hi_lo_375};
  wire [7:0]    dataGroup_55_5 = dataGroup_lo_375[1343:1336];
  wire [2047:0] dataGroup_lo_376 = {dataGroup_lo_hi_376, dataGroup_lo_lo_376};
  wire [2047:0] dataGroup_hi_376 = {dataGroup_hi_hi_376, dataGroup_hi_lo_376};
  wire [7:0]    dataGroup_56_5 = dataGroup_lo_376[1367:1360];
  wire [2047:0] dataGroup_lo_377 = {dataGroup_lo_hi_377, dataGroup_lo_lo_377};
  wire [2047:0] dataGroup_hi_377 = {dataGroup_hi_hi_377, dataGroup_hi_lo_377};
  wire [7:0]    dataGroup_57_5 = dataGroup_lo_377[1391:1384];
  wire [2047:0] dataGroup_lo_378 = {dataGroup_lo_hi_378, dataGroup_lo_lo_378};
  wire [2047:0] dataGroup_hi_378 = {dataGroup_hi_hi_378, dataGroup_hi_lo_378};
  wire [7:0]    dataGroup_58_5 = dataGroup_lo_378[1415:1408];
  wire [2047:0] dataGroup_lo_379 = {dataGroup_lo_hi_379, dataGroup_lo_lo_379};
  wire [2047:0] dataGroup_hi_379 = {dataGroup_hi_hi_379, dataGroup_hi_lo_379};
  wire [7:0]    dataGroup_59_5 = dataGroup_lo_379[1439:1432];
  wire [2047:0] dataGroup_lo_380 = {dataGroup_lo_hi_380, dataGroup_lo_lo_380};
  wire [2047:0] dataGroup_hi_380 = {dataGroup_hi_hi_380, dataGroup_hi_lo_380};
  wire [7:0]    dataGroup_60_5 = dataGroup_lo_380[1463:1456];
  wire [2047:0] dataGroup_lo_381 = {dataGroup_lo_hi_381, dataGroup_lo_lo_381};
  wire [2047:0] dataGroup_hi_381 = {dataGroup_hi_hi_381, dataGroup_hi_lo_381};
  wire [7:0]    dataGroup_61_5 = dataGroup_lo_381[1487:1480];
  wire [2047:0] dataGroup_lo_382 = {dataGroup_lo_hi_382, dataGroup_lo_lo_382};
  wire [2047:0] dataGroup_hi_382 = {dataGroup_hi_hi_382, dataGroup_hi_lo_382};
  wire [7:0]    dataGroup_62_5 = dataGroup_lo_382[1511:1504];
  wire [2047:0] dataGroup_lo_383 = {dataGroup_lo_hi_383, dataGroup_lo_lo_383};
  wire [2047:0] dataGroup_hi_383 = {dataGroup_hi_hi_383, dataGroup_hi_lo_383};
  wire [7:0]    dataGroup_63_5 = dataGroup_lo_383[1535:1528];
  wire [15:0]   res_lo_lo_lo_lo_lo_5 = {dataGroup_1_5, dataGroup_0_5};
  wire [15:0]   res_lo_lo_lo_lo_hi_5 = {dataGroup_3_5, dataGroup_2_5};
  wire [31:0]   res_lo_lo_lo_lo_5 = {res_lo_lo_lo_lo_hi_5, res_lo_lo_lo_lo_lo_5};
  wire [15:0]   res_lo_lo_lo_hi_lo_5 = {dataGroup_5_5, dataGroup_4_5};
  wire [15:0]   res_lo_lo_lo_hi_hi_5 = {dataGroup_7_5, dataGroup_6_5};
  wire [31:0]   res_lo_lo_lo_hi_5 = {res_lo_lo_lo_hi_hi_5, res_lo_lo_lo_hi_lo_5};
  wire [63:0]   res_lo_lo_lo_5 = {res_lo_lo_lo_hi_5, res_lo_lo_lo_lo_5};
  wire [15:0]   res_lo_lo_hi_lo_lo_5 = {dataGroup_9_5, dataGroup_8_5};
  wire [15:0]   res_lo_lo_hi_lo_hi_5 = {dataGroup_11_5, dataGroup_10_5};
  wire [31:0]   res_lo_lo_hi_lo_5 = {res_lo_lo_hi_lo_hi_5, res_lo_lo_hi_lo_lo_5};
  wire [15:0]   res_lo_lo_hi_hi_lo_5 = {dataGroup_13_5, dataGroup_12_5};
  wire [15:0]   res_lo_lo_hi_hi_hi_5 = {dataGroup_15_5, dataGroup_14_5};
  wire [31:0]   res_lo_lo_hi_hi_5 = {res_lo_lo_hi_hi_hi_5, res_lo_lo_hi_hi_lo_5};
  wire [63:0]   res_lo_lo_hi_5 = {res_lo_lo_hi_hi_5, res_lo_lo_hi_lo_5};
  wire [127:0]  res_lo_lo_5 = {res_lo_lo_hi_5, res_lo_lo_lo_5};
  wire [15:0]   res_lo_hi_lo_lo_lo_5 = {dataGroup_17_5, dataGroup_16_5};
  wire [15:0]   res_lo_hi_lo_lo_hi_5 = {dataGroup_19_5, dataGroup_18_5};
  wire [31:0]   res_lo_hi_lo_lo_5 = {res_lo_hi_lo_lo_hi_5, res_lo_hi_lo_lo_lo_5};
  wire [15:0]   res_lo_hi_lo_hi_lo_5 = {dataGroup_21_5, dataGroup_20_5};
  wire [15:0]   res_lo_hi_lo_hi_hi_5 = {dataGroup_23_5, dataGroup_22_5};
  wire [31:0]   res_lo_hi_lo_hi_5 = {res_lo_hi_lo_hi_hi_5, res_lo_hi_lo_hi_lo_5};
  wire [63:0]   res_lo_hi_lo_5 = {res_lo_hi_lo_hi_5, res_lo_hi_lo_lo_5};
  wire [15:0]   res_lo_hi_hi_lo_lo_5 = {dataGroup_25_5, dataGroup_24_5};
  wire [15:0]   res_lo_hi_hi_lo_hi_5 = {dataGroup_27_5, dataGroup_26_5};
  wire [31:0]   res_lo_hi_hi_lo_5 = {res_lo_hi_hi_lo_hi_5, res_lo_hi_hi_lo_lo_5};
  wire [15:0]   res_lo_hi_hi_hi_lo_5 = {dataGroup_29_5, dataGroup_28_5};
  wire [15:0]   res_lo_hi_hi_hi_hi_5 = {dataGroup_31_5, dataGroup_30_5};
  wire [31:0]   res_lo_hi_hi_hi_5 = {res_lo_hi_hi_hi_hi_5, res_lo_hi_hi_hi_lo_5};
  wire [63:0]   res_lo_hi_hi_5 = {res_lo_hi_hi_hi_5, res_lo_hi_hi_lo_5};
  wire [127:0]  res_lo_hi_5 = {res_lo_hi_hi_5, res_lo_hi_lo_5};
  wire [255:0]  res_lo_5 = {res_lo_hi_5, res_lo_lo_5};
  wire [15:0]   res_hi_lo_lo_lo_lo_5 = {dataGroup_33_5, dataGroup_32_5};
  wire [15:0]   res_hi_lo_lo_lo_hi_5 = {dataGroup_35_5, dataGroup_34_5};
  wire [31:0]   res_hi_lo_lo_lo_5 = {res_hi_lo_lo_lo_hi_5, res_hi_lo_lo_lo_lo_5};
  wire [15:0]   res_hi_lo_lo_hi_lo_5 = {dataGroup_37_5, dataGroup_36_5};
  wire [15:0]   res_hi_lo_lo_hi_hi_5 = {dataGroup_39_5, dataGroup_38_5};
  wire [31:0]   res_hi_lo_lo_hi_5 = {res_hi_lo_lo_hi_hi_5, res_hi_lo_lo_hi_lo_5};
  wire [63:0]   res_hi_lo_lo_5 = {res_hi_lo_lo_hi_5, res_hi_lo_lo_lo_5};
  wire [15:0]   res_hi_lo_hi_lo_lo_5 = {dataGroup_41_5, dataGroup_40_5};
  wire [15:0]   res_hi_lo_hi_lo_hi_5 = {dataGroup_43_5, dataGroup_42_5};
  wire [31:0]   res_hi_lo_hi_lo_5 = {res_hi_lo_hi_lo_hi_5, res_hi_lo_hi_lo_lo_5};
  wire [15:0]   res_hi_lo_hi_hi_lo_5 = {dataGroup_45_5, dataGroup_44_5};
  wire [15:0]   res_hi_lo_hi_hi_hi_5 = {dataGroup_47_5, dataGroup_46_5};
  wire [31:0]   res_hi_lo_hi_hi_5 = {res_hi_lo_hi_hi_hi_5, res_hi_lo_hi_hi_lo_5};
  wire [63:0]   res_hi_lo_hi_5 = {res_hi_lo_hi_hi_5, res_hi_lo_hi_lo_5};
  wire [127:0]  res_hi_lo_5 = {res_hi_lo_hi_5, res_hi_lo_lo_5};
  wire [15:0]   res_hi_hi_lo_lo_lo_5 = {dataGroup_49_5, dataGroup_48_5};
  wire [15:0]   res_hi_hi_lo_lo_hi_5 = {dataGroup_51_5, dataGroup_50_5};
  wire [31:0]   res_hi_hi_lo_lo_5 = {res_hi_hi_lo_lo_hi_5, res_hi_hi_lo_lo_lo_5};
  wire [15:0]   res_hi_hi_lo_hi_lo_5 = {dataGroup_53_5, dataGroup_52_5};
  wire [15:0]   res_hi_hi_lo_hi_hi_5 = {dataGroup_55_5, dataGroup_54_5};
  wire [31:0]   res_hi_hi_lo_hi_5 = {res_hi_hi_lo_hi_hi_5, res_hi_hi_lo_hi_lo_5};
  wire [63:0]   res_hi_hi_lo_5 = {res_hi_hi_lo_hi_5, res_hi_hi_lo_lo_5};
  wire [15:0]   res_hi_hi_hi_lo_lo_5 = {dataGroup_57_5, dataGroup_56_5};
  wire [15:0]   res_hi_hi_hi_lo_hi_5 = {dataGroup_59_5, dataGroup_58_5};
  wire [31:0]   res_hi_hi_hi_lo_5 = {res_hi_hi_hi_lo_hi_5, res_hi_hi_hi_lo_lo_5};
  wire [15:0]   res_hi_hi_hi_hi_lo_5 = {dataGroup_61_5, dataGroup_60_5};
  wire [15:0]   res_hi_hi_hi_hi_hi_5 = {dataGroup_63_5, dataGroup_62_5};
  wire [31:0]   res_hi_hi_hi_hi_5 = {res_hi_hi_hi_hi_hi_5, res_hi_hi_hi_hi_lo_5};
  wire [63:0]   res_hi_hi_hi_5 = {res_hi_hi_hi_hi_5, res_hi_hi_hi_lo_5};
  wire [127:0]  res_hi_hi_5 = {res_hi_hi_hi_5, res_hi_hi_lo_5};
  wire [255:0]  res_hi_5 = {res_hi_hi_5, res_hi_lo_5};
  wire [511:0]  res_18 = {res_hi_5, res_lo_5};
  wire [1023:0] lo_lo_2 = {res_17, res_16};
  wire [1023:0] lo_hi_2 = {512'h0, res_18};
  wire [2047:0] lo_2 = {lo_hi_2, lo_lo_2};
  wire [4095:0] regroupLoadData_0_2 = {2048'h0, lo_2};
  wire [2047:0] dataGroup_lo_384 = {dataGroup_lo_hi_384, dataGroup_lo_lo_384};
  wire [2047:0] dataGroup_hi_384 = {dataGroup_hi_hi_384, dataGroup_hi_lo_384};
  wire [7:0]    dataGroup_0_6 = dataGroup_lo_384[7:0];
  wire [2047:0] dataGroup_lo_385 = {dataGroup_lo_hi_385, dataGroup_lo_lo_385};
  wire [2047:0] dataGroup_hi_385 = {dataGroup_hi_hi_385, dataGroup_hi_lo_385};
  wire [7:0]    dataGroup_1_6 = dataGroup_lo_385[39:32];
  wire [2047:0] dataGroup_lo_386 = {dataGroup_lo_hi_386, dataGroup_lo_lo_386};
  wire [2047:0] dataGroup_hi_386 = {dataGroup_hi_hi_386, dataGroup_hi_lo_386};
  wire [7:0]    dataGroup_2_6 = dataGroup_lo_386[71:64];
  wire [2047:0] dataGroup_lo_387 = {dataGroup_lo_hi_387, dataGroup_lo_lo_387};
  wire [2047:0] dataGroup_hi_387 = {dataGroup_hi_hi_387, dataGroup_hi_lo_387};
  wire [7:0]    dataGroup_3_6 = dataGroup_lo_387[103:96];
  wire [2047:0] dataGroup_lo_388 = {dataGroup_lo_hi_388, dataGroup_lo_lo_388};
  wire [2047:0] dataGroup_hi_388 = {dataGroup_hi_hi_388, dataGroup_hi_lo_388};
  wire [7:0]    dataGroup_4_6 = dataGroup_lo_388[135:128];
  wire [2047:0] dataGroup_lo_389 = {dataGroup_lo_hi_389, dataGroup_lo_lo_389};
  wire [2047:0] dataGroup_hi_389 = {dataGroup_hi_hi_389, dataGroup_hi_lo_389};
  wire [7:0]    dataGroup_5_6 = dataGroup_lo_389[167:160];
  wire [2047:0] dataGroup_lo_390 = {dataGroup_lo_hi_390, dataGroup_lo_lo_390};
  wire [2047:0] dataGroup_hi_390 = {dataGroup_hi_hi_390, dataGroup_hi_lo_390};
  wire [7:0]    dataGroup_6_6 = dataGroup_lo_390[199:192];
  wire [2047:0] dataGroup_lo_391 = {dataGroup_lo_hi_391, dataGroup_lo_lo_391};
  wire [2047:0] dataGroup_hi_391 = {dataGroup_hi_hi_391, dataGroup_hi_lo_391};
  wire [7:0]    dataGroup_7_6 = dataGroup_lo_391[231:224];
  wire [2047:0] dataGroup_lo_392 = {dataGroup_lo_hi_392, dataGroup_lo_lo_392};
  wire [2047:0] dataGroup_hi_392 = {dataGroup_hi_hi_392, dataGroup_hi_lo_392};
  wire [7:0]    dataGroup_8_6 = dataGroup_lo_392[263:256];
  wire [2047:0] dataGroup_lo_393 = {dataGroup_lo_hi_393, dataGroup_lo_lo_393};
  wire [2047:0] dataGroup_hi_393 = {dataGroup_hi_hi_393, dataGroup_hi_lo_393};
  wire [7:0]    dataGroup_9_6 = dataGroup_lo_393[295:288];
  wire [2047:0] dataGroup_lo_394 = {dataGroup_lo_hi_394, dataGroup_lo_lo_394};
  wire [2047:0] dataGroup_hi_394 = {dataGroup_hi_hi_394, dataGroup_hi_lo_394};
  wire [7:0]    dataGroup_10_6 = dataGroup_lo_394[327:320];
  wire [2047:0] dataGroup_lo_395 = {dataGroup_lo_hi_395, dataGroup_lo_lo_395};
  wire [2047:0] dataGroup_hi_395 = {dataGroup_hi_hi_395, dataGroup_hi_lo_395};
  wire [7:0]    dataGroup_11_6 = dataGroup_lo_395[359:352];
  wire [2047:0] dataGroup_lo_396 = {dataGroup_lo_hi_396, dataGroup_lo_lo_396};
  wire [2047:0] dataGroup_hi_396 = {dataGroup_hi_hi_396, dataGroup_hi_lo_396};
  wire [7:0]    dataGroup_12_6 = dataGroup_lo_396[391:384];
  wire [2047:0] dataGroup_lo_397 = {dataGroup_lo_hi_397, dataGroup_lo_lo_397};
  wire [2047:0] dataGroup_hi_397 = {dataGroup_hi_hi_397, dataGroup_hi_lo_397};
  wire [7:0]    dataGroup_13_6 = dataGroup_lo_397[423:416];
  wire [2047:0] dataGroup_lo_398 = {dataGroup_lo_hi_398, dataGroup_lo_lo_398};
  wire [2047:0] dataGroup_hi_398 = {dataGroup_hi_hi_398, dataGroup_hi_lo_398};
  wire [7:0]    dataGroup_14_6 = dataGroup_lo_398[455:448];
  wire [2047:0] dataGroup_lo_399 = {dataGroup_lo_hi_399, dataGroup_lo_lo_399};
  wire [2047:0] dataGroup_hi_399 = {dataGroup_hi_hi_399, dataGroup_hi_lo_399};
  wire [7:0]    dataGroup_15_6 = dataGroup_lo_399[487:480];
  wire [2047:0] dataGroup_lo_400 = {dataGroup_lo_hi_400, dataGroup_lo_lo_400};
  wire [2047:0] dataGroup_hi_400 = {dataGroup_hi_hi_400, dataGroup_hi_lo_400};
  wire [7:0]    dataGroup_16_6 = dataGroup_lo_400[519:512];
  wire [2047:0] dataGroup_lo_401 = {dataGroup_lo_hi_401, dataGroup_lo_lo_401};
  wire [2047:0] dataGroup_hi_401 = {dataGroup_hi_hi_401, dataGroup_hi_lo_401};
  wire [7:0]    dataGroup_17_6 = dataGroup_lo_401[551:544];
  wire [2047:0] dataGroup_lo_402 = {dataGroup_lo_hi_402, dataGroup_lo_lo_402};
  wire [2047:0] dataGroup_hi_402 = {dataGroup_hi_hi_402, dataGroup_hi_lo_402};
  wire [7:0]    dataGroup_18_6 = dataGroup_lo_402[583:576];
  wire [2047:0] dataGroup_lo_403 = {dataGroup_lo_hi_403, dataGroup_lo_lo_403};
  wire [2047:0] dataGroup_hi_403 = {dataGroup_hi_hi_403, dataGroup_hi_lo_403};
  wire [7:0]    dataGroup_19_6 = dataGroup_lo_403[615:608];
  wire [2047:0] dataGroup_lo_404 = {dataGroup_lo_hi_404, dataGroup_lo_lo_404};
  wire [2047:0] dataGroup_hi_404 = {dataGroup_hi_hi_404, dataGroup_hi_lo_404};
  wire [7:0]    dataGroup_20_6 = dataGroup_lo_404[647:640];
  wire [2047:0] dataGroup_lo_405 = {dataGroup_lo_hi_405, dataGroup_lo_lo_405};
  wire [2047:0] dataGroup_hi_405 = {dataGroup_hi_hi_405, dataGroup_hi_lo_405};
  wire [7:0]    dataGroup_21_6 = dataGroup_lo_405[679:672];
  wire [2047:0] dataGroup_lo_406 = {dataGroup_lo_hi_406, dataGroup_lo_lo_406};
  wire [2047:0] dataGroup_hi_406 = {dataGroup_hi_hi_406, dataGroup_hi_lo_406};
  wire [7:0]    dataGroup_22_6 = dataGroup_lo_406[711:704];
  wire [2047:0] dataGroup_lo_407 = {dataGroup_lo_hi_407, dataGroup_lo_lo_407};
  wire [2047:0] dataGroup_hi_407 = {dataGroup_hi_hi_407, dataGroup_hi_lo_407};
  wire [7:0]    dataGroup_23_6 = dataGroup_lo_407[743:736];
  wire [2047:0] dataGroup_lo_408 = {dataGroup_lo_hi_408, dataGroup_lo_lo_408};
  wire [2047:0] dataGroup_hi_408 = {dataGroup_hi_hi_408, dataGroup_hi_lo_408};
  wire [7:0]    dataGroup_24_6 = dataGroup_lo_408[775:768];
  wire [2047:0] dataGroup_lo_409 = {dataGroup_lo_hi_409, dataGroup_lo_lo_409};
  wire [2047:0] dataGroup_hi_409 = {dataGroup_hi_hi_409, dataGroup_hi_lo_409};
  wire [7:0]    dataGroup_25_6 = dataGroup_lo_409[807:800];
  wire [2047:0] dataGroup_lo_410 = {dataGroup_lo_hi_410, dataGroup_lo_lo_410};
  wire [2047:0] dataGroup_hi_410 = {dataGroup_hi_hi_410, dataGroup_hi_lo_410};
  wire [7:0]    dataGroup_26_6 = dataGroup_lo_410[839:832];
  wire [2047:0] dataGroup_lo_411 = {dataGroup_lo_hi_411, dataGroup_lo_lo_411};
  wire [2047:0] dataGroup_hi_411 = {dataGroup_hi_hi_411, dataGroup_hi_lo_411};
  wire [7:0]    dataGroup_27_6 = dataGroup_lo_411[871:864];
  wire [2047:0] dataGroup_lo_412 = {dataGroup_lo_hi_412, dataGroup_lo_lo_412};
  wire [2047:0] dataGroup_hi_412 = {dataGroup_hi_hi_412, dataGroup_hi_lo_412};
  wire [7:0]    dataGroup_28_6 = dataGroup_lo_412[903:896];
  wire [2047:0] dataGroup_lo_413 = {dataGroup_lo_hi_413, dataGroup_lo_lo_413};
  wire [2047:0] dataGroup_hi_413 = {dataGroup_hi_hi_413, dataGroup_hi_lo_413};
  wire [7:0]    dataGroup_29_6 = dataGroup_lo_413[935:928];
  wire [2047:0] dataGroup_lo_414 = {dataGroup_lo_hi_414, dataGroup_lo_lo_414};
  wire [2047:0] dataGroup_hi_414 = {dataGroup_hi_hi_414, dataGroup_hi_lo_414};
  wire [7:0]    dataGroup_30_6 = dataGroup_lo_414[967:960];
  wire [2047:0] dataGroup_lo_415 = {dataGroup_lo_hi_415, dataGroup_lo_lo_415};
  wire [2047:0] dataGroup_hi_415 = {dataGroup_hi_hi_415, dataGroup_hi_lo_415};
  wire [7:0]    dataGroup_31_6 = dataGroup_lo_415[999:992];
  wire [2047:0] dataGroup_lo_416 = {dataGroup_lo_hi_416, dataGroup_lo_lo_416};
  wire [2047:0] dataGroup_hi_416 = {dataGroup_hi_hi_416, dataGroup_hi_lo_416};
  wire [7:0]    dataGroup_32_6 = dataGroup_lo_416[1031:1024];
  wire [2047:0] dataGroup_lo_417 = {dataGroup_lo_hi_417, dataGroup_lo_lo_417};
  wire [2047:0] dataGroup_hi_417 = {dataGroup_hi_hi_417, dataGroup_hi_lo_417};
  wire [7:0]    dataGroup_33_6 = dataGroup_lo_417[1063:1056];
  wire [2047:0] dataGroup_lo_418 = {dataGroup_lo_hi_418, dataGroup_lo_lo_418};
  wire [2047:0] dataGroup_hi_418 = {dataGroup_hi_hi_418, dataGroup_hi_lo_418};
  wire [7:0]    dataGroup_34_6 = dataGroup_lo_418[1095:1088];
  wire [2047:0] dataGroup_lo_419 = {dataGroup_lo_hi_419, dataGroup_lo_lo_419};
  wire [2047:0] dataGroup_hi_419 = {dataGroup_hi_hi_419, dataGroup_hi_lo_419};
  wire [7:0]    dataGroup_35_6 = dataGroup_lo_419[1127:1120];
  wire [2047:0] dataGroup_lo_420 = {dataGroup_lo_hi_420, dataGroup_lo_lo_420};
  wire [2047:0] dataGroup_hi_420 = {dataGroup_hi_hi_420, dataGroup_hi_lo_420};
  wire [7:0]    dataGroup_36_6 = dataGroup_lo_420[1159:1152];
  wire [2047:0] dataGroup_lo_421 = {dataGroup_lo_hi_421, dataGroup_lo_lo_421};
  wire [2047:0] dataGroup_hi_421 = {dataGroup_hi_hi_421, dataGroup_hi_lo_421};
  wire [7:0]    dataGroup_37_6 = dataGroup_lo_421[1191:1184];
  wire [2047:0] dataGroup_lo_422 = {dataGroup_lo_hi_422, dataGroup_lo_lo_422};
  wire [2047:0] dataGroup_hi_422 = {dataGroup_hi_hi_422, dataGroup_hi_lo_422};
  wire [7:0]    dataGroup_38_6 = dataGroup_lo_422[1223:1216];
  wire [2047:0] dataGroup_lo_423 = {dataGroup_lo_hi_423, dataGroup_lo_lo_423};
  wire [2047:0] dataGroup_hi_423 = {dataGroup_hi_hi_423, dataGroup_hi_lo_423};
  wire [7:0]    dataGroup_39_6 = dataGroup_lo_423[1255:1248];
  wire [2047:0] dataGroup_lo_424 = {dataGroup_lo_hi_424, dataGroup_lo_lo_424};
  wire [2047:0] dataGroup_hi_424 = {dataGroup_hi_hi_424, dataGroup_hi_lo_424};
  wire [7:0]    dataGroup_40_6 = dataGroup_lo_424[1287:1280];
  wire [2047:0] dataGroup_lo_425 = {dataGroup_lo_hi_425, dataGroup_lo_lo_425};
  wire [2047:0] dataGroup_hi_425 = {dataGroup_hi_hi_425, dataGroup_hi_lo_425};
  wire [7:0]    dataGroup_41_6 = dataGroup_lo_425[1319:1312];
  wire [2047:0] dataGroup_lo_426 = {dataGroup_lo_hi_426, dataGroup_lo_lo_426};
  wire [2047:0] dataGroup_hi_426 = {dataGroup_hi_hi_426, dataGroup_hi_lo_426};
  wire [7:0]    dataGroup_42_6 = dataGroup_lo_426[1351:1344];
  wire [2047:0] dataGroup_lo_427 = {dataGroup_lo_hi_427, dataGroup_lo_lo_427};
  wire [2047:0] dataGroup_hi_427 = {dataGroup_hi_hi_427, dataGroup_hi_lo_427};
  wire [7:0]    dataGroup_43_6 = dataGroup_lo_427[1383:1376];
  wire [2047:0] dataGroup_lo_428 = {dataGroup_lo_hi_428, dataGroup_lo_lo_428};
  wire [2047:0] dataGroup_hi_428 = {dataGroup_hi_hi_428, dataGroup_hi_lo_428};
  wire [7:0]    dataGroup_44_6 = dataGroup_lo_428[1415:1408];
  wire [2047:0] dataGroup_lo_429 = {dataGroup_lo_hi_429, dataGroup_lo_lo_429};
  wire [2047:0] dataGroup_hi_429 = {dataGroup_hi_hi_429, dataGroup_hi_lo_429};
  wire [7:0]    dataGroup_45_6 = dataGroup_lo_429[1447:1440];
  wire [2047:0] dataGroup_lo_430 = {dataGroup_lo_hi_430, dataGroup_lo_lo_430};
  wire [2047:0] dataGroup_hi_430 = {dataGroup_hi_hi_430, dataGroup_hi_lo_430};
  wire [7:0]    dataGroup_46_6 = dataGroup_lo_430[1479:1472];
  wire [2047:0] dataGroup_lo_431 = {dataGroup_lo_hi_431, dataGroup_lo_lo_431};
  wire [2047:0] dataGroup_hi_431 = {dataGroup_hi_hi_431, dataGroup_hi_lo_431};
  wire [7:0]    dataGroup_47_6 = dataGroup_lo_431[1511:1504];
  wire [2047:0] dataGroup_lo_432 = {dataGroup_lo_hi_432, dataGroup_lo_lo_432};
  wire [2047:0] dataGroup_hi_432 = {dataGroup_hi_hi_432, dataGroup_hi_lo_432};
  wire [7:0]    dataGroup_48_6 = dataGroup_lo_432[1543:1536];
  wire [2047:0] dataGroup_lo_433 = {dataGroup_lo_hi_433, dataGroup_lo_lo_433};
  wire [2047:0] dataGroup_hi_433 = {dataGroup_hi_hi_433, dataGroup_hi_lo_433};
  wire [7:0]    dataGroup_49_6 = dataGroup_lo_433[1575:1568];
  wire [2047:0] dataGroup_lo_434 = {dataGroup_lo_hi_434, dataGroup_lo_lo_434};
  wire [2047:0] dataGroup_hi_434 = {dataGroup_hi_hi_434, dataGroup_hi_lo_434};
  wire [7:0]    dataGroup_50_6 = dataGroup_lo_434[1607:1600];
  wire [2047:0] dataGroup_lo_435 = {dataGroup_lo_hi_435, dataGroup_lo_lo_435};
  wire [2047:0] dataGroup_hi_435 = {dataGroup_hi_hi_435, dataGroup_hi_lo_435};
  wire [7:0]    dataGroup_51_6 = dataGroup_lo_435[1639:1632];
  wire [2047:0] dataGroup_lo_436 = {dataGroup_lo_hi_436, dataGroup_lo_lo_436};
  wire [2047:0] dataGroup_hi_436 = {dataGroup_hi_hi_436, dataGroup_hi_lo_436};
  wire [7:0]    dataGroup_52_6 = dataGroup_lo_436[1671:1664];
  wire [2047:0] dataGroup_lo_437 = {dataGroup_lo_hi_437, dataGroup_lo_lo_437};
  wire [2047:0] dataGroup_hi_437 = {dataGroup_hi_hi_437, dataGroup_hi_lo_437};
  wire [7:0]    dataGroup_53_6 = dataGroup_lo_437[1703:1696];
  wire [2047:0] dataGroup_lo_438 = {dataGroup_lo_hi_438, dataGroup_lo_lo_438};
  wire [2047:0] dataGroup_hi_438 = {dataGroup_hi_hi_438, dataGroup_hi_lo_438};
  wire [7:0]    dataGroup_54_6 = dataGroup_lo_438[1735:1728];
  wire [2047:0] dataGroup_lo_439 = {dataGroup_lo_hi_439, dataGroup_lo_lo_439};
  wire [2047:0] dataGroup_hi_439 = {dataGroup_hi_hi_439, dataGroup_hi_lo_439};
  wire [7:0]    dataGroup_55_6 = dataGroup_lo_439[1767:1760];
  wire [2047:0] dataGroup_lo_440 = {dataGroup_lo_hi_440, dataGroup_lo_lo_440};
  wire [2047:0] dataGroup_hi_440 = {dataGroup_hi_hi_440, dataGroup_hi_lo_440};
  wire [7:0]    dataGroup_56_6 = dataGroup_lo_440[1799:1792];
  wire [2047:0] dataGroup_lo_441 = {dataGroup_lo_hi_441, dataGroup_lo_lo_441};
  wire [2047:0] dataGroup_hi_441 = {dataGroup_hi_hi_441, dataGroup_hi_lo_441};
  wire [7:0]    dataGroup_57_6 = dataGroup_lo_441[1831:1824];
  wire [2047:0] dataGroup_lo_442 = {dataGroup_lo_hi_442, dataGroup_lo_lo_442};
  wire [2047:0] dataGroup_hi_442 = {dataGroup_hi_hi_442, dataGroup_hi_lo_442};
  wire [7:0]    dataGroup_58_6 = dataGroup_lo_442[1863:1856];
  wire [2047:0] dataGroup_lo_443 = {dataGroup_lo_hi_443, dataGroup_lo_lo_443};
  wire [2047:0] dataGroup_hi_443 = {dataGroup_hi_hi_443, dataGroup_hi_lo_443};
  wire [7:0]    dataGroup_59_6 = dataGroup_lo_443[1895:1888];
  wire [2047:0] dataGroup_lo_444 = {dataGroup_lo_hi_444, dataGroup_lo_lo_444};
  wire [2047:0] dataGroup_hi_444 = {dataGroup_hi_hi_444, dataGroup_hi_lo_444};
  wire [7:0]    dataGroup_60_6 = dataGroup_lo_444[1927:1920];
  wire [2047:0] dataGroup_lo_445 = {dataGroup_lo_hi_445, dataGroup_lo_lo_445};
  wire [2047:0] dataGroup_hi_445 = {dataGroup_hi_hi_445, dataGroup_hi_lo_445};
  wire [7:0]    dataGroup_61_6 = dataGroup_lo_445[1959:1952];
  wire [2047:0] dataGroup_lo_446 = {dataGroup_lo_hi_446, dataGroup_lo_lo_446};
  wire [2047:0] dataGroup_hi_446 = {dataGroup_hi_hi_446, dataGroup_hi_lo_446};
  wire [7:0]    dataGroup_62_6 = dataGroup_lo_446[1991:1984];
  wire [2047:0] dataGroup_lo_447 = {dataGroup_lo_hi_447, dataGroup_lo_lo_447};
  wire [2047:0] dataGroup_hi_447 = {dataGroup_hi_hi_447, dataGroup_hi_lo_447};
  wire [7:0]    dataGroup_63_6 = dataGroup_lo_447[2023:2016];
  wire [15:0]   res_lo_lo_lo_lo_lo_6 = {dataGroup_1_6, dataGroup_0_6};
  wire [15:0]   res_lo_lo_lo_lo_hi_6 = {dataGroup_3_6, dataGroup_2_6};
  wire [31:0]   res_lo_lo_lo_lo_6 = {res_lo_lo_lo_lo_hi_6, res_lo_lo_lo_lo_lo_6};
  wire [15:0]   res_lo_lo_lo_hi_lo_6 = {dataGroup_5_6, dataGroup_4_6};
  wire [15:0]   res_lo_lo_lo_hi_hi_6 = {dataGroup_7_6, dataGroup_6_6};
  wire [31:0]   res_lo_lo_lo_hi_6 = {res_lo_lo_lo_hi_hi_6, res_lo_lo_lo_hi_lo_6};
  wire [63:0]   res_lo_lo_lo_6 = {res_lo_lo_lo_hi_6, res_lo_lo_lo_lo_6};
  wire [15:0]   res_lo_lo_hi_lo_lo_6 = {dataGroup_9_6, dataGroup_8_6};
  wire [15:0]   res_lo_lo_hi_lo_hi_6 = {dataGroup_11_6, dataGroup_10_6};
  wire [31:0]   res_lo_lo_hi_lo_6 = {res_lo_lo_hi_lo_hi_6, res_lo_lo_hi_lo_lo_6};
  wire [15:0]   res_lo_lo_hi_hi_lo_6 = {dataGroup_13_6, dataGroup_12_6};
  wire [15:0]   res_lo_lo_hi_hi_hi_6 = {dataGroup_15_6, dataGroup_14_6};
  wire [31:0]   res_lo_lo_hi_hi_6 = {res_lo_lo_hi_hi_hi_6, res_lo_lo_hi_hi_lo_6};
  wire [63:0]   res_lo_lo_hi_6 = {res_lo_lo_hi_hi_6, res_lo_lo_hi_lo_6};
  wire [127:0]  res_lo_lo_6 = {res_lo_lo_hi_6, res_lo_lo_lo_6};
  wire [15:0]   res_lo_hi_lo_lo_lo_6 = {dataGroup_17_6, dataGroup_16_6};
  wire [15:0]   res_lo_hi_lo_lo_hi_6 = {dataGroup_19_6, dataGroup_18_6};
  wire [31:0]   res_lo_hi_lo_lo_6 = {res_lo_hi_lo_lo_hi_6, res_lo_hi_lo_lo_lo_6};
  wire [15:0]   res_lo_hi_lo_hi_lo_6 = {dataGroup_21_6, dataGroup_20_6};
  wire [15:0]   res_lo_hi_lo_hi_hi_6 = {dataGroup_23_6, dataGroup_22_6};
  wire [31:0]   res_lo_hi_lo_hi_6 = {res_lo_hi_lo_hi_hi_6, res_lo_hi_lo_hi_lo_6};
  wire [63:0]   res_lo_hi_lo_6 = {res_lo_hi_lo_hi_6, res_lo_hi_lo_lo_6};
  wire [15:0]   res_lo_hi_hi_lo_lo_6 = {dataGroup_25_6, dataGroup_24_6};
  wire [15:0]   res_lo_hi_hi_lo_hi_6 = {dataGroup_27_6, dataGroup_26_6};
  wire [31:0]   res_lo_hi_hi_lo_6 = {res_lo_hi_hi_lo_hi_6, res_lo_hi_hi_lo_lo_6};
  wire [15:0]   res_lo_hi_hi_hi_lo_6 = {dataGroup_29_6, dataGroup_28_6};
  wire [15:0]   res_lo_hi_hi_hi_hi_6 = {dataGroup_31_6, dataGroup_30_6};
  wire [31:0]   res_lo_hi_hi_hi_6 = {res_lo_hi_hi_hi_hi_6, res_lo_hi_hi_hi_lo_6};
  wire [63:0]   res_lo_hi_hi_6 = {res_lo_hi_hi_hi_6, res_lo_hi_hi_lo_6};
  wire [127:0]  res_lo_hi_6 = {res_lo_hi_hi_6, res_lo_hi_lo_6};
  wire [255:0]  res_lo_6 = {res_lo_hi_6, res_lo_lo_6};
  wire [15:0]   res_hi_lo_lo_lo_lo_6 = {dataGroup_33_6, dataGroup_32_6};
  wire [15:0]   res_hi_lo_lo_lo_hi_6 = {dataGroup_35_6, dataGroup_34_6};
  wire [31:0]   res_hi_lo_lo_lo_6 = {res_hi_lo_lo_lo_hi_6, res_hi_lo_lo_lo_lo_6};
  wire [15:0]   res_hi_lo_lo_hi_lo_6 = {dataGroup_37_6, dataGroup_36_6};
  wire [15:0]   res_hi_lo_lo_hi_hi_6 = {dataGroup_39_6, dataGroup_38_6};
  wire [31:0]   res_hi_lo_lo_hi_6 = {res_hi_lo_lo_hi_hi_6, res_hi_lo_lo_hi_lo_6};
  wire [63:0]   res_hi_lo_lo_6 = {res_hi_lo_lo_hi_6, res_hi_lo_lo_lo_6};
  wire [15:0]   res_hi_lo_hi_lo_lo_6 = {dataGroup_41_6, dataGroup_40_6};
  wire [15:0]   res_hi_lo_hi_lo_hi_6 = {dataGroup_43_6, dataGroup_42_6};
  wire [31:0]   res_hi_lo_hi_lo_6 = {res_hi_lo_hi_lo_hi_6, res_hi_lo_hi_lo_lo_6};
  wire [15:0]   res_hi_lo_hi_hi_lo_6 = {dataGroup_45_6, dataGroup_44_6};
  wire [15:0]   res_hi_lo_hi_hi_hi_6 = {dataGroup_47_6, dataGroup_46_6};
  wire [31:0]   res_hi_lo_hi_hi_6 = {res_hi_lo_hi_hi_hi_6, res_hi_lo_hi_hi_lo_6};
  wire [63:0]   res_hi_lo_hi_6 = {res_hi_lo_hi_hi_6, res_hi_lo_hi_lo_6};
  wire [127:0]  res_hi_lo_6 = {res_hi_lo_hi_6, res_hi_lo_lo_6};
  wire [15:0]   res_hi_hi_lo_lo_lo_6 = {dataGroup_49_6, dataGroup_48_6};
  wire [15:0]   res_hi_hi_lo_lo_hi_6 = {dataGroup_51_6, dataGroup_50_6};
  wire [31:0]   res_hi_hi_lo_lo_6 = {res_hi_hi_lo_lo_hi_6, res_hi_hi_lo_lo_lo_6};
  wire [15:0]   res_hi_hi_lo_hi_lo_6 = {dataGroup_53_6, dataGroup_52_6};
  wire [15:0]   res_hi_hi_lo_hi_hi_6 = {dataGroup_55_6, dataGroup_54_6};
  wire [31:0]   res_hi_hi_lo_hi_6 = {res_hi_hi_lo_hi_hi_6, res_hi_hi_lo_hi_lo_6};
  wire [63:0]   res_hi_hi_lo_6 = {res_hi_hi_lo_hi_6, res_hi_hi_lo_lo_6};
  wire [15:0]   res_hi_hi_hi_lo_lo_6 = {dataGroup_57_6, dataGroup_56_6};
  wire [15:0]   res_hi_hi_hi_lo_hi_6 = {dataGroup_59_6, dataGroup_58_6};
  wire [31:0]   res_hi_hi_hi_lo_6 = {res_hi_hi_hi_lo_hi_6, res_hi_hi_hi_lo_lo_6};
  wire [15:0]   res_hi_hi_hi_hi_lo_6 = {dataGroup_61_6, dataGroup_60_6};
  wire [15:0]   res_hi_hi_hi_hi_hi_6 = {dataGroup_63_6, dataGroup_62_6};
  wire [31:0]   res_hi_hi_hi_hi_6 = {res_hi_hi_hi_hi_hi_6, res_hi_hi_hi_hi_lo_6};
  wire [63:0]   res_hi_hi_hi_6 = {res_hi_hi_hi_hi_6, res_hi_hi_hi_lo_6};
  wire [127:0]  res_hi_hi_6 = {res_hi_hi_hi_6, res_hi_hi_lo_6};
  wire [255:0]  res_hi_6 = {res_hi_hi_6, res_hi_lo_6};
  wire [511:0]  res_24 = {res_hi_6, res_lo_6};
  wire [2047:0] dataGroup_lo_448 = {dataGroup_lo_hi_448, dataGroup_lo_lo_448};
  wire [2047:0] dataGroup_hi_448 = {dataGroup_hi_hi_448, dataGroup_hi_lo_448};
  wire [7:0]    dataGroup_0_7 = dataGroup_lo_448[15:8];
  wire [2047:0] dataGroup_lo_449 = {dataGroup_lo_hi_449, dataGroup_lo_lo_449};
  wire [2047:0] dataGroup_hi_449 = {dataGroup_hi_hi_449, dataGroup_hi_lo_449};
  wire [7:0]    dataGroup_1_7 = dataGroup_lo_449[47:40];
  wire [2047:0] dataGroup_lo_450 = {dataGroup_lo_hi_450, dataGroup_lo_lo_450};
  wire [2047:0] dataGroup_hi_450 = {dataGroup_hi_hi_450, dataGroup_hi_lo_450};
  wire [7:0]    dataGroup_2_7 = dataGroup_lo_450[79:72];
  wire [2047:0] dataGroup_lo_451 = {dataGroup_lo_hi_451, dataGroup_lo_lo_451};
  wire [2047:0] dataGroup_hi_451 = {dataGroup_hi_hi_451, dataGroup_hi_lo_451};
  wire [7:0]    dataGroup_3_7 = dataGroup_lo_451[111:104];
  wire [2047:0] dataGroup_lo_452 = {dataGroup_lo_hi_452, dataGroup_lo_lo_452};
  wire [2047:0] dataGroup_hi_452 = {dataGroup_hi_hi_452, dataGroup_hi_lo_452};
  wire [7:0]    dataGroup_4_7 = dataGroup_lo_452[143:136];
  wire [2047:0] dataGroup_lo_453 = {dataGroup_lo_hi_453, dataGroup_lo_lo_453};
  wire [2047:0] dataGroup_hi_453 = {dataGroup_hi_hi_453, dataGroup_hi_lo_453};
  wire [7:0]    dataGroup_5_7 = dataGroup_lo_453[175:168];
  wire [2047:0] dataGroup_lo_454 = {dataGroup_lo_hi_454, dataGroup_lo_lo_454};
  wire [2047:0] dataGroup_hi_454 = {dataGroup_hi_hi_454, dataGroup_hi_lo_454};
  wire [7:0]    dataGroup_6_7 = dataGroup_lo_454[207:200];
  wire [2047:0] dataGroup_lo_455 = {dataGroup_lo_hi_455, dataGroup_lo_lo_455};
  wire [2047:0] dataGroup_hi_455 = {dataGroup_hi_hi_455, dataGroup_hi_lo_455};
  wire [7:0]    dataGroup_7_7 = dataGroup_lo_455[239:232];
  wire [2047:0] dataGroup_lo_456 = {dataGroup_lo_hi_456, dataGroup_lo_lo_456};
  wire [2047:0] dataGroup_hi_456 = {dataGroup_hi_hi_456, dataGroup_hi_lo_456};
  wire [7:0]    dataGroup_8_7 = dataGroup_lo_456[271:264];
  wire [2047:0] dataGroup_lo_457 = {dataGroup_lo_hi_457, dataGroup_lo_lo_457};
  wire [2047:0] dataGroup_hi_457 = {dataGroup_hi_hi_457, dataGroup_hi_lo_457};
  wire [7:0]    dataGroup_9_7 = dataGroup_lo_457[303:296];
  wire [2047:0] dataGroup_lo_458 = {dataGroup_lo_hi_458, dataGroup_lo_lo_458};
  wire [2047:0] dataGroup_hi_458 = {dataGroup_hi_hi_458, dataGroup_hi_lo_458};
  wire [7:0]    dataGroup_10_7 = dataGroup_lo_458[335:328];
  wire [2047:0] dataGroup_lo_459 = {dataGroup_lo_hi_459, dataGroup_lo_lo_459};
  wire [2047:0] dataGroup_hi_459 = {dataGroup_hi_hi_459, dataGroup_hi_lo_459};
  wire [7:0]    dataGroup_11_7 = dataGroup_lo_459[367:360];
  wire [2047:0] dataGroup_lo_460 = {dataGroup_lo_hi_460, dataGroup_lo_lo_460};
  wire [2047:0] dataGroup_hi_460 = {dataGroup_hi_hi_460, dataGroup_hi_lo_460};
  wire [7:0]    dataGroup_12_7 = dataGroup_lo_460[399:392];
  wire [2047:0] dataGroup_lo_461 = {dataGroup_lo_hi_461, dataGroup_lo_lo_461};
  wire [2047:0] dataGroup_hi_461 = {dataGroup_hi_hi_461, dataGroup_hi_lo_461};
  wire [7:0]    dataGroup_13_7 = dataGroup_lo_461[431:424];
  wire [2047:0] dataGroup_lo_462 = {dataGroup_lo_hi_462, dataGroup_lo_lo_462};
  wire [2047:0] dataGroup_hi_462 = {dataGroup_hi_hi_462, dataGroup_hi_lo_462};
  wire [7:0]    dataGroup_14_7 = dataGroup_lo_462[463:456];
  wire [2047:0] dataGroup_lo_463 = {dataGroup_lo_hi_463, dataGroup_lo_lo_463};
  wire [2047:0] dataGroup_hi_463 = {dataGroup_hi_hi_463, dataGroup_hi_lo_463};
  wire [7:0]    dataGroup_15_7 = dataGroup_lo_463[495:488];
  wire [2047:0] dataGroup_lo_464 = {dataGroup_lo_hi_464, dataGroup_lo_lo_464};
  wire [2047:0] dataGroup_hi_464 = {dataGroup_hi_hi_464, dataGroup_hi_lo_464};
  wire [7:0]    dataGroup_16_7 = dataGroup_lo_464[527:520];
  wire [2047:0] dataGroup_lo_465 = {dataGroup_lo_hi_465, dataGroup_lo_lo_465};
  wire [2047:0] dataGroup_hi_465 = {dataGroup_hi_hi_465, dataGroup_hi_lo_465};
  wire [7:0]    dataGroup_17_7 = dataGroup_lo_465[559:552];
  wire [2047:0] dataGroup_lo_466 = {dataGroup_lo_hi_466, dataGroup_lo_lo_466};
  wire [2047:0] dataGroup_hi_466 = {dataGroup_hi_hi_466, dataGroup_hi_lo_466};
  wire [7:0]    dataGroup_18_7 = dataGroup_lo_466[591:584];
  wire [2047:0] dataGroup_lo_467 = {dataGroup_lo_hi_467, dataGroup_lo_lo_467};
  wire [2047:0] dataGroup_hi_467 = {dataGroup_hi_hi_467, dataGroup_hi_lo_467};
  wire [7:0]    dataGroup_19_7 = dataGroup_lo_467[623:616];
  wire [2047:0] dataGroup_lo_468 = {dataGroup_lo_hi_468, dataGroup_lo_lo_468};
  wire [2047:0] dataGroup_hi_468 = {dataGroup_hi_hi_468, dataGroup_hi_lo_468};
  wire [7:0]    dataGroup_20_7 = dataGroup_lo_468[655:648];
  wire [2047:0] dataGroup_lo_469 = {dataGroup_lo_hi_469, dataGroup_lo_lo_469};
  wire [2047:0] dataGroup_hi_469 = {dataGroup_hi_hi_469, dataGroup_hi_lo_469};
  wire [7:0]    dataGroup_21_7 = dataGroup_lo_469[687:680];
  wire [2047:0] dataGroup_lo_470 = {dataGroup_lo_hi_470, dataGroup_lo_lo_470};
  wire [2047:0] dataGroup_hi_470 = {dataGroup_hi_hi_470, dataGroup_hi_lo_470};
  wire [7:0]    dataGroup_22_7 = dataGroup_lo_470[719:712];
  wire [2047:0] dataGroup_lo_471 = {dataGroup_lo_hi_471, dataGroup_lo_lo_471};
  wire [2047:0] dataGroup_hi_471 = {dataGroup_hi_hi_471, dataGroup_hi_lo_471};
  wire [7:0]    dataGroup_23_7 = dataGroup_lo_471[751:744];
  wire [2047:0] dataGroup_lo_472 = {dataGroup_lo_hi_472, dataGroup_lo_lo_472};
  wire [2047:0] dataGroup_hi_472 = {dataGroup_hi_hi_472, dataGroup_hi_lo_472};
  wire [7:0]    dataGroup_24_7 = dataGroup_lo_472[783:776];
  wire [2047:0] dataGroup_lo_473 = {dataGroup_lo_hi_473, dataGroup_lo_lo_473};
  wire [2047:0] dataGroup_hi_473 = {dataGroup_hi_hi_473, dataGroup_hi_lo_473};
  wire [7:0]    dataGroup_25_7 = dataGroup_lo_473[815:808];
  wire [2047:0] dataGroup_lo_474 = {dataGroup_lo_hi_474, dataGroup_lo_lo_474};
  wire [2047:0] dataGroup_hi_474 = {dataGroup_hi_hi_474, dataGroup_hi_lo_474};
  wire [7:0]    dataGroup_26_7 = dataGroup_lo_474[847:840];
  wire [2047:0] dataGroup_lo_475 = {dataGroup_lo_hi_475, dataGroup_lo_lo_475};
  wire [2047:0] dataGroup_hi_475 = {dataGroup_hi_hi_475, dataGroup_hi_lo_475};
  wire [7:0]    dataGroup_27_7 = dataGroup_lo_475[879:872];
  wire [2047:0] dataGroup_lo_476 = {dataGroup_lo_hi_476, dataGroup_lo_lo_476};
  wire [2047:0] dataGroup_hi_476 = {dataGroup_hi_hi_476, dataGroup_hi_lo_476};
  wire [7:0]    dataGroup_28_7 = dataGroup_lo_476[911:904];
  wire [2047:0] dataGroup_lo_477 = {dataGroup_lo_hi_477, dataGroup_lo_lo_477};
  wire [2047:0] dataGroup_hi_477 = {dataGroup_hi_hi_477, dataGroup_hi_lo_477};
  wire [7:0]    dataGroup_29_7 = dataGroup_lo_477[943:936];
  wire [2047:0] dataGroup_lo_478 = {dataGroup_lo_hi_478, dataGroup_lo_lo_478};
  wire [2047:0] dataGroup_hi_478 = {dataGroup_hi_hi_478, dataGroup_hi_lo_478};
  wire [7:0]    dataGroup_30_7 = dataGroup_lo_478[975:968];
  wire [2047:0] dataGroup_lo_479 = {dataGroup_lo_hi_479, dataGroup_lo_lo_479};
  wire [2047:0] dataGroup_hi_479 = {dataGroup_hi_hi_479, dataGroup_hi_lo_479};
  wire [7:0]    dataGroup_31_7 = dataGroup_lo_479[1007:1000];
  wire [2047:0] dataGroup_lo_480 = {dataGroup_lo_hi_480, dataGroup_lo_lo_480};
  wire [2047:0] dataGroup_hi_480 = {dataGroup_hi_hi_480, dataGroup_hi_lo_480};
  wire [7:0]    dataGroup_32_7 = dataGroup_lo_480[1039:1032];
  wire [2047:0] dataGroup_lo_481 = {dataGroup_lo_hi_481, dataGroup_lo_lo_481};
  wire [2047:0] dataGroup_hi_481 = {dataGroup_hi_hi_481, dataGroup_hi_lo_481};
  wire [7:0]    dataGroup_33_7 = dataGroup_lo_481[1071:1064];
  wire [2047:0] dataGroup_lo_482 = {dataGroup_lo_hi_482, dataGroup_lo_lo_482};
  wire [2047:0] dataGroup_hi_482 = {dataGroup_hi_hi_482, dataGroup_hi_lo_482};
  wire [7:0]    dataGroup_34_7 = dataGroup_lo_482[1103:1096];
  wire [2047:0] dataGroup_lo_483 = {dataGroup_lo_hi_483, dataGroup_lo_lo_483};
  wire [2047:0] dataGroup_hi_483 = {dataGroup_hi_hi_483, dataGroup_hi_lo_483};
  wire [7:0]    dataGroup_35_7 = dataGroup_lo_483[1135:1128];
  wire [2047:0] dataGroup_lo_484 = {dataGroup_lo_hi_484, dataGroup_lo_lo_484};
  wire [2047:0] dataGroup_hi_484 = {dataGroup_hi_hi_484, dataGroup_hi_lo_484};
  wire [7:0]    dataGroup_36_7 = dataGroup_lo_484[1167:1160];
  wire [2047:0] dataGroup_lo_485 = {dataGroup_lo_hi_485, dataGroup_lo_lo_485};
  wire [2047:0] dataGroup_hi_485 = {dataGroup_hi_hi_485, dataGroup_hi_lo_485};
  wire [7:0]    dataGroup_37_7 = dataGroup_lo_485[1199:1192];
  wire [2047:0] dataGroup_lo_486 = {dataGroup_lo_hi_486, dataGroup_lo_lo_486};
  wire [2047:0] dataGroup_hi_486 = {dataGroup_hi_hi_486, dataGroup_hi_lo_486};
  wire [7:0]    dataGroup_38_7 = dataGroup_lo_486[1231:1224];
  wire [2047:0] dataGroup_lo_487 = {dataGroup_lo_hi_487, dataGroup_lo_lo_487};
  wire [2047:0] dataGroup_hi_487 = {dataGroup_hi_hi_487, dataGroup_hi_lo_487};
  wire [7:0]    dataGroup_39_7 = dataGroup_lo_487[1263:1256];
  wire [2047:0] dataGroup_lo_488 = {dataGroup_lo_hi_488, dataGroup_lo_lo_488};
  wire [2047:0] dataGroup_hi_488 = {dataGroup_hi_hi_488, dataGroup_hi_lo_488};
  wire [7:0]    dataGroup_40_7 = dataGroup_lo_488[1295:1288];
  wire [2047:0] dataGroup_lo_489 = {dataGroup_lo_hi_489, dataGroup_lo_lo_489};
  wire [2047:0] dataGroup_hi_489 = {dataGroup_hi_hi_489, dataGroup_hi_lo_489};
  wire [7:0]    dataGroup_41_7 = dataGroup_lo_489[1327:1320];
  wire [2047:0] dataGroup_lo_490 = {dataGroup_lo_hi_490, dataGroup_lo_lo_490};
  wire [2047:0] dataGroup_hi_490 = {dataGroup_hi_hi_490, dataGroup_hi_lo_490};
  wire [7:0]    dataGroup_42_7 = dataGroup_lo_490[1359:1352];
  wire [2047:0] dataGroup_lo_491 = {dataGroup_lo_hi_491, dataGroup_lo_lo_491};
  wire [2047:0] dataGroup_hi_491 = {dataGroup_hi_hi_491, dataGroup_hi_lo_491};
  wire [7:0]    dataGroup_43_7 = dataGroup_lo_491[1391:1384];
  wire [2047:0] dataGroup_lo_492 = {dataGroup_lo_hi_492, dataGroup_lo_lo_492};
  wire [2047:0] dataGroup_hi_492 = {dataGroup_hi_hi_492, dataGroup_hi_lo_492};
  wire [7:0]    dataGroup_44_7 = dataGroup_lo_492[1423:1416];
  wire [2047:0] dataGroup_lo_493 = {dataGroup_lo_hi_493, dataGroup_lo_lo_493};
  wire [2047:0] dataGroup_hi_493 = {dataGroup_hi_hi_493, dataGroup_hi_lo_493};
  wire [7:0]    dataGroup_45_7 = dataGroup_lo_493[1455:1448];
  wire [2047:0] dataGroup_lo_494 = {dataGroup_lo_hi_494, dataGroup_lo_lo_494};
  wire [2047:0] dataGroup_hi_494 = {dataGroup_hi_hi_494, dataGroup_hi_lo_494};
  wire [7:0]    dataGroup_46_7 = dataGroup_lo_494[1487:1480];
  wire [2047:0] dataGroup_lo_495 = {dataGroup_lo_hi_495, dataGroup_lo_lo_495};
  wire [2047:0] dataGroup_hi_495 = {dataGroup_hi_hi_495, dataGroup_hi_lo_495};
  wire [7:0]    dataGroup_47_7 = dataGroup_lo_495[1519:1512];
  wire [2047:0] dataGroup_lo_496 = {dataGroup_lo_hi_496, dataGroup_lo_lo_496};
  wire [2047:0] dataGroup_hi_496 = {dataGroup_hi_hi_496, dataGroup_hi_lo_496};
  wire [7:0]    dataGroup_48_7 = dataGroup_lo_496[1551:1544];
  wire [2047:0] dataGroup_lo_497 = {dataGroup_lo_hi_497, dataGroup_lo_lo_497};
  wire [2047:0] dataGroup_hi_497 = {dataGroup_hi_hi_497, dataGroup_hi_lo_497};
  wire [7:0]    dataGroup_49_7 = dataGroup_lo_497[1583:1576];
  wire [2047:0] dataGroup_lo_498 = {dataGroup_lo_hi_498, dataGroup_lo_lo_498};
  wire [2047:0] dataGroup_hi_498 = {dataGroup_hi_hi_498, dataGroup_hi_lo_498};
  wire [7:0]    dataGroup_50_7 = dataGroup_lo_498[1615:1608];
  wire [2047:0] dataGroup_lo_499 = {dataGroup_lo_hi_499, dataGroup_lo_lo_499};
  wire [2047:0] dataGroup_hi_499 = {dataGroup_hi_hi_499, dataGroup_hi_lo_499};
  wire [7:0]    dataGroup_51_7 = dataGroup_lo_499[1647:1640];
  wire [2047:0] dataGroup_lo_500 = {dataGroup_lo_hi_500, dataGroup_lo_lo_500};
  wire [2047:0] dataGroup_hi_500 = {dataGroup_hi_hi_500, dataGroup_hi_lo_500};
  wire [7:0]    dataGroup_52_7 = dataGroup_lo_500[1679:1672];
  wire [2047:0] dataGroup_lo_501 = {dataGroup_lo_hi_501, dataGroup_lo_lo_501};
  wire [2047:0] dataGroup_hi_501 = {dataGroup_hi_hi_501, dataGroup_hi_lo_501};
  wire [7:0]    dataGroup_53_7 = dataGroup_lo_501[1711:1704];
  wire [2047:0] dataGroup_lo_502 = {dataGroup_lo_hi_502, dataGroup_lo_lo_502};
  wire [2047:0] dataGroup_hi_502 = {dataGroup_hi_hi_502, dataGroup_hi_lo_502};
  wire [7:0]    dataGroup_54_7 = dataGroup_lo_502[1743:1736];
  wire [2047:0] dataGroup_lo_503 = {dataGroup_lo_hi_503, dataGroup_lo_lo_503};
  wire [2047:0] dataGroup_hi_503 = {dataGroup_hi_hi_503, dataGroup_hi_lo_503};
  wire [7:0]    dataGroup_55_7 = dataGroup_lo_503[1775:1768];
  wire [2047:0] dataGroup_lo_504 = {dataGroup_lo_hi_504, dataGroup_lo_lo_504};
  wire [2047:0] dataGroup_hi_504 = {dataGroup_hi_hi_504, dataGroup_hi_lo_504};
  wire [7:0]    dataGroup_56_7 = dataGroup_lo_504[1807:1800];
  wire [2047:0] dataGroup_lo_505 = {dataGroup_lo_hi_505, dataGroup_lo_lo_505};
  wire [2047:0] dataGroup_hi_505 = {dataGroup_hi_hi_505, dataGroup_hi_lo_505};
  wire [7:0]    dataGroup_57_7 = dataGroup_lo_505[1839:1832];
  wire [2047:0] dataGroup_lo_506 = {dataGroup_lo_hi_506, dataGroup_lo_lo_506};
  wire [2047:0] dataGroup_hi_506 = {dataGroup_hi_hi_506, dataGroup_hi_lo_506};
  wire [7:0]    dataGroup_58_7 = dataGroup_lo_506[1871:1864];
  wire [2047:0] dataGroup_lo_507 = {dataGroup_lo_hi_507, dataGroup_lo_lo_507};
  wire [2047:0] dataGroup_hi_507 = {dataGroup_hi_hi_507, dataGroup_hi_lo_507};
  wire [7:0]    dataGroup_59_7 = dataGroup_lo_507[1903:1896];
  wire [2047:0] dataGroup_lo_508 = {dataGroup_lo_hi_508, dataGroup_lo_lo_508};
  wire [2047:0] dataGroup_hi_508 = {dataGroup_hi_hi_508, dataGroup_hi_lo_508};
  wire [7:0]    dataGroup_60_7 = dataGroup_lo_508[1935:1928];
  wire [2047:0] dataGroup_lo_509 = {dataGroup_lo_hi_509, dataGroup_lo_lo_509};
  wire [2047:0] dataGroup_hi_509 = {dataGroup_hi_hi_509, dataGroup_hi_lo_509};
  wire [7:0]    dataGroup_61_7 = dataGroup_lo_509[1967:1960];
  wire [2047:0] dataGroup_lo_510 = {dataGroup_lo_hi_510, dataGroup_lo_lo_510};
  wire [2047:0] dataGroup_hi_510 = {dataGroup_hi_hi_510, dataGroup_hi_lo_510};
  wire [7:0]    dataGroup_62_7 = dataGroup_lo_510[1999:1992];
  wire [2047:0] dataGroup_lo_511 = {dataGroup_lo_hi_511, dataGroup_lo_lo_511};
  wire [2047:0] dataGroup_hi_511 = {dataGroup_hi_hi_511, dataGroup_hi_lo_511};
  wire [7:0]    dataGroup_63_7 = dataGroup_lo_511[2031:2024];
  wire [15:0]   res_lo_lo_lo_lo_lo_7 = {dataGroup_1_7, dataGroup_0_7};
  wire [15:0]   res_lo_lo_lo_lo_hi_7 = {dataGroup_3_7, dataGroup_2_7};
  wire [31:0]   res_lo_lo_lo_lo_7 = {res_lo_lo_lo_lo_hi_7, res_lo_lo_lo_lo_lo_7};
  wire [15:0]   res_lo_lo_lo_hi_lo_7 = {dataGroup_5_7, dataGroup_4_7};
  wire [15:0]   res_lo_lo_lo_hi_hi_7 = {dataGroup_7_7, dataGroup_6_7};
  wire [31:0]   res_lo_lo_lo_hi_7 = {res_lo_lo_lo_hi_hi_7, res_lo_lo_lo_hi_lo_7};
  wire [63:0]   res_lo_lo_lo_7 = {res_lo_lo_lo_hi_7, res_lo_lo_lo_lo_7};
  wire [15:0]   res_lo_lo_hi_lo_lo_7 = {dataGroup_9_7, dataGroup_8_7};
  wire [15:0]   res_lo_lo_hi_lo_hi_7 = {dataGroup_11_7, dataGroup_10_7};
  wire [31:0]   res_lo_lo_hi_lo_7 = {res_lo_lo_hi_lo_hi_7, res_lo_lo_hi_lo_lo_7};
  wire [15:0]   res_lo_lo_hi_hi_lo_7 = {dataGroup_13_7, dataGroup_12_7};
  wire [15:0]   res_lo_lo_hi_hi_hi_7 = {dataGroup_15_7, dataGroup_14_7};
  wire [31:0]   res_lo_lo_hi_hi_7 = {res_lo_lo_hi_hi_hi_7, res_lo_lo_hi_hi_lo_7};
  wire [63:0]   res_lo_lo_hi_7 = {res_lo_lo_hi_hi_7, res_lo_lo_hi_lo_7};
  wire [127:0]  res_lo_lo_7 = {res_lo_lo_hi_7, res_lo_lo_lo_7};
  wire [15:0]   res_lo_hi_lo_lo_lo_7 = {dataGroup_17_7, dataGroup_16_7};
  wire [15:0]   res_lo_hi_lo_lo_hi_7 = {dataGroup_19_7, dataGroup_18_7};
  wire [31:0]   res_lo_hi_lo_lo_7 = {res_lo_hi_lo_lo_hi_7, res_lo_hi_lo_lo_lo_7};
  wire [15:0]   res_lo_hi_lo_hi_lo_7 = {dataGroup_21_7, dataGroup_20_7};
  wire [15:0]   res_lo_hi_lo_hi_hi_7 = {dataGroup_23_7, dataGroup_22_7};
  wire [31:0]   res_lo_hi_lo_hi_7 = {res_lo_hi_lo_hi_hi_7, res_lo_hi_lo_hi_lo_7};
  wire [63:0]   res_lo_hi_lo_7 = {res_lo_hi_lo_hi_7, res_lo_hi_lo_lo_7};
  wire [15:0]   res_lo_hi_hi_lo_lo_7 = {dataGroup_25_7, dataGroup_24_7};
  wire [15:0]   res_lo_hi_hi_lo_hi_7 = {dataGroup_27_7, dataGroup_26_7};
  wire [31:0]   res_lo_hi_hi_lo_7 = {res_lo_hi_hi_lo_hi_7, res_lo_hi_hi_lo_lo_7};
  wire [15:0]   res_lo_hi_hi_hi_lo_7 = {dataGroup_29_7, dataGroup_28_7};
  wire [15:0]   res_lo_hi_hi_hi_hi_7 = {dataGroup_31_7, dataGroup_30_7};
  wire [31:0]   res_lo_hi_hi_hi_7 = {res_lo_hi_hi_hi_hi_7, res_lo_hi_hi_hi_lo_7};
  wire [63:0]   res_lo_hi_hi_7 = {res_lo_hi_hi_hi_7, res_lo_hi_hi_lo_7};
  wire [127:0]  res_lo_hi_7 = {res_lo_hi_hi_7, res_lo_hi_lo_7};
  wire [255:0]  res_lo_7 = {res_lo_hi_7, res_lo_lo_7};
  wire [15:0]   res_hi_lo_lo_lo_lo_7 = {dataGroup_33_7, dataGroup_32_7};
  wire [15:0]   res_hi_lo_lo_lo_hi_7 = {dataGroup_35_7, dataGroup_34_7};
  wire [31:0]   res_hi_lo_lo_lo_7 = {res_hi_lo_lo_lo_hi_7, res_hi_lo_lo_lo_lo_7};
  wire [15:0]   res_hi_lo_lo_hi_lo_7 = {dataGroup_37_7, dataGroup_36_7};
  wire [15:0]   res_hi_lo_lo_hi_hi_7 = {dataGroup_39_7, dataGroup_38_7};
  wire [31:0]   res_hi_lo_lo_hi_7 = {res_hi_lo_lo_hi_hi_7, res_hi_lo_lo_hi_lo_7};
  wire [63:0]   res_hi_lo_lo_7 = {res_hi_lo_lo_hi_7, res_hi_lo_lo_lo_7};
  wire [15:0]   res_hi_lo_hi_lo_lo_7 = {dataGroup_41_7, dataGroup_40_7};
  wire [15:0]   res_hi_lo_hi_lo_hi_7 = {dataGroup_43_7, dataGroup_42_7};
  wire [31:0]   res_hi_lo_hi_lo_7 = {res_hi_lo_hi_lo_hi_7, res_hi_lo_hi_lo_lo_7};
  wire [15:0]   res_hi_lo_hi_hi_lo_7 = {dataGroup_45_7, dataGroup_44_7};
  wire [15:0]   res_hi_lo_hi_hi_hi_7 = {dataGroup_47_7, dataGroup_46_7};
  wire [31:0]   res_hi_lo_hi_hi_7 = {res_hi_lo_hi_hi_hi_7, res_hi_lo_hi_hi_lo_7};
  wire [63:0]   res_hi_lo_hi_7 = {res_hi_lo_hi_hi_7, res_hi_lo_hi_lo_7};
  wire [127:0]  res_hi_lo_7 = {res_hi_lo_hi_7, res_hi_lo_lo_7};
  wire [15:0]   res_hi_hi_lo_lo_lo_7 = {dataGroup_49_7, dataGroup_48_7};
  wire [15:0]   res_hi_hi_lo_lo_hi_7 = {dataGroup_51_7, dataGroup_50_7};
  wire [31:0]   res_hi_hi_lo_lo_7 = {res_hi_hi_lo_lo_hi_7, res_hi_hi_lo_lo_lo_7};
  wire [15:0]   res_hi_hi_lo_hi_lo_7 = {dataGroup_53_7, dataGroup_52_7};
  wire [15:0]   res_hi_hi_lo_hi_hi_7 = {dataGroup_55_7, dataGroup_54_7};
  wire [31:0]   res_hi_hi_lo_hi_7 = {res_hi_hi_lo_hi_hi_7, res_hi_hi_lo_hi_lo_7};
  wire [63:0]   res_hi_hi_lo_7 = {res_hi_hi_lo_hi_7, res_hi_hi_lo_lo_7};
  wire [15:0]   res_hi_hi_hi_lo_lo_7 = {dataGroup_57_7, dataGroup_56_7};
  wire [15:0]   res_hi_hi_hi_lo_hi_7 = {dataGroup_59_7, dataGroup_58_7};
  wire [31:0]   res_hi_hi_hi_lo_7 = {res_hi_hi_hi_lo_hi_7, res_hi_hi_hi_lo_lo_7};
  wire [15:0]   res_hi_hi_hi_hi_lo_7 = {dataGroup_61_7, dataGroup_60_7};
  wire [15:0]   res_hi_hi_hi_hi_hi_7 = {dataGroup_63_7, dataGroup_62_7};
  wire [31:0]   res_hi_hi_hi_hi_7 = {res_hi_hi_hi_hi_hi_7, res_hi_hi_hi_hi_lo_7};
  wire [63:0]   res_hi_hi_hi_7 = {res_hi_hi_hi_hi_7, res_hi_hi_hi_lo_7};
  wire [127:0]  res_hi_hi_7 = {res_hi_hi_hi_7, res_hi_hi_lo_7};
  wire [255:0]  res_hi_7 = {res_hi_hi_7, res_hi_lo_7};
  wire [511:0]  res_25 = {res_hi_7, res_lo_7};
  wire [2047:0] dataGroup_lo_512 = {dataGroup_lo_hi_512, dataGroup_lo_lo_512};
  wire [2047:0] dataGroup_hi_512 = {dataGroup_hi_hi_512, dataGroup_hi_lo_512};
  wire [7:0]    dataGroup_0_8 = dataGroup_lo_512[23:16];
  wire [2047:0] dataGroup_lo_513 = {dataGroup_lo_hi_513, dataGroup_lo_lo_513};
  wire [2047:0] dataGroup_hi_513 = {dataGroup_hi_hi_513, dataGroup_hi_lo_513};
  wire [7:0]    dataGroup_1_8 = dataGroup_lo_513[55:48];
  wire [2047:0] dataGroup_lo_514 = {dataGroup_lo_hi_514, dataGroup_lo_lo_514};
  wire [2047:0] dataGroup_hi_514 = {dataGroup_hi_hi_514, dataGroup_hi_lo_514};
  wire [7:0]    dataGroup_2_8 = dataGroup_lo_514[87:80];
  wire [2047:0] dataGroup_lo_515 = {dataGroup_lo_hi_515, dataGroup_lo_lo_515};
  wire [2047:0] dataGroup_hi_515 = {dataGroup_hi_hi_515, dataGroup_hi_lo_515};
  wire [7:0]    dataGroup_3_8 = dataGroup_lo_515[119:112];
  wire [2047:0] dataGroup_lo_516 = {dataGroup_lo_hi_516, dataGroup_lo_lo_516};
  wire [2047:0] dataGroup_hi_516 = {dataGroup_hi_hi_516, dataGroup_hi_lo_516};
  wire [7:0]    dataGroup_4_8 = dataGroup_lo_516[151:144];
  wire [2047:0] dataGroup_lo_517 = {dataGroup_lo_hi_517, dataGroup_lo_lo_517};
  wire [2047:0] dataGroup_hi_517 = {dataGroup_hi_hi_517, dataGroup_hi_lo_517};
  wire [7:0]    dataGroup_5_8 = dataGroup_lo_517[183:176];
  wire [2047:0] dataGroup_lo_518 = {dataGroup_lo_hi_518, dataGroup_lo_lo_518};
  wire [2047:0] dataGroup_hi_518 = {dataGroup_hi_hi_518, dataGroup_hi_lo_518};
  wire [7:0]    dataGroup_6_8 = dataGroup_lo_518[215:208];
  wire [2047:0] dataGroup_lo_519 = {dataGroup_lo_hi_519, dataGroup_lo_lo_519};
  wire [2047:0] dataGroup_hi_519 = {dataGroup_hi_hi_519, dataGroup_hi_lo_519};
  wire [7:0]    dataGroup_7_8 = dataGroup_lo_519[247:240];
  wire [2047:0] dataGroup_lo_520 = {dataGroup_lo_hi_520, dataGroup_lo_lo_520};
  wire [2047:0] dataGroup_hi_520 = {dataGroup_hi_hi_520, dataGroup_hi_lo_520};
  wire [7:0]    dataGroup_8_8 = dataGroup_lo_520[279:272];
  wire [2047:0] dataGroup_lo_521 = {dataGroup_lo_hi_521, dataGroup_lo_lo_521};
  wire [2047:0] dataGroup_hi_521 = {dataGroup_hi_hi_521, dataGroup_hi_lo_521};
  wire [7:0]    dataGroup_9_8 = dataGroup_lo_521[311:304];
  wire [2047:0] dataGroup_lo_522 = {dataGroup_lo_hi_522, dataGroup_lo_lo_522};
  wire [2047:0] dataGroup_hi_522 = {dataGroup_hi_hi_522, dataGroup_hi_lo_522};
  wire [7:0]    dataGroup_10_8 = dataGroup_lo_522[343:336];
  wire [2047:0] dataGroup_lo_523 = {dataGroup_lo_hi_523, dataGroup_lo_lo_523};
  wire [2047:0] dataGroup_hi_523 = {dataGroup_hi_hi_523, dataGroup_hi_lo_523};
  wire [7:0]    dataGroup_11_8 = dataGroup_lo_523[375:368];
  wire [2047:0] dataGroup_lo_524 = {dataGroup_lo_hi_524, dataGroup_lo_lo_524};
  wire [2047:0] dataGroup_hi_524 = {dataGroup_hi_hi_524, dataGroup_hi_lo_524};
  wire [7:0]    dataGroup_12_8 = dataGroup_lo_524[407:400];
  wire [2047:0] dataGroup_lo_525 = {dataGroup_lo_hi_525, dataGroup_lo_lo_525};
  wire [2047:0] dataGroup_hi_525 = {dataGroup_hi_hi_525, dataGroup_hi_lo_525};
  wire [7:0]    dataGroup_13_8 = dataGroup_lo_525[439:432];
  wire [2047:0] dataGroup_lo_526 = {dataGroup_lo_hi_526, dataGroup_lo_lo_526};
  wire [2047:0] dataGroup_hi_526 = {dataGroup_hi_hi_526, dataGroup_hi_lo_526};
  wire [7:0]    dataGroup_14_8 = dataGroup_lo_526[471:464];
  wire [2047:0] dataGroup_lo_527 = {dataGroup_lo_hi_527, dataGroup_lo_lo_527};
  wire [2047:0] dataGroup_hi_527 = {dataGroup_hi_hi_527, dataGroup_hi_lo_527};
  wire [7:0]    dataGroup_15_8 = dataGroup_lo_527[503:496];
  wire [2047:0] dataGroup_lo_528 = {dataGroup_lo_hi_528, dataGroup_lo_lo_528};
  wire [2047:0] dataGroup_hi_528 = {dataGroup_hi_hi_528, dataGroup_hi_lo_528};
  wire [7:0]    dataGroup_16_8 = dataGroup_lo_528[535:528];
  wire [2047:0] dataGroup_lo_529 = {dataGroup_lo_hi_529, dataGroup_lo_lo_529};
  wire [2047:0] dataGroup_hi_529 = {dataGroup_hi_hi_529, dataGroup_hi_lo_529};
  wire [7:0]    dataGroup_17_8 = dataGroup_lo_529[567:560];
  wire [2047:0] dataGroup_lo_530 = {dataGroup_lo_hi_530, dataGroup_lo_lo_530};
  wire [2047:0] dataGroup_hi_530 = {dataGroup_hi_hi_530, dataGroup_hi_lo_530};
  wire [7:0]    dataGroup_18_8 = dataGroup_lo_530[599:592];
  wire [2047:0] dataGroup_lo_531 = {dataGroup_lo_hi_531, dataGroup_lo_lo_531};
  wire [2047:0] dataGroup_hi_531 = {dataGroup_hi_hi_531, dataGroup_hi_lo_531};
  wire [7:0]    dataGroup_19_8 = dataGroup_lo_531[631:624];
  wire [2047:0] dataGroup_lo_532 = {dataGroup_lo_hi_532, dataGroup_lo_lo_532};
  wire [2047:0] dataGroup_hi_532 = {dataGroup_hi_hi_532, dataGroup_hi_lo_532};
  wire [7:0]    dataGroup_20_8 = dataGroup_lo_532[663:656];
  wire [2047:0] dataGroup_lo_533 = {dataGroup_lo_hi_533, dataGroup_lo_lo_533};
  wire [2047:0] dataGroup_hi_533 = {dataGroup_hi_hi_533, dataGroup_hi_lo_533};
  wire [7:0]    dataGroup_21_8 = dataGroup_lo_533[695:688];
  wire [2047:0] dataGroup_lo_534 = {dataGroup_lo_hi_534, dataGroup_lo_lo_534};
  wire [2047:0] dataGroup_hi_534 = {dataGroup_hi_hi_534, dataGroup_hi_lo_534};
  wire [7:0]    dataGroup_22_8 = dataGroup_lo_534[727:720];
  wire [2047:0] dataGroup_lo_535 = {dataGroup_lo_hi_535, dataGroup_lo_lo_535};
  wire [2047:0] dataGroup_hi_535 = {dataGroup_hi_hi_535, dataGroup_hi_lo_535};
  wire [7:0]    dataGroup_23_8 = dataGroup_lo_535[759:752];
  wire [2047:0] dataGroup_lo_536 = {dataGroup_lo_hi_536, dataGroup_lo_lo_536};
  wire [2047:0] dataGroup_hi_536 = {dataGroup_hi_hi_536, dataGroup_hi_lo_536};
  wire [7:0]    dataGroup_24_8 = dataGroup_lo_536[791:784];
  wire [2047:0] dataGroup_lo_537 = {dataGroup_lo_hi_537, dataGroup_lo_lo_537};
  wire [2047:0] dataGroup_hi_537 = {dataGroup_hi_hi_537, dataGroup_hi_lo_537};
  wire [7:0]    dataGroup_25_8 = dataGroup_lo_537[823:816];
  wire [2047:0] dataGroup_lo_538 = {dataGroup_lo_hi_538, dataGroup_lo_lo_538};
  wire [2047:0] dataGroup_hi_538 = {dataGroup_hi_hi_538, dataGroup_hi_lo_538};
  wire [7:0]    dataGroup_26_8 = dataGroup_lo_538[855:848];
  wire [2047:0] dataGroup_lo_539 = {dataGroup_lo_hi_539, dataGroup_lo_lo_539};
  wire [2047:0] dataGroup_hi_539 = {dataGroup_hi_hi_539, dataGroup_hi_lo_539};
  wire [7:0]    dataGroup_27_8 = dataGroup_lo_539[887:880];
  wire [2047:0] dataGroup_lo_540 = {dataGroup_lo_hi_540, dataGroup_lo_lo_540};
  wire [2047:0] dataGroup_hi_540 = {dataGroup_hi_hi_540, dataGroup_hi_lo_540};
  wire [7:0]    dataGroup_28_8 = dataGroup_lo_540[919:912];
  wire [2047:0] dataGroup_lo_541 = {dataGroup_lo_hi_541, dataGroup_lo_lo_541};
  wire [2047:0] dataGroup_hi_541 = {dataGroup_hi_hi_541, dataGroup_hi_lo_541};
  wire [7:0]    dataGroup_29_8 = dataGroup_lo_541[951:944];
  wire [2047:0] dataGroup_lo_542 = {dataGroup_lo_hi_542, dataGroup_lo_lo_542};
  wire [2047:0] dataGroup_hi_542 = {dataGroup_hi_hi_542, dataGroup_hi_lo_542};
  wire [7:0]    dataGroup_30_8 = dataGroup_lo_542[983:976];
  wire [2047:0] dataGroup_lo_543 = {dataGroup_lo_hi_543, dataGroup_lo_lo_543};
  wire [2047:0] dataGroup_hi_543 = {dataGroup_hi_hi_543, dataGroup_hi_lo_543};
  wire [7:0]    dataGroup_31_8 = dataGroup_lo_543[1015:1008];
  wire [2047:0] dataGroup_lo_544 = {dataGroup_lo_hi_544, dataGroup_lo_lo_544};
  wire [2047:0] dataGroup_hi_544 = {dataGroup_hi_hi_544, dataGroup_hi_lo_544};
  wire [7:0]    dataGroup_32_8 = dataGroup_lo_544[1047:1040];
  wire [2047:0] dataGroup_lo_545 = {dataGroup_lo_hi_545, dataGroup_lo_lo_545};
  wire [2047:0] dataGroup_hi_545 = {dataGroup_hi_hi_545, dataGroup_hi_lo_545};
  wire [7:0]    dataGroup_33_8 = dataGroup_lo_545[1079:1072];
  wire [2047:0] dataGroup_lo_546 = {dataGroup_lo_hi_546, dataGroup_lo_lo_546};
  wire [2047:0] dataGroup_hi_546 = {dataGroup_hi_hi_546, dataGroup_hi_lo_546};
  wire [7:0]    dataGroup_34_8 = dataGroup_lo_546[1111:1104];
  wire [2047:0] dataGroup_lo_547 = {dataGroup_lo_hi_547, dataGroup_lo_lo_547};
  wire [2047:0] dataGroup_hi_547 = {dataGroup_hi_hi_547, dataGroup_hi_lo_547};
  wire [7:0]    dataGroup_35_8 = dataGroup_lo_547[1143:1136];
  wire [2047:0] dataGroup_lo_548 = {dataGroup_lo_hi_548, dataGroup_lo_lo_548};
  wire [2047:0] dataGroup_hi_548 = {dataGroup_hi_hi_548, dataGroup_hi_lo_548};
  wire [7:0]    dataGroup_36_8 = dataGroup_lo_548[1175:1168];
  wire [2047:0] dataGroup_lo_549 = {dataGroup_lo_hi_549, dataGroup_lo_lo_549};
  wire [2047:0] dataGroup_hi_549 = {dataGroup_hi_hi_549, dataGroup_hi_lo_549};
  wire [7:0]    dataGroup_37_8 = dataGroup_lo_549[1207:1200];
  wire [2047:0] dataGroup_lo_550 = {dataGroup_lo_hi_550, dataGroup_lo_lo_550};
  wire [2047:0] dataGroup_hi_550 = {dataGroup_hi_hi_550, dataGroup_hi_lo_550};
  wire [7:0]    dataGroup_38_8 = dataGroup_lo_550[1239:1232];
  wire [2047:0] dataGroup_lo_551 = {dataGroup_lo_hi_551, dataGroup_lo_lo_551};
  wire [2047:0] dataGroup_hi_551 = {dataGroup_hi_hi_551, dataGroup_hi_lo_551};
  wire [7:0]    dataGroup_39_8 = dataGroup_lo_551[1271:1264];
  wire [2047:0] dataGroup_lo_552 = {dataGroup_lo_hi_552, dataGroup_lo_lo_552};
  wire [2047:0] dataGroup_hi_552 = {dataGroup_hi_hi_552, dataGroup_hi_lo_552};
  wire [7:0]    dataGroup_40_8 = dataGroup_lo_552[1303:1296];
  wire [2047:0] dataGroup_lo_553 = {dataGroup_lo_hi_553, dataGroup_lo_lo_553};
  wire [2047:0] dataGroup_hi_553 = {dataGroup_hi_hi_553, dataGroup_hi_lo_553};
  wire [7:0]    dataGroup_41_8 = dataGroup_lo_553[1335:1328];
  wire [2047:0] dataGroup_lo_554 = {dataGroup_lo_hi_554, dataGroup_lo_lo_554};
  wire [2047:0] dataGroup_hi_554 = {dataGroup_hi_hi_554, dataGroup_hi_lo_554};
  wire [7:0]    dataGroup_42_8 = dataGroup_lo_554[1367:1360];
  wire [2047:0] dataGroup_lo_555 = {dataGroup_lo_hi_555, dataGroup_lo_lo_555};
  wire [2047:0] dataGroup_hi_555 = {dataGroup_hi_hi_555, dataGroup_hi_lo_555};
  wire [7:0]    dataGroup_43_8 = dataGroup_lo_555[1399:1392];
  wire [2047:0] dataGroup_lo_556 = {dataGroup_lo_hi_556, dataGroup_lo_lo_556};
  wire [2047:0] dataGroup_hi_556 = {dataGroup_hi_hi_556, dataGroup_hi_lo_556};
  wire [7:0]    dataGroup_44_8 = dataGroup_lo_556[1431:1424];
  wire [2047:0] dataGroup_lo_557 = {dataGroup_lo_hi_557, dataGroup_lo_lo_557};
  wire [2047:0] dataGroup_hi_557 = {dataGroup_hi_hi_557, dataGroup_hi_lo_557};
  wire [7:0]    dataGroup_45_8 = dataGroup_lo_557[1463:1456];
  wire [2047:0] dataGroup_lo_558 = {dataGroup_lo_hi_558, dataGroup_lo_lo_558};
  wire [2047:0] dataGroup_hi_558 = {dataGroup_hi_hi_558, dataGroup_hi_lo_558};
  wire [7:0]    dataGroup_46_8 = dataGroup_lo_558[1495:1488];
  wire [2047:0] dataGroup_lo_559 = {dataGroup_lo_hi_559, dataGroup_lo_lo_559};
  wire [2047:0] dataGroup_hi_559 = {dataGroup_hi_hi_559, dataGroup_hi_lo_559};
  wire [7:0]    dataGroup_47_8 = dataGroup_lo_559[1527:1520];
  wire [2047:0] dataGroup_lo_560 = {dataGroup_lo_hi_560, dataGroup_lo_lo_560};
  wire [2047:0] dataGroup_hi_560 = {dataGroup_hi_hi_560, dataGroup_hi_lo_560};
  wire [7:0]    dataGroup_48_8 = dataGroup_lo_560[1559:1552];
  wire [2047:0] dataGroup_lo_561 = {dataGroup_lo_hi_561, dataGroup_lo_lo_561};
  wire [2047:0] dataGroup_hi_561 = {dataGroup_hi_hi_561, dataGroup_hi_lo_561};
  wire [7:0]    dataGroup_49_8 = dataGroup_lo_561[1591:1584];
  wire [2047:0] dataGroup_lo_562 = {dataGroup_lo_hi_562, dataGroup_lo_lo_562};
  wire [2047:0] dataGroup_hi_562 = {dataGroup_hi_hi_562, dataGroup_hi_lo_562};
  wire [7:0]    dataGroup_50_8 = dataGroup_lo_562[1623:1616];
  wire [2047:0] dataGroup_lo_563 = {dataGroup_lo_hi_563, dataGroup_lo_lo_563};
  wire [2047:0] dataGroup_hi_563 = {dataGroup_hi_hi_563, dataGroup_hi_lo_563};
  wire [7:0]    dataGroup_51_8 = dataGroup_lo_563[1655:1648];
  wire [2047:0] dataGroup_lo_564 = {dataGroup_lo_hi_564, dataGroup_lo_lo_564};
  wire [2047:0] dataGroup_hi_564 = {dataGroup_hi_hi_564, dataGroup_hi_lo_564};
  wire [7:0]    dataGroup_52_8 = dataGroup_lo_564[1687:1680];
  wire [2047:0] dataGroup_lo_565 = {dataGroup_lo_hi_565, dataGroup_lo_lo_565};
  wire [2047:0] dataGroup_hi_565 = {dataGroup_hi_hi_565, dataGroup_hi_lo_565};
  wire [7:0]    dataGroup_53_8 = dataGroup_lo_565[1719:1712];
  wire [2047:0] dataGroup_lo_566 = {dataGroup_lo_hi_566, dataGroup_lo_lo_566};
  wire [2047:0] dataGroup_hi_566 = {dataGroup_hi_hi_566, dataGroup_hi_lo_566};
  wire [7:0]    dataGroup_54_8 = dataGroup_lo_566[1751:1744];
  wire [2047:0] dataGroup_lo_567 = {dataGroup_lo_hi_567, dataGroup_lo_lo_567};
  wire [2047:0] dataGroup_hi_567 = {dataGroup_hi_hi_567, dataGroup_hi_lo_567};
  wire [7:0]    dataGroup_55_8 = dataGroup_lo_567[1783:1776];
  wire [2047:0] dataGroup_lo_568 = {dataGroup_lo_hi_568, dataGroup_lo_lo_568};
  wire [2047:0] dataGroup_hi_568 = {dataGroup_hi_hi_568, dataGroup_hi_lo_568};
  wire [7:0]    dataGroup_56_8 = dataGroup_lo_568[1815:1808];
  wire [2047:0] dataGroup_lo_569 = {dataGroup_lo_hi_569, dataGroup_lo_lo_569};
  wire [2047:0] dataGroup_hi_569 = {dataGroup_hi_hi_569, dataGroup_hi_lo_569};
  wire [7:0]    dataGroup_57_8 = dataGroup_lo_569[1847:1840];
  wire [2047:0] dataGroup_lo_570 = {dataGroup_lo_hi_570, dataGroup_lo_lo_570};
  wire [2047:0] dataGroup_hi_570 = {dataGroup_hi_hi_570, dataGroup_hi_lo_570};
  wire [7:0]    dataGroup_58_8 = dataGroup_lo_570[1879:1872];
  wire [2047:0] dataGroup_lo_571 = {dataGroup_lo_hi_571, dataGroup_lo_lo_571};
  wire [2047:0] dataGroup_hi_571 = {dataGroup_hi_hi_571, dataGroup_hi_lo_571};
  wire [7:0]    dataGroup_59_8 = dataGroup_lo_571[1911:1904];
  wire [2047:0] dataGroup_lo_572 = {dataGroup_lo_hi_572, dataGroup_lo_lo_572};
  wire [2047:0] dataGroup_hi_572 = {dataGroup_hi_hi_572, dataGroup_hi_lo_572};
  wire [7:0]    dataGroup_60_8 = dataGroup_lo_572[1943:1936];
  wire [2047:0] dataGroup_lo_573 = {dataGroup_lo_hi_573, dataGroup_lo_lo_573};
  wire [2047:0] dataGroup_hi_573 = {dataGroup_hi_hi_573, dataGroup_hi_lo_573};
  wire [7:0]    dataGroup_61_8 = dataGroup_lo_573[1975:1968];
  wire [2047:0] dataGroup_lo_574 = {dataGroup_lo_hi_574, dataGroup_lo_lo_574};
  wire [2047:0] dataGroup_hi_574 = {dataGroup_hi_hi_574, dataGroup_hi_lo_574};
  wire [7:0]    dataGroup_62_8 = dataGroup_lo_574[2007:2000];
  wire [2047:0] dataGroup_lo_575 = {dataGroup_lo_hi_575, dataGroup_lo_lo_575};
  wire [2047:0] dataGroup_hi_575 = {dataGroup_hi_hi_575, dataGroup_hi_lo_575};
  wire [7:0]    dataGroup_63_8 = dataGroup_lo_575[2039:2032];
  wire [15:0]   res_lo_lo_lo_lo_lo_8 = {dataGroup_1_8, dataGroup_0_8};
  wire [15:0]   res_lo_lo_lo_lo_hi_8 = {dataGroup_3_8, dataGroup_2_8};
  wire [31:0]   res_lo_lo_lo_lo_8 = {res_lo_lo_lo_lo_hi_8, res_lo_lo_lo_lo_lo_8};
  wire [15:0]   res_lo_lo_lo_hi_lo_8 = {dataGroup_5_8, dataGroup_4_8};
  wire [15:0]   res_lo_lo_lo_hi_hi_8 = {dataGroup_7_8, dataGroup_6_8};
  wire [31:0]   res_lo_lo_lo_hi_8 = {res_lo_lo_lo_hi_hi_8, res_lo_lo_lo_hi_lo_8};
  wire [63:0]   res_lo_lo_lo_8 = {res_lo_lo_lo_hi_8, res_lo_lo_lo_lo_8};
  wire [15:0]   res_lo_lo_hi_lo_lo_8 = {dataGroup_9_8, dataGroup_8_8};
  wire [15:0]   res_lo_lo_hi_lo_hi_8 = {dataGroup_11_8, dataGroup_10_8};
  wire [31:0]   res_lo_lo_hi_lo_8 = {res_lo_lo_hi_lo_hi_8, res_lo_lo_hi_lo_lo_8};
  wire [15:0]   res_lo_lo_hi_hi_lo_8 = {dataGroup_13_8, dataGroup_12_8};
  wire [15:0]   res_lo_lo_hi_hi_hi_8 = {dataGroup_15_8, dataGroup_14_8};
  wire [31:0]   res_lo_lo_hi_hi_8 = {res_lo_lo_hi_hi_hi_8, res_lo_lo_hi_hi_lo_8};
  wire [63:0]   res_lo_lo_hi_8 = {res_lo_lo_hi_hi_8, res_lo_lo_hi_lo_8};
  wire [127:0]  res_lo_lo_8 = {res_lo_lo_hi_8, res_lo_lo_lo_8};
  wire [15:0]   res_lo_hi_lo_lo_lo_8 = {dataGroup_17_8, dataGroup_16_8};
  wire [15:0]   res_lo_hi_lo_lo_hi_8 = {dataGroup_19_8, dataGroup_18_8};
  wire [31:0]   res_lo_hi_lo_lo_8 = {res_lo_hi_lo_lo_hi_8, res_lo_hi_lo_lo_lo_8};
  wire [15:0]   res_lo_hi_lo_hi_lo_8 = {dataGroup_21_8, dataGroup_20_8};
  wire [15:0]   res_lo_hi_lo_hi_hi_8 = {dataGroup_23_8, dataGroup_22_8};
  wire [31:0]   res_lo_hi_lo_hi_8 = {res_lo_hi_lo_hi_hi_8, res_lo_hi_lo_hi_lo_8};
  wire [63:0]   res_lo_hi_lo_8 = {res_lo_hi_lo_hi_8, res_lo_hi_lo_lo_8};
  wire [15:0]   res_lo_hi_hi_lo_lo_8 = {dataGroup_25_8, dataGroup_24_8};
  wire [15:0]   res_lo_hi_hi_lo_hi_8 = {dataGroup_27_8, dataGroup_26_8};
  wire [31:0]   res_lo_hi_hi_lo_8 = {res_lo_hi_hi_lo_hi_8, res_lo_hi_hi_lo_lo_8};
  wire [15:0]   res_lo_hi_hi_hi_lo_8 = {dataGroup_29_8, dataGroup_28_8};
  wire [15:0]   res_lo_hi_hi_hi_hi_8 = {dataGroup_31_8, dataGroup_30_8};
  wire [31:0]   res_lo_hi_hi_hi_8 = {res_lo_hi_hi_hi_hi_8, res_lo_hi_hi_hi_lo_8};
  wire [63:0]   res_lo_hi_hi_8 = {res_lo_hi_hi_hi_8, res_lo_hi_hi_lo_8};
  wire [127:0]  res_lo_hi_8 = {res_lo_hi_hi_8, res_lo_hi_lo_8};
  wire [255:0]  res_lo_8 = {res_lo_hi_8, res_lo_lo_8};
  wire [15:0]   res_hi_lo_lo_lo_lo_8 = {dataGroup_33_8, dataGroup_32_8};
  wire [15:0]   res_hi_lo_lo_lo_hi_8 = {dataGroup_35_8, dataGroup_34_8};
  wire [31:0]   res_hi_lo_lo_lo_8 = {res_hi_lo_lo_lo_hi_8, res_hi_lo_lo_lo_lo_8};
  wire [15:0]   res_hi_lo_lo_hi_lo_8 = {dataGroup_37_8, dataGroup_36_8};
  wire [15:0]   res_hi_lo_lo_hi_hi_8 = {dataGroup_39_8, dataGroup_38_8};
  wire [31:0]   res_hi_lo_lo_hi_8 = {res_hi_lo_lo_hi_hi_8, res_hi_lo_lo_hi_lo_8};
  wire [63:0]   res_hi_lo_lo_8 = {res_hi_lo_lo_hi_8, res_hi_lo_lo_lo_8};
  wire [15:0]   res_hi_lo_hi_lo_lo_8 = {dataGroup_41_8, dataGroup_40_8};
  wire [15:0]   res_hi_lo_hi_lo_hi_8 = {dataGroup_43_8, dataGroup_42_8};
  wire [31:0]   res_hi_lo_hi_lo_8 = {res_hi_lo_hi_lo_hi_8, res_hi_lo_hi_lo_lo_8};
  wire [15:0]   res_hi_lo_hi_hi_lo_8 = {dataGroup_45_8, dataGroup_44_8};
  wire [15:0]   res_hi_lo_hi_hi_hi_8 = {dataGroup_47_8, dataGroup_46_8};
  wire [31:0]   res_hi_lo_hi_hi_8 = {res_hi_lo_hi_hi_hi_8, res_hi_lo_hi_hi_lo_8};
  wire [63:0]   res_hi_lo_hi_8 = {res_hi_lo_hi_hi_8, res_hi_lo_hi_lo_8};
  wire [127:0]  res_hi_lo_8 = {res_hi_lo_hi_8, res_hi_lo_lo_8};
  wire [15:0]   res_hi_hi_lo_lo_lo_8 = {dataGroup_49_8, dataGroup_48_8};
  wire [15:0]   res_hi_hi_lo_lo_hi_8 = {dataGroup_51_8, dataGroup_50_8};
  wire [31:0]   res_hi_hi_lo_lo_8 = {res_hi_hi_lo_lo_hi_8, res_hi_hi_lo_lo_lo_8};
  wire [15:0]   res_hi_hi_lo_hi_lo_8 = {dataGroup_53_8, dataGroup_52_8};
  wire [15:0]   res_hi_hi_lo_hi_hi_8 = {dataGroup_55_8, dataGroup_54_8};
  wire [31:0]   res_hi_hi_lo_hi_8 = {res_hi_hi_lo_hi_hi_8, res_hi_hi_lo_hi_lo_8};
  wire [63:0]   res_hi_hi_lo_8 = {res_hi_hi_lo_hi_8, res_hi_hi_lo_lo_8};
  wire [15:0]   res_hi_hi_hi_lo_lo_8 = {dataGroup_57_8, dataGroup_56_8};
  wire [15:0]   res_hi_hi_hi_lo_hi_8 = {dataGroup_59_8, dataGroup_58_8};
  wire [31:0]   res_hi_hi_hi_lo_8 = {res_hi_hi_hi_lo_hi_8, res_hi_hi_hi_lo_lo_8};
  wire [15:0]   res_hi_hi_hi_hi_lo_8 = {dataGroup_61_8, dataGroup_60_8};
  wire [15:0]   res_hi_hi_hi_hi_hi_8 = {dataGroup_63_8, dataGroup_62_8};
  wire [31:0]   res_hi_hi_hi_hi_8 = {res_hi_hi_hi_hi_hi_8, res_hi_hi_hi_hi_lo_8};
  wire [63:0]   res_hi_hi_hi_8 = {res_hi_hi_hi_hi_8, res_hi_hi_hi_lo_8};
  wire [127:0]  res_hi_hi_8 = {res_hi_hi_hi_8, res_hi_hi_lo_8};
  wire [255:0]  res_hi_8 = {res_hi_hi_8, res_hi_lo_8};
  wire [511:0]  res_26 = {res_hi_8, res_lo_8};
  wire [2047:0] dataGroup_lo_576 = {dataGroup_lo_hi_576, dataGroup_lo_lo_576};
  wire [2047:0] dataGroup_hi_576 = {dataGroup_hi_hi_576, dataGroup_hi_lo_576};
  wire [7:0]    dataGroup_0_9 = dataGroup_lo_576[31:24];
  wire [2047:0] dataGroup_lo_577 = {dataGroup_lo_hi_577, dataGroup_lo_lo_577};
  wire [2047:0] dataGroup_hi_577 = {dataGroup_hi_hi_577, dataGroup_hi_lo_577};
  wire [7:0]    dataGroup_1_9 = dataGroup_lo_577[63:56];
  wire [2047:0] dataGroup_lo_578 = {dataGroup_lo_hi_578, dataGroup_lo_lo_578};
  wire [2047:0] dataGroup_hi_578 = {dataGroup_hi_hi_578, dataGroup_hi_lo_578};
  wire [7:0]    dataGroup_2_9 = dataGroup_lo_578[95:88];
  wire [2047:0] dataGroup_lo_579 = {dataGroup_lo_hi_579, dataGroup_lo_lo_579};
  wire [2047:0] dataGroup_hi_579 = {dataGroup_hi_hi_579, dataGroup_hi_lo_579};
  wire [7:0]    dataGroup_3_9 = dataGroup_lo_579[127:120];
  wire [2047:0] dataGroup_lo_580 = {dataGroup_lo_hi_580, dataGroup_lo_lo_580};
  wire [2047:0] dataGroup_hi_580 = {dataGroup_hi_hi_580, dataGroup_hi_lo_580};
  wire [7:0]    dataGroup_4_9 = dataGroup_lo_580[159:152];
  wire [2047:0] dataGroup_lo_581 = {dataGroup_lo_hi_581, dataGroup_lo_lo_581};
  wire [2047:0] dataGroup_hi_581 = {dataGroup_hi_hi_581, dataGroup_hi_lo_581};
  wire [7:0]    dataGroup_5_9 = dataGroup_lo_581[191:184];
  wire [2047:0] dataGroup_lo_582 = {dataGroup_lo_hi_582, dataGroup_lo_lo_582};
  wire [2047:0] dataGroup_hi_582 = {dataGroup_hi_hi_582, dataGroup_hi_lo_582};
  wire [7:0]    dataGroup_6_9 = dataGroup_lo_582[223:216];
  wire [2047:0] dataGroup_lo_583 = {dataGroup_lo_hi_583, dataGroup_lo_lo_583};
  wire [2047:0] dataGroup_hi_583 = {dataGroup_hi_hi_583, dataGroup_hi_lo_583};
  wire [7:0]    dataGroup_7_9 = dataGroup_lo_583[255:248];
  wire [2047:0] dataGroup_lo_584 = {dataGroup_lo_hi_584, dataGroup_lo_lo_584};
  wire [2047:0] dataGroup_hi_584 = {dataGroup_hi_hi_584, dataGroup_hi_lo_584};
  wire [7:0]    dataGroup_8_9 = dataGroup_lo_584[287:280];
  wire [2047:0] dataGroup_lo_585 = {dataGroup_lo_hi_585, dataGroup_lo_lo_585};
  wire [2047:0] dataGroup_hi_585 = {dataGroup_hi_hi_585, dataGroup_hi_lo_585};
  wire [7:0]    dataGroup_9_9 = dataGroup_lo_585[319:312];
  wire [2047:0] dataGroup_lo_586 = {dataGroup_lo_hi_586, dataGroup_lo_lo_586};
  wire [2047:0] dataGroup_hi_586 = {dataGroup_hi_hi_586, dataGroup_hi_lo_586};
  wire [7:0]    dataGroup_10_9 = dataGroup_lo_586[351:344];
  wire [2047:0] dataGroup_lo_587 = {dataGroup_lo_hi_587, dataGroup_lo_lo_587};
  wire [2047:0] dataGroup_hi_587 = {dataGroup_hi_hi_587, dataGroup_hi_lo_587};
  wire [7:0]    dataGroup_11_9 = dataGroup_lo_587[383:376];
  wire [2047:0] dataGroup_lo_588 = {dataGroup_lo_hi_588, dataGroup_lo_lo_588};
  wire [2047:0] dataGroup_hi_588 = {dataGroup_hi_hi_588, dataGroup_hi_lo_588};
  wire [7:0]    dataGroup_12_9 = dataGroup_lo_588[415:408];
  wire [2047:0] dataGroup_lo_589 = {dataGroup_lo_hi_589, dataGroup_lo_lo_589};
  wire [2047:0] dataGroup_hi_589 = {dataGroup_hi_hi_589, dataGroup_hi_lo_589};
  wire [7:0]    dataGroup_13_9 = dataGroup_lo_589[447:440];
  wire [2047:0] dataGroup_lo_590 = {dataGroup_lo_hi_590, dataGroup_lo_lo_590};
  wire [2047:0] dataGroup_hi_590 = {dataGroup_hi_hi_590, dataGroup_hi_lo_590};
  wire [7:0]    dataGroup_14_9 = dataGroup_lo_590[479:472];
  wire [2047:0] dataGroup_lo_591 = {dataGroup_lo_hi_591, dataGroup_lo_lo_591};
  wire [2047:0] dataGroup_hi_591 = {dataGroup_hi_hi_591, dataGroup_hi_lo_591};
  wire [7:0]    dataGroup_15_9 = dataGroup_lo_591[511:504];
  wire [2047:0] dataGroup_lo_592 = {dataGroup_lo_hi_592, dataGroup_lo_lo_592};
  wire [2047:0] dataGroup_hi_592 = {dataGroup_hi_hi_592, dataGroup_hi_lo_592};
  wire [7:0]    dataGroup_16_9 = dataGroup_lo_592[543:536];
  wire [2047:0] dataGroup_lo_593 = {dataGroup_lo_hi_593, dataGroup_lo_lo_593};
  wire [2047:0] dataGroup_hi_593 = {dataGroup_hi_hi_593, dataGroup_hi_lo_593};
  wire [7:0]    dataGroup_17_9 = dataGroup_lo_593[575:568];
  wire [2047:0] dataGroup_lo_594 = {dataGroup_lo_hi_594, dataGroup_lo_lo_594};
  wire [2047:0] dataGroup_hi_594 = {dataGroup_hi_hi_594, dataGroup_hi_lo_594};
  wire [7:0]    dataGroup_18_9 = dataGroup_lo_594[607:600];
  wire [2047:0] dataGroup_lo_595 = {dataGroup_lo_hi_595, dataGroup_lo_lo_595};
  wire [2047:0] dataGroup_hi_595 = {dataGroup_hi_hi_595, dataGroup_hi_lo_595};
  wire [7:0]    dataGroup_19_9 = dataGroup_lo_595[639:632];
  wire [2047:0] dataGroup_lo_596 = {dataGroup_lo_hi_596, dataGroup_lo_lo_596};
  wire [2047:0] dataGroup_hi_596 = {dataGroup_hi_hi_596, dataGroup_hi_lo_596};
  wire [7:0]    dataGroup_20_9 = dataGroup_lo_596[671:664];
  wire [2047:0] dataGroup_lo_597 = {dataGroup_lo_hi_597, dataGroup_lo_lo_597};
  wire [2047:0] dataGroup_hi_597 = {dataGroup_hi_hi_597, dataGroup_hi_lo_597};
  wire [7:0]    dataGroup_21_9 = dataGroup_lo_597[703:696];
  wire [2047:0] dataGroup_lo_598 = {dataGroup_lo_hi_598, dataGroup_lo_lo_598};
  wire [2047:0] dataGroup_hi_598 = {dataGroup_hi_hi_598, dataGroup_hi_lo_598};
  wire [7:0]    dataGroup_22_9 = dataGroup_lo_598[735:728];
  wire [2047:0] dataGroup_lo_599 = {dataGroup_lo_hi_599, dataGroup_lo_lo_599};
  wire [2047:0] dataGroup_hi_599 = {dataGroup_hi_hi_599, dataGroup_hi_lo_599};
  wire [7:0]    dataGroup_23_9 = dataGroup_lo_599[767:760];
  wire [2047:0] dataGroup_lo_600 = {dataGroup_lo_hi_600, dataGroup_lo_lo_600};
  wire [2047:0] dataGroup_hi_600 = {dataGroup_hi_hi_600, dataGroup_hi_lo_600};
  wire [7:0]    dataGroup_24_9 = dataGroup_lo_600[799:792];
  wire [2047:0] dataGroup_lo_601 = {dataGroup_lo_hi_601, dataGroup_lo_lo_601};
  wire [2047:0] dataGroup_hi_601 = {dataGroup_hi_hi_601, dataGroup_hi_lo_601};
  wire [7:0]    dataGroup_25_9 = dataGroup_lo_601[831:824];
  wire [2047:0] dataGroup_lo_602 = {dataGroup_lo_hi_602, dataGroup_lo_lo_602};
  wire [2047:0] dataGroup_hi_602 = {dataGroup_hi_hi_602, dataGroup_hi_lo_602};
  wire [7:0]    dataGroup_26_9 = dataGroup_lo_602[863:856];
  wire [2047:0] dataGroup_lo_603 = {dataGroup_lo_hi_603, dataGroup_lo_lo_603};
  wire [2047:0] dataGroup_hi_603 = {dataGroup_hi_hi_603, dataGroup_hi_lo_603};
  wire [7:0]    dataGroup_27_9 = dataGroup_lo_603[895:888];
  wire [2047:0] dataGroup_lo_604 = {dataGroup_lo_hi_604, dataGroup_lo_lo_604};
  wire [2047:0] dataGroup_hi_604 = {dataGroup_hi_hi_604, dataGroup_hi_lo_604};
  wire [7:0]    dataGroup_28_9 = dataGroup_lo_604[927:920];
  wire [2047:0] dataGroup_lo_605 = {dataGroup_lo_hi_605, dataGroup_lo_lo_605};
  wire [2047:0] dataGroup_hi_605 = {dataGroup_hi_hi_605, dataGroup_hi_lo_605};
  wire [7:0]    dataGroup_29_9 = dataGroup_lo_605[959:952];
  wire [2047:0] dataGroup_lo_606 = {dataGroup_lo_hi_606, dataGroup_lo_lo_606};
  wire [2047:0] dataGroup_hi_606 = {dataGroup_hi_hi_606, dataGroup_hi_lo_606};
  wire [7:0]    dataGroup_30_9 = dataGroup_lo_606[991:984];
  wire [2047:0] dataGroup_lo_607 = {dataGroup_lo_hi_607, dataGroup_lo_lo_607};
  wire [2047:0] dataGroup_hi_607 = {dataGroup_hi_hi_607, dataGroup_hi_lo_607};
  wire [7:0]    dataGroup_31_9 = dataGroup_lo_607[1023:1016];
  wire [2047:0] dataGroup_lo_608 = {dataGroup_lo_hi_608, dataGroup_lo_lo_608};
  wire [2047:0] dataGroup_hi_608 = {dataGroup_hi_hi_608, dataGroup_hi_lo_608};
  wire [7:0]    dataGroup_32_9 = dataGroup_lo_608[1055:1048];
  wire [2047:0] dataGroup_lo_609 = {dataGroup_lo_hi_609, dataGroup_lo_lo_609};
  wire [2047:0] dataGroup_hi_609 = {dataGroup_hi_hi_609, dataGroup_hi_lo_609};
  wire [7:0]    dataGroup_33_9 = dataGroup_lo_609[1087:1080];
  wire [2047:0] dataGroup_lo_610 = {dataGroup_lo_hi_610, dataGroup_lo_lo_610};
  wire [2047:0] dataGroup_hi_610 = {dataGroup_hi_hi_610, dataGroup_hi_lo_610};
  wire [7:0]    dataGroup_34_9 = dataGroup_lo_610[1119:1112];
  wire [2047:0] dataGroup_lo_611 = {dataGroup_lo_hi_611, dataGroup_lo_lo_611};
  wire [2047:0] dataGroup_hi_611 = {dataGroup_hi_hi_611, dataGroup_hi_lo_611};
  wire [7:0]    dataGroup_35_9 = dataGroup_lo_611[1151:1144];
  wire [2047:0] dataGroup_lo_612 = {dataGroup_lo_hi_612, dataGroup_lo_lo_612};
  wire [2047:0] dataGroup_hi_612 = {dataGroup_hi_hi_612, dataGroup_hi_lo_612};
  wire [7:0]    dataGroup_36_9 = dataGroup_lo_612[1183:1176];
  wire [2047:0] dataGroup_lo_613 = {dataGroup_lo_hi_613, dataGroup_lo_lo_613};
  wire [2047:0] dataGroup_hi_613 = {dataGroup_hi_hi_613, dataGroup_hi_lo_613};
  wire [7:0]    dataGroup_37_9 = dataGroup_lo_613[1215:1208];
  wire [2047:0] dataGroup_lo_614 = {dataGroup_lo_hi_614, dataGroup_lo_lo_614};
  wire [2047:0] dataGroup_hi_614 = {dataGroup_hi_hi_614, dataGroup_hi_lo_614};
  wire [7:0]    dataGroup_38_9 = dataGroup_lo_614[1247:1240];
  wire [2047:0] dataGroup_lo_615 = {dataGroup_lo_hi_615, dataGroup_lo_lo_615};
  wire [2047:0] dataGroup_hi_615 = {dataGroup_hi_hi_615, dataGroup_hi_lo_615};
  wire [7:0]    dataGroup_39_9 = dataGroup_lo_615[1279:1272];
  wire [2047:0] dataGroup_lo_616 = {dataGroup_lo_hi_616, dataGroup_lo_lo_616};
  wire [2047:0] dataGroup_hi_616 = {dataGroup_hi_hi_616, dataGroup_hi_lo_616};
  wire [7:0]    dataGroup_40_9 = dataGroup_lo_616[1311:1304];
  wire [2047:0] dataGroup_lo_617 = {dataGroup_lo_hi_617, dataGroup_lo_lo_617};
  wire [2047:0] dataGroup_hi_617 = {dataGroup_hi_hi_617, dataGroup_hi_lo_617};
  wire [7:0]    dataGroup_41_9 = dataGroup_lo_617[1343:1336];
  wire [2047:0] dataGroup_lo_618 = {dataGroup_lo_hi_618, dataGroup_lo_lo_618};
  wire [2047:0] dataGroup_hi_618 = {dataGroup_hi_hi_618, dataGroup_hi_lo_618};
  wire [7:0]    dataGroup_42_9 = dataGroup_lo_618[1375:1368];
  wire [2047:0] dataGroup_lo_619 = {dataGroup_lo_hi_619, dataGroup_lo_lo_619};
  wire [2047:0] dataGroup_hi_619 = {dataGroup_hi_hi_619, dataGroup_hi_lo_619};
  wire [7:0]    dataGroup_43_9 = dataGroup_lo_619[1407:1400];
  wire [2047:0] dataGroup_lo_620 = {dataGroup_lo_hi_620, dataGroup_lo_lo_620};
  wire [2047:0] dataGroup_hi_620 = {dataGroup_hi_hi_620, dataGroup_hi_lo_620};
  wire [7:0]    dataGroup_44_9 = dataGroup_lo_620[1439:1432];
  wire [2047:0] dataGroup_lo_621 = {dataGroup_lo_hi_621, dataGroup_lo_lo_621};
  wire [2047:0] dataGroup_hi_621 = {dataGroup_hi_hi_621, dataGroup_hi_lo_621};
  wire [7:0]    dataGroup_45_9 = dataGroup_lo_621[1471:1464];
  wire [2047:0] dataGroup_lo_622 = {dataGroup_lo_hi_622, dataGroup_lo_lo_622};
  wire [2047:0] dataGroup_hi_622 = {dataGroup_hi_hi_622, dataGroup_hi_lo_622};
  wire [7:0]    dataGroup_46_9 = dataGroup_lo_622[1503:1496];
  wire [2047:0] dataGroup_lo_623 = {dataGroup_lo_hi_623, dataGroup_lo_lo_623};
  wire [2047:0] dataGroup_hi_623 = {dataGroup_hi_hi_623, dataGroup_hi_lo_623};
  wire [7:0]    dataGroup_47_9 = dataGroup_lo_623[1535:1528];
  wire [2047:0] dataGroup_lo_624 = {dataGroup_lo_hi_624, dataGroup_lo_lo_624};
  wire [2047:0] dataGroup_hi_624 = {dataGroup_hi_hi_624, dataGroup_hi_lo_624};
  wire [7:0]    dataGroup_48_9 = dataGroup_lo_624[1567:1560];
  wire [2047:0] dataGroup_lo_625 = {dataGroup_lo_hi_625, dataGroup_lo_lo_625};
  wire [2047:0] dataGroup_hi_625 = {dataGroup_hi_hi_625, dataGroup_hi_lo_625};
  wire [7:0]    dataGroup_49_9 = dataGroup_lo_625[1599:1592];
  wire [2047:0] dataGroup_lo_626 = {dataGroup_lo_hi_626, dataGroup_lo_lo_626};
  wire [2047:0] dataGroup_hi_626 = {dataGroup_hi_hi_626, dataGroup_hi_lo_626};
  wire [7:0]    dataGroup_50_9 = dataGroup_lo_626[1631:1624];
  wire [2047:0] dataGroup_lo_627 = {dataGroup_lo_hi_627, dataGroup_lo_lo_627};
  wire [2047:0] dataGroup_hi_627 = {dataGroup_hi_hi_627, dataGroup_hi_lo_627};
  wire [7:0]    dataGroup_51_9 = dataGroup_lo_627[1663:1656];
  wire [2047:0] dataGroup_lo_628 = {dataGroup_lo_hi_628, dataGroup_lo_lo_628};
  wire [2047:0] dataGroup_hi_628 = {dataGroup_hi_hi_628, dataGroup_hi_lo_628};
  wire [7:0]    dataGroup_52_9 = dataGroup_lo_628[1695:1688];
  wire [2047:0] dataGroup_lo_629 = {dataGroup_lo_hi_629, dataGroup_lo_lo_629};
  wire [2047:0] dataGroup_hi_629 = {dataGroup_hi_hi_629, dataGroup_hi_lo_629};
  wire [7:0]    dataGroup_53_9 = dataGroup_lo_629[1727:1720];
  wire [2047:0] dataGroup_lo_630 = {dataGroup_lo_hi_630, dataGroup_lo_lo_630};
  wire [2047:0] dataGroup_hi_630 = {dataGroup_hi_hi_630, dataGroup_hi_lo_630};
  wire [7:0]    dataGroup_54_9 = dataGroup_lo_630[1759:1752];
  wire [2047:0] dataGroup_lo_631 = {dataGroup_lo_hi_631, dataGroup_lo_lo_631};
  wire [2047:0] dataGroup_hi_631 = {dataGroup_hi_hi_631, dataGroup_hi_lo_631};
  wire [7:0]    dataGroup_55_9 = dataGroup_lo_631[1791:1784];
  wire [2047:0] dataGroup_lo_632 = {dataGroup_lo_hi_632, dataGroup_lo_lo_632};
  wire [2047:0] dataGroup_hi_632 = {dataGroup_hi_hi_632, dataGroup_hi_lo_632};
  wire [7:0]    dataGroup_56_9 = dataGroup_lo_632[1823:1816];
  wire [2047:0] dataGroup_lo_633 = {dataGroup_lo_hi_633, dataGroup_lo_lo_633};
  wire [2047:0] dataGroup_hi_633 = {dataGroup_hi_hi_633, dataGroup_hi_lo_633};
  wire [7:0]    dataGroup_57_9 = dataGroup_lo_633[1855:1848];
  wire [2047:0] dataGroup_lo_634 = {dataGroup_lo_hi_634, dataGroup_lo_lo_634};
  wire [2047:0] dataGroup_hi_634 = {dataGroup_hi_hi_634, dataGroup_hi_lo_634};
  wire [7:0]    dataGroup_58_9 = dataGroup_lo_634[1887:1880];
  wire [2047:0] dataGroup_lo_635 = {dataGroup_lo_hi_635, dataGroup_lo_lo_635};
  wire [2047:0] dataGroup_hi_635 = {dataGroup_hi_hi_635, dataGroup_hi_lo_635};
  wire [7:0]    dataGroup_59_9 = dataGroup_lo_635[1919:1912];
  wire [2047:0] dataGroup_lo_636 = {dataGroup_lo_hi_636, dataGroup_lo_lo_636};
  wire [2047:0] dataGroup_hi_636 = {dataGroup_hi_hi_636, dataGroup_hi_lo_636};
  wire [7:0]    dataGroup_60_9 = dataGroup_lo_636[1951:1944];
  wire [2047:0] dataGroup_lo_637 = {dataGroup_lo_hi_637, dataGroup_lo_lo_637};
  wire [2047:0] dataGroup_hi_637 = {dataGroup_hi_hi_637, dataGroup_hi_lo_637};
  wire [7:0]    dataGroup_61_9 = dataGroup_lo_637[1983:1976];
  wire [2047:0] dataGroup_lo_638 = {dataGroup_lo_hi_638, dataGroup_lo_lo_638};
  wire [2047:0] dataGroup_hi_638 = {dataGroup_hi_hi_638, dataGroup_hi_lo_638};
  wire [7:0]    dataGroup_62_9 = dataGroup_lo_638[2015:2008];
  wire [2047:0] dataGroup_lo_639 = {dataGroup_lo_hi_639, dataGroup_lo_lo_639};
  wire [2047:0] dataGroup_hi_639 = {dataGroup_hi_hi_639, dataGroup_hi_lo_639};
  wire [7:0]    dataGroup_63_9 = dataGroup_lo_639[2047:2040];
  wire [15:0]   res_lo_lo_lo_lo_lo_9 = {dataGroup_1_9, dataGroup_0_9};
  wire [15:0]   res_lo_lo_lo_lo_hi_9 = {dataGroup_3_9, dataGroup_2_9};
  wire [31:0]   res_lo_lo_lo_lo_9 = {res_lo_lo_lo_lo_hi_9, res_lo_lo_lo_lo_lo_9};
  wire [15:0]   res_lo_lo_lo_hi_lo_9 = {dataGroup_5_9, dataGroup_4_9};
  wire [15:0]   res_lo_lo_lo_hi_hi_9 = {dataGroup_7_9, dataGroup_6_9};
  wire [31:0]   res_lo_lo_lo_hi_9 = {res_lo_lo_lo_hi_hi_9, res_lo_lo_lo_hi_lo_9};
  wire [63:0]   res_lo_lo_lo_9 = {res_lo_lo_lo_hi_9, res_lo_lo_lo_lo_9};
  wire [15:0]   res_lo_lo_hi_lo_lo_9 = {dataGroup_9_9, dataGroup_8_9};
  wire [15:0]   res_lo_lo_hi_lo_hi_9 = {dataGroup_11_9, dataGroup_10_9};
  wire [31:0]   res_lo_lo_hi_lo_9 = {res_lo_lo_hi_lo_hi_9, res_lo_lo_hi_lo_lo_9};
  wire [15:0]   res_lo_lo_hi_hi_lo_9 = {dataGroup_13_9, dataGroup_12_9};
  wire [15:0]   res_lo_lo_hi_hi_hi_9 = {dataGroup_15_9, dataGroup_14_9};
  wire [31:0]   res_lo_lo_hi_hi_9 = {res_lo_lo_hi_hi_hi_9, res_lo_lo_hi_hi_lo_9};
  wire [63:0]   res_lo_lo_hi_9 = {res_lo_lo_hi_hi_9, res_lo_lo_hi_lo_9};
  wire [127:0]  res_lo_lo_9 = {res_lo_lo_hi_9, res_lo_lo_lo_9};
  wire [15:0]   res_lo_hi_lo_lo_lo_9 = {dataGroup_17_9, dataGroup_16_9};
  wire [15:0]   res_lo_hi_lo_lo_hi_9 = {dataGroup_19_9, dataGroup_18_9};
  wire [31:0]   res_lo_hi_lo_lo_9 = {res_lo_hi_lo_lo_hi_9, res_lo_hi_lo_lo_lo_9};
  wire [15:0]   res_lo_hi_lo_hi_lo_9 = {dataGroup_21_9, dataGroup_20_9};
  wire [15:0]   res_lo_hi_lo_hi_hi_9 = {dataGroup_23_9, dataGroup_22_9};
  wire [31:0]   res_lo_hi_lo_hi_9 = {res_lo_hi_lo_hi_hi_9, res_lo_hi_lo_hi_lo_9};
  wire [63:0]   res_lo_hi_lo_9 = {res_lo_hi_lo_hi_9, res_lo_hi_lo_lo_9};
  wire [15:0]   res_lo_hi_hi_lo_lo_9 = {dataGroup_25_9, dataGroup_24_9};
  wire [15:0]   res_lo_hi_hi_lo_hi_9 = {dataGroup_27_9, dataGroup_26_9};
  wire [31:0]   res_lo_hi_hi_lo_9 = {res_lo_hi_hi_lo_hi_9, res_lo_hi_hi_lo_lo_9};
  wire [15:0]   res_lo_hi_hi_hi_lo_9 = {dataGroup_29_9, dataGroup_28_9};
  wire [15:0]   res_lo_hi_hi_hi_hi_9 = {dataGroup_31_9, dataGroup_30_9};
  wire [31:0]   res_lo_hi_hi_hi_9 = {res_lo_hi_hi_hi_hi_9, res_lo_hi_hi_hi_lo_9};
  wire [63:0]   res_lo_hi_hi_9 = {res_lo_hi_hi_hi_9, res_lo_hi_hi_lo_9};
  wire [127:0]  res_lo_hi_9 = {res_lo_hi_hi_9, res_lo_hi_lo_9};
  wire [255:0]  res_lo_9 = {res_lo_hi_9, res_lo_lo_9};
  wire [15:0]   res_hi_lo_lo_lo_lo_9 = {dataGroup_33_9, dataGroup_32_9};
  wire [15:0]   res_hi_lo_lo_lo_hi_9 = {dataGroup_35_9, dataGroup_34_9};
  wire [31:0]   res_hi_lo_lo_lo_9 = {res_hi_lo_lo_lo_hi_9, res_hi_lo_lo_lo_lo_9};
  wire [15:0]   res_hi_lo_lo_hi_lo_9 = {dataGroup_37_9, dataGroup_36_9};
  wire [15:0]   res_hi_lo_lo_hi_hi_9 = {dataGroup_39_9, dataGroup_38_9};
  wire [31:0]   res_hi_lo_lo_hi_9 = {res_hi_lo_lo_hi_hi_9, res_hi_lo_lo_hi_lo_9};
  wire [63:0]   res_hi_lo_lo_9 = {res_hi_lo_lo_hi_9, res_hi_lo_lo_lo_9};
  wire [15:0]   res_hi_lo_hi_lo_lo_9 = {dataGroup_41_9, dataGroup_40_9};
  wire [15:0]   res_hi_lo_hi_lo_hi_9 = {dataGroup_43_9, dataGroup_42_9};
  wire [31:0]   res_hi_lo_hi_lo_9 = {res_hi_lo_hi_lo_hi_9, res_hi_lo_hi_lo_lo_9};
  wire [15:0]   res_hi_lo_hi_hi_lo_9 = {dataGroup_45_9, dataGroup_44_9};
  wire [15:0]   res_hi_lo_hi_hi_hi_9 = {dataGroup_47_9, dataGroup_46_9};
  wire [31:0]   res_hi_lo_hi_hi_9 = {res_hi_lo_hi_hi_hi_9, res_hi_lo_hi_hi_lo_9};
  wire [63:0]   res_hi_lo_hi_9 = {res_hi_lo_hi_hi_9, res_hi_lo_hi_lo_9};
  wire [127:0]  res_hi_lo_9 = {res_hi_lo_hi_9, res_hi_lo_lo_9};
  wire [15:0]   res_hi_hi_lo_lo_lo_9 = {dataGroup_49_9, dataGroup_48_9};
  wire [15:0]   res_hi_hi_lo_lo_hi_9 = {dataGroup_51_9, dataGroup_50_9};
  wire [31:0]   res_hi_hi_lo_lo_9 = {res_hi_hi_lo_lo_hi_9, res_hi_hi_lo_lo_lo_9};
  wire [15:0]   res_hi_hi_lo_hi_lo_9 = {dataGroup_53_9, dataGroup_52_9};
  wire [15:0]   res_hi_hi_lo_hi_hi_9 = {dataGroup_55_9, dataGroup_54_9};
  wire [31:0]   res_hi_hi_lo_hi_9 = {res_hi_hi_lo_hi_hi_9, res_hi_hi_lo_hi_lo_9};
  wire [63:0]   res_hi_hi_lo_9 = {res_hi_hi_lo_hi_9, res_hi_hi_lo_lo_9};
  wire [15:0]   res_hi_hi_hi_lo_lo_9 = {dataGroup_57_9, dataGroup_56_9};
  wire [15:0]   res_hi_hi_hi_lo_hi_9 = {dataGroup_59_9, dataGroup_58_9};
  wire [31:0]   res_hi_hi_hi_lo_9 = {res_hi_hi_hi_lo_hi_9, res_hi_hi_hi_lo_lo_9};
  wire [15:0]   res_hi_hi_hi_hi_lo_9 = {dataGroup_61_9, dataGroup_60_9};
  wire [15:0]   res_hi_hi_hi_hi_hi_9 = {dataGroup_63_9, dataGroup_62_9};
  wire [31:0]   res_hi_hi_hi_hi_9 = {res_hi_hi_hi_hi_hi_9, res_hi_hi_hi_hi_lo_9};
  wire [63:0]   res_hi_hi_hi_9 = {res_hi_hi_hi_hi_9, res_hi_hi_hi_lo_9};
  wire [127:0]  res_hi_hi_9 = {res_hi_hi_hi_9, res_hi_hi_lo_9};
  wire [255:0]  res_hi_9 = {res_hi_hi_9, res_hi_lo_9};
  wire [511:0]  res_27 = {res_hi_9, res_lo_9};
  wire [1023:0] lo_lo_3 = {res_25, res_24};
  wire [1023:0] lo_hi_3 = {res_27, res_26};
  wire [2047:0] lo_3 = {lo_hi_3, lo_lo_3};
  wire [4095:0] regroupLoadData_0_3 = {2048'h0, lo_3};
  wire [2047:0] dataGroup_lo_640 = {dataGroup_lo_hi_640, dataGroup_lo_lo_640};
  wire [2047:0] dataGroup_hi_640 = {dataGroup_hi_hi_640, dataGroup_hi_lo_640};
  wire [7:0]    dataGroup_0_10 = dataGroup_lo_640[7:0];
  wire [2047:0] dataGroup_lo_641 = {dataGroup_lo_hi_641, dataGroup_lo_lo_641};
  wire [2047:0] dataGroup_hi_641 = {dataGroup_hi_hi_641, dataGroup_hi_lo_641};
  wire [7:0]    dataGroup_1_10 = dataGroup_lo_641[47:40];
  wire [2047:0] dataGroup_lo_642 = {dataGroup_lo_hi_642, dataGroup_lo_lo_642};
  wire [2047:0] dataGroup_hi_642 = {dataGroup_hi_hi_642, dataGroup_hi_lo_642};
  wire [7:0]    dataGroup_2_10 = dataGroup_lo_642[87:80];
  wire [2047:0] dataGroup_lo_643 = {dataGroup_lo_hi_643, dataGroup_lo_lo_643};
  wire [2047:0] dataGroup_hi_643 = {dataGroup_hi_hi_643, dataGroup_hi_lo_643};
  wire [7:0]    dataGroup_3_10 = dataGroup_lo_643[127:120];
  wire [2047:0] dataGroup_lo_644 = {dataGroup_lo_hi_644, dataGroup_lo_lo_644};
  wire [2047:0] dataGroup_hi_644 = {dataGroup_hi_hi_644, dataGroup_hi_lo_644};
  wire [7:0]    dataGroup_4_10 = dataGroup_lo_644[167:160];
  wire [2047:0] dataGroup_lo_645 = {dataGroup_lo_hi_645, dataGroup_lo_lo_645};
  wire [2047:0] dataGroup_hi_645 = {dataGroup_hi_hi_645, dataGroup_hi_lo_645};
  wire [7:0]    dataGroup_5_10 = dataGroup_lo_645[207:200];
  wire [2047:0] dataGroup_lo_646 = {dataGroup_lo_hi_646, dataGroup_lo_lo_646};
  wire [2047:0] dataGroup_hi_646 = {dataGroup_hi_hi_646, dataGroup_hi_lo_646};
  wire [7:0]    dataGroup_6_10 = dataGroup_lo_646[247:240];
  wire [2047:0] dataGroup_lo_647 = {dataGroup_lo_hi_647, dataGroup_lo_lo_647};
  wire [2047:0] dataGroup_hi_647 = {dataGroup_hi_hi_647, dataGroup_hi_lo_647};
  wire [7:0]    dataGroup_7_10 = dataGroup_lo_647[287:280];
  wire [2047:0] dataGroup_lo_648 = {dataGroup_lo_hi_648, dataGroup_lo_lo_648};
  wire [2047:0] dataGroup_hi_648 = {dataGroup_hi_hi_648, dataGroup_hi_lo_648};
  wire [7:0]    dataGroup_8_10 = dataGroup_lo_648[327:320];
  wire [2047:0] dataGroup_lo_649 = {dataGroup_lo_hi_649, dataGroup_lo_lo_649};
  wire [2047:0] dataGroup_hi_649 = {dataGroup_hi_hi_649, dataGroup_hi_lo_649};
  wire [7:0]    dataGroup_9_10 = dataGroup_lo_649[367:360];
  wire [2047:0] dataGroup_lo_650 = {dataGroup_lo_hi_650, dataGroup_lo_lo_650};
  wire [2047:0] dataGroup_hi_650 = {dataGroup_hi_hi_650, dataGroup_hi_lo_650};
  wire [7:0]    dataGroup_10_10 = dataGroup_lo_650[407:400];
  wire [2047:0] dataGroup_lo_651 = {dataGroup_lo_hi_651, dataGroup_lo_lo_651};
  wire [2047:0] dataGroup_hi_651 = {dataGroup_hi_hi_651, dataGroup_hi_lo_651};
  wire [7:0]    dataGroup_11_10 = dataGroup_lo_651[447:440];
  wire [2047:0] dataGroup_lo_652 = {dataGroup_lo_hi_652, dataGroup_lo_lo_652};
  wire [2047:0] dataGroup_hi_652 = {dataGroup_hi_hi_652, dataGroup_hi_lo_652};
  wire [7:0]    dataGroup_12_10 = dataGroup_lo_652[487:480];
  wire [2047:0] dataGroup_lo_653 = {dataGroup_lo_hi_653, dataGroup_lo_lo_653};
  wire [2047:0] dataGroup_hi_653 = {dataGroup_hi_hi_653, dataGroup_hi_lo_653};
  wire [7:0]    dataGroup_13_10 = dataGroup_lo_653[527:520];
  wire [2047:0] dataGroup_lo_654 = {dataGroup_lo_hi_654, dataGroup_lo_lo_654};
  wire [2047:0] dataGroup_hi_654 = {dataGroup_hi_hi_654, dataGroup_hi_lo_654};
  wire [7:0]    dataGroup_14_10 = dataGroup_lo_654[567:560];
  wire [2047:0] dataGroup_lo_655 = {dataGroup_lo_hi_655, dataGroup_lo_lo_655};
  wire [2047:0] dataGroup_hi_655 = {dataGroup_hi_hi_655, dataGroup_hi_lo_655};
  wire [7:0]    dataGroup_15_10 = dataGroup_lo_655[607:600];
  wire [2047:0] dataGroup_lo_656 = {dataGroup_lo_hi_656, dataGroup_lo_lo_656};
  wire [2047:0] dataGroup_hi_656 = {dataGroup_hi_hi_656, dataGroup_hi_lo_656};
  wire [7:0]    dataGroup_16_10 = dataGroup_lo_656[647:640];
  wire [2047:0] dataGroup_lo_657 = {dataGroup_lo_hi_657, dataGroup_lo_lo_657};
  wire [2047:0] dataGroup_hi_657 = {dataGroup_hi_hi_657, dataGroup_hi_lo_657};
  wire [7:0]    dataGroup_17_10 = dataGroup_lo_657[687:680];
  wire [2047:0] dataGroup_lo_658 = {dataGroup_lo_hi_658, dataGroup_lo_lo_658};
  wire [2047:0] dataGroup_hi_658 = {dataGroup_hi_hi_658, dataGroup_hi_lo_658};
  wire [7:0]    dataGroup_18_10 = dataGroup_lo_658[727:720];
  wire [2047:0] dataGroup_lo_659 = {dataGroup_lo_hi_659, dataGroup_lo_lo_659};
  wire [2047:0] dataGroup_hi_659 = {dataGroup_hi_hi_659, dataGroup_hi_lo_659};
  wire [7:0]    dataGroup_19_10 = dataGroup_lo_659[767:760];
  wire [2047:0] dataGroup_lo_660 = {dataGroup_lo_hi_660, dataGroup_lo_lo_660};
  wire [2047:0] dataGroup_hi_660 = {dataGroup_hi_hi_660, dataGroup_hi_lo_660};
  wire [7:0]    dataGroup_20_10 = dataGroup_lo_660[807:800];
  wire [2047:0] dataGroup_lo_661 = {dataGroup_lo_hi_661, dataGroup_lo_lo_661};
  wire [2047:0] dataGroup_hi_661 = {dataGroup_hi_hi_661, dataGroup_hi_lo_661};
  wire [7:0]    dataGroup_21_10 = dataGroup_lo_661[847:840];
  wire [2047:0] dataGroup_lo_662 = {dataGroup_lo_hi_662, dataGroup_lo_lo_662};
  wire [2047:0] dataGroup_hi_662 = {dataGroup_hi_hi_662, dataGroup_hi_lo_662};
  wire [7:0]    dataGroup_22_10 = dataGroup_lo_662[887:880];
  wire [2047:0] dataGroup_lo_663 = {dataGroup_lo_hi_663, dataGroup_lo_lo_663};
  wire [2047:0] dataGroup_hi_663 = {dataGroup_hi_hi_663, dataGroup_hi_lo_663};
  wire [7:0]    dataGroup_23_10 = dataGroup_lo_663[927:920];
  wire [2047:0] dataGroup_lo_664 = {dataGroup_lo_hi_664, dataGroup_lo_lo_664};
  wire [2047:0] dataGroup_hi_664 = {dataGroup_hi_hi_664, dataGroup_hi_lo_664};
  wire [7:0]    dataGroup_24_10 = dataGroup_lo_664[967:960];
  wire [2047:0] dataGroup_lo_665 = {dataGroup_lo_hi_665, dataGroup_lo_lo_665};
  wire [2047:0] dataGroup_hi_665 = {dataGroup_hi_hi_665, dataGroup_hi_lo_665};
  wire [7:0]    dataGroup_25_10 = dataGroup_lo_665[1007:1000];
  wire [2047:0] dataGroup_lo_666 = {dataGroup_lo_hi_666, dataGroup_lo_lo_666};
  wire [2047:0] dataGroup_hi_666 = {dataGroup_hi_hi_666, dataGroup_hi_lo_666};
  wire [7:0]    dataGroup_26_10 = dataGroup_lo_666[1047:1040];
  wire [2047:0] dataGroup_lo_667 = {dataGroup_lo_hi_667, dataGroup_lo_lo_667};
  wire [2047:0] dataGroup_hi_667 = {dataGroup_hi_hi_667, dataGroup_hi_lo_667};
  wire [7:0]    dataGroup_27_10 = dataGroup_lo_667[1087:1080];
  wire [2047:0] dataGroup_lo_668 = {dataGroup_lo_hi_668, dataGroup_lo_lo_668};
  wire [2047:0] dataGroup_hi_668 = {dataGroup_hi_hi_668, dataGroup_hi_lo_668};
  wire [7:0]    dataGroup_28_10 = dataGroup_lo_668[1127:1120];
  wire [2047:0] dataGroup_lo_669 = {dataGroup_lo_hi_669, dataGroup_lo_lo_669};
  wire [2047:0] dataGroup_hi_669 = {dataGroup_hi_hi_669, dataGroup_hi_lo_669};
  wire [7:0]    dataGroup_29_10 = dataGroup_lo_669[1167:1160];
  wire [2047:0] dataGroup_lo_670 = {dataGroup_lo_hi_670, dataGroup_lo_lo_670};
  wire [2047:0] dataGroup_hi_670 = {dataGroup_hi_hi_670, dataGroup_hi_lo_670};
  wire [7:0]    dataGroup_30_10 = dataGroup_lo_670[1207:1200];
  wire [2047:0] dataGroup_lo_671 = {dataGroup_lo_hi_671, dataGroup_lo_lo_671};
  wire [2047:0] dataGroup_hi_671 = {dataGroup_hi_hi_671, dataGroup_hi_lo_671};
  wire [7:0]    dataGroup_31_10 = dataGroup_lo_671[1247:1240];
  wire [2047:0] dataGroup_lo_672 = {dataGroup_lo_hi_672, dataGroup_lo_lo_672};
  wire [2047:0] dataGroup_hi_672 = {dataGroup_hi_hi_672, dataGroup_hi_lo_672};
  wire [7:0]    dataGroup_32_10 = dataGroup_lo_672[1287:1280];
  wire [2047:0] dataGroup_lo_673 = {dataGroup_lo_hi_673, dataGroup_lo_lo_673};
  wire [2047:0] dataGroup_hi_673 = {dataGroup_hi_hi_673, dataGroup_hi_lo_673};
  wire [7:0]    dataGroup_33_10 = dataGroup_lo_673[1327:1320];
  wire [2047:0] dataGroup_lo_674 = {dataGroup_lo_hi_674, dataGroup_lo_lo_674};
  wire [2047:0] dataGroup_hi_674 = {dataGroup_hi_hi_674, dataGroup_hi_lo_674};
  wire [7:0]    dataGroup_34_10 = dataGroup_lo_674[1367:1360];
  wire [2047:0] dataGroup_lo_675 = {dataGroup_lo_hi_675, dataGroup_lo_lo_675};
  wire [2047:0] dataGroup_hi_675 = {dataGroup_hi_hi_675, dataGroup_hi_lo_675};
  wire [7:0]    dataGroup_35_10 = dataGroup_lo_675[1407:1400];
  wire [2047:0] dataGroup_lo_676 = {dataGroup_lo_hi_676, dataGroup_lo_lo_676};
  wire [2047:0] dataGroup_hi_676 = {dataGroup_hi_hi_676, dataGroup_hi_lo_676};
  wire [7:0]    dataGroup_36_10 = dataGroup_lo_676[1447:1440];
  wire [2047:0] dataGroup_lo_677 = {dataGroup_lo_hi_677, dataGroup_lo_lo_677};
  wire [2047:0] dataGroup_hi_677 = {dataGroup_hi_hi_677, dataGroup_hi_lo_677};
  wire [7:0]    dataGroup_37_10 = dataGroup_lo_677[1487:1480];
  wire [2047:0] dataGroup_lo_678 = {dataGroup_lo_hi_678, dataGroup_lo_lo_678};
  wire [2047:0] dataGroup_hi_678 = {dataGroup_hi_hi_678, dataGroup_hi_lo_678};
  wire [7:0]    dataGroup_38_10 = dataGroup_lo_678[1527:1520];
  wire [2047:0] dataGroup_lo_679 = {dataGroup_lo_hi_679, dataGroup_lo_lo_679};
  wire [2047:0] dataGroup_hi_679 = {dataGroup_hi_hi_679, dataGroup_hi_lo_679};
  wire [7:0]    dataGroup_39_10 = dataGroup_lo_679[1567:1560];
  wire [2047:0] dataGroup_lo_680 = {dataGroup_lo_hi_680, dataGroup_lo_lo_680};
  wire [2047:0] dataGroup_hi_680 = {dataGroup_hi_hi_680, dataGroup_hi_lo_680};
  wire [7:0]    dataGroup_40_10 = dataGroup_lo_680[1607:1600];
  wire [2047:0] dataGroup_lo_681 = {dataGroup_lo_hi_681, dataGroup_lo_lo_681};
  wire [2047:0] dataGroup_hi_681 = {dataGroup_hi_hi_681, dataGroup_hi_lo_681};
  wire [7:0]    dataGroup_41_10 = dataGroup_lo_681[1647:1640];
  wire [2047:0] dataGroup_lo_682 = {dataGroup_lo_hi_682, dataGroup_lo_lo_682};
  wire [2047:0] dataGroup_hi_682 = {dataGroup_hi_hi_682, dataGroup_hi_lo_682};
  wire [7:0]    dataGroup_42_10 = dataGroup_lo_682[1687:1680];
  wire [2047:0] dataGroup_lo_683 = {dataGroup_lo_hi_683, dataGroup_lo_lo_683};
  wire [2047:0] dataGroup_hi_683 = {dataGroup_hi_hi_683, dataGroup_hi_lo_683};
  wire [7:0]    dataGroup_43_10 = dataGroup_lo_683[1727:1720];
  wire [2047:0] dataGroup_lo_684 = {dataGroup_lo_hi_684, dataGroup_lo_lo_684};
  wire [2047:0] dataGroup_hi_684 = {dataGroup_hi_hi_684, dataGroup_hi_lo_684};
  wire [7:0]    dataGroup_44_10 = dataGroup_lo_684[1767:1760];
  wire [2047:0] dataGroup_lo_685 = {dataGroup_lo_hi_685, dataGroup_lo_lo_685};
  wire [2047:0] dataGroup_hi_685 = {dataGroup_hi_hi_685, dataGroup_hi_lo_685};
  wire [7:0]    dataGroup_45_10 = dataGroup_lo_685[1807:1800];
  wire [2047:0] dataGroup_lo_686 = {dataGroup_lo_hi_686, dataGroup_lo_lo_686};
  wire [2047:0] dataGroup_hi_686 = {dataGroup_hi_hi_686, dataGroup_hi_lo_686};
  wire [7:0]    dataGroup_46_10 = dataGroup_lo_686[1847:1840];
  wire [2047:0] dataGroup_lo_687 = {dataGroup_lo_hi_687, dataGroup_lo_lo_687};
  wire [2047:0] dataGroup_hi_687 = {dataGroup_hi_hi_687, dataGroup_hi_lo_687};
  wire [7:0]    dataGroup_47_10 = dataGroup_lo_687[1887:1880];
  wire [2047:0] dataGroup_lo_688 = {dataGroup_lo_hi_688, dataGroup_lo_lo_688};
  wire [2047:0] dataGroup_hi_688 = {dataGroup_hi_hi_688, dataGroup_hi_lo_688};
  wire [7:0]    dataGroup_48_10 = dataGroup_lo_688[1927:1920];
  wire [2047:0] dataGroup_lo_689 = {dataGroup_lo_hi_689, dataGroup_lo_lo_689};
  wire [2047:0] dataGroup_hi_689 = {dataGroup_hi_hi_689, dataGroup_hi_lo_689};
  wire [7:0]    dataGroup_49_10 = dataGroup_lo_689[1967:1960];
  wire [2047:0] dataGroup_lo_690 = {dataGroup_lo_hi_690, dataGroup_lo_lo_690};
  wire [2047:0] dataGroup_hi_690 = {dataGroup_hi_hi_690, dataGroup_hi_lo_690};
  wire [7:0]    dataGroup_50_10 = dataGroup_lo_690[2007:2000];
  wire [2047:0] dataGroup_lo_691 = {dataGroup_lo_hi_691, dataGroup_lo_lo_691};
  wire [2047:0] dataGroup_hi_691 = {dataGroup_hi_hi_691, dataGroup_hi_lo_691};
  wire [7:0]    dataGroup_51_10 = dataGroup_lo_691[2047:2040];
  wire [2047:0] dataGroup_lo_692 = {dataGroup_lo_hi_692, dataGroup_lo_lo_692};
  wire [2047:0] dataGroup_hi_692 = {dataGroup_hi_hi_692, dataGroup_hi_lo_692};
  wire [7:0]    dataGroup_52_10 = dataGroup_hi_692[39:32];
  wire [2047:0] dataGroup_lo_693 = {dataGroup_lo_hi_693, dataGroup_lo_lo_693};
  wire [2047:0] dataGroup_hi_693 = {dataGroup_hi_hi_693, dataGroup_hi_lo_693};
  wire [7:0]    dataGroup_53_10 = dataGroup_hi_693[79:72];
  wire [2047:0] dataGroup_lo_694 = {dataGroup_lo_hi_694, dataGroup_lo_lo_694};
  wire [2047:0] dataGroup_hi_694 = {dataGroup_hi_hi_694, dataGroup_hi_lo_694};
  wire [7:0]    dataGroup_54_10 = dataGroup_hi_694[119:112];
  wire [2047:0] dataGroup_lo_695 = {dataGroup_lo_hi_695, dataGroup_lo_lo_695};
  wire [2047:0] dataGroup_hi_695 = {dataGroup_hi_hi_695, dataGroup_hi_lo_695};
  wire [7:0]    dataGroup_55_10 = dataGroup_hi_695[159:152];
  wire [2047:0] dataGroup_lo_696 = {dataGroup_lo_hi_696, dataGroup_lo_lo_696};
  wire [2047:0] dataGroup_hi_696 = {dataGroup_hi_hi_696, dataGroup_hi_lo_696};
  wire [7:0]    dataGroup_56_10 = dataGroup_hi_696[199:192];
  wire [2047:0] dataGroup_lo_697 = {dataGroup_lo_hi_697, dataGroup_lo_lo_697};
  wire [2047:0] dataGroup_hi_697 = {dataGroup_hi_hi_697, dataGroup_hi_lo_697};
  wire [7:0]    dataGroup_57_10 = dataGroup_hi_697[239:232];
  wire [2047:0] dataGroup_lo_698 = {dataGroup_lo_hi_698, dataGroup_lo_lo_698};
  wire [2047:0] dataGroup_hi_698 = {dataGroup_hi_hi_698, dataGroup_hi_lo_698};
  wire [7:0]    dataGroup_58_10 = dataGroup_hi_698[279:272];
  wire [2047:0] dataGroup_lo_699 = {dataGroup_lo_hi_699, dataGroup_lo_lo_699};
  wire [2047:0] dataGroup_hi_699 = {dataGroup_hi_hi_699, dataGroup_hi_lo_699};
  wire [7:0]    dataGroup_59_10 = dataGroup_hi_699[319:312];
  wire [2047:0] dataGroup_lo_700 = {dataGroup_lo_hi_700, dataGroup_lo_lo_700};
  wire [2047:0] dataGroup_hi_700 = {dataGroup_hi_hi_700, dataGroup_hi_lo_700};
  wire [7:0]    dataGroup_60_10 = dataGroup_hi_700[359:352];
  wire [2047:0] dataGroup_lo_701 = {dataGroup_lo_hi_701, dataGroup_lo_lo_701};
  wire [2047:0] dataGroup_hi_701 = {dataGroup_hi_hi_701, dataGroup_hi_lo_701};
  wire [7:0]    dataGroup_61_10 = dataGroup_hi_701[399:392];
  wire [2047:0] dataGroup_lo_702 = {dataGroup_lo_hi_702, dataGroup_lo_lo_702};
  wire [2047:0] dataGroup_hi_702 = {dataGroup_hi_hi_702, dataGroup_hi_lo_702};
  wire [7:0]    dataGroup_62_10 = dataGroup_hi_702[439:432];
  wire [2047:0] dataGroup_lo_703 = {dataGroup_lo_hi_703, dataGroup_lo_lo_703};
  wire [2047:0] dataGroup_hi_703 = {dataGroup_hi_hi_703, dataGroup_hi_lo_703};
  wire [7:0]    dataGroup_63_10 = dataGroup_hi_703[479:472];
  wire [15:0]   res_lo_lo_lo_lo_lo_10 = {dataGroup_1_10, dataGroup_0_10};
  wire [15:0]   res_lo_lo_lo_lo_hi_10 = {dataGroup_3_10, dataGroup_2_10};
  wire [31:0]   res_lo_lo_lo_lo_10 = {res_lo_lo_lo_lo_hi_10, res_lo_lo_lo_lo_lo_10};
  wire [15:0]   res_lo_lo_lo_hi_lo_10 = {dataGroup_5_10, dataGroup_4_10};
  wire [15:0]   res_lo_lo_lo_hi_hi_10 = {dataGroup_7_10, dataGroup_6_10};
  wire [31:0]   res_lo_lo_lo_hi_10 = {res_lo_lo_lo_hi_hi_10, res_lo_lo_lo_hi_lo_10};
  wire [63:0]   res_lo_lo_lo_10 = {res_lo_lo_lo_hi_10, res_lo_lo_lo_lo_10};
  wire [15:0]   res_lo_lo_hi_lo_lo_10 = {dataGroup_9_10, dataGroup_8_10};
  wire [15:0]   res_lo_lo_hi_lo_hi_10 = {dataGroup_11_10, dataGroup_10_10};
  wire [31:0]   res_lo_lo_hi_lo_10 = {res_lo_lo_hi_lo_hi_10, res_lo_lo_hi_lo_lo_10};
  wire [15:0]   res_lo_lo_hi_hi_lo_10 = {dataGroup_13_10, dataGroup_12_10};
  wire [15:0]   res_lo_lo_hi_hi_hi_10 = {dataGroup_15_10, dataGroup_14_10};
  wire [31:0]   res_lo_lo_hi_hi_10 = {res_lo_lo_hi_hi_hi_10, res_lo_lo_hi_hi_lo_10};
  wire [63:0]   res_lo_lo_hi_10 = {res_lo_lo_hi_hi_10, res_lo_lo_hi_lo_10};
  wire [127:0]  res_lo_lo_10 = {res_lo_lo_hi_10, res_lo_lo_lo_10};
  wire [15:0]   res_lo_hi_lo_lo_lo_10 = {dataGroup_17_10, dataGroup_16_10};
  wire [15:0]   res_lo_hi_lo_lo_hi_10 = {dataGroup_19_10, dataGroup_18_10};
  wire [31:0]   res_lo_hi_lo_lo_10 = {res_lo_hi_lo_lo_hi_10, res_lo_hi_lo_lo_lo_10};
  wire [15:0]   res_lo_hi_lo_hi_lo_10 = {dataGroup_21_10, dataGroup_20_10};
  wire [15:0]   res_lo_hi_lo_hi_hi_10 = {dataGroup_23_10, dataGroup_22_10};
  wire [31:0]   res_lo_hi_lo_hi_10 = {res_lo_hi_lo_hi_hi_10, res_lo_hi_lo_hi_lo_10};
  wire [63:0]   res_lo_hi_lo_10 = {res_lo_hi_lo_hi_10, res_lo_hi_lo_lo_10};
  wire [15:0]   res_lo_hi_hi_lo_lo_10 = {dataGroup_25_10, dataGroup_24_10};
  wire [15:0]   res_lo_hi_hi_lo_hi_10 = {dataGroup_27_10, dataGroup_26_10};
  wire [31:0]   res_lo_hi_hi_lo_10 = {res_lo_hi_hi_lo_hi_10, res_lo_hi_hi_lo_lo_10};
  wire [15:0]   res_lo_hi_hi_hi_lo_10 = {dataGroup_29_10, dataGroup_28_10};
  wire [15:0]   res_lo_hi_hi_hi_hi_10 = {dataGroup_31_10, dataGroup_30_10};
  wire [31:0]   res_lo_hi_hi_hi_10 = {res_lo_hi_hi_hi_hi_10, res_lo_hi_hi_hi_lo_10};
  wire [63:0]   res_lo_hi_hi_10 = {res_lo_hi_hi_hi_10, res_lo_hi_hi_lo_10};
  wire [127:0]  res_lo_hi_10 = {res_lo_hi_hi_10, res_lo_hi_lo_10};
  wire [255:0]  res_lo_10 = {res_lo_hi_10, res_lo_lo_10};
  wire [15:0]   res_hi_lo_lo_lo_lo_10 = {dataGroup_33_10, dataGroup_32_10};
  wire [15:0]   res_hi_lo_lo_lo_hi_10 = {dataGroup_35_10, dataGroup_34_10};
  wire [31:0]   res_hi_lo_lo_lo_10 = {res_hi_lo_lo_lo_hi_10, res_hi_lo_lo_lo_lo_10};
  wire [15:0]   res_hi_lo_lo_hi_lo_10 = {dataGroup_37_10, dataGroup_36_10};
  wire [15:0]   res_hi_lo_lo_hi_hi_10 = {dataGroup_39_10, dataGroup_38_10};
  wire [31:0]   res_hi_lo_lo_hi_10 = {res_hi_lo_lo_hi_hi_10, res_hi_lo_lo_hi_lo_10};
  wire [63:0]   res_hi_lo_lo_10 = {res_hi_lo_lo_hi_10, res_hi_lo_lo_lo_10};
  wire [15:0]   res_hi_lo_hi_lo_lo_10 = {dataGroup_41_10, dataGroup_40_10};
  wire [15:0]   res_hi_lo_hi_lo_hi_10 = {dataGroup_43_10, dataGroup_42_10};
  wire [31:0]   res_hi_lo_hi_lo_10 = {res_hi_lo_hi_lo_hi_10, res_hi_lo_hi_lo_lo_10};
  wire [15:0]   res_hi_lo_hi_hi_lo_10 = {dataGroup_45_10, dataGroup_44_10};
  wire [15:0]   res_hi_lo_hi_hi_hi_10 = {dataGroup_47_10, dataGroup_46_10};
  wire [31:0]   res_hi_lo_hi_hi_10 = {res_hi_lo_hi_hi_hi_10, res_hi_lo_hi_hi_lo_10};
  wire [63:0]   res_hi_lo_hi_10 = {res_hi_lo_hi_hi_10, res_hi_lo_hi_lo_10};
  wire [127:0]  res_hi_lo_10 = {res_hi_lo_hi_10, res_hi_lo_lo_10};
  wire [15:0]   res_hi_hi_lo_lo_lo_10 = {dataGroup_49_10, dataGroup_48_10};
  wire [15:0]   res_hi_hi_lo_lo_hi_10 = {dataGroup_51_10, dataGroup_50_10};
  wire [31:0]   res_hi_hi_lo_lo_10 = {res_hi_hi_lo_lo_hi_10, res_hi_hi_lo_lo_lo_10};
  wire [15:0]   res_hi_hi_lo_hi_lo_10 = {dataGroup_53_10, dataGroup_52_10};
  wire [15:0]   res_hi_hi_lo_hi_hi_10 = {dataGroup_55_10, dataGroup_54_10};
  wire [31:0]   res_hi_hi_lo_hi_10 = {res_hi_hi_lo_hi_hi_10, res_hi_hi_lo_hi_lo_10};
  wire [63:0]   res_hi_hi_lo_10 = {res_hi_hi_lo_hi_10, res_hi_hi_lo_lo_10};
  wire [15:0]   res_hi_hi_hi_lo_lo_10 = {dataGroup_57_10, dataGroup_56_10};
  wire [15:0]   res_hi_hi_hi_lo_hi_10 = {dataGroup_59_10, dataGroup_58_10};
  wire [31:0]   res_hi_hi_hi_lo_10 = {res_hi_hi_hi_lo_hi_10, res_hi_hi_hi_lo_lo_10};
  wire [15:0]   res_hi_hi_hi_hi_lo_10 = {dataGroup_61_10, dataGroup_60_10};
  wire [15:0]   res_hi_hi_hi_hi_hi_10 = {dataGroup_63_10, dataGroup_62_10};
  wire [31:0]   res_hi_hi_hi_hi_10 = {res_hi_hi_hi_hi_hi_10, res_hi_hi_hi_hi_lo_10};
  wire [63:0]   res_hi_hi_hi_10 = {res_hi_hi_hi_hi_10, res_hi_hi_hi_lo_10};
  wire [127:0]  res_hi_hi_10 = {res_hi_hi_hi_10, res_hi_hi_lo_10};
  wire [255:0]  res_hi_10 = {res_hi_hi_10, res_hi_lo_10};
  wire [511:0]  res_32 = {res_hi_10, res_lo_10};
  wire [2047:0] dataGroup_lo_704 = {dataGroup_lo_hi_704, dataGroup_lo_lo_704};
  wire [2047:0] dataGroup_hi_704 = {dataGroup_hi_hi_704, dataGroup_hi_lo_704};
  wire [7:0]    dataGroup_0_11 = dataGroup_lo_704[15:8];
  wire [2047:0] dataGroup_lo_705 = {dataGroup_lo_hi_705, dataGroup_lo_lo_705};
  wire [2047:0] dataGroup_hi_705 = {dataGroup_hi_hi_705, dataGroup_hi_lo_705};
  wire [7:0]    dataGroup_1_11 = dataGroup_lo_705[55:48];
  wire [2047:0] dataGroup_lo_706 = {dataGroup_lo_hi_706, dataGroup_lo_lo_706};
  wire [2047:0] dataGroup_hi_706 = {dataGroup_hi_hi_706, dataGroup_hi_lo_706};
  wire [7:0]    dataGroup_2_11 = dataGroup_lo_706[95:88];
  wire [2047:0] dataGroup_lo_707 = {dataGroup_lo_hi_707, dataGroup_lo_lo_707};
  wire [2047:0] dataGroup_hi_707 = {dataGroup_hi_hi_707, dataGroup_hi_lo_707};
  wire [7:0]    dataGroup_3_11 = dataGroup_lo_707[135:128];
  wire [2047:0] dataGroup_lo_708 = {dataGroup_lo_hi_708, dataGroup_lo_lo_708};
  wire [2047:0] dataGroup_hi_708 = {dataGroup_hi_hi_708, dataGroup_hi_lo_708};
  wire [7:0]    dataGroup_4_11 = dataGroup_lo_708[175:168];
  wire [2047:0] dataGroup_lo_709 = {dataGroup_lo_hi_709, dataGroup_lo_lo_709};
  wire [2047:0] dataGroup_hi_709 = {dataGroup_hi_hi_709, dataGroup_hi_lo_709};
  wire [7:0]    dataGroup_5_11 = dataGroup_lo_709[215:208];
  wire [2047:0] dataGroup_lo_710 = {dataGroup_lo_hi_710, dataGroup_lo_lo_710};
  wire [2047:0] dataGroup_hi_710 = {dataGroup_hi_hi_710, dataGroup_hi_lo_710};
  wire [7:0]    dataGroup_6_11 = dataGroup_lo_710[255:248];
  wire [2047:0] dataGroup_lo_711 = {dataGroup_lo_hi_711, dataGroup_lo_lo_711};
  wire [2047:0] dataGroup_hi_711 = {dataGroup_hi_hi_711, dataGroup_hi_lo_711};
  wire [7:0]    dataGroup_7_11 = dataGroup_lo_711[295:288];
  wire [2047:0] dataGroup_lo_712 = {dataGroup_lo_hi_712, dataGroup_lo_lo_712};
  wire [2047:0] dataGroup_hi_712 = {dataGroup_hi_hi_712, dataGroup_hi_lo_712};
  wire [7:0]    dataGroup_8_11 = dataGroup_lo_712[335:328];
  wire [2047:0] dataGroup_lo_713 = {dataGroup_lo_hi_713, dataGroup_lo_lo_713};
  wire [2047:0] dataGroup_hi_713 = {dataGroup_hi_hi_713, dataGroup_hi_lo_713};
  wire [7:0]    dataGroup_9_11 = dataGroup_lo_713[375:368];
  wire [2047:0] dataGroup_lo_714 = {dataGroup_lo_hi_714, dataGroup_lo_lo_714};
  wire [2047:0] dataGroup_hi_714 = {dataGroup_hi_hi_714, dataGroup_hi_lo_714};
  wire [7:0]    dataGroup_10_11 = dataGroup_lo_714[415:408];
  wire [2047:0] dataGroup_lo_715 = {dataGroup_lo_hi_715, dataGroup_lo_lo_715};
  wire [2047:0] dataGroup_hi_715 = {dataGroup_hi_hi_715, dataGroup_hi_lo_715};
  wire [7:0]    dataGroup_11_11 = dataGroup_lo_715[455:448];
  wire [2047:0] dataGroup_lo_716 = {dataGroup_lo_hi_716, dataGroup_lo_lo_716};
  wire [2047:0] dataGroup_hi_716 = {dataGroup_hi_hi_716, dataGroup_hi_lo_716};
  wire [7:0]    dataGroup_12_11 = dataGroup_lo_716[495:488];
  wire [2047:0] dataGroup_lo_717 = {dataGroup_lo_hi_717, dataGroup_lo_lo_717};
  wire [2047:0] dataGroup_hi_717 = {dataGroup_hi_hi_717, dataGroup_hi_lo_717};
  wire [7:0]    dataGroup_13_11 = dataGroup_lo_717[535:528];
  wire [2047:0] dataGroup_lo_718 = {dataGroup_lo_hi_718, dataGroup_lo_lo_718};
  wire [2047:0] dataGroup_hi_718 = {dataGroup_hi_hi_718, dataGroup_hi_lo_718};
  wire [7:0]    dataGroup_14_11 = dataGroup_lo_718[575:568];
  wire [2047:0] dataGroup_lo_719 = {dataGroup_lo_hi_719, dataGroup_lo_lo_719};
  wire [2047:0] dataGroup_hi_719 = {dataGroup_hi_hi_719, dataGroup_hi_lo_719};
  wire [7:0]    dataGroup_15_11 = dataGroup_lo_719[615:608];
  wire [2047:0] dataGroup_lo_720 = {dataGroup_lo_hi_720, dataGroup_lo_lo_720};
  wire [2047:0] dataGroup_hi_720 = {dataGroup_hi_hi_720, dataGroup_hi_lo_720};
  wire [7:0]    dataGroup_16_11 = dataGroup_lo_720[655:648];
  wire [2047:0] dataGroup_lo_721 = {dataGroup_lo_hi_721, dataGroup_lo_lo_721};
  wire [2047:0] dataGroup_hi_721 = {dataGroup_hi_hi_721, dataGroup_hi_lo_721};
  wire [7:0]    dataGroup_17_11 = dataGroup_lo_721[695:688];
  wire [2047:0] dataGroup_lo_722 = {dataGroup_lo_hi_722, dataGroup_lo_lo_722};
  wire [2047:0] dataGroup_hi_722 = {dataGroup_hi_hi_722, dataGroup_hi_lo_722};
  wire [7:0]    dataGroup_18_11 = dataGroup_lo_722[735:728];
  wire [2047:0] dataGroup_lo_723 = {dataGroup_lo_hi_723, dataGroup_lo_lo_723};
  wire [2047:0] dataGroup_hi_723 = {dataGroup_hi_hi_723, dataGroup_hi_lo_723};
  wire [7:0]    dataGroup_19_11 = dataGroup_lo_723[775:768];
  wire [2047:0] dataGroup_lo_724 = {dataGroup_lo_hi_724, dataGroup_lo_lo_724};
  wire [2047:0] dataGroup_hi_724 = {dataGroup_hi_hi_724, dataGroup_hi_lo_724};
  wire [7:0]    dataGroup_20_11 = dataGroup_lo_724[815:808];
  wire [2047:0] dataGroup_lo_725 = {dataGroup_lo_hi_725, dataGroup_lo_lo_725};
  wire [2047:0] dataGroup_hi_725 = {dataGroup_hi_hi_725, dataGroup_hi_lo_725};
  wire [7:0]    dataGroup_21_11 = dataGroup_lo_725[855:848];
  wire [2047:0] dataGroup_lo_726 = {dataGroup_lo_hi_726, dataGroup_lo_lo_726};
  wire [2047:0] dataGroup_hi_726 = {dataGroup_hi_hi_726, dataGroup_hi_lo_726};
  wire [7:0]    dataGroup_22_11 = dataGroup_lo_726[895:888];
  wire [2047:0] dataGroup_lo_727 = {dataGroup_lo_hi_727, dataGroup_lo_lo_727};
  wire [2047:0] dataGroup_hi_727 = {dataGroup_hi_hi_727, dataGroup_hi_lo_727};
  wire [7:0]    dataGroup_23_11 = dataGroup_lo_727[935:928];
  wire [2047:0] dataGroup_lo_728 = {dataGroup_lo_hi_728, dataGroup_lo_lo_728};
  wire [2047:0] dataGroup_hi_728 = {dataGroup_hi_hi_728, dataGroup_hi_lo_728};
  wire [7:0]    dataGroup_24_11 = dataGroup_lo_728[975:968];
  wire [2047:0] dataGroup_lo_729 = {dataGroup_lo_hi_729, dataGroup_lo_lo_729};
  wire [2047:0] dataGroup_hi_729 = {dataGroup_hi_hi_729, dataGroup_hi_lo_729};
  wire [7:0]    dataGroup_25_11 = dataGroup_lo_729[1015:1008];
  wire [2047:0] dataGroup_lo_730 = {dataGroup_lo_hi_730, dataGroup_lo_lo_730};
  wire [2047:0] dataGroup_hi_730 = {dataGroup_hi_hi_730, dataGroup_hi_lo_730};
  wire [7:0]    dataGroup_26_11 = dataGroup_lo_730[1055:1048];
  wire [2047:0] dataGroup_lo_731 = {dataGroup_lo_hi_731, dataGroup_lo_lo_731};
  wire [2047:0] dataGroup_hi_731 = {dataGroup_hi_hi_731, dataGroup_hi_lo_731};
  wire [7:0]    dataGroup_27_11 = dataGroup_lo_731[1095:1088];
  wire [2047:0] dataGroup_lo_732 = {dataGroup_lo_hi_732, dataGroup_lo_lo_732};
  wire [2047:0] dataGroup_hi_732 = {dataGroup_hi_hi_732, dataGroup_hi_lo_732};
  wire [7:0]    dataGroup_28_11 = dataGroup_lo_732[1135:1128];
  wire [2047:0] dataGroup_lo_733 = {dataGroup_lo_hi_733, dataGroup_lo_lo_733};
  wire [2047:0] dataGroup_hi_733 = {dataGroup_hi_hi_733, dataGroup_hi_lo_733};
  wire [7:0]    dataGroup_29_11 = dataGroup_lo_733[1175:1168];
  wire [2047:0] dataGroup_lo_734 = {dataGroup_lo_hi_734, dataGroup_lo_lo_734};
  wire [2047:0] dataGroup_hi_734 = {dataGroup_hi_hi_734, dataGroup_hi_lo_734};
  wire [7:0]    dataGroup_30_11 = dataGroup_lo_734[1215:1208];
  wire [2047:0] dataGroup_lo_735 = {dataGroup_lo_hi_735, dataGroup_lo_lo_735};
  wire [2047:0] dataGroup_hi_735 = {dataGroup_hi_hi_735, dataGroup_hi_lo_735};
  wire [7:0]    dataGroup_31_11 = dataGroup_lo_735[1255:1248];
  wire [2047:0] dataGroup_lo_736 = {dataGroup_lo_hi_736, dataGroup_lo_lo_736};
  wire [2047:0] dataGroup_hi_736 = {dataGroup_hi_hi_736, dataGroup_hi_lo_736};
  wire [7:0]    dataGroup_32_11 = dataGroup_lo_736[1295:1288];
  wire [2047:0] dataGroup_lo_737 = {dataGroup_lo_hi_737, dataGroup_lo_lo_737};
  wire [2047:0] dataGroup_hi_737 = {dataGroup_hi_hi_737, dataGroup_hi_lo_737};
  wire [7:0]    dataGroup_33_11 = dataGroup_lo_737[1335:1328];
  wire [2047:0] dataGroup_lo_738 = {dataGroup_lo_hi_738, dataGroup_lo_lo_738};
  wire [2047:0] dataGroup_hi_738 = {dataGroup_hi_hi_738, dataGroup_hi_lo_738};
  wire [7:0]    dataGroup_34_11 = dataGroup_lo_738[1375:1368];
  wire [2047:0] dataGroup_lo_739 = {dataGroup_lo_hi_739, dataGroup_lo_lo_739};
  wire [2047:0] dataGroup_hi_739 = {dataGroup_hi_hi_739, dataGroup_hi_lo_739};
  wire [7:0]    dataGroup_35_11 = dataGroup_lo_739[1415:1408];
  wire [2047:0] dataGroup_lo_740 = {dataGroup_lo_hi_740, dataGroup_lo_lo_740};
  wire [2047:0] dataGroup_hi_740 = {dataGroup_hi_hi_740, dataGroup_hi_lo_740};
  wire [7:0]    dataGroup_36_11 = dataGroup_lo_740[1455:1448];
  wire [2047:0] dataGroup_lo_741 = {dataGroup_lo_hi_741, dataGroup_lo_lo_741};
  wire [2047:0] dataGroup_hi_741 = {dataGroup_hi_hi_741, dataGroup_hi_lo_741};
  wire [7:0]    dataGroup_37_11 = dataGroup_lo_741[1495:1488];
  wire [2047:0] dataGroup_lo_742 = {dataGroup_lo_hi_742, dataGroup_lo_lo_742};
  wire [2047:0] dataGroup_hi_742 = {dataGroup_hi_hi_742, dataGroup_hi_lo_742};
  wire [7:0]    dataGroup_38_11 = dataGroup_lo_742[1535:1528];
  wire [2047:0] dataGroup_lo_743 = {dataGroup_lo_hi_743, dataGroup_lo_lo_743};
  wire [2047:0] dataGroup_hi_743 = {dataGroup_hi_hi_743, dataGroup_hi_lo_743};
  wire [7:0]    dataGroup_39_11 = dataGroup_lo_743[1575:1568];
  wire [2047:0] dataGroup_lo_744 = {dataGroup_lo_hi_744, dataGroup_lo_lo_744};
  wire [2047:0] dataGroup_hi_744 = {dataGroup_hi_hi_744, dataGroup_hi_lo_744};
  wire [7:0]    dataGroup_40_11 = dataGroup_lo_744[1615:1608];
  wire [2047:0] dataGroup_lo_745 = {dataGroup_lo_hi_745, dataGroup_lo_lo_745};
  wire [2047:0] dataGroup_hi_745 = {dataGroup_hi_hi_745, dataGroup_hi_lo_745};
  wire [7:0]    dataGroup_41_11 = dataGroup_lo_745[1655:1648];
  wire [2047:0] dataGroup_lo_746 = {dataGroup_lo_hi_746, dataGroup_lo_lo_746};
  wire [2047:0] dataGroup_hi_746 = {dataGroup_hi_hi_746, dataGroup_hi_lo_746};
  wire [7:0]    dataGroup_42_11 = dataGroup_lo_746[1695:1688];
  wire [2047:0] dataGroup_lo_747 = {dataGroup_lo_hi_747, dataGroup_lo_lo_747};
  wire [2047:0] dataGroup_hi_747 = {dataGroup_hi_hi_747, dataGroup_hi_lo_747};
  wire [7:0]    dataGroup_43_11 = dataGroup_lo_747[1735:1728];
  wire [2047:0] dataGroup_lo_748 = {dataGroup_lo_hi_748, dataGroup_lo_lo_748};
  wire [2047:0] dataGroup_hi_748 = {dataGroup_hi_hi_748, dataGroup_hi_lo_748};
  wire [7:0]    dataGroup_44_11 = dataGroup_lo_748[1775:1768];
  wire [2047:0] dataGroup_lo_749 = {dataGroup_lo_hi_749, dataGroup_lo_lo_749};
  wire [2047:0] dataGroup_hi_749 = {dataGroup_hi_hi_749, dataGroup_hi_lo_749};
  wire [7:0]    dataGroup_45_11 = dataGroup_lo_749[1815:1808];
  wire [2047:0] dataGroup_lo_750 = {dataGroup_lo_hi_750, dataGroup_lo_lo_750};
  wire [2047:0] dataGroup_hi_750 = {dataGroup_hi_hi_750, dataGroup_hi_lo_750};
  wire [7:0]    dataGroup_46_11 = dataGroup_lo_750[1855:1848];
  wire [2047:0] dataGroup_lo_751 = {dataGroup_lo_hi_751, dataGroup_lo_lo_751};
  wire [2047:0] dataGroup_hi_751 = {dataGroup_hi_hi_751, dataGroup_hi_lo_751};
  wire [7:0]    dataGroup_47_11 = dataGroup_lo_751[1895:1888];
  wire [2047:0] dataGroup_lo_752 = {dataGroup_lo_hi_752, dataGroup_lo_lo_752};
  wire [2047:0] dataGroup_hi_752 = {dataGroup_hi_hi_752, dataGroup_hi_lo_752};
  wire [7:0]    dataGroup_48_11 = dataGroup_lo_752[1935:1928];
  wire [2047:0] dataGroup_lo_753 = {dataGroup_lo_hi_753, dataGroup_lo_lo_753};
  wire [2047:0] dataGroup_hi_753 = {dataGroup_hi_hi_753, dataGroup_hi_lo_753};
  wire [7:0]    dataGroup_49_11 = dataGroup_lo_753[1975:1968];
  wire [2047:0] dataGroup_lo_754 = {dataGroup_lo_hi_754, dataGroup_lo_lo_754};
  wire [2047:0] dataGroup_hi_754 = {dataGroup_hi_hi_754, dataGroup_hi_lo_754};
  wire [7:0]    dataGroup_50_11 = dataGroup_lo_754[2015:2008];
  wire [2047:0] dataGroup_lo_755 = {dataGroup_lo_hi_755, dataGroup_lo_lo_755};
  wire [2047:0] dataGroup_hi_755 = {dataGroup_hi_hi_755, dataGroup_hi_lo_755};
  wire [7:0]    dataGroup_51_11 = dataGroup_hi_755[7:0];
  wire [2047:0] dataGroup_lo_756 = {dataGroup_lo_hi_756, dataGroup_lo_lo_756};
  wire [2047:0] dataGroup_hi_756 = {dataGroup_hi_hi_756, dataGroup_hi_lo_756};
  wire [7:0]    dataGroup_52_11 = dataGroup_hi_756[47:40];
  wire [2047:0] dataGroup_lo_757 = {dataGroup_lo_hi_757, dataGroup_lo_lo_757};
  wire [2047:0] dataGroup_hi_757 = {dataGroup_hi_hi_757, dataGroup_hi_lo_757};
  wire [7:0]    dataGroup_53_11 = dataGroup_hi_757[87:80];
  wire [2047:0] dataGroup_lo_758 = {dataGroup_lo_hi_758, dataGroup_lo_lo_758};
  wire [2047:0] dataGroup_hi_758 = {dataGroup_hi_hi_758, dataGroup_hi_lo_758};
  wire [7:0]    dataGroup_54_11 = dataGroup_hi_758[127:120];
  wire [2047:0] dataGroup_lo_759 = {dataGroup_lo_hi_759, dataGroup_lo_lo_759};
  wire [2047:0] dataGroup_hi_759 = {dataGroup_hi_hi_759, dataGroup_hi_lo_759};
  wire [7:0]    dataGroup_55_11 = dataGroup_hi_759[167:160];
  wire [2047:0] dataGroup_lo_760 = {dataGroup_lo_hi_760, dataGroup_lo_lo_760};
  wire [2047:0] dataGroup_hi_760 = {dataGroup_hi_hi_760, dataGroup_hi_lo_760};
  wire [7:0]    dataGroup_56_11 = dataGroup_hi_760[207:200];
  wire [2047:0] dataGroup_lo_761 = {dataGroup_lo_hi_761, dataGroup_lo_lo_761};
  wire [2047:0] dataGroup_hi_761 = {dataGroup_hi_hi_761, dataGroup_hi_lo_761};
  wire [7:0]    dataGroup_57_11 = dataGroup_hi_761[247:240];
  wire [2047:0] dataGroup_lo_762 = {dataGroup_lo_hi_762, dataGroup_lo_lo_762};
  wire [2047:0] dataGroup_hi_762 = {dataGroup_hi_hi_762, dataGroup_hi_lo_762};
  wire [7:0]    dataGroup_58_11 = dataGroup_hi_762[287:280];
  wire [2047:0] dataGroup_lo_763 = {dataGroup_lo_hi_763, dataGroup_lo_lo_763};
  wire [2047:0] dataGroup_hi_763 = {dataGroup_hi_hi_763, dataGroup_hi_lo_763};
  wire [7:0]    dataGroup_59_11 = dataGroup_hi_763[327:320];
  wire [2047:0] dataGroup_lo_764 = {dataGroup_lo_hi_764, dataGroup_lo_lo_764};
  wire [2047:0] dataGroup_hi_764 = {dataGroup_hi_hi_764, dataGroup_hi_lo_764};
  wire [7:0]    dataGroup_60_11 = dataGroup_hi_764[367:360];
  wire [2047:0] dataGroup_lo_765 = {dataGroup_lo_hi_765, dataGroup_lo_lo_765};
  wire [2047:0] dataGroup_hi_765 = {dataGroup_hi_hi_765, dataGroup_hi_lo_765};
  wire [7:0]    dataGroup_61_11 = dataGroup_hi_765[407:400];
  wire [2047:0] dataGroup_lo_766 = {dataGroup_lo_hi_766, dataGroup_lo_lo_766};
  wire [2047:0] dataGroup_hi_766 = {dataGroup_hi_hi_766, dataGroup_hi_lo_766};
  wire [7:0]    dataGroup_62_11 = dataGroup_hi_766[447:440];
  wire [2047:0] dataGroup_lo_767 = {dataGroup_lo_hi_767, dataGroup_lo_lo_767};
  wire [2047:0] dataGroup_hi_767 = {dataGroup_hi_hi_767, dataGroup_hi_lo_767};
  wire [7:0]    dataGroup_63_11 = dataGroup_hi_767[487:480];
  wire [15:0]   res_lo_lo_lo_lo_lo_11 = {dataGroup_1_11, dataGroup_0_11};
  wire [15:0]   res_lo_lo_lo_lo_hi_11 = {dataGroup_3_11, dataGroup_2_11};
  wire [31:0]   res_lo_lo_lo_lo_11 = {res_lo_lo_lo_lo_hi_11, res_lo_lo_lo_lo_lo_11};
  wire [15:0]   res_lo_lo_lo_hi_lo_11 = {dataGroup_5_11, dataGroup_4_11};
  wire [15:0]   res_lo_lo_lo_hi_hi_11 = {dataGroup_7_11, dataGroup_6_11};
  wire [31:0]   res_lo_lo_lo_hi_11 = {res_lo_lo_lo_hi_hi_11, res_lo_lo_lo_hi_lo_11};
  wire [63:0]   res_lo_lo_lo_11 = {res_lo_lo_lo_hi_11, res_lo_lo_lo_lo_11};
  wire [15:0]   res_lo_lo_hi_lo_lo_11 = {dataGroup_9_11, dataGroup_8_11};
  wire [15:0]   res_lo_lo_hi_lo_hi_11 = {dataGroup_11_11, dataGroup_10_11};
  wire [31:0]   res_lo_lo_hi_lo_11 = {res_lo_lo_hi_lo_hi_11, res_lo_lo_hi_lo_lo_11};
  wire [15:0]   res_lo_lo_hi_hi_lo_11 = {dataGroup_13_11, dataGroup_12_11};
  wire [15:0]   res_lo_lo_hi_hi_hi_11 = {dataGroup_15_11, dataGroup_14_11};
  wire [31:0]   res_lo_lo_hi_hi_11 = {res_lo_lo_hi_hi_hi_11, res_lo_lo_hi_hi_lo_11};
  wire [63:0]   res_lo_lo_hi_11 = {res_lo_lo_hi_hi_11, res_lo_lo_hi_lo_11};
  wire [127:0]  res_lo_lo_11 = {res_lo_lo_hi_11, res_lo_lo_lo_11};
  wire [15:0]   res_lo_hi_lo_lo_lo_11 = {dataGroup_17_11, dataGroup_16_11};
  wire [15:0]   res_lo_hi_lo_lo_hi_11 = {dataGroup_19_11, dataGroup_18_11};
  wire [31:0]   res_lo_hi_lo_lo_11 = {res_lo_hi_lo_lo_hi_11, res_lo_hi_lo_lo_lo_11};
  wire [15:0]   res_lo_hi_lo_hi_lo_11 = {dataGroup_21_11, dataGroup_20_11};
  wire [15:0]   res_lo_hi_lo_hi_hi_11 = {dataGroup_23_11, dataGroup_22_11};
  wire [31:0]   res_lo_hi_lo_hi_11 = {res_lo_hi_lo_hi_hi_11, res_lo_hi_lo_hi_lo_11};
  wire [63:0]   res_lo_hi_lo_11 = {res_lo_hi_lo_hi_11, res_lo_hi_lo_lo_11};
  wire [15:0]   res_lo_hi_hi_lo_lo_11 = {dataGroup_25_11, dataGroup_24_11};
  wire [15:0]   res_lo_hi_hi_lo_hi_11 = {dataGroup_27_11, dataGroup_26_11};
  wire [31:0]   res_lo_hi_hi_lo_11 = {res_lo_hi_hi_lo_hi_11, res_lo_hi_hi_lo_lo_11};
  wire [15:0]   res_lo_hi_hi_hi_lo_11 = {dataGroup_29_11, dataGroup_28_11};
  wire [15:0]   res_lo_hi_hi_hi_hi_11 = {dataGroup_31_11, dataGroup_30_11};
  wire [31:0]   res_lo_hi_hi_hi_11 = {res_lo_hi_hi_hi_hi_11, res_lo_hi_hi_hi_lo_11};
  wire [63:0]   res_lo_hi_hi_11 = {res_lo_hi_hi_hi_11, res_lo_hi_hi_lo_11};
  wire [127:0]  res_lo_hi_11 = {res_lo_hi_hi_11, res_lo_hi_lo_11};
  wire [255:0]  res_lo_11 = {res_lo_hi_11, res_lo_lo_11};
  wire [15:0]   res_hi_lo_lo_lo_lo_11 = {dataGroup_33_11, dataGroup_32_11};
  wire [15:0]   res_hi_lo_lo_lo_hi_11 = {dataGroup_35_11, dataGroup_34_11};
  wire [31:0]   res_hi_lo_lo_lo_11 = {res_hi_lo_lo_lo_hi_11, res_hi_lo_lo_lo_lo_11};
  wire [15:0]   res_hi_lo_lo_hi_lo_11 = {dataGroup_37_11, dataGroup_36_11};
  wire [15:0]   res_hi_lo_lo_hi_hi_11 = {dataGroup_39_11, dataGroup_38_11};
  wire [31:0]   res_hi_lo_lo_hi_11 = {res_hi_lo_lo_hi_hi_11, res_hi_lo_lo_hi_lo_11};
  wire [63:0]   res_hi_lo_lo_11 = {res_hi_lo_lo_hi_11, res_hi_lo_lo_lo_11};
  wire [15:0]   res_hi_lo_hi_lo_lo_11 = {dataGroup_41_11, dataGroup_40_11};
  wire [15:0]   res_hi_lo_hi_lo_hi_11 = {dataGroup_43_11, dataGroup_42_11};
  wire [31:0]   res_hi_lo_hi_lo_11 = {res_hi_lo_hi_lo_hi_11, res_hi_lo_hi_lo_lo_11};
  wire [15:0]   res_hi_lo_hi_hi_lo_11 = {dataGroup_45_11, dataGroup_44_11};
  wire [15:0]   res_hi_lo_hi_hi_hi_11 = {dataGroup_47_11, dataGroup_46_11};
  wire [31:0]   res_hi_lo_hi_hi_11 = {res_hi_lo_hi_hi_hi_11, res_hi_lo_hi_hi_lo_11};
  wire [63:0]   res_hi_lo_hi_11 = {res_hi_lo_hi_hi_11, res_hi_lo_hi_lo_11};
  wire [127:0]  res_hi_lo_11 = {res_hi_lo_hi_11, res_hi_lo_lo_11};
  wire [15:0]   res_hi_hi_lo_lo_lo_11 = {dataGroup_49_11, dataGroup_48_11};
  wire [15:0]   res_hi_hi_lo_lo_hi_11 = {dataGroup_51_11, dataGroup_50_11};
  wire [31:0]   res_hi_hi_lo_lo_11 = {res_hi_hi_lo_lo_hi_11, res_hi_hi_lo_lo_lo_11};
  wire [15:0]   res_hi_hi_lo_hi_lo_11 = {dataGroup_53_11, dataGroup_52_11};
  wire [15:0]   res_hi_hi_lo_hi_hi_11 = {dataGroup_55_11, dataGroup_54_11};
  wire [31:0]   res_hi_hi_lo_hi_11 = {res_hi_hi_lo_hi_hi_11, res_hi_hi_lo_hi_lo_11};
  wire [63:0]   res_hi_hi_lo_11 = {res_hi_hi_lo_hi_11, res_hi_hi_lo_lo_11};
  wire [15:0]   res_hi_hi_hi_lo_lo_11 = {dataGroup_57_11, dataGroup_56_11};
  wire [15:0]   res_hi_hi_hi_lo_hi_11 = {dataGroup_59_11, dataGroup_58_11};
  wire [31:0]   res_hi_hi_hi_lo_11 = {res_hi_hi_hi_lo_hi_11, res_hi_hi_hi_lo_lo_11};
  wire [15:0]   res_hi_hi_hi_hi_lo_11 = {dataGroup_61_11, dataGroup_60_11};
  wire [15:0]   res_hi_hi_hi_hi_hi_11 = {dataGroup_63_11, dataGroup_62_11};
  wire [31:0]   res_hi_hi_hi_hi_11 = {res_hi_hi_hi_hi_hi_11, res_hi_hi_hi_hi_lo_11};
  wire [63:0]   res_hi_hi_hi_11 = {res_hi_hi_hi_hi_11, res_hi_hi_hi_lo_11};
  wire [127:0]  res_hi_hi_11 = {res_hi_hi_hi_11, res_hi_hi_lo_11};
  wire [255:0]  res_hi_11 = {res_hi_hi_11, res_hi_lo_11};
  wire [511:0]  res_33 = {res_hi_11, res_lo_11};
  wire [2047:0] dataGroup_lo_768 = {dataGroup_lo_hi_768, dataGroup_lo_lo_768};
  wire [2047:0] dataGroup_hi_768 = {dataGroup_hi_hi_768, dataGroup_hi_lo_768};
  wire [7:0]    dataGroup_0_12 = dataGroup_lo_768[23:16];
  wire [2047:0] dataGroup_lo_769 = {dataGroup_lo_hi_769, dataGroup_lo_lo_769};
  wire [2047:0] dataGroup_hi_769 = {dataGroup_hi_hi_769, dataGroup_hi_lo_769};
  wire [7:0]    dataGroup_1_12 = dataGroup_lo_769[63:56];
  wire [2047:0] dataGroup_lo_770 = {dataGroup_lo_hi_770, dataGroup_lo_lo_770};
  wire [2047:0] dataGroup_hi_770 = {dataGroup_hi_hi_770, dataGroup_hi_lo_770};
  wire [7:0]    dataGroup_2_12 = dataGroup_lo_770[103:96];
  wire [2047:0] dataGroup_lo_771 = {dataGroup_lo_hi_771, dataGroup_lo_lo_771};
  wire [2047:0] dataGroup_hi_771 = {dataGroup_hi_hi_771, dataGroup_hi_lo_771};
  wire [7:0]    dataGroup_3_12 = dataGroup_lo_771[143:136];
  wire [2047:0] dataGroup_lo_772 = {dataGroup_lo_hi_772, dataGroup_lo_lo_772};
  wire [2047:0] dataGroup_hi_772 = {dataGroup_hi_hi_772, dataGroup_hi_lo_772};
  wire [7:0]    dataGroup_4_12 = dataGroup_lo_772[183:176];
  wire [2047:0] dataGroup_lo_773 = {dataGroup_lo_hi_773, dataGroup_lo_lo_773};
  wire [2047:0] dataGroup_hi_773 = {dataGroup_hi_hi_773, dataGroup_hi_lo_773};
  wire [7:0]    dataGroup_5_12 = dataGroup_lo_773[223:216];
  wire [2047:0] dataGroup_lo_774 = {dataGroup_lo_hi_774, dataGroup_lo_lo_774};
  wire [2047:0] dataGroup_hi_774 = {dataGroup_hi_hi_774, dataGroup_hi_lo_774};
  wire [7:0]    dataGroup_6_12 = dataGroup_lo_774[263:256];
  wire [2047:0] dataGroup_lo_775 = {dataGroup_lo_hi_775, dataGroup_lo_lo_775};
  wire [2047:0] dataGroup_hi_775 = {dataGroup_hi_hi_775, dataGroup_hi_lo_775};
  wire [7:0]    dataGroup_7_12 = dataGroup_lo_775[303:296];
  wire [2047:0] dataGroup_lo_776 = {dataGroup_lo_hi_776, dataGroup_lo_lo_776};
  wire [2047:0] dataGroup_hi_776 = {dataGroup_hi_hi_776, dataGroup_hi_lo_776};
  wire [7:0]    dataGroup_8_12 = dataGroup_lo_776[343:336];
  wire [2047:0] dataGroup_lo_777 = {dataGroup_lo_hi_777, dataGroup_lo_lo_777};
  wire [2047:0] dataGroup_hi_777 = {dataGroup_hi_hi_777, dataGroup_hi_lo_777};
  wire [7:0]    dataGroup_9_12 = dataGroup_lo_777[383:376];
  wire [2047:0] dataGroup_lo_778 = {dataGroup_lo_hi_778, dataGroup_lo_lo_778};
  wire [2047:0] dataGroup_hi_778 = {dataGroup_hi_hi_778, dataGroup_hi_lo_778};
  wire [7:0]    dataGroup_10_12 = dataGroup_lo_778[423:416];
  wire [2047:0] dataGroup_lo_779 = {dataGroup_lo_hi_779, dataGroup_lo_lo_779};
  wire [2047:0] dataGroup_hi_779 = {dataGroup_hi_hi_779, dataGroup_hi_lo_779};
  wire [7:0]    dataGroup_11_12 = dataGroup_lo_779[463:456];
  wire [2047:0] dataGroup_lo_780 = {dataGroup_lo_hi_780, dataGroup_lo_lo_780};
  wire [2047:0] dataGroup_hi_780 = {dataGroup_hi_hi_780, dataGroup_hi_lo_780};
  wire [7:0]    dataGroup_12_12 = dataGroup_lo_780[503:496];
  wire [2047:0] dataGroup_lo_781 = {dataGroup_lo_hi_781, dataGroup_lo_lo_781};
  wire [2047:0] dataGroup_hi_781 = {dataGroup_hi_hi_781, dataGroup_hi_lo_781};
  wire [7:0]    dataGroup_13_12 = dataGroup_lo_781[543:536];
  wire [2047:0] dataGroup_lo_782 = {dataGroup_lo_hi_782, dataGroup_lo_lo_782};
  wire [2047:0] dataGroup_hi_782 = {dataGroup_hi_hi_782, dataGroup_hi_lo_782};
  wire [7:0]    dataGroup_14_12 = dataGroup_lo_782[583:576];
  wire [2047:0] dataGroup_lo_783 = {dataGroup_lo_hi_783, dataGroup_lo_lo_783};
  wire [2047:0] dataGroup_hi_783 = {dataGroup_hi_hi_783, dataGroup_hi_lo_783};
  wire [7:0]    dataGroup_15_12 = dataGroup_lo_783[623:616];
  wire [2047:0] dataGroup_lo_784 = {dataGroup_lo_hi_784, dataGroup_lo_lo_784};
  wire [2047:0] dataGroup_hi_784 = {dataGroup_hi_hi_784, dataGroup_hi_lo_784};
  wire [7:0]    dataGroup_16_12 = dataGroup_lo_784[663:656];
  wire [2047:0] dataGroup_lo_785 = {dataGroup_lo_hi_785, dataGroup_lo_lo_785};
  wire [2047:0] dataGroup_hi_785 = {dataGroup_hi_hi_785, dataGroup_hi_lo_785};
  wire [7:0]    dataGroup_17_12 = dataGroup_lo_785[703:696];
  wire [2047:0] dataGroup_lo_786 = {dataGroup_lo_hi_786, dataGroup_lo_lo_786};
  wire [2047:0] dataGroup_hi_786 = {dataGroup_hi_hi_786, dataGroup_hi_lo_786};
  wire [7:0]    dataGroup_18_12 = dataGroup_lo_786[743:736];
  wire [2047:0] dataGroup_lo_787 = {dataGroup_lo_hi_787, dataGroup_lo_lo_787};
  wire [2047:0] dataGroup_hi_787 = {dataGroup_hi_hi_787, dataGroup_hi_lo_787};
  wire [7:0]    dataGroup_19_12 = dataGroup_lo_787[783:776];
  wire [2047:0] dataGroup_lo_788 = {dataGroup_lo_hi_788, dataGroup_lo_lo_788};
  wire [2047:0] dataGroup_hi_788 = {dataGroup_hi_hi_788, dataGroup_hi_lo_788};
  wire [7:0]    dataGroup_20_12 = dataGroup_lo_788[823:816];
  wire [2047:0] dataGroup_lo_789 = {dataGroup_lo_hi_789, dataGroup_lo_lo_789};
  wire [2047:0] dataGroup_hi_789 = {dataGroup_hi_hi_789, dataGroup_hi_lo_789};
  wire [7:0]    dataGroup_21_12 = dataGroup_lo_789[863:856];
  wire [2047:0] dataGroup_lo_790 = {dataGroup_lo_hi_790, dataGroup_lo_lo_790};
  wire [2047:0] dataGroup_hi_790 = {dataGroup_hi_hi_790, dataGroup_hi_lo_790};
  wire [7:0]    dataGroup_22_12 = dataGroup_lo_790[903:896];
  wire [2047:0] dataGroup_lo_791 = {dataGroup_lo_hi_791, dataGroup_lo_lo_791};
  wire [2047:0] dataGroup_hi_791 = {dataGroup_hi_hi_791, dataGroup_hi_lo_791};
  wire [7:0]    dataGroup_23_12 = dataGroup_lo_791[943:936];
  wire [2047:0] dataGroup_lo_792 = {dataGroup_lo_hi_792, dataGroup_lo_lo_792};
  wire [2047:0] dataGroup_hi_792 = {dataGroup_hi_hi_792, dataGroup_hi_lo_792};
  wire [7:0]    dataGroup_24_12 = dataGroup_lo_792[983:976];
  wire [2047:0] dataGroup_lo_793 = {dataGroup_lo_hi_793, dataGroup_lo_lo_793};
  wire [2047:0] dataGroup_hi_793 = {dataGroup_hi_hi_793, dataGroup_hi_lo_793};
  wire [7:0]    dataGroup_25_12 = dataGroup_lo_793[1023:1016];
  wire [2047:0] dataGroup_lo_794 = {dataGroup_lo_hi_794, dataGroup_lo_lo_794};
  wire [2047:0] dataGroup_hi_794 = {dataGroup_hi_hi_794, dataGroup_hi_lo_794};
  wire [7:0]    dataGroup_26_12 = dataGroup_lo_794[1063:1056];
  wire [2047:0] dataGroup_lo_795 = {dataGroup_lo_hi_795, dataGroup_lo_lo_795};
  wire [2047:0] dataGroup_hi_795 = {dataGroup_hi_hi_795, dataGroup_hi_lo_795};
  wire [7:0]    dataGroup_27_12 = dataGroup_lo_795[1103:1096];
  wire [2047:0] dataGroup_lo_796 = {dataGroup_lo_hi_796, dataGroup_lo_lo_796};
  wire [2047:0] dataGroup_hi_796 = {dataGroup_hi_hi_796, dataGroup_hi_lo_796};
  wire [7:0]    dataGroup_28_12 = dataGroup_lo_796[1143:1136];
  wire [2047:0] dataGroup_lo_797 = {dataGroup_lo_hi_797, dataGroup_lo_lo_797};
  wire [2047:0] dataGroup_hi_797 = {dataGroup_hi_hi_797, dataGroup_hi_lo_797};
  wire [7:0]    dataGroup_29_12 = dataGroup_lo_797[1183:1176];
  wire [2047:0] dataGroup_lo_798 = {dataGroup_lo_hi_798, dataGroup_lo_lo_798};
  wire [2047:0] dataGroup_hi_798 = {dataGroup_hi_hi_798, dataGroup_hi_lo_798};
  wire [7:0]    dataGroup_30_12 = dataGroup_lo_798[1223:1216];
  wire [2047:0] dataGroup_lo_799 = {dataGroup_lo_hi_799, dataGroup_lo_lo_799};
  wire [2047:0] dataGroup_hi_799 = {dataGroup_hi_hi_799, dataGroup_hi_lo_799};
  wire [7:0]    dataGroup_31_12 = dataGroup_lo_799[1263:1256];
  wire [2047:0] dataGroup_lo_800 = {dataGroup_lo_hi_800, dataGroup_lo_lo_800};
  wire [2047:0] dataGroup_hi_800 = {dataGroup_hi_hi_800, dataGroup_hi_lo_800};
  wire [7:0]    dataGroup_32_12 = dataGroup_lo_800[1303:1296];
  wire [2047:0] dataGroup_lo_801 = {dataGroup_lo_hi_801, dataGroup_lo_lo_801};
  wire [2047:0] dataGroup_hi_801 = {dataGroup_hi_hi_801, dataGroup_hi_lo_801};
  wire [7:0]    dataGroup_33_12 = dataGroup_lo_801[1343:1336];
  wire [2047:0] dataGroup_lo_802 = {dataGroup_lo_hi_802, dataGroup_lo_lo_802};
  wire [2047:0] dataGroup_hi_802 = {dataGroup_hi_hi_802, dataGroup_hi_lo_802};
  wire [7:0]    dataGroup_34_12 = dataGroup_lo_802[1383:1376];
  wire [2047:0] dataGroup_lo_803 = {dataGroup_lo_hi_803, dataGroup_lo_lo_803};
  wire [2047:0] dataGroup_hi_803 = {dataGroup_hi_hi_803, dataGroup_hi_lo_803};
  wire [7:0]    dataGroup_35_12 = dataGroup_lo_803[1423:1416];
  wire [2047:0] dataGroup_lo_804 = {dataGroup_lo_hi_804, dataGroup_lo_lo_804};
  wire [2047:0] dataGroup_hi_804 = {dataGroup_hi_hi_804, dataGroup_hi_lo_804};
  wire [7:0]    dataGroup_36_12 = dataGroup_lo_804[1463:1456];
  wire [2047:0] dataGroup_lo_805 = {dataGroup_lo_hi_805, dataGroup_lo_lo_805};
  wire [2047:0] dataGroup_hi_805 = {dataGroup_hi_hi_805, dataGroup_hi_lo_805};
  wire [7:0]    dataGroup_37_12 = dataGroup_lo_805[1503:1496];
  wire [2047:0] dataGroup_lo_806 = {dataGroup_lo_hi_806, dataGroup_lo_lo_806};
  wire [2047:0] dataGroup_hi_806 = {dataGroup_hi_hi_806, dataGroup_hi_lo_806};
  wire [7:0]    dataGroup_38_12 = dataGroup_lo_806[1543:1536];
  wire [2047:0] dataGroup_lo_807 = {dataGroup_lo_hi_807, dataGroup_lo_lo_807};
  wire [2047:0] dataGroup_hi_807 = {dataGroup_hi_hi_807, dataGroup_hi_lo_807};
  wire [7:0]    dataGroup_39_12 = dataGroup_lo_807[1583:1576];
  wire [2047:0] dataGroup_lo_808 = {dataGroup_lo_hi_808, dataGroup_lo_lo_808};
  wire [2047:0] dataGroup_hi_808 = {dataGroup_hi_hi_808, dataGroup_hi_lo_808};
  wire [7:0]    dataGroup_40_12 = dataGroup_lo_808[1623:1616];
  wire [2047:0] dataGroup_lo_809 = {dataGroup_lo_hi_809, dataGroup_lo_lo_809};
  wire [2047:0] dataGroup_hi_809 = {dataGroup_hi_hi_809, dataGroup_hi_lo_809};
  wire [7:0]    dataGroup_41_12 = dataGroup_lo_809[1663:1656];
  wire [2047:0] dataGroup_lo_810 = {dataGroup_lo_hi_810, dataGroup_lo_lo_810};
  wire [2047:0] dataGroup_hi_810 = {dataGroup_hi_hi_810, dataGroup_hi_lo_810};
  wire [7:0]    dataGroup_42_12 = dataGroup_lo_810[1703:1696];
  wire [2047:0] dataGroup_lo_811 = {dataGroup_lo_hi_811, dataGroup_lo_lo_811};
  wire [2047:0] dataGroup_hi_811 = {dataGroup_hi_hi_811, dataGroup_hi_lo_811};
  wire [7:0]    dataGroup_43_12 = dataGroup_lo_811[1743:1736];
  wire [2047:0] dataGroup_lo_812 = {dataGroup_lo_hi_812, dataGroup_lo_lo_812};
  wire [2047:0] dataGroup_hi_812 = {dataGroup_hi_hi_812, dataGroup_hi_lo_812};
  wire [7:0]    dataGroup_44_12 = dataGroup_lo_812[1783:1776];
  wire [2047:0] dataGroup_lo_813 = {dataGroup_lo_hi_813, dataGroup_lo_lo_813};
  wire [2047:0] dataGroup_hi_813 = {dataGroup_hi_hi_813, dataGroup_hi_lo_813};
  wire [7:0]    dataGroup_45_12 = dataGroup_lo_813[1823:1816];
  wire [2047:0] dataGroup_lo_814 = {dataGroup_lo_hi_814, dataGroup_lo_lo_814};
  wire [2047:0] dataGroup_hi_814 = {dataGroup_hi_hi_814, dataGroup_hi_lo_814};
  wire [7:0]    dataGroup_46_12 = dataGroup_lo_814[1863:1856];
  wire [2047:0] dataGroup_lo_815 = {dataGroup_lo_hi_815, dataGroup_lo_lo_815};
  wire [2047:0] dataGroup_hi_815 = {dataGroup_hi_hi_815, dataGroup_hi_lo_815};
  wire [7:0]    dataGroup_47_12 = dataGroup_lo_815[1903:1896];
  wire [2047:0] dataGroup_lo_816 = {dataGroup_lo_hi_816, dataGroup_lo_lo_816};
  wire [2047:0] dataGroup_hi_816 = {dataGroup_hi_hi_816, dataGroup_hi_lo_816};
  wire [7:0]    dataGroup_48_12 = dataGroup_lo_816[1943:1936];
  wire [2047:0] dataGroup_lo_817 = {dataGroup_lo_hi_817, dataGroup_lo_lo_817};
  wire [2047:0] dataGroup_hi_817 = {dataGroup_hi_hi_817, dataGroup_hi_lo_817};
  wire [7:0]    dataGroup_49_12 = dataGroup_lo_817[1983:1976];
  wire [2047:0] dataGroup_lo_818 = {dataGroup_lo_hi_818, dataGroup_lo_lo_818};
  wire [2047:0] dataGroup_hi_818 = {dataGroup_hi_hi_818, dataGroup_hi_lo_818};
  wire [7:0]    dataGroup_50_12 = dataGroup_lo_818[2023:2016];
  wire [2047:0] dataGroup_lo_819 = {dataGroup_lo_hi_819, dataGroup_lo_lo_819};
  wire [2047:0] dataGroup_hi_819 = {dataGroup_hi_hi_819, dataGroup_hi_lo_819};
  wire [7:0]    dataGroup_51_12 = dataGroup_hi_819[15:8];
  wire [2047:0] dataGroup_lo_820 = {dataGroup_lo_hi_820, dataGroup_lo_lo_820};
  wire [2047:0] dataGroup_hi_820 = {dataGroup_hi_hi_820, dataGroup_hi_lo_820};
  wire [7:0]    dataGroup_52_12 = dataGroup_hi_820[55:48];
  wire [2047:0] dataGroup_lo_821 = {dataGroup_lo_hi_821, dataGroup_lo_lo_821};
  wire [2047:0] dataGroup_hi_821 = {dataGroup_hi_hi_821, dataGroup_hi_lo_821};
  wire [7:0]    dataGroup_53_12 = dataGroup_hi_821[95:88];
  wire [2047:0] dataGroup_lo_822 = {dataGroup_lo_hi_822, dataGroup_lo_lo_822};
  wire [2047:0] dataGroup_hi_822 = {dataGroup_hi_hi_822, dataGroup_hi_lo_822};
  wire [7:0]    dataGroup_54_12 = dataGroup_hi_822[135:128];
  wire [2047:0] dataGroup_lo_823 = {dataGroup_lo_hi_823, dataGroup_lo_lo_823};
  wire [2047:0] dataGroup_hi_823 = {dataGroup_hi_hi_823, dataGroup_hi_lo_823};
  wire [7:0]    dataGroup_55_12 = dataGroup_hi_823[175:168];
  wire [2047:0] dataGroup_lo_824 = {dataGroup_lo_hi_824, dataGroup_lo_lo_824};
  wire [2047:0] dataGroup_hi_824 = {dataGroup_hi_hi_824, dataGroup_hi_lo_824};
  wire [7:0]    dataGroup_56_12 = dataGroup_hi_824[215:208];
  wire [2047:0] dataGroup_lo_825 = {dataGroup_lo_hi_825, dataGroup_lo_lo_825};
  wire [2047:0] dataGroup_hi_825 = {dataGroup_hi_hi_825, dataGroup_hi_lo_825};
  wire [7:0]    dataGroup_57_12 = dataGroup_hi_825[255:248];
  wire [2047:0] dataGroup_lo_826 = {dataGroup_lo_hi_826, dataGroup_lo_lo_826};
  wire [2047:0] dataGroup_hi_826 = {dataGroup_hi_hi_826, dataGroup_hi_lo_826};
  wire [7:0]    dataGroup_58_12 = dataGroup_hi_826[295:288];
  wire [2047:0] dataGroup_lo_827 = {dataGroup_lo_hi_827, dataGroup_lo_lo_827};
  wire [2047:0] dataGroup_hi_827 = {dataGroup_hi_hi_827, dataGroup_hi_lo_827};
  wire [7:0]    dataGroup_59_12 = dataGroup_hi_827[335:328];
  wire [2047:0] dataGroup_lo_828 = {dataGroup_lo_hi_828, dataGroup_lo_lo_828};
  wire [2047:0] dataGroup_hi_828 = {dataGroup_hi_hi_828, dataGroup_hi_lo_828};
  wire [7:0]    dataGroup_60_12 = dataGroup_hi_828[375:368];
  wire [2047:0] dataGroup_lo_829 = {dataGroup_lo_hi_829, dataGroup_lo_lo_829};
  wire [2047:0] dataGroup_hi_829 = {dataGroup_hi_hi_829, dataGroup_hi_lo_829};
  wire [7:0]    dataGroup_61_12 = dataGroup_hi_829[415:408];
  wire [2047:0] dataGroup_lo_830 = {dataGroup_lo_hi_830, dataGroup_lo_lo_830};
  wire [2047:0] dataGroup_hi_830 = {dataGroup_hi_hi_830, dataGroup_hi_lo_830};
  wire [7:0]    dataGroup_62_12 = dataGroup_hi_830[455:448];
  wire [2047:0] dataGroup_lo_831 = {dataGroup_lo_hi_831, dataGroup_lo_lo_831};
  wire [2047:0] dataGroup_hi_831 = {dataGroup_hi_hi_831, dataGroup_hi_lo_831};
  wire [7:0]    dataGroup_63_12 = dataGroup_hi_831[495:488];
  wire [15:0]   res_lo_lo_lo_lo_lo_12 = {dataGroup_1_12, dataGroup_0_12};
  wire [15:0]   res_lo_lo_lo_lo_hi_12 = {dataGroup_3_12, dataGroup_2_12};
  wire [31:0]   res_lo_lo_lo_lo_12 = {res_lo_lo_lo_lo_hi_12, res_lo_lo_lo_lo_lo_12};
  wire [15:0]   res_lo_lo_lo_hi_lo_12 = {dataGroup_5_12, dataGroup_4_12};
  wire [15:0]   res_lo_lo_lo_hi_hi_12 = {dataGroup_7_12, dataGroup_6_12};
  wire [31:0]   res_lo_lo_lo_hi_12 = {res_lo_lo_lo_hi_hi_12, res_lo_lo_lo_hi_lo_12};
  wire [63:0]   res_lo_lo_lo_12 = {res_lo_lo_lo_hi_12, res_lo_lo_lo_lo_12};
  wire [15:0]   res_lo_lo_hi_lo_lo_12 = {dataGroup_9_12, dataGroup_8_12};
  wire [15:0]   res_lo_lo_hi_lo_hi_12 = {dataGroup_11_12, dataGroup_10_12};
  wire [31:0]   res_lo_lo_hi_lo_12 = {res_lo_lo_hi_lo_hi_12, res_lo_lo_hi_lo_lo_12};
  wire [15:0]   res_lo_lo_hi_hi_lo_12 = {dataGroup_13_12, dataGroup_12_12};
  wire [15:0]   res_lo_lo_hi_hi_hi_12 = {dataGroup_15_12, dataGroup_14_12};
  wire [31:0]   res_lo_lo_hi_hi_12 = {res_lo_lo_hi_hi_hi_12, res_lo_lo_hi_hi_lo_12};
  wire [63:0]   res_lo_lo_hi_12 = {res_lo_lo_hi_hi_12, res_lo_lo_hi_lo_12};
  wire [127:0]  res_lo_lo_12 = {res_lo_lo_hi_12, res_lo_lo_lo_12};
  wire [15:0]   res_lo_hi_lo_lo_lo_12 = {dataGroup_17_12, dataGroup_16_12};
  wire [15:0]   res_lo_hi_lo_lo_hi_12 = {dataGroup_19_12, dataGroup_18_12};
  wire [31:0]   res_lo_hi_lo_lo_12 = {res_lo_hi_lo_lo_hi_12, res_lo_hi_lo_lo_lo_12};
  wire [15:0]   res_lo_hi_lo_hi_lo_12 = {dataGroup_21_12, dataGroup_20_12};
  wire [15:0]   res_lo_hi_lo_hi_hi_12 = {dataGroup_23_12, dataGroup_22_12};
  wire [31:0]   res_lo_hi_lo_hi_12 = {res_lo_hi_lo_hi_hi_12, res_lo_hi_lo_hi_lo_12};
  wire [63:0]   res_lo_hi_lo_12 = {res_lo_hi_lo_hi_12, res_lo_hi_lo_lo_12};
  wire [15:0]   res_lo_hi_hi_lo_lo_12 = {dataGroup_25_12, dataGroup_24_12};
  wire [15:0]   res_lo_hi_hi_lo_hi_12 = {dataGroup_27_12, dataGroup_26_12};
  wire [31:0]   res_lo_hi_hi_lo_12 = {res_lo_hi_hi_lo_hi_12, res_lo_hi_hi_lo_lo_12};
  wire [15:0]   res_lo_hi_hi_hi_lo_12 = {dataGroup_29_12, dataGroup_28_12};
  wire [15:0]   res_lo_hi_hi_hi_hi_12 = {dataGroup_31_12, dataGroup_30_12};
  wire [31:0]   res_lo_hi_hi_hi_12 = {res_lo_hi_hi_hi_hi_12, res_lo_hi_hi_hi_lo_12};
  wire [63:0]   res_lo_hi_hi_12 = {res_lo_hi_hi_hi_12, res_lo_hi_hi_lo_12};
  wire [127:0]  res_lo_hi_12 = {res_lo_hi_hi_12, res_lo_hi_lo_12};
  wire [255:0]  res_lo_12 = {res_lo_hi_12, res_lo_lo_12};
  wire [15:0]   res_hi_lo_lo_lo_lo_12 = {dataGroup_33_12, dataGroup_32_12};
  wire [15:0]   res_hi_lo_lo_lo_hi_12 = {dataGroup_35_12, dataGroup_34_12};
  wire [31:0]   res_hi_lo_lo_lo_12 = {res_hi_lo_lo_lo_hi_12, res_hi_lo_lo_lo_lo_12};
  wire [15:0]   res_hi_lo_lo_hi_lo_12 = {dataGroup_37_12, dataGroup_36_12};
  wire [15:0]   res_hi_lo_lo_hi_hi_12 = {dataGroup_39_12, dataGroup_38_12};
  wire [31:0]   res_hi_lo_lo_hi_12 = {res_hi_lo_lo_hi_hi_12, res_hi_lo_lo_hi_lo_12};
  wire [63:0]   res_hi_lo_lo_12 = {res_hi_lo_lo_hi_12, res_hi_lo_lo_lo_12};
  wire [15:0]   res_hi_lo_hi_lo_lo_12 = {dataGroup_41_12, dataGroup_40_12};
  wire [15:0]   res_hi_lo_hi_lo_hi_12 = {dataGroup_43_12, dataGroup_42_12};
  wire [31:0]   res_hi_lo_hi_lo_12 = {res_hi_lo_hi_lo_hi_12, res_hi_lo_hi_lo_lo_12};
  wire [15:0]   res_hi_lo_hi_hi_lo_12 = {dataGroup_45_12, dataGroup_44_12};
  wire [15:0]   res_hi_lo_hi_hi_hi_12 = {dataGroup_47_12, dataGroup_46_12};
  wire [31:0]   res_hi_lo_hi_hi_12 = {res_hi_lo_hi_hi_hi_12, res_hi_lo_hi_hi_lo_12};
  wire [63:0]   res_hi_lo_hi_12 = {res_hi_lo_hi_hi_12, res_hi_lo_hi_lo_12};
  wire [127:0]  res_hi_lo_12 = {res_hi_lo_hi_12, res_hi_lo_lo_12};
  wire [15:0]   res_hi_hi_lo_lo_lo_12 = {dataGroup_49_12, dataGroup_48_12};
  wire [15:0]   res_hi_hi_lo_lo_hi_12 = {dataGroup_51_12, dataGroup_50_12};
  wire [31:0]   res_hi_hi_lo_lo_12 = {res_hi_hi_lo_lo_hi_12, res_hi_hi_lo_lo_lo_12};
  wire [15:0]   res_hi_hi_lo_hi_lo_12 = {dataGroup_53_12, dataGroup_52_12};
  wire [15:0]   res_hi_hi_lo_hi_hi_12 = {dataGroup_55_12, dataGroup_54_12};
  wire [31:0]   res_hi_hi_lo_hi_12 = {res_hi_hi_lo_hi_hi_12, res_hi_hi_lo_hi_lo_12};
  wire [63:0]   res_hi_hi_lo_12 = {res_hi_hi_lo_hi_12, res_hi_hi_lo_lo_12};
  wire [15:0]   res_hi_hi_hi_lo_lo_12 = {dataGroup_57_12, dataGroup_56_12};
  wire [15:0]   res_hi_hi_hi_lo_hi_12 = {dataGroup_59_12, dataGroup_58_12};
  wire [31:0]   res_hi_hi_hi_lo_12 = {res_hi_hi_hi_lo_hi_12, res_hi_hi_hi_lo_lo_12};
  wire [15:0]   res_hi_hi_hi_hi_lo_12 = {dataGroup_61_12, dataGroup_60_12};
  wire [15:0]   res_hi_hi_hi_hi_hi_12 = {dataGroup_63_12, dataGroup_62_12};
  wire [31:0]   res_hi_hi_hi_hi_12 = {res_hi_hi_hi_hi_hi_12, res_hi_hi_hi_hi_lo_12};
  wire [63:0]   res_hi_hi_hi_12 = {res_hi_hi_hi_hi_12, res_hi_hi_hi_lo_12};
  wire [127:0]  res_hi_hi_12 = {res_hi_hi_hi_12, res_hi_hi_lo_12};
  wire [255:0]  res_hi_12 = {res_hi_hi_12, res_hi_lo_12};
  wire [511:0]  res_34 = {res_hi_12, res_lo_12};
  wire [2047:0] dataGroup_lo_832 = {dataGroup_lo_hi_832, dataGroup_lo_lo_832};
  wire [2047:0] dataGroup_hi_832 = {dataGroup_hi_hi_832, dataGroup_hi_lo_832};
  wire [7:0]    dataGroup_0_13 = dataGroup_lo_832[31:24];
  wire [2047:0] dataGroup_lo_833 = {dataGroup_lo_hi_833, dataGroup_lo_lo_833};
  wire [2047:0] dataGroup_hi_833 = {dataGroup_hi_hi_833, dataGroup_hi_lo_833};
  wire [7:0]    dataGroup_1_13 = dataGroup_lo_833[71:64];
  wire [2047:0] dataGroup_lo_834 = {dataGroup_lo_hi_834, dataGroup_lo_lo_834};
  wire [2047:0] dataGroup_hi_834 = {dataGroup_hi_hi_834, dataGroup_hi_lo_834};
  wire [7:0]    dataGroup_2_13 = dataGroup_lo_834[111:104];
  wire [2047:0] dataGroup_lo_835 = {dataGroup_lo_hi_835, dataGroup_lo_lo_835};
  wire [2047:0] dataGroup_hi_835 = {dataGroup_hi_hi_835, dataGroup_hi_lo_835};
  wire [7:0]    dataGroup_3_13 = dataGroup_lo_835[151:144];
  wire [2047:0] dataGroup_lo_836 = {dataGroup_lo_hi_836, dataGroup_lo_lo_836};
  wire [2047:0] dataGroup_hi_836 = {dataGroup_hi_hi_836, dataGroup_hi_lo_836};
  wire [7:0]    dataGroup_4_13 = dataGroup_lo_836[191:184];
  wire [2047:0] dataGroup_lo_837 = {dataGroup_lo_hi_837, dataGroup_lo_lo_837};
  wire [2047:0] dataGroup_hi_837 = {dataGroup_hi_hi_837, dataGroup_hi_lo_837};
  wire [7:0]    dataGroup_5_13 = dataGroup_lo_837[231:224];
  wire [2047:0] dataGroup_lo_838 = {dataGroup_lo_hi_838, dataGroup_lo_lo_838};
  wire [2047:0] dataGroup_hi_838 = {dataGroup_hi_hi_838, dataGroup_hi_lo_838};
  wire [7:0]    dataGroup_6_13 = dataGroup_lo_838[271:264];
  wire [2047:0] dataGroup_lo_839 = {dataGroup_lo_hi_839, dataGroup_lo_lo_839};
  wire [2047:0] dataGroup_hi_839 = {dataGroup_hi_hi_839, dataGroup_hi_lo_839};
  wire [7:0]    dataGroup_7_13 = dataGroup_lo_839[311:304];
  wire [2047:0] dataGroup_lo_840 = {dataGroup_lo_hi_840, dataGroup_lo_lo_840};
  wire [2047:0] dataGroup_hi_840 = {dataGroup_hi_hi_840, dataGroup_hi_lo_840};
  wire [7:0]    dataGroup_8_13 = dataGroup_lo_840[351:344];
  wire [2047:0] dataGroup_lo_841 = {dataGroup_lo_hi_841, dataGroup_lo_lo_841};
  wire [2047:0] dataGroup_hi_841 = {dataGroup_hi_hi_841, dataGroup_hi_lo_841};
  wire [7:0]    dataGroup_9_13 = dataGroup_lo_841[391:384];
  wire [2047:0] dataGroup_lo_842 = {dataGroup_lo_hi_842, dataGroup_lo_lo_842};
  wire [2047:0] dataGroup_hi_842 = {dataGroup_hi_hi_842, dataGroup_hi_lo_842};
  wire [7:0]    dataGroup_10_13 = dataGroup_lo_842[431:424];
  wire [2047:0] dataGroup_lo_843 = {dataGroup_lo_hi_843, dataGroup_lo_lo_843};
  wire [2047:0] dataGroup_hi_843 = {dataGroup_hi_hi_843, dataGroup_hi_lo_843};
  wire [7:0]    dataGroup_11_13 = dataGroup_lo_843[471:464];
  wire [2047:0] dataGroup_lo_844 = {dataGroup_lo_hi_844, dataGroup_lo_lo_844};
  wire [2047:0] dataGroup_hi_844 = {dataGroup_hi_hi_844, dataGroup_hi_lo_844};
  wire [7:0]    dataGroup_12_13 = dataGroup_lo_844[511:504];
  wire [2047:0] dataGroup_lo_845 = {dataGroup_lo_hi_845, dataGroup_lo_lo_845};
  wire [2047:0] dataGroup_hi_845 = {dataGroup_hi_hi_845, dataGroup_hi_lo_845};
  wire [7:0]    dataGroup_13_13 = dataGroup_lo_845[551:544];
  wire [2047:0] dataGroup_lo_846 = {dataGroup_lo_hi_846, dataGroup_lo_lo_846};
  wire [2047:0] dataGroup_hi_846 = {dataGroup_hi_hi_846, dataGroup_hi_lo_846};
  wire [7:0]    dataGroup_14_13 = dataGroup_lo_846[591:584];
  wire [2047:0] dataGroup_lo_847 = {dataGroup_lo_hi_847, dataGroup_lo_lo_847};
  wire [2047:0] dataGroup_hi_847 = {dataGroup_hi_hi_847, dataGroup_hi_lo_847};
  wire [7:0]    dataGroup_15_13 = dataGroup_lo_847[631:624];
  wire [2047:0] dataGroup_lo_848 = {dataGroup_lo_hi_848, dataGroup_lo_lo_848};
  wire [2047:0] dataGroup_hi_848 = {dataGroup_hi_hi_848, dataGroup_hi_lo_848};
  wire [7:0]    dataGroup_16_13 = dataGroup_lo_848[671:664];
  wire [2047:0] dataGroup_lo_849 = {dataGroup_lo_hi_849, dataGroup_lo_lo_849};
  wire [2047:0] dataGroup_hi_849 = {dataGroup_hi_hi_849, dataGroup_hi_lo_849};
  wire [7:0]    dataGroup_17_13 = dataGroup_lo_849[711:704];
  wire [2047:0] dataGroup_lo_850 = {dataGroup_lo_hi_850, dataGroup_lo_lo_850};
  wire [2047:0] dataGroup_hi_850 = {dataGroup_hi_hi_850, dataGroup_hi_lo_850};
  wire [7:0]    dataGroup_18_13 = dataGroup_lo_850[751:744];
  wire [2047:0] dataGroup_lo_851 = {dataGroup_lo_hi_851, dataGroup_lo_lo_851};
  wire [2047:0] dataGroup_hi_851 = {dataGroup_hi_hi_851, dataGroup_hi_lo_851};
  wire [7:0]    dataGroup_19_13 = dataGroup_lo_851[791:784];
  wire [2047:0] dataGroup_lo_852 = {dataGroup_lo_hi_852, dataGroup_lo_lo_852};
  wire [2047:0] dataGroup_hi_852 = {dataGroup_hi_hi_852, dataGroup_hi_lo_852};
  wire [7:0]    dataGroup_20_13 = dataGroup_lo_852[831:824];
  wire [2047:0] dataGroup_lo_853 = {dataGroup_lo_hi_853, dataGroup_lo_lo_853};
  wire [2047:0] dataGroup_hi_853 = {dataGroup_hi_hi_853, dataGroup_hi_lo_853};
  wire [7:0]    dataGroup_21_13 = dataGroup_lo_853[871:864];
  wire [2047:0] dataGroup_lo_854 = {dataGroup_lo_hi_854, dataGroup_lo_lo_854};
  wire [2047:0] dataGroup_hi_854 = {dataGroup_hi_hi_854, dataGroup_hi_lo_854};
  wire [7:0]    dataGroup_22_13 = dataGroup_lo_854[911:904];
  wire [2047:0] dataGroup_lo_855 = {dataGroup_lo_hi_855, dataGroup_lo_lo_855};
  wire [2047:0] dataGroup_hi_855 = {dataGroup_hi_hi_855, dataGroup_hi_lo_855};
  wire [7:0]    dataGroup_23_13 = dataGroup_lo_855[951:944];
  wire [2047:0] dataGroup_lo_856 = {dataGroup_lo_hi_856, dataGroup_lo_lo_856};
  wire [2047:0] dataGroup_hi_856 = {dataGroup_hi_hi_856, dataGroup_hi_lo_856};
  wire [7:0]    dataGroup_24_13 = dataGroup_lo_856[991:984];
  wire [2047:0] dataGroup_lo_857 = {dataGroup_lo_hi_857, dataGroup_lo_lo_857};
  wire [2047:0] dataGroup_hi_857 = {dataGroup_hi_hi_857, dataGroup_hi_lo_857};
  wire [7:0]    dataGroup_25_13 = dataGroup_lo_857[1031:1024];
  wire [2047:0] dataGroup_lo_858 = {dataGroup_lo_hi_858, dataGroup_lo_lo_858};
  wire [2047:0] dataGroup_hi_858 = {dataGroup_hi_hi_858, dataGroup_hi_lo_858};
  wire [7:0]    dataGroup_26_13 = dataGroup_lo_858[1071:1064];
  wire [2047:0] dataGroup_lo_859 = {dataGroup_lo_hi_859, dataGroup_lo_lo_859};
  wire [2047:0] dataGroup_hi_859 = {dataGroup_hi_hi_859, dataGroup_hi_lo_859};
  wire [7:0]    dataGroup_27_13 = dataGroup_lo_859[1111:1104];
  wire [2047:0] dataGroup_lo_860 = {dataGroup_lo_hi_860, dataGroup_lo_lo_860};
  wire [2047:0] dataGroup_hi_860 = {dataGroup_hi_hi_860, dataGroup_hi_lo_860};
  wire [7:0]    dataGroup_28_13 = dataGroup_lo_860[1151:1144];
  wire [2047:0] dataGroup_lo_861 = {dataGroup_lo_hi_861, dataGroup_lo_lo_861};
  wire [2047:0] dataGroup_hi_861 = {dataGroup_hi_hi_861, dataGroup_hi_lo_861};
  wire [7:0]    dataGroup_29_13 = dataGroup_lo_861[1191:1184];
  wire [2047:0] dataGroup_lo_862 = {dataGroup_lo_hi_862, dataGroup_lo_lo_862};
  wire [2047:0] dataGroup_hi_862 = {dataGroup_hi_hi_862, dataGroup_hi_lo_862};
  wire [7:0]    dataGroup_30_13 = dataGroup_lo_862[1231:1224];
  wire [2047:0] dataGroup_lo_863 = {dataGroup_lo_hi_863, dataGroup_lo_lo_863};
  wire [2047:0] dataGroup_hi_863 = {dataGroup_hi_hi_863, dataGroup_hi_lo_863};
  wire [7:0]    dataGroup_31_13 = dataGroup_lo_863[1271:1264];
  wire [2047:0] dataGroup_lo_864 = {dataGroup_lo_hi_864, dataGroup_lo_lo_864};
  wire [2047:0] dataGroup_hi_864 = {dataGroup_hi_hi_864, dataGroup_hi_lo_864};
  wire [7:0]    dataGroup_32_13 = dataGroup_lo_864[1311:1304];
  wire [2047:0] dataGroup_lo_865 = {dataGroup_lo_hi_865, dataGroup_lo_lo_865};
  wire [2047:0] dataGroup_hi_865 = {dataGroup_hi_hi_865, dataGroup_hi_lo_865};
  wire [7:0]    dataGroup_33_13 = dataGroup_lo_865[1351:1344];
  wire [2047:0] dataGroup_lo_866 = {dataGroup_lo_hi_866, dataGroup_lo_lo_866};
  wire [2047:0] dataGroup_hi_866 = {dataGroup_hi_hi_866, dataGroup_hi_lo_866};
  wire [7:0]    dataGroup_34_13 = dataGroup_lo_866[1391:1384];
  wire [2047:0] dataGroup_lo_867 = {dataGroup_lo_hi_867, dataGroup_lo_lo_867};
  wire [2047:0] dataGroup_hi_867 = {dataGroup_hi_hi_867, dataGroup_hi_lo_867};
  wire [7:0]    dataGroup_35_13 = dataGroup_lo_867[1431:1424];
  wire [2047:0] dataGroup_lo_868 = {dataGroup_lo_hi_868, dataGroup_lo_lo_868};
  wire [2047:0] dataGroup_hi_868 = {dataGroup_hi_hi_868, dataGroup_hi_lo_868};
  wire [7:0]    dataGroup_36_13 = dataGroup_lo_868[1471:1464];
  wire [2047:0] dataGroup_lo_869 = {dataGroup_lo_hi_869, dataGroup_lo_lo_869};
  wire [2047:0] dataGroup_hi_869 = {dataGroup_hi_hi_869, dataGroup_hi_lo_869};
  wire [7:0]    dataGroup_37_13 = dataGroup_lo_869[1511:1504];
  wire [2047:0] dataGroup_lo_870 = {dataGroup_lo_hi_870, dataGroup_lo_lo_870};
  wire [2047:0] dataGroup_hi_870 = {dataGroup_hi_hi_870, dataGroup_hi_lo_870};
  wire [7:0]    dataGroup_38_13 = dataGroup_lo_870[1551:1544];
  wire [2047:0] dataGroup_lo_871 = {dataGroup_lo_hi_871, dataGroup_lo_lo_871};
  wire [2047:0] dataGroup_hi_871 = {dataGroup_hi_hi_871, dataGroup_hi_lo_871};
  wire [7:0]    dataGroup_39_13 = dataGroup_lo_871[1591:1584];
  wire [2047:0] dataGroup_lo_872 = {dataGroup_lo_hi_872, dataGroup_lo_lo_872};
  wire [2047:0] dataGroup_hi_872 = {dataGroup_hi_hi_872, dataGroup_hi_lo_872};
  wire [7:0]    dataGroup_40_13 = dataGroup_lo_872[1631:1624];
  wire [2047:0] dataGroup_lo_873 = {dataGroup_lo_hi_873, dataGroup_lo_lo_873};
  wire [2047:0] dataGroup_hi_873 = {dataGroup_hi_hi_873, dataGroup_hi_lo_873};
  wire [7:0]    dataGroup_41_13 = dataGroup_lo_873[1671:1664];
  wire [2047:0] dataGroup_lo_874 = {dataGroup_lo_hi_874, dataGroup_lo_lo_874};
  wire [2047:0] dataGroup_hi_874 = {dataGroup_hi_hi_874, dataGroup_hi_lo_874};
  wire [7:0]    dataGroup_42_13 = dataGroup_lo_874[1711:1704];
  wire [2047:0] dataGroup_lo_875 = {dataGroup_lo_hi_875, dataGroup_lo_lo_875};
  wire [2047:0] dataGroup_hi_875 = {dataGroup_hi_hi_875, dataGroup_hi_lo_875};
  wire [7:0]    dataGroup_43_13 = dataGroup_lo_875[1751:1744];
  wire [2047:0] dataGroup_lo_876 = {dataGroup_lo_hi_876, dataGroup_lo_lo_876};
  wire [2047:0] dataGroup_hi_876 = {dataGroup_hi_hi_876, dataGroup_hi_lo_876};
  wire [7:0]    dataGroup_44_13 = dataGroup_lo_876[1791:1784];
  wire [2047:0] dataGroup_lo_877 = {dataGroup_lo_hi_877, dataGroup_lo_lo_877};
  wire [2047:0] dataGroup_hi_877 = {dataGroup_hi_hi_877, dataGroup_hi_lo_877};
  wire [7:0]    dataGroup_45_13 = dataGroup_lo_877[1831:1824];
  wire [2047:0] dataGroup_lo_878 = {dataGroup_lo_hi_878, dataGroup_lo_lo_878};
  wire [2047:0] dataGroup_hi_878 = {dataGroup_hi_hi_878, dataGroup_hi_lo_878};
  wire [7:0]    dataGroup_46_13 = dataGroup_lo_878[1871:1864];
  wire [2047:0] dataGroup_lo_879 = {dataGroup_lo_hi_879, dataGroup_lo_lo_879};
  wire [2047:0] dataGroup_hi_879 = {dataGroup_hi_hi_879, dataGroup_hi_lo_879};
  wire [7:0]    dataGroup_47_13 = dataGroup_lo_879[1911:1904];
  wire [2047:0] dataGroup_lo_880 = {dataGroup_lo_hi_880, dataGroup_lo_lo_880};
  wire [2047:0] dataGroup_hi_880 = {dataGroup_hi_hi_880, dataGroup_hi_lo_880};
  wire [7:0]    dataGroup_48_13 = dataGroup_lo_880[1951:1944];
  wire [2047:0] dataGroup_lo_881 = {dataGroup_lo_hi_881, dataGroup_lo_lo_881};
  wire [2047:0] dataGroup_hi_881 = {dataGroup_hi_hi_881, dataGroup_hi_lo_881};
  wire [7:0]    dataGroup_49_13 = dataGroup_lo_881[1991:1984];
  wire [2047:0] dataGroup_lo_882 = {dataGroup_lo_hi_882, dataGroup_lo_lo_882};
  wire [2047:0] dataGroup_hi_882 = {dataGroup_hi_hi_882, dataGroup_hi_lo_882};
  wire [7:0]    dataGroup_50_13 = dataGroup_lo_882[2031:2024];
  wire [2047:0] dataGroup_lo_883 = {dataGroup_lo_hi_883, dataGroup_lo_lo_883};
  wire [2047:0] dataGroup_hi_883 = {dataGroup_hi_hi_883, dataGroup_hi_lo_883};
  wire [7:0]    dataGroup_51_13 = dataGroup_hi_883[23:16];
  wire [2047:0] dataGroup_lo_884 = {dataGroup_lo_hi_884, dataGroup_lo_lo_884};
  wire [2047:0] dataGroup_hi_884 = {dataGroup_hi_hi_884, dataGroup_hi_lo_884};
  wire [7:0]    dataGroup_52_13 = dataGroup_hi_884[63:56];
  wire [2047:0] dataGroup_lo_885 = {dataGroup_lo_hi_885, dataGroup_lo_lo_885};
  wire [2047:0] dataGroup_hi_885 = {dataGroup_hi_hi_885, dataGroup_hi_lo_885};
  wire [7:0]    dataGroup_53_13 = dataGroup_hi_885[103:96];
  wire [2047:0] dataGroup_lo_886 = {dataGroup_lo_hi_886, dataGroup_lo_lo_886};
  wire [2047:0] dataGroup_hi_886 = {dataGroup_hi_hi_886, dataGroup_hi_lo_886};
  wire [7:0]    dataGroup_54_13 = dataGroup_hi_886[143:136];
  wire [2047:0] dataGroup_lo_887 = {dataGroup_lo_hi_887, dataGroup_lo_lo_887};
  wire [2047:0] dataGroup_hi_887 = {dataGroup_hi_hi_887, dataGroup_hi_lo_887};
  wire [7:0]    dataGroup_55_13 = dataGroup_hi_887[183:176];
  wire [2047:0] dataGroup_lo_888 = {dataGroup_lo_hi_888, dataGroup_lo_lo_888};
  wire [2047:0] dataGroup_hi_888 = {dataGroup_hi_hi_888, dataGroup_hi_lo_888};
  wire [7:0]    dataGroup_56_13 = dataGroup_hi_888[223:216];
  wire [2047:0] dataGroup_lo_889 = {dataGroup_lo_hi_889, dataGroup_lo_lo_889};
  wire [2047:0] dataGroup_hi_889 = {dataGroup_hi_hi_889, dataGroup_hi_lo_889};
  wire [7:0]    dataGroup_57_13 = dataGroup_hi_889[263:256];
  wire [2047:0] dataGroup_lo_890 = {dataGroup_lo_hi_890, dataGroup_lo_lo_890};
  wire [2047:0] dataGroup_hi_890 = {dataGroup_hi_hi_890, dataGroup_hi_lo_890};
  wire [7:0]    dataGroup_58_13 = dataGroup_hi_890[303:296];
  wire [2047:0] dataGroup_lo_891 = {dataGroup_lo_hi_891, dataGroup_lo_lo_891};
  wire [2047:0] dataGroup_hi_891 = {dataGroup_hi_hi_891, dataGroup_hi_lo_891};
  wire [7:0]    dataGroup_59_13 = dataGroup_hi_891[343:336];
  wire [2047:0] dataGroup_lo_892 = {dataGroup_lo_hi_892, dataGroup_lo_lo_892};
  wire [2047:0] dataGroup_hi_892 = {dataGroup_hi_hi_892, dataGroup_hi_lo_892};
  wire [7:0]    dataGroup_60_13 = dataGroup_hi_892[383:376];
  wire [2047:0] dataGroup_lo_893 = {dataGroup_lo_hi_893, dataGroup_lo_lo_893};
  wire [2047:0] dataGroup_hi_893 = {dataGroup_hi_hi_893, dataGroup_hi_lo_893};
  wire [7:0]    dataGroup_61_13 = dataGroup_hi_893[423:416];
  wire [2047:0] dataGroup_lo_894 = {dataGroup_lo_hi_894, dataGroup_lo_lo_894};
  wire [2047:0] dataGroup_hi_894 = {dataGroup_hi_hi_894, dataGroup_hi_lo_894};
  wire [7:0]    dataGroup_62_13 = dataGroup_hi_894[463:456];
  wire [2047:0] dataGroup_lo_895 = {dataGroup_lo_hi_895, dataGroup_lo_lo_895};
  wire [2047:0] dataGroup_hi_895 = {dataGroup_hi_hi_895, dataGroup_hi_lo_895};
  wire [7:0]    dataGroup_63_13 = dataGroup_hi_895[503:496];
  wire [15:0]   res_lo_lo_lo_lo_lo_13 = {dataGroup_1_13, dataGroup_0_13};
  wire [15:0]   res_lo_lo_lo_lo_hi_13 = {dataGroup_3_13, dataGroup_2_13};
  wire [31:0]   res_lo_lo_lo_lo_13 = {res_lo_lo_lo_lo_hi_13, res_lo_lo_lo_lo_lo_13};
  wire [15:0]   res_lo_lo_lo_hi_lo_13 = {dataGroup_5_13, dataGroup_4_13};
  wire [15:0]   res_lo_lo_lo_hi_hi_13 = {dataGroup_7_13, dataGroup_6_13};
  wire [31:0]   res_lo_lo_lo_hi_13 = {res_lo_lo_lo_hi_hi_13, res_lo_lo_lo_hi_lo_13};
  wire [63:0]   res_lo_lo_lo_13 = {res_lo_lo_lo_hi_13, res_lo_lo_lo_lo_13};
  wire [15:0]   res_lo_lo_hi_lo_lo_13 = {dataGroup_9_13, dataGroup_8_13};
  wire [15:0]   res_lo_lo_hi_lo_hi_13 = {dataGroup_11_13, dataGroup_10_13};
  wire [31:0]   res_lo_lo_hi_lo_13 = {res_lo_lo_hi_lo_hi_13, res_lo_lo_hi_lo_lo_13};
  wire [15:0]   res_lo_lo_hi_hi_lo_13 = {dataGroup_13_13, dataGroup_12_13};
  wire [15:0]   res_lo_lo_hi_hi_hi_13 = {dataGroup_15_13, dataGroup_14_13};
  wire [31:0]   res_lo_lo_hi_hi_13 = {res_lo_lo_hi_hi_hi_13, res_lo_lo_hi_hi_lo_13};
  wire [63:0]   res_lo_lo_hi_13 = {res_lo_lo_hi_hi_13, res_lo_lo_hi_lo_13};
  wire [127:0]  res_lo_lo_13 = {res_lo_lo_hi_13, res_lo_lo_lo_13};
  wire [15:0]   res_lo_hi_lo_lo_lo_13 = {dataGroup_17_13, dataGroup_16_13};
  wire [15:0]   res_lo_hi_lo_lo_hi_13 = {dataGroup_19_13, dataGroup_18_13};
  wire [31:0]   res_lo_hi_lo_lo_13 = {res_lo_hi_lo_lo_hi_13, res_lo_hi_lo_lo_lo_13};
  wire [15:0]   res_lo_hi_lo_hi_lo_13 = {dataGroup_21_13, dataGroup_20_13};
  wire [15:0]   res_lo_hi_lo_hi_hi_13 = {dataGroup_23_13, dataGroup_22_13};
  wire [31:0]   res_lo_hi_lo_hi_13 = {res_lo_hi_lo_hi_hi_13, res_lo_hi_lo_hi_lo_13};
  wire [63:0]   res_lo_hi_lo_13 = {res_lo_hi_lo_hi_13, res_lo_hi_lo_lo_13};
  wire [15:0]   res_lo_hi_hi_lo_lo_13 = {dataGroup_25_13, dataGroup_24_13};
  wire [15:0]   res_lo_hi_hi_lo_hi_13 = {dataGroup_27_13, dataGroup_26_13};
  wire [31:0]   res_lo_hi_hi_lo_13 = {res_lo_hi_hi_lo_hi_13, res_lo_hi_hi_lo_lo_13};
  wire [15:0]   res_lo_hi_hi_hi_lo_13 = {dataGroup_29_13, dataGroup_28_13};
  wire [15:0]   res_lo_hi_hi_hi_hi_13 = {dataGroup_31_13, dataGroup_30_13};
  wire [31:0]   res_lo_hi_hi_hi_13 = {res_lo_hi_hi_hi_hi_13, res_lo_hi_hi_hi_lo_13};
  wire [63:0]   res_lo_hi_hi_13 = {res_lo_hi_hi_hi_13, res_lo_hi_hi_lo_13};
  wire [127:0]  res_lo_hi_13 = {res_lo_hi_hi_13, res_lo_hi_lo_13};
  wire [255:0]  res_lo_13 = {res_lo_hi_13, res_lo_lo_13};
  wire [15:0]   res_hi_lo_lo_lo_lo_13 = {dataGroup_33_13, dataGroup_32_13};
  wire [15:0]   res_hi_lo_lo_lo_hi_13 = {dataGroup_35_13, dataGroup_34_13};
  wire [31:0]   res_hi_lo_lo_lo_13 = {res_hi_lo_lo_lo_hi_13, res_hi_lo_lo_lo_lo_13};
  wire [15:0]   res_hi_lo_lo_hi_lo_13 = {dataGroup_37_13, dataGroup_36_13};
  wire [15:0]   res_hi_lo_lo_hi_hi_13 = {dataGroup_39_13, dataGroup_38_13};
  wire [31:0]   res_hi_lo_lo_hi_13 = {res_hi_lo_lo_hi_hi_13, res_hi_lo_lo_hi_lo_13};
  wire [63:0]   res_hi_lo_lo_13 = {res_hi_lo_lo_hi_13, res_hi_lo_lo_lo_13};
  wire [15:0]   res_hi_lo_hi_lo_lo_13 = {dataGroup_41_13, dataGroup_40_13};
  wire [15:0]   res_hi_lo_hi_lo_hi_13 = {dataGroup_43_13, dataGroup_42_13};
  wire [31:0]   res_hi_lo_hi_lo_13 = {res_hi_lo_hi_lo_hi_13, res_hi_lo_hi_lo_lo_13};
  wire [15:0]   res_hi_lo_hi_hi_lo_13 = {dataGroup_45_13, dataGroup_44_13};
  wire [15:0]   res_hi_lo_hi_hi_hi_13 = {dataGroup_47_13, dataGroup_46_13};
  wire [31:0]   res_hi_lo_hi_hi_13 = {res_hi_lo_hi_hi_hi_13, res_hi_lo_hi_hi_lo_13};
  wire [63:0]   res_hi_lo_hi_13 = {res_hi_lo_hi_hi_13, res_hi_lo_hi_lo_13};
  wire [127:0]  res_hi_lo_13 = {res_hi_lo_hi_13, res_hi_lo_lo_13};
  wire [15:0]   res_hi_hi_lo_lo_lo_13 = {dataGroup_49_13, dataGroup_48_13};
  wire [15:0]   res_hi_hi_lo_lo_hi_13 = {dataGroup_51_13, dataGroup_50_13};
  wire [31:0]   res_hi_hi_lo_lo_13 = {res_hi_hi_lo_lo_hi_13, res_hi_hi_lo_lo_lo_13};
  wire [15:0]   res_hi_hi_lo_hi_lo_13 = {dataGroup_53_13, dataGroup_52_13};
  wire [15:0]   res_hi_hi_lo_hi_hi_13 = {dataGroup_55_13, dataGroup_54_13};
  wire [31:0]   res_hi_hi_lo_hi_13 = {res_hi_hi_lo_hi_hi_13, res_hi_hi_lo_hi_lo_13};
  wire [63:0]   res_hi_hi_lo_13 = {res_hi_hi_lo_hi_13, res_hi_hi_lo_lo_13};
  wire [15:0]   res_hi_hi_hi_lo_lo_13 = {dataGroup_57_13, dataGroup_56_13};
  wire [15:0]   res_hi_hi_hi_lo_hi_13 = {dataGroup_59_13, dataGroup_58_13};
  wire [31:0]   res_hi_hi_hi_lo_13 = {res_hi_hi_hi_lo_hi_13, res_hi_hi_hi_lo_lo_13};
  wire [15:0]   res_hi_hi_hi_hi_lo_13 = {dataGroup_61_13, dataGroup_60_13};
  wire [15:0]   res_hi_hi_hi_hi_hi_13 = {dataGroup_63_13, dataGroup_62_13};
  wire [31:0]   res_hi_hi_hi_hi_13 = {res_hi_hi_hi_hi_hi_13, res_hi_hi_hi_hi_lo_13};
  wire [63:0]   res_hi_hi_hi_13 = {res_hi_hi_hi_hi_13, res_hi_hi_hi_lo_13};
  wire [127:0]  res_hi_hi_13 = {res_hi_hi_hi_13, res_hi_hi_lo_13};
  wire [255:0]  res_hi_13 = {res_hi_hi_13, res_hi_lo_13};
  wire [511:0]  res_35 = {res_hi_13, res_lo_13};
  wire [2047:0] dataGroup_lo_896 = {dataGroup_lo_hi_896, dataGroup_lo_lo_896};
  wire [2047:0] dataGroup_hi_896 = {dataGroup_hi_hi_896, dataGroup_hi_lo_896};
  wire [7:0]    dataGroup_0_14 = dataGroup_lo_896[39:32];
  wire [2047:0] dataGroup_lo_897 = {dataGroup_lo_hi_897, dataGroup_lo_lo_897};
  wire [2047:0] dataGroup_hi_897 = {dataGroup_hi_hi_897, dataGroup_hi_lo_897};
  wire [7:0]    dataGroup_1_14 = dataGroup_lo_897[79:72];
  wire [2047:0] dataGroup_lo_898 = {dataGroup_lo_hi_898, dataGroup_lo_lo_898};
  wire [2047:0] dataGroup_hi_898 = {dataGroup_hi_hi_898, dataGroup_hi_lo_898};
  wire [7:0]    dataGroup_2_14 = dataGroup_lo_898[119:112];
  wire [2047:0] dataGroup_lo_899 = {dataGroup_lo_hi_899, dataGroup_lo_lo_899};
  wire [2047:0] dataGroup_hi_899 = {dataGroup_hi_hi_899, dataGroup_hi_lo_899};
  wire [7:0]    dataGroup_3_14 = dataGroup_lo_899[159:152];
  wire [2047:0] dataGroup_lo_900 = {dataGroup_lo_hi_900, dataGroup_lo_lo_900};
  wire [2047:0] dataGroup_hi_900 = {dataGroup_hi_hi_900, dataGroup_hi_lo_900};
  wire [7:0]    dataGroup_4_14 = dataGroup_lo_900[199:192];
  wire [2047:0] dataGroup_lo_901 = {dataGroup_lo_hi_901, dataGroup_lo_lo_901};
  wire [2047:0] dataGroup_hi_901 = {dataGroup_hi_hi_901, dataGroup_hi_lo_901};
  wire [7:0]    dataGroup_5_14 = dataGroup_lo_901[239:232];
  wire [2047:0] dataGroup_lo_902 = {dataGroup_lo_hi_902, dataGroup_lo_lo_902};
  wire [2047:0] dataGroup_hi_902 = {dataGroup_hi_hi_902, dataGroup_hi_lo_902};
  wire [7:0]    dataGroup_6_14 = dataGroup_lo_902[279:272];
  wire [2047:0] dataGroup_lo_903 = {dataGroup_lo_hi_903, dataGroup_lo_lo_903};
  wire [2047:0] dataGroup_hi_903 = {dataGroup_hi_hi_903, dataGroup_hi_lo_903};
  wire [7:0]    dataGroup_7_14 = dataGroup_lo_903[319:312];
  wire [2047:0] dataGroup_lo_904 = {dataGroup_lo_hi_904, dataGroup_lo_lo_904};
  wire [2047:0] dataGroup_hi_904 = {dataGroup_hi_hi_904, dataGroup_hi_lo_904};
  wire [7:0]    dataGroup_8_14 = dataGroup_lo_904[359:352];
  wire [2047:0] dataGroup_lo_905 = {dataGroup_lo_hi_905, dataGroup_lo_lo_905};
  wire [2047:0] dataGroup_hi_905 = {dataGroup_hi_hi_905, dataGroup_hi_lo_905};
  wire [7:0]    dataGroup_9_14 = dataGroup_lo_905[399:392];
  wire [2047:0] dataGroup_lo_906 = {dataGroup_lo_hi_906, dataGroup_lo_lo_906};
  wire [2047:0] dataGroup_hi_906 = {dataGroup_hi_hi_906, dataGroup_hi_lo_906};
  wire [7:0]    dataGroup_10_14 = dataGroup_lo_906[439:432];
  wire [2047:0] dataGroup_lo_907 = {dataGroup_lo_hi_907, dataGroup_lo_lo_907};
  wire [2047:0] dataGroup_hi_907 = {dataGroup_hi_hi_907, dataGroup_hi_lo_907};
  wire [7:0]    dataGroup_11_14 = dataGroup_lo_907[479:472];
  wire [2047:0] dataGroup_lo_908 = {dataGroup_lo_hi_908, dataGroup_lo_lo_908};
  wire [2047:0] dataGroup_hi_908 = {dataGroup_hi_hi_908, dataGroup_hi_lo_908};
  wire [7:0]    dataGroup_12_14 = dataGroup_lo_908[519:512];
  wire [2047:0] dataGroup_lo_909 = {dataGroup_lo_hi_909, dataGroup_lo_lo_909};
  wire [2047:0] dataGroup_hi_909 = {dataGroup_hi_hi_909, dataGroup_hi_lo_909};
  wire [7:0]    dataGroup_13_14 = dataGroup_lo_909[559:552];
  wire [2047:0] dataGroup_lo_910 = {dataGroup_lo_hi_910, dataGroup_lo_lo_910};
  wire [2047:0] dataGroup_hi_910 = {dataGroup_hi_hi_910, dataGroup_hi_lo_910};
  wire [7:0]    dataGroup_14_14 = dataGroup_lo_910[599:592];
  wire [2047:0] dataGroup_lo_911 = {dataGroup_lo_hi_911, dataGroup_lo_lo_911};
  wire [2047:0] dataGroup_hi_911 = {dataGroup_hi_hi_911, dataGroup_hi_lo_911};
  wire [7:0]    dataGroup_15_14 = dataGroup_lo_911[639:632];
  wire [2047:0] dataGroup_lo_912 = {dataGroup_lo_hi_912, dataGroup_lo_lo_912};
  wire [2047:0] dataGroup_hi_912 = {dataGroup_hi_hi_912, dataGroup_hi_lo_912};
  wire [7:0]    dataGroup_16_14 = dataGroup_lo_912[679:672];
  wire [2047:0] dataGroup_lo_913 = {dataGroup_lo_hi_913, dataGroup_lo_lo_913};
  wire [2047:0] dataGroup_hi_913 = {dataGroup_hi_hi_913, dataGroup_hi_lo_913};
  wire [7:0]    dataGroup_17_14 = dataGroup_lo_913[719:712];
  wire [2047:0] dataGroup_lo_914 = {dataGroup_lo_hi_914, dataGroup_lo_lo_914};
  wire [2047:0] dataGroup_hi_914 = {dataGroup_hi_hi_914, dataGroup_hi_lo_914};
  wire [7:0]    dataGroup_18_14 = dataGroup_lo_914[759:752];
  wire [2047:0] dataGroup_lo_915 = {dataGroup_lo_hi_915, dataGroup_lo_lo_915};
  wire [2047:0] dataGroup_hi_915 = {dataGroup_hi_hi_915, dataGroup_hi_lo_915};
  wire [7:0]    dataGroup_19_14 = dataGroup_lo_915[799:792];
  wire [2047:0] dataGroup_lo_916 = {dataGroup_lo_hi_916, dataGroup_lo_lo_916};
  wire [2047:0] dataGroup_hi_916 = {dataGroup_hi_hi_916, dataGroup_hi_lo_916};
  wire [7:0]    dataGroup_20_14 = dataGroup_lo_916[839:832];
  wire [2047:0] dataGroup_lo_917 = {dataGroup_lo_hi_917, dataGroup_lo_lo_917};
  wire [2047:0] dataGroup_hi_917 = {dataGroup_hi_hi_917, dataGroup_hi_lo_917};
  wire [7:0]    dataGroup_21_14 = dataGroup_lo_917[879:872];
  wire [2047:0] dataGroup_lo_918 = {dataGroup_lo_hi_918, dataGroup_lo_lo_918};
  wire [2047:0] dataGroup_hi_918 = {dataGroup_hi_hi_918, dataGroup_hi_lo_918};
  wire [7:0]    dataGroup_22_14 = dataGroup_lo_918[919:912];
  wire [2047:0] dataGroup_lo_919 = {dataGroup_lo_hi_919, dataGroup_lo_lo_919};
  wire [2047:0] dataGroup_hi_919 = {dataGroup_hi_hi_919, dataGroup_hi_lo_919};
  wire [7:0]    dataGroup_23_14 = dataGroup_lo_919[959:952];
  wire [2047:0] dataGroup_lo_920 = {dataGroup_lo_hi_920, dataGroup_lo_lo_920};
  wire [2047:0] dataGroup_hi_920 = {dataGroup_hi_hi_920, dataGroup_hi_lo_920};
  wire [7:0]    dataGroup_24_14 = dataGroup_lo_920[999:992];
  wire [2047:0] dataGroup_lo_921 = {dataGroup_lo_hi_921, dataGroup_lo_lo_921};
  wire [2047:0] dataGroup_hi_921 = {dataGroup_hi_hi_921, dataGroup_hi_lo_921};
  wire [7:0]    dataGroup_25_14 = dataGroup_lo_921[1039:1032];
  wire [2047:0] dataGroup_lo_922 = {dataGroup_lo_hi_922, dataGroup_lo_lo_922};
  wire [2047:0] dataGroup_hi_922 = {dataGroup_hi_hi_922, dataGroup_hi_lo_922};
  wire [7:0]    dataGroup_26_14 = dataGroup_lo_922[1079:1072];
  wire [2047:0] dataGroup_lo_923 = {dataGroup_lo_hi_923, dataGroup_lo_lo_923};
  wire [2047:0] dataGroup_hi_923 = {dataGroup_hi_hi_923, dataGroup_hi_lo_923};
  wire [7:0]    dataGroup_27_14 = dataGroup_lo_923[1119:1112];
  wire [2047:0] dataGroup_lo_924 = {dataGroup_lo_hi_924, dataGroup_lo_lo_924};
  wire [2047:0] dataGroup_hi_924 = {dataGroup_hi_hi_924, dataGroup_hi_lo_924};
  wire [7:0]    dataGroup_28_14 = dataGroup_lo_924[1159:1152];
  wire [2047:0] dataGroup_lo_925 = {dataGroup_lo_hi_925, dataGroup_lo_lo_925};
  wire [2047:0] dataGroup_hi_925 = {dataGroup_hi_hi_925, dataGroup_hi_lo_925};
  wire [7:0]    dataGroup_29_14 = dataGroup_lo_925[1199:1192];
  wire [2047:0] dataGroup_lo_926 = {dataGroup_lo_hi_926, dataGroup_lo_lo_926};
  wire [2047:0] dataGroup_hi_926 = {dataGroup_hi_hi_926, dataGroup_hi_lo_926};
  wire [7:0]    dataGroup_30_14 = dataGroup_lo_926[1239:1232];
  wire [2047:0] dataGroup_lo_927 = {dataGroup_lo_hi_927, dataGroup_lo_lo_927};
  wire [2047:0] dataGroup_hi_927 = {dataGroup_hi_hi_927, dataGroup_hi_lo_927};
  wire [7:0]    dataGroup_31_14 = dataGroup_lo_927[1279:1272];
  wire [2047:0] dataGroup_lo_928 = {dataGroup_lo_hi_928, dataGroup_lo_lo_928};
  wire [2047:0] dataGroup_hi_928 = {dataGroup_hi_hi_928, dataGroup_hi_lo_928};
  wire [7:0]    dataGroup_32_14 = dataGroup_lo_928[1319:1312];
  wire [2047:0] dataGroup_lo_929 = {dataGroup_lo_hi_929, dataGroup_lo_lo_929};
  wire [2047:0] dataGroup_hi_929 = {dataGroup_hi_hi_929, dataGroup_hi_lo_929};
  wire [7:0]    dataGroup_33_14 = dataGroup_lo_929[1359:1352];
  wire [2047:0] dataGroup_lo_930 = {dataGroup_lo_hi_930, dataGroup_lo_lo_930};
  wire [2047:0] dataGroup_hi_930 = {dataGroup_hi_hi_930, dataGroup_hi_lo_930};
  wire [7:0]    dataGroup_34_14 = dataGroup_lo_930[1399:1392];
  wire [2047:0] dataGroup_lo_931 = {dataGroup_lo_hi_931, dataGroup_lo_lo_931};
  wire [2047:0] dataGroup_hi_931 = {dataGroup_hi_hi_931, dataGroup_hi_lo_931};
  wire [7:0]    dataGroup_35_14 = dataGroup_lo_931[1439:1432];
  wire [2047:0] dataGroup_lo_932 = {dataGroup_lo_hi_932, dataGroup_lo_lo_932};
  wire [2047:0] dataGroup_hi_932 = {dataGroup_hi_hi_932, dataGroup_hi_lo_932};
  wire [7:0]    dataGroup_36_14 = dataGroup_lo_932[1479:1472];
  wire [2047:0] dataGroup_lo_933 = {dataGroup_lo_hi_933, dataGroup_lo_lo_933};
  wire [2047:0] dataGroup_hi_933 = {dataGroup_hi_hi_933, dataGroup_hi_lo_933};
  wire [7:0]    dataGroup_37_14 = dataGroup_lo_933[1519:1512];
  wire [2047:0] dataGroup_lo_934 = {dataGroup_lo_hi_934, dataGroup_lo_lo_934};
  wire [2047:0] dataGroup_hi_934 = {dataGroup_hi_hi_934, dataGroup_hi_lo_934};
  wire [7:0]    dataGroup_38_14 = dataGroup_lo_934[1559:1552];
  wire [2047:0] dataGroup_lo_935 = {dataGroup_lo_hi_935, dataGroup_lo_lo_935};
  wire [2047:0] dataGroup_hi_935 = {dataGroup_hi_hi_935, dataGroup_hi_lo_935};
  wire [7:0]    dataGroup_39_14 = dataGroup_lo_935[1599:1592];
  wire [2047:0] dataGroup_lo_936 = {dataGroup_lo_hi_936, dataGroup_lo_lo_936};
  wire [2047:0] dataGroup_hi_936 = {dataGroup_hi_hi_936, dataGroup_hi_lo_936};
  wire [7:0]    dataGroup_40_14 = dataGroup_lo_936[1639:1632];
  wire [2047:0] dataGroup_lo_937 = {dataGroup_lo_hi_937, dataGroup_lo_lo_937};
  wire [2047:0] dataGroup_hi_937 = {dataGroup_hi_hi_937, dataGroup_hi_lo_937};
  wire [7:0]    dataGroup_41_14 = dataGroup_lo_937[1679:1672];
  wire [2047:0] dataGroup_lo_938 = {dataGroup_lo_hi_938, dataGroup_lo_lo_938};
  wire [2047:0] dataGroup_hi_938 = {dataGroup_hi_hi_938, dataGroup_hi_lo_938};
  wire [7:0]    dataGroup_42_14 = dataGroup_lo_938[1719:1712];
  wire [2047:0] dataGroup_lo_939 = {dataGroup_lo_hi_939, dataGroup_lo_lo_939};
  wire [2047:0] dataGroup_hi_939 = {dataGroup_hi_hi_939, dataGroup_hi_lo_939};
  wire [7:0]    dataGroup_43_14 = dataGroup_lo_939[1759:1752];
  wire [2047:0] dataGroup_lo_940 = {dataGroup_lo_hi_940, dataGroup_lo_lo_940};
  wire [2047:0] dataGroup_hi_940 = {dataGroup_hi_hi_940, dataGroup_hi_lo_940};
  wire [7:0]    dataGroup_44_14 = dataGroup_lo_940[1799:1792];
  wire [2047:0] dataGroup_lo_941 = {dataGroup_lo_hi_941, dataGroup_lo_lo_941};
  wire [2047:0] dataGroup_hi_941 = {dataGroup_hi_hi_941, dataGroup_hi_lo_941};
  wire [7:0]    dataGroup_45_14 = dataGroup_lo_941[1839:1832];
  wire [2047:0] dataGroup_lo_942 = {dataGroup_lo_hi_942, dataGroup_lo_lo_942};
  wire [2047:0] dataGroup_hi_942 = {dataGroup_hi_hi_942, dataGroup_hi_lo_942};
  wire [7:0]    dataGroup_46_14 = dataGroup_lo_942[1879:1872];
  wire [2047:0] dataGroup_lo_943 = {dataGroup_lo_hi_943, dataGroup_lo_lo_943};
  wire [2047:0] dataGroup_hi_943 = {dataGroup_hi_hi_943, dataGroup_hi_lo_943};
  wire [7:0]    dataGroup_47_14 = dataGroup_lo_943[1919:1912];
  wire [2047:0] dataGroup_lo_944 = {dataGroup_lo_hi_944, dataGroup_lo_lo_944};
  wire [2047:0] dataGroup_hi_944 = {dataGroup_hi_hi_944, dataGroup_hi_lo_944};
  wire [7:0]    dataGroup_48_14 = dataGroup_lo_944[1959:1952];
  wire [2047:0] dataGroup_lo_945 = {dataGroup_lo_hi_945, dataGroup_lo_lo_945};
  wire [2047:0] dataGroup_hi_945 = {dataGroup_hi_hi_945, dataGroup_hi_lo_945};
  wire [7:0]    dataGroup_49_14 = dataGroup_lo_945[1999:1992];
  wire [2047:0] dataGroup_lo_946 = {dataGroup_lo_hi_946, dataGroup_lo_lo_946};
  wire [2047:0] dataGroup_hi_946 = {dataGroup_hi_hi_946, dataGroup_hi_lo_946};
  wire [7:0]    dataGroup_50_14 = dataGroup_lo_946[2039:2032];
  wire [2047:0] dataGroup_lo_947 = {dataGroup_lo_hi_947, dataGroup_lo_lo_947};
  wire [2047:0] dataGroup_hi_947 = {dataGroup_hi_hi_947, dataGroup_hi_lo_947};
  wire [7:0]    dataGroup_51_14 = dataGroup_hi_947[31:24];
  wire [2047:0] dataGroup_lo_948 = {dataGroup_lo_hi_948, dataGroup_lo_lo_948};
  wire [2047:0] dataGroup_hi_948 = {dataGroup_hi_hi_948, dataGroup_hi_lo_948};
  wire [7:0]    dataGroup_52_14 = dataGroup_hi_948[71:64];
  wire [2047:0] dataGroup_lo_949 = {dataGroup_lo_hi_949, dataGroup_lo_lo_949};
  wire [2047:0] dataGroup_hi_949 = {dataGroup_hi_hi_949, dataGroup_hi_lo_949};
  wire [7:0]    dataGroup_53_14 = dataGroup_hi_949[111:104];
  wire [2047:0] dataGroup_lo_950 = {dataGroup_lo_hi_950, dataGroup_lo_lo_950};
  wire [2047:0] dataGroup_hi_950 = {dataGroup_hi_hi_950, dataGroup_hi_lo_950};
  wire [7:0]    dataGroup_54_14 = dataGroup_hi_950[151:144];
  wire [2047:0] dataGroup_lo_951 = {dataGroup_lo_hi_951, dataGroup_lo_lo_951};
  wire [2047:0] dataGroup_hi_951 = {dataGroup_hi_hi_951, dataGroup_hi_lo_951};
  wire [7:0]    dataGroup_55_14 = dataGroup_hi_951[191:184];
  wire [2047:0] dataGroup_lo_952 = {dataGroup_lo_hi_952, dataGroup_lo_lo_952};
  wire [2047:0] dataGroup_hi_952 = {dataGroup_hi_hi_952, dataGroup_hi_lo_952};
  wire [7:0]    dataGroup_56_14 = dataGroup_hi_952[231:224];
  wire [2047:0] dataGroup_lo_953 = {dataGroup_lo_hi_953, dataGroup_lo_lo_953};
  wire [2047:0] dataGroup_hi_953 = {dataGroup_hi_hi_953, dataGroup_hi_lo_953};
  wire [7:0]    dataGroup_57_14 = dataGroup_hi_953[271:264];
  wire [2047:0] dataGroup_lo_954 = {dataGroup_lo_hi_954, dataGroup_lo_lo_954};
  wire [2047:0] dataGroup_hi_954 = {dataGroup_hi_hi_954, dataGroup_hi_lo_954};
  wire [7:0]    dataGroup_58_14 = dataGroup_hi_954[311:304];
  wire [2047:0] dataGroup_lo_955 = {dataGroup_lo_hi_955, dataGroup_lo_lo_955};
  wire [2047:0] dataGroup_hi_955 = {dataGroup_hi_hi_955, dataGroup_hi_lo_955};
  wire [7:0]    dataGroup_59_14 = dataGroup_hi_955[351:344];
  wire [2047:0] dataGroup_lo_956 = {dataGroup_lo_hi_956, dataGroup_lo_lo_956};
  wire [2047:0] dataGroup_hi_956 = {dataGroup_hi_hi_956, dataGroup_hi_lo_956};
  wire [7:0]    dataGroup_60_14 = dataGroup_hi_956[391:384];
  wire [2047:0] dataGroup_lo_957 = {dataGroup_lo_hi_957, dataGroup_lo_lo_957};
  wire [2047:0] dataGroup_hi_957 = {dataGroup_hi_hi_957, dataGroup_hi_lo_957};
  wire [7:0]    dataGroup_61_14 = dataGroup_hi_957[431:424];
  wire [2047:0] dataGroup_lo_958 = {dataGroup_lo_hi_958, dataGroup_lo_lo_958};
  wire [2047:0] dataGroup_hi_958 = {dataGroup_hi_hi_958, dataGroup_hi_lo_958};
  wire [7:0]    dataGroup_62_14 = dataGroup_hi_958[471:464];
  wire [2047:0] dataGroup_lo_959 = {dataGroup_lo_hi_959, dataGroup_lo_lo_959};
  wire [2047:0] dataGroup_hi_959 = {dataGroup_hi_hi_959, dataGroup_hi_lo_959};
  wire [7:0]    dataGroup_63_14 = dataGroup_hi_959[511:504];
  wire [15:0]   res_lo_lo_lo_lo_lo_14 = {dataGroup_1_14, dataGroup_0_14};
  wire [15:0]   res_lo_lo_lo_lo_hi_14 = {dataGroup_3_14, dataGroup_2_14};
  wire [31:0]   res_lo_lo_lo_lo_14 = {res_lo_lo_lo_lo_hi_14, res_lo_lo_lo_lo_lo_14};
  wire [15:0]   res_lo_lo_lo_hi_lo_14 = {dataGroup_5_14, dataGroup_4_14};
  wire [15:0]   res_lo_lo_lo_hi_hi_14 = {dataGroup_7_14, dataGroup_6_14};
  wire [31:0]   res_lo_lo_lo_hi_14 = {res_lo_lo_lo_hi_hi_14, res_lo_lo_lo_hi_lo_14};
  wire [63:0]   res_lo_lo_lo_14 = {res_lo_lo_lo_hi_14, res_lo_lo_lo_lo_14};
  wire [15:0]   res_lo_lo_hi_lo_lo_14 = {dataGroup_9_14, dataGroup_8_14};
  wire [15:0]   res_lo_lo_hi_lo_hi_14 = {dataGroup_11_14, dataGroup_10_14};
  wire [31:0]   res_lo_lo_hi_lo_14 = {res_lo_lo_hi_lo_hi_14, res_lo_lo_hi_lo_lo_14};
  wire [15:0]   res_lo_lo_hi_hi_lo_14 = {dataGroup_13_14, dataGroup_12_14};
  wire [15:0]   res_lo_lo_hi_hi_hi_14 = {dataGroup_15_14, dataGroup_14_14};
  wire [31:0]   res_lo_lo_hi_hi_14 = {res_lo_lo_hi_hi_hi_14, res_lo_lo_hi_hi_lo_14};
  wire [63:0]   res_lo_lo_hi_14 = {res_lo_lo_hi_hi_14, res_lo_lo_hi_lo_14};
  wire [127:0]  res_lo_lo_14 = {res_lo_lo_hi_14, res_lo_lo_lo_14};
  wire [15:0]   res_lo_hi_lo_lo_lo_14 = {dataGroup_17_14, dataGroup_16_14};
  wire [15:0]   res_lo_hi_lo_lo_hi_14 = {dataGroup_19_14, dataGroup_18_14};
  wire [31:0]   res_lo_hi_lo_lo_14 = {res_lo_hi_lo_lo_hi_14, res_lo_hi_lo_lo_lo_14};
  wire [15:0]   res_lo_hi_lo_hi_lo_14 = {dataGroup_21_14, dataGroup_20_14};
  wire [15:0]   res_lo_hi_lo_hi_hi_14 = {dataGroup_23_14, dataGroup_22_14};
  wire [31:0]   res_lo_hi_lo_hi_14 = {res_lo_hi_lo_hi_hi_14, res_lo_hi_lo_hi_lo_14};
  wire [63:0]   res_lo_hi_lo_14 = {res_lo_hi_lo_hi_14, res_lo_hi_lo_lo_14};
  wire [15:0]   res_lo_hi_hi_lo_lo_14 = {dataGroup_25_14, dataGroup_24_14};
  wire [15:0]   res_lo_hi_hi_lo_hi_14 = {dataGroup_27_14, dataGroup_26_14};
  wire [31:0]   res_lo_hi_hi_lo_14 = {res_lo_hi_hi_lo_hi_14, res_lo_hi_hi_lo_lo_14};
  wire [15:0]   res_lo_hi_hi_hi_lo_14 = {dataGroup_29_14, dataGroup_28_14};
  wire [15:0]   res_lo_hi_hi_hi_hi_14 = {dataGroup_31_14, dataGroup_30_14};
  wire [31:0]   res_lo_hi_hi_hi_14 = {res_lo_hi_hi_hi_hi_14, res_lo_hi_hi_hi_lo_14};
  wire [63:0]   res_lo_hi_hi_14 = {res_lo_hi_hi_hi_14, res_lo_hi_hi_lo_14};
  wire [127:0]  res_lo_hi_14 = {res_lo_hi_hi_14, res_lo_hi_lo_14};
  wire [255:0]  res_lo_14 = {res_lo_hi_14, res_lo_lo_14};
  wire [15:0]   res_hi_lo_lo_lo_lo_14 = {dataGroup_33_14, dataGroup_32_14};
  wire [15:0]   res_hi_lo_lo_lo_hi_14 = {dataGroup_35_14, dataGroup_34_14};
  wire [31:0]   res_hi_lo_lo_lo_14 = {res_hi_lo_lo_lo_hi_14, res_hi_lo_lo_lo_lo_14};
  wire [15:0]   res_hi_lo_lo_hi_lo_14 = {dataGroup_37_14, dataGroup_36_14};
  wire [15:0]   res_hi_lo_lo_hi_hi_14 = {dataGroup_39_14, dataGroup_38_14};
  wire [31:0]   res_hi_lo_lo_hi_14 = {res_hi_lo_lo_hi_hi_14, res_hi_lo_lo_hi_lo_14};
  wire [63:0]   res_hi_lo_lo_14 = {res_hi_lo_lo_hi_14, res_hi_lo_lo_lo_14};
  wire [15:0]   res_hi_lo_hi_lo_lo_14 = {dataGroup_41_14, dataGroup_40_14};
  wire [15:0]   res_hi_lo_hi_lo_hi_14 = {dataGroup_43_14, dataGroup_42_14};
  wire [31:0]   res_hi_lo_hi_lo_14 = {res_hi_lo_hi_lo_hi_14, res_hi_lo_hi_lo_lo_14};
  wire [15:0]   res_hi_lo_hi_hi_lo_14 = {dataGroup_45_14, dataGroup_44_14};
  wire [15:0]   res_hi_lo_hi_hi_hi_14 = {dataGroup_47_14, dataGroup_46_14};
  wire [31:0]   res_hi_lo_hi_hi_14 = {res_hi_lo_hi_hi_hi_14, res_hi_lo_hi_hi_lo_14};
  wire [63:0]   res_hi_lo_hi_14 = {res_hi_lo_hi_hi_14, res_hi_lo_hi_lo_14};
  wire [127:0]  res_hi_lo_14 = {res_hi_lo_hi_14, res_hi_lo_lo_14};
  wire [15:0]   res_hi_hi_lo_lo_lo_14 = {dataGroup_49_14, dataGroup_48_14};
  wire [15:0]   res_hi_hi_lo_lo_hi_14 = {dataGroup_51_14, dataGroup_50_14};
  wire [31:0]   res_hi_hi_lo_lo_14 = {res_hi_hi_lo_lo_hi_14, res_hi_hi_lo_lo_lo_14};
  wire [15:0]   res_hi_hi_lo_hi_lo_14 = {dataGroup_53_14, dataGroup_52_14};
  wire [15:0]   res_hi_hi_lo_hi_hi_14 = {dataGroup_55_14, dataGroup_54_14};
  wire [31:0]   res_hi_hi_lo_hi_14 = {res_hi_hi_lo_hi_hi_14, res_hi_hi_lo_hi_lo_14};
  wire [63:0]   res_hi_hi_lo_14 = {res_hi_hi_lo_hi_14, res_hi_hi_lo_lo_14};
  wire [15:0]   res_hi_hi_hi_lo_lo_14 = {dataGroup_57_14, dataGroup_56_14};
  wire [15:0]   res_hi_hi_hi_lo_hi_14 = {dataGroup_59_14, dataGroup_58_14};
  wire [31:0]   res_hi_hi_hi_lo_14 = {res_hi_hi_hi_lo_hi_14, res_hi_hi_hi_lo_lo_14};
  wire [15:0]   res_hi_hi_hi_hi_lo_14 = {dataGroup_61_14, dataGroup_60_14};
  wire [15:0]   res_hi_hi_hi_hi_hi_14 = {dataGroup_63_14, dataGroup_62_14};
  wire [31:0]   res_hi_hi_hi_hi_14 = {res_hi_hi_hi_hi_hi_14, res_hi_hi_hi_hi_lo_14};
  wire [63:0]   res_hi_hi_hi_14 = {res_hi_hi_hi_hi_14, res_hi_hi_hi_lo_14};
  wire [127:0]  res_hi_hi_14 = {res_hi_hi_hi_14, res_hi_hi_lo_14};
  wire [255:0]  res_hi_14 = {res_hi_hi_14, res_hi_lo_14};
  wire [511:0]  res_36 = {res_hi_14, res_lo_14};
  wire [1023:0] lo_lo_4 = {res_33, res_32};
  wire [1023:0] lo_hi_4 = {res_35, res_34};
  wire [2047:0] lo_4 = {lo_hi_4, lo_lo_4};
  wire [1023:0] hi_lo_4 = {512'h0, res_36};
  wire [2047:0] hi_4 = {1024'h0, hi_lo_4};
  wire [4095:0] regroupLoadData_0_4 = {hi_4, lo_4};
  wire [2047:0] dataGroup_lo_960 = {dataGroup_lo_hi_960, dataGroup_lo_lo_960};
  wire [2047:0] dataGroup_hi_960 = {dataGroup_hi_hi_960, dataGroup_hi_lo_960};
  wire [7:0]    dataGroup_0_15 = dataGroup_lo_960[7:0];
  wire [2047:0] dataGroup_lo_961 = {dataGroup_lo_hi_961, dataGroup_lo_lo_961};
  wire [2047:0] dataGroup_hi_961 = {dataGroup_hi_hi_961, dataGroup_hi_lo_961};
  wire [7:0]    dataGroup_1_15 = dataGroup_lo_961[55:48];
  wire [2047:0] dataGroup_lo_962 = {dataGroup_lo_hi_962, dataGroup_lo_lo_962};
  wire [2047:0] dataGroup_hi_962 = {dataGroup_hi_hi_962, dataGroup_hi_lo_962};
  wire [7:0]    dataGroup_2_15 = dataGroup_lo_962[103:96];
  wire [2047:0] dataGroup_lo_963 = {dataGroup_lo_hi_963, dataGroup_lo_lo_963};
  wire [2047:0] dataGroup_hi_963 = {dataGroup_hi_hi_963, dataGroup_hi_lo_963};
  wire [7:0]    dataGroup_3_15 = dataGroup_lo_963[151:144];
  wire [2047:0] dataGroup_lo_964 = {dataGroup_lo_hi_964, dataGroup_lo_lo_964};
  wire [2047:0] dataGroup_hi_964 = {dataGroup_hi_hi_964, dataGroup_hi_lo_964};
  wire [7:0]    dataGroup_4_15 = dataGroup_lo_964[199:192];
  wire [2047:0] dataGroup_lo_965 = {dataGroup_lo_hi_965, dataGroup_lo_lo_965};
  wire [2047:0] dataGroup_hi_965 = {dataGroup_hi_hi_965, dataGroup_hi_lo_965};
  wire [7:0]    dataGroup_5_15 = dataGroup_lo_965[247:240];
  wire [2047:0] dataGroup_lo_966 = {dataGroup_lo_hi_966, dataGroup_lo_lo_966};
  wire [2047:0] dataGroup_hi_966 = {dataGroup_hi_hi_966, dataGroup_hi_lo_966};
  wire [7:0]    dataGroup_6_15 = dataGroup_lo_966[295:288];
  wire [2047:0] dataGroup_lo_967 = {dataGroup_lo_hi_967, dataGroup_lo_lo_967};
  wire [2047:0] dataGroup_hi_967 = {dataGroup_hi_hi_967, dataGroup_hi_lo_967};
  wire [7:0]    dataGroup_7_15 = dataGroup_lo_967[343:336];
  wire [2047:0] dataGroup_lo_968 = {dataGroup_lo_hi_968, dataGroup_lo_lo_968};
  wire [2047:0] dataGroup_hi_968 = {dataGroup_hi_hi_968, dataGroup_hi_lo_968};
  wire [7:0]    dataGroup_8_15 = dataGroup_lo_968[391:384];
  wire [2047:0] dataGroup_lo_969 = {dataGroup_lo_hi_969, dataGroup_lo_lo_969};
  wire [2047:0] dataGroup_hi_969 = {dataGroup_hi_hi_969, dataGroup_hi_lo_969};
  wire [7:0]    dataGroup_9_15 = dataGroup_lo_969[439:432];
  wire [2047:0] dataGroup_lo_970 = {dataGroup_lo_hi_970, dataGroup_lo_lo_970};
  wire [2047:0] dataGroup_hi_970 = {dataGroup_hi_hi_970, dataGroup_hi_lo_970};
  wire [7:0]    dataGroup_10_15 = dataGroup_lo_970[487:480];
  wire [2047:0] dataGroup_lo_971 = {dataGroup_lo_hi_971, dataGroup_lo_lo_971};
  wire [2047:0] dataGroup_hi_971 = {dataGroup_hi_hi_971, dataGroup_hi_lo_971};
  wire [7:0]    dataGroup_11_15 = dataGroup_lo_971[535:528];
  wire [2047:0] dataGroup_lo_972 = {dataGroup_lo_hi_972, dataGroup_lo_lo_972};
  wire [2047:0] dataGroup_hi_972 = {dataGroup_hi_hi_972, dataGroup_hi_lo_972};
  wire [7:0]    dataGroup_12_15 = dataGroup_lo_972[583:576];
  wire [2047:0] dataGroup_lo_973 = {dataGroup_lo_hi_973, dataGroup_lo_lo_973};
  wire [2047:0] dataGroup_hi_973 = {dataGroup_hi_hi_973, dataGroup_hi_lo_973};
  wire [7:0]    dataGroup_13_15 = dataGroup_lo_973[631:624];
  wire [2047:0] dataGroup_lo_974 = {dataGroup_lo_hi_974, dataGroup_lo_lo_974};
  wire [2047:0] dataGroup_hi_974 = {dataGroup_hi_hi_974, dataGroup_hi_lo_974};
  wire [7:0]    dataGroup_14_15 = dataGroup_lo_974[679:672];
  wire [2047:0] dataGroup_lo_975 = {dataGroup_lo_hi_975, dataGroup_lo_lo_975};
  wire [2047:0] dataGroup_hi_975 = {dataGroup_hi_hi_975, dataGroup_hi_lo_975};
  wire [7:0]    dataGroup_15_15 = dataGroup_lo_975[727:720];
  wire [2047:0] dataGroup_lo_976 = {dataGroup_lo_hi_976, dataGroup_lo_lo_976};
  wire [2047:0] dataGroup_hi_976 = {dataGroup_hi_hi_976, dataGroup_hi_lo_976};
  wire [7:0]    dataGroup_16_15 = dataGroup_lo_976[775:768];
  wire [2047:0] dataGroup_lo_977 = {dataGroup_lo_hi_977, dataGroup_lo_lo_977};
  wire [2047:0] dataGroup_hi_977 = {dataGroup_hi_hi_977, dataGroup_hi_lo_977};
  wire [7:0]    dataGroup_17_15 = dataGroup_lo_977[823:816];
  wire [2047:0] dataGroup_lo_978 = {dataGroup_lo_hi_978, dataGroup_lo_lo_978};
  wire [2047:0] dataGroup_hi_978 = {dataGroup_hi_hi_978, dataGroup_hi_lo_978};
  wire [7:0]    dataGroup_18_15 = dataGroup_lo_978[871:864];
  wire [2047:0] dataGroup_lo_979 = {dataGroup_lo_hi_979, dataGroup_lo_lo_979};
  wire [2047:0] dataGroup_hi_979 = {dataGroup_hi_hi_979, dataGroup_hi_lo_979};
  wire [7:0]    dataGroup_19_15 = dataGroup_lo_979[919:912];
  wire [2047:0] dataGroup_lo_980 = {dataGroup_lo_hi_980, dataGroup_lo_lo_980};
  wire [2047:0] dataGroup_hi_980 = {dataGroup_hi_hi_980, dataGroup_hi_lo_980};
  wire [7:0]    dataGroup_20_15 = dataGroup_lo_980[967:960];
  wire [2047:0] dataGroup_lo_981 = {dataGroup_lo_hi_981, dataGroup_lo_lo_981};
  wire [2047:0] dataGroup_hi_981 = {dataGroup_hi_hi_981, dataGroup_hi_lo_981};
  wire [7:0]    dataGroup_21_15 = dataGroup_lo_981[1015:1008];
  wire [2047:0] dataGroup_lo_982 = {dataGroup_lo_hi_982, dataGroup_lo_lo_982};
  wire [2047:0] dataGroup_hi_982 = {dataGroup_hi_hi_982, dataGroup_hi_lo_982};
  wire [7:0]    dataGroup_22_15 = dataGroup_lo_982[1063:1056];
  wire [2047:0] dataGroup_lo_983 = {dataGroup_lo_hi_983, dataGroup_lo_lo_983};
  wire [2047:0] dataGroup_hi_983 = {dataGroup_hi_hi_983, dataGroup_hi_lo_983};
  wire [7:0]    dataGroup_23_15 = dataGroup_lo_983[1111:1104];
  wire [2047:0] dataGroup_lo_984 = {dataGroup_lo_hi_984, dataGroup_lo_lo_984};
  wire [2047:0] dataGroup_hi_984 = {dataGroup_hi_hi_984, dataGroup_hi_lo_984};
  wire [7:0]    dataGroup_24_15 = dataGroup_lo_984[1159:1152];
  wire [2047:0] dataGroup_lo_985 = {dataGroup_lo_hi_985, dataGroup_lo_lo_985};
  wire [2047:0] dataGroup_hi_985 = {dataGroup_hi_hi_985, dataGroup_hi_lo_985};
  wire [7:0]    dataGroup_25_15 = dataGroup_lo_985[1207:1200];
  wire [2047:0] dataGroup_lo_986 = {dataGroup_lo_hi_986, dataGroup_lo_lo_986};
  wire [2047:0] dataGroup_hi_986 = {dataGroup_hi_hi_986, dataGroup_hi_lo_986};
  wire [7:0]    dataGroup_26_15 = dataGroup_lo_986[1255:1248];
  wire [2047:0] dataGroup_lo_987 = {dataGroup_lo_hi_987, dataGroup_lo_lo_987};
  wire [2047:0] dataGroup_hi_987 = {dataGroup_hi_hi_987, dataGroup_hi_lo_987};
  wire [7:0]    dataGroup_27_15 = dataGroup_lo_987[1303:1296];
  wire [2047:0] dataGroup_lo_988 = {dataGroup_lo_hi_988, dataGroup_lo_lo_988};
  wire [2047:0] dataGroup_hi_988 = {dataGroup_hi_hi_988, dataGroup_hi_lo_988};
  wire [7:0]    dataGroup_28_15 = dataGroup_lo_988[1351:1344];
  wire [2047:0] dataGroup_lo_989 = {dataGroup_lo_hi_989, dataGroup_lo_lo_989};
  wire [2047:0] dataGroup_hi_989 = {dataGroup_hi_hi_989, dataGroup_hi_lo_989};
  wire [7:0]    dataGroup_29_15 = dataGroup_lo_989[1399:1392];
  wire [2047:0] dataGroup_lo_990 = {dataGroup_lo_hi_990, dataGroup_lo_lo_990};
  wire [2047:0] dataGroup_hi_990 = {dataGroup_hi_hi_990, dataGroup_hi_lo_990};
  wire [7:0]    dataGroup_30_15 = dataGroup_lo_990[1447:1440];
  wire [2047:0] dataGroup_lo_991 = {dataGroup_lo_hi_991, dataGroup_lo_lo_991};
  wire [2047:0] dataGroup_hi_991 = {dataGroup_hi_hi_991, dataGroup_hi_lo_991};
  wire [7:0]    dataGroup_31_15 = dataGroup_lo_991[1495:1488];
  wire [2047:0] dataGroup_lo_992 = {dataGroup_lo_hi_992, dataGroup_lo_lo_992};
  wire [2047:0] dataGroup_hi_992 = {dataGroup_hi_hi_992, dataGroup_hi_lo_992};
  wire [7:0]    dataGroup_32_15 = dataGroup_lo_992[1543:1536];
  wire [2047:0] dataGroup_lo_993 = {dataGroup_lo_hi_993, dataGroup_lo_lo_993};
  wire [2047:0] dataGroup_hi_993 = {dataGroup_hi_hi_993, dataGroup_hi_lo_993};
  wire [7:0]    dataGroup_33_15 = dataGroup_lo_993[1591:1584];
  wire [2047:0] dataGroup_lo_994 = {dataGroup_lo_hi_994, dataGroup_lo_lo_994};
  wire [2047:0] dataGroup_hi_994 = {dataGroup_hi_hi_994, dataGroup_hi_lo_994};
  wire [7:0]    dataGroup_34_15 = dataGroup_lo_994[1639:1632];
  wire [2047:0] dataGroup_lo_995 = {dataGroup_lo_hi_995, dataGroup_lo_lo_995};
  wire [2047:0] dataGroup_hi_995 = {dataGroup_hi_hi_995, dataGroup_hi_lo_995};
  wire [7:0]    dataGroup_35_15 = dataGroup_lo_995[1687:1680];
  wire [2047:0] dataGroup_lo_996 = {dataGroup_lo_hi_996, dataGroup_lo_lo_996};
  wire [2047:0] dataGroup_hi_996 = {dataGroup_hi_hi_996, dataGroup_hi_lo_996};
  wire [7:0]    dataGroup_36_15 = dataGroup_lo_996[1735:1728];
  wire [2047:0] dataGroup_lo_997 = {dataGroup_lo_hi_997, dataGroup_lo_lo_997};
  wire [2047:0] dataGroup_hi_997 = {dataGroup_hi_hi_997, dataGroup_hi_lo_997};
  wire [7:0]    dataGroup_37_15 = dataGroup_lo_997[1783:1776];
  wire [2047:0] dataGroup_lo_998 = {dataGroup_lo_hi_998, dataGroup_lo_lo_998};
  wire [2047:0] dataGroup_hi_998 = {dataGroup_hi_hi_998, dataGroup_hi_lo_998};
  wire [7:0]    dataGroup_38_15 = dataGroup_lo_998[1831:1824];
  wire [2047:0] dataGroup_lo_999 = {dataGroup_lo_hi_999, dataGroup_lo_lo_999};
  wire [2047:0] dataGroup_hi_999 = {dataGroup_hi_hi_999, dataGroup_hi_lo_999};
  wire [7:0]    dataGroup_39_15 = dataGroup_lo_999[1879:1872];
  wire [2047:0] dataGroup_lo_1000 = {dataGroup_lo_hi_1000, dataGroup_lo_lo_1000};
  wire [2047:0] dataGroup_hi_1000 = {dataGroup_hi_hi_1000, dataGroup_hi_lo_1000};
  wire [7:0]    dataGroup_40_15 = dataGroup_lo_1000[1927:1920];
  wire [2047:0] dataGroup_lo_1001 = {dataGroup_lo_hi_1001, dataGroup_lo_lo_1001};
  wire [2047:0] dataGroup_hi_1001 = {dataGroup_hi_hi_1001, dataGroup_hi_lo_1001};
  wire [7:0]    dataGroup_41_15 = dataGroup_lo_1001[1975:1968];
  wire [2047:0] dataGroup_lo_1002 = {dataGroup_lo_hi_1002, dataGroup_lo_lo_1002};
  wire [2047:0] dataGroup_hi_1002 = {dataGroup_hi_hi_1002, dataGroup_hi_lo_1002};
  wire [7:0]    dataGroup_42_15 = dataGroup_lo_1002[2023:2016];
  wire [2047:0] dataGroup_lo_1003 = {dataGroup_lo_hi_1003, dataGroup_lo_lo_1003};
  wire [2047:0] dataGroup_hi_1003 = {dataGroup_hi_hi_1003, dataGroup_hi_lo_1003};
  wire [7:0]    dataGroup_43_15 = dataGroup_hi_1003[23:16];
  wire [2047:0] dataGroup_lo_1004 = {dataGroup_lo_hi_1004, dataGroup_lo_lo_1004};
  wire [2047:0] dataGroup_hi_1004 = {dataGroup_hi_hi_1004, dataGroup_hi_lo_1004};
  wire [7:0]    dataGroup_44_15 = dataGroup_hi_1004[71:64];
  wire [2047:0] dataGroup_lo_1005 = {dataGroup_lo_hi_1005, dataGroup_lo_lo_1005};
  wire [2047:0] dataGroup_hi_1005 = {dataGroup_hi_hi_1005, dataGroup_hi_lo_1005};
  wire [7:0]    dataGroup_45_15 = dataGroup_hi_1005[119:112];
  wire [2047:0] dataGroup_lo_1006 = {dataGroup_lo_hi_1006, dataGroup_lo_lo_1006};
  wire [2047:0] dataGroup_hi_1006 = {dataGroup_hi_hi_1006, dataGroup_hi_lo_1006};
  wire [7:0]    dataGroup_46_15 = dataGroup_hi_1006[167:160];
  wire [2047:0] dataGroup_lo_1007 = {dataGroup_lo_hi_1007, dataGroup_lo_lo_1007};
  wire [2047:0] dataGroup_hi_1007 = {dataGroup_hi_hi_1007, dataGroup_hi_lo_1007};
  wire [7:0]    dataGroup_47_15 = dataGroup_hi_1007[215:208];
  wire [2047:0] dataGroup_lo_1008 = {dataGroup_lo_hi_1008, dataGroup_lo_lo_1008};
  wire [2047:0] dataGroup_hi_1008 = {dataGroup_hi_hi_1008, dataGroup_hi_lo_1008};
  wire [7:0]    dataGroup_48_15 = dataGroup_hi_1008[263:256];
  wire [2047:0] dataGroup_lo_1009 = {dataGroup_lo_hi_1009, dataGroup_lo_lo_1009};
  wire [2047:0] dataGroup_hi_1009 = {dataGroup_hi_hi_1009, dataGroup_hi_lo_1009};
  wire [7:0]    dataGroup_49_15 = dataGroup_hi_1009[311:304];
  wire [2047:0] dataGroup_lo_1010 = {dataGroup_lo_hi_1010, dataGroup_lo_lo_1010};
  wire [2047:0] dataGroup_hi_1010 = {dataGroup_hi_hi_1010, dataGroup_hi_lo_1010};
  wire [7:0]    dataGroup_50_15 = dataGroup_hi_1010[359:352];
  wire [2047:0] dataGroup_lo_1011 = {dataGroup_lo_hi_1011, dataGroup_lo_lo_1011};
  wire [2047:0] dataGroup_hi_1011 = {dataGroup_hi_hi_1011, dataGroup_hi_lo_1011};
  wire [7:0]    dataGroup_51_15 = dataGroup_hi_1011[407:400];
  wire [2047:0] dataGroup_lo_1012 = {dataGroup_lo_hi_1012, dataGroup_lo_lo_1012};
  wire [2047:0] dataGroup_hi_1012 = {dataGroup_hi_hi_1012, dataGroup_hi_lo_1012};
  wire [7:0]    dataGroup_52_15 = dataGroup_hi_1012[455:448];
  wire [2047:0] dataGroup_lo_1013 = {dataGroup_lo_hi_1013, dataGroup_lo_lo_1013};
  wire [2047:0] dataGroup_hi_1013 = {dataGroup_hi_hi_1013, dataGroup_hi_lo_1013};
  wire [7:0]    dataGroup_53_15 = dataGroup_hi_1013[503:496];
  wire [2047:0] dataGroup_lo_1014 = {dataGroup_lo_hi_1014, dataGroup_lo_lo_1014};
  wire [2047:0] dataGroup_hi_1014 = {dataGroup_hi_hi_1014, dataGroup_hi_lo_1014};
  wire [7:0]    dataGroup_54_15 = dataGroup_hi_1014[551:544];
  wire [2047:0] dataGroup_lo_1015 = {dataGroup_lo_hi_1015, dataGroup_lo_lo_1015};
  wire [2047:0] dataGroup_hi_1015 = {dataGroup_hi_hi_1015, dataGroup_hi_lo_1015};
  wire [7:0]    dataGroup_55_15 = dataGroup_hi_1015[599:592];
  wire [2047:0] dataGroup_lo_1016 = {dataGroup_lo_hi_1016, dataGroup_lo_lo_1016};
  wire [2047:0] dataGroup_hi_1016 = {dataGroup_hi_hi_1016, dataGroup_hi_lo_1016};
  wire [7:0]    dataGroup_56_15 = dataGroup_hi_1016[647:640];
  wire [2047:0] dataGroup_lo_1017 = {dataGroup_lo_hi_1017, dataGroup_lo_lo_1017};
  wire [2047:0] dataGroup_hi_1017 = {dataGroup_hi_hi_1017, dataGroup_hi_lo_1017};
  wire [7:0]    dataGroup_57_15 = dataGroup_hi_1017[695:688];
  wire [2047:0] dataGroup_lo_1018 = {dataGroup_lo_hi_1018, dataGroup_lo_lo_1018};
  wire [2047:0] dataGroup_hi_1018 = {dataGroup_hi_hi_1018, dataGroup_hi_lo_1018};
  wire [7:0]    dataGroup_58_15 = dataGroup_hi_1018[743:736];
  wire [2047:0] dataGroup_lo_1019 = {dataGroup_lo_hi_1019, dataGroup_lo_lo_1019};
  wire [2047:0] dataGroup_hi_1019 = {dataGroup_hi_hi_1019, dataGroup_hi_lo_1019};
  wire [7:0]    dataGroup_59_15 = dataGroup_hi_1019[791:784];
  wire [2047:0] dataGroup_lo_1020 = {dataGroup_lo_hi_1020, dataGroup_lo_lo_1020};
  wire [2047:0] dataGroup_hi_1020 = {dataGroup_hi_hi_1020, dataGroup_hi_lo_1020};
  wire [7:0]    dataGroup_60_15 = dataGroup_hi_1020[839:832];
  wire [2047:0] dataGroup_lo_1021 = {dataGroup_lo_hi_1021, dataGroup_lo_lo_1021};
  wire [2047:0] dataGroup_hi_1021 = {dataGroup_hi_hi_1021, dataGroup_hi_lo_1021};
  wire [7:0]    dataGroup_61_15 = dataGroup_hi_1021[887:880];
  wire [2047:0] dataGroup_lo_1022 = {dataGroup_lo_hi_1022, dataGroup_lo_lo_1022};
  wire [2047:0] dataGroup_hi_1022 = {dataGroup_hi_hi_1022, dataGroup_hi_lo_1022};
  wire [7:0]    dataGroup_62_15 = dataGroup_hi_1022[935:928];
  wire [2047:0] dataGroup_lo_1023 = {dataGroup_lo_hi_1023, dataGroup_lo_lo_1023};
  wire [2047:0] dataGroup_hi_1023 = {dataGroup_hi_hi_1023, dataGroup_hi_lo_1023};
  wire [7:0]    dataGroup_63_15 = dataGroup_hi_1023[983:976];
  wire [15:0]   res_lo_lo_lo_lo_lo_15 = {dataGroup_1_15, dataGroup_0_15};
  wire [15:0]   res_lo_lo_lo_lo_hi_15 = {dataGroup_3_15, dataGroup_2_15};
  wire [31:0]   res_lo_lo_lo_lo_15 = {res_lo_lo_lo_lo_hi_15, res_lo_lo_lo_lo_lo_15};
  wire [15:0]   res_lo_lo_lo_hi_lo_15 = {dataGroup_5_15, dataGroup_4_15};
  wire [15:0]   res_lo_lo_lo_hi_hi_15 = {dataGroup_7_15, dataGroup_6_15};
  wire [31:0]   res_lo_lo_lo_hi_15 = {res_lo_lo_lo_hi_hi_15, res_lo_lo_lo_hi_lo_15};
  wire [63:0]   res_lo_lo_lo_15 = {res_lo_lo_lo_hi_15, res_lo_lo_lo_lo_15};
  wire [15:0]   res_lo_lo_hi_lo_lo_15 = {dataGroup_9_15, dataGroup_8_15};
  wire [15:0]   res_lo_lo_hi_lo_hi_15 = {dataGroup_11_15, dataGroup_10_15};
  wire [31:0]   res_lo_lo_hi_lo_15 = {res_lo_lo_hi_lo_hi_15, res_lo_lo_hi_lo_lo_15};
  wire [15:0]   res_lo_lo_hi_hi_lo_15 = {dataGroup_13_15, dataGroup_12_15};
  wire [15:0]   res_lo_lo_hi_hi_hi_15 = {dataGroup_15_15, dataGroup_14_15};
  wire [31:0]   res_lo_lo_hi_hi_15 = {res_lo_lo_hi_hi_hi_15, res_lo_lo_hi_hi_lo_15};
  wire [63:0]   res_lo_lo_hi_15 = {res_lo_lo_hi_hi_15, res_lo_lo_hi_lo_15};
  wire [127:0]  res_lo_lo_15 = {res_lo_lo_hi_15, res_lo_lo_lo_15};
  wire [15:0]   res_lo_hi_lo_lo_lo_15 = {dataGroup_17_15, dataGroup_16_15};
  wire [15:0]   res_lo_hi_lo_lo_hi_15 = {dataGroup_19_15, dataGroup_18_15};
  wire [31:0]   res_lo_hi_lo_lo_15 = {res_lo_hi_lo_lo_hi_15, res_lo_hi_lo_lo_lo_15};
  wire [15:0]   res_lo_hi_lo_hi_lo_15 = {dataGroup_21_15, dataGroup_20_15};
  wire [15:0]   res_lo_hi_lo_hi_hi_15 = {dataGroup_23_15, dataGroup_22_15};
  wire [31:0]   res_lo_hi_lo_hi_15 = {res_lo_hi_lo_hi_hi_15, res_lo_hi_lo_hi_lo_15};
  wire [63:0]   res_lo_hi_lo_15 = {res_lo_hi_lo_hi_15, res_lo_hi_lo_lo_15};
  wire [15:0]   res_lo_hi_hi_lo_lo_15 = {dataGroup_25_15, dataGroup_24_15};
  wire [15:0]   res_lo_hi_hi_lo_hi_15 = {dataGroup_27_15, dataGroup_26_15};
  wire [31:0]   res_lo_hi_hi_lo_15 = {res_lo_hi_hi_lo_hi_15, res_lo_hi_hi_lo_lo_15};
  wire [15:0]   res_lo_hi_hi_hi_lo_15 = {dataGroup_29_15, dataGroup_28_15};
  wire [15:0]   res_lo_hi_hi_hi_hi_15 = {dataGroup_31_15, dataGroup_30_15};
  wire [31:0]   res_lo_hi_hi_hi_15 = {res_lo_hi_hi_hi_hi_15, res_lo_hi_hi_hi_lo_15};
  wire [63:0]   res_lo_hi_hi_15 = {res_lo_hi_hi_hi_15, res_lo_hi_hi_lo_15};
  wire [127:0]  res_lo_hi_15 = {res_lo_hi_hi_15, res_lo_hi_lo_15};
  wire [255:0]  res_lo_15 = {res_lo_hi_15, res_lo_lo_15};
  wire [15:0]   res_hi_lo_lo_lo_lo_15 = {dataGroup_33_15, dataGroup_32_15};
  wire [15:0]   res_hi_lo_lo_lo_hi_15 = {dataGroup_35_15, dataGroup_34_15};
  wire [31:0]   res_hi_lo_lo_lo_15 = {res_hi_lo_lo_lo_hi_15, res_hi_lo_lo_lo_lo_15};
  wire [15:0]   res_hi_lo_lo_hi_lo_15 = {dataGroup_37_15, dataGroup_36_15};
  wire [15:0]   res_hi_lo_lo_hi_hi_15 = {dataGroup_39_15, dataGroup_38_15};
  wire [31:0]   res_hi_lo_lo_hi_15 = {res_hi_lo_lo_hi_hi_15, res_hi_lo_lo_hi_lo_15};
  wire [63:0]   res_hi_lo_lo_15 = {res_hi_lo_lo_hi_15, res_hi_lo_lo_lo_15};
  wire [15:0]   res_hi_lo_hi_lo_lo_15 = {dataGroup_41_15, dataGroup_40_15};
  wire [15:0]   res_hi_lo_hi_lo_hi_15 = {dataGroup_43_15, dataGroup_42_15};
  wire [31:0]   res_hi_lo_hi_lo_15 = {res_hi_lo_hi_lo_hi_15, res_hi_lo_hi_lo_lo_15};
  wire [15:0]   res_hi_lo_hi_hi_lo_15 = {dataGroup_45_15, dataGroup_44_15};
  wire [15:0]   res_hi_lo_hi_hi_hi_15 = {dataGroup_47_15, dataGroup_46_15};
  wire [31:0]   res_hi_lo_hi_hi_15 = {res_hi_lo_hi_hi_hi_15, res_hi_lo_hi_hi_lo_15};
  wire [63:0]   res_hi_lo_hi_15 = {res_hi_lo_hi_hi_15, res_hi_lo_hi_lo_15};
  wire [127:0]  res_hi_lo_15 = {res_hi_lo_hi_15, res_hi_lo_lo_15};
  wire [15:0]   res_hi_hi_lo_lo_lo_15 = {dataGroup_49_15, dataGroup_48_15};
  wire [15:0]   res_hi_hi_lo_lo_hi_15 = {dataGroup_51_15, dataGroup_50_15};
  wire [31:0]   res_hi_hi_lo_lo_15 = {res_hi_hi_lo_lo_hi_15, res_hi_hi_lo_lo_lo_15};
  wire [15:0]   res_hi_hi_lo_hi_lo_15 = {dataGroup_53_15, dataGroup_52_15};
  wire [15:0]   res_hi_hi_lo_hi_hi_15 = {dataGroup_55_15, dataGroup_54_15};
  wire [31:0]   res_hi_hi_lo_hi_15 = {res_hi_hi_lo_hi_hi_15, res_hi_hi_lo_hi_lo_15};
  wire [63:0]   res_hi_hi_lo_15 = {res_hi_hi_lo_hi_15, res_hi_hi_lo_lo_15};
  wire [15:0]   res_hi_hi_hi_lo_lo_15 = {dataGroup_57_15, dataGroup_56_15};
  wire [15:0]   res_hi_hi_hi_lo_hi_15 = {dataGroup_59_15, dataGroup_58_15};
  wire [31:0]   res_hi_hi_hi_lo_15 = {res_hi_hi_hi_lo_hi_15, res_hi_hi_hi_lo_lo_15};
  wire [15:0]   res_hi_hi_hi_hi_lo_15 = {dataGroup_61_15, dataGroup_60_15};
  wire [15:0]   res_hi_hi_hi_hi_hi_15 = {dataGroup_63_15, dataGroup_62_15};
  wire [31:0]   res_hi_hi_hi_hi_15 = {res_hi_hi_hi_hi_hi_15, res_hi_hi_hi_hi_lo_15};
  wire [63:0]   res_hi_hi_hi_15 = {res_hi_hi_hi_hi_15, res_hi_hi_hi_lo_15};
  wire [127:0]  res_hi_hi_15 = {res_hi_hi_hi_15, res_hi_hi_lo_15};
  wire [255:0]  res_hi_15 = {res_hi_hi_15, res_hi_lo_15};
  wire [511:0]  res_40 = {res_hi_15, res_lo_15};
  wire [2047:0] dataGroup_lo_1024 = {dataGroup_lo_hi_1024, dataGroup_lo_lo_1024};
  wire [2047:0] dataGroup_hi_1024 = {dataGroup_hi_hi_1024, dataGroup_hi_lo_1024};
  wire [7:0]    dataGroup_0_16 = dataGroup_lo_1024[15:8];
  wire [2047:0] dataGroup_lo_1025 = {dataGroup_lo_hi_1025, dataGroup_lo_lo_1025};
  wire [2047:0] dataGroup_hi_1025 = {dataGroup_hi_hi_1025, dataGroup_hi_lo_1025};
  wire [7:0]    dataGroup_1_16 = dataGroup_lo_1025[63:56];
  wire [2047:0] dataGroup_lo_1026 = {dataGroup_lo_hi_1026, dataGroup_lo_lo_1026};
  wire [2047:0] dataGroup_hi_1026 = {dataGroup_hi_hi_1026, dataGroup_hi_lo_1026};
  wire [7:0]    dataGroup_2_16 = dataGroup_lo_1026[111:104];
  wire [2047:0] dataGroup_lo_1027 = {dataGroup_lo_hi_1027, dataGroup_lo_lo_1027};
  wire [2047:0] dataGroup_hi_1027 = {dataGroup_hi_hi_1027, dataGroup_hi_lo_1027};
  wire [7:0]    dataGroup_3_16 = dataGroup_lo_1027[159:152];
  wire [2047:0] dataGroup_lo_1028 = {dataGroup_lo_hi_1028, dataGroup_lo_lo_1028};
  wire [2047:0] dataGroup_hi_1028 = {dataGroup_hi_hi_1028, dataGroup_hi_lo_1028};
  wire [7:0]    dataGroup_4_16 = dataGroup_lo_1028[207:200];
  wire [2047:0] dataGroup_lo_1029 = {dataGroup_lo_hi_1029, dataGroup_lo_lo_1029};
  wire [2047:0] dataGroup_hi_1029 = {dataGroup_hi_hi_1029, dataGroup_hi_lo_1029};
  wire [7:0]    dataGroup_5_16 = dataGroup_lo_1029[255:248];
  wire [2047:0] dataGroup_lo_1030 = {dataGroup_lo_hi_1030, dataGroup_lo_lo_1030};
  wire [2047:0] dataGroup_hi_1030 = {dataGroup_hi_hi_1030, dataGroup_hi_lo_1030};
  wire [7:0]    dataGroup_6_16 = dataGroup_lo_1030[303:296];
  wire [2047:0] dataGroup_lo_1031 = {dataGroup_lo_hi_1031, dataGroup_lo_lo_1031};
  wire [2047:0] dataGroup_hi_1031 = {dataGroup_hi_hi_1031, dataGroup_hi_lo_1031};
  wire [7:0]    dataGroup_7_16 = dataGroup_lo_1031[351:344];
  wire [2047:0] dataGroup_lo_1032 = {dataGroup_lo_hi_1032, dataGroup_lo_lo_1032};
  wire [2047:0] dataGroup_hi_1032 = {dataGroup_hi_hi_1032, dataGroup_hi_lo_1032};
  wire [7:0]    dataGroup_8_16 = dataGroup_lo_1032[399:392];
  wire [2047:0] dataGroup_lo_1033 = {dataGroup_lo_hi_1033, dataGroup_lo_lo_1033};
  wire [2047:0] dataGroup_hi_1033 = {dataGroup_hi_hi_1033, dataGroup_hi_lo_1033};
  wire [7:0]    dataGroup_9_16 = dataGroup_lo_1033[447:440];
  wire [2047:0] dataGroup_lo_1034 = {dataGroup_lo_hi_1034, dataGroup_lo_lo_1034};
  wire [2047:0] dataGroup_hi_1034 = {dataGroup_hi_hi_1034, dataGroup_hi_lo_1034};
  wire [7:0]    dataGroup_10_16 = dataGroup_lo_1034[495:488];
  wire [2047:0] dataGroup_lo_1035 = {dataGroup_lo_hi_1035, dataGroup_lo_lo_1035};
  wire [2047:0] dataGroup_hi_1035 = {dataGroup_hi_hi_1035, dataGroup_hi_lo_1035};
  wire [7:0]    dataGroup_11_16 = dataGroup_lo_1035[543:536];
  wire [2047:0] dataGroup_lo_1036 = {dataGroup_lo_hi_1036, dataGroup_lo_lo_1036};
  wire [2047:0] dataGroup_hi_1036 = {dataGroup_hi_hi_1036, dataGroup_hi_lo_1036};
  wire [7:0]    dataGroup_12_16 = dataGroup_lo_1036[591:584];
  wire [2047:0] dataGroup_lo_1037 = {dataGroup_lo_hi_1037, dataGroup_lo_lo_1037};
  wire [2047:0] dataGroup_hi_1037 = {dataGroup_hi_hi_1037, dataGroup_hi_lo_1037};
  wire [7:0]    dataGroup_13_16 = dataGroup_lo_1037[639:632];
  wire [2047:0] dataGroup_lo_1038 = {dataGroup_lo_hi_1038, dataGroup_lo_lo_1038};
  wire [2047:0] dataGroup_hi_1038 = {dataGroup_hi_hi_1038, dataGroup_hi_lo_1038};
  wire [7:0]    dataGroup_14_16 = dataGroup_lo_1038[687:680];
  wire [2047:0] dataGroup_lo_1039 = {dataGroup_lo_hi_1039, dataGroup_lo_lo_1039};
  wire [2047:0] dataGroup_hi_1039 = {dataGroup_hi_hi_1039, dataGroup_hi_lo_1039};
  wire [7:0]    dataGroup_15_16 = dataGroup_lo_1039[735:728];
  wire [2047:0] dataGroup_lo_1040 = {dataGroup_lo_hi_1040, dataGroup_lo_lo_1040};
  wire [2047:0] dataGroup_hi_1040 = {dataGroup_hi_hi_1040, dataGroup_hi_lo_1040};
  wire [7:0]    dataGroup_16_16 = dataGroup_lo_1040[783:776];
  wire [2047:0] dataGroup_lo_1041 = {dataGroup_lo_hi_1041, dataGroup_lo_lo_1041};
  wire [2047:0] dataGroup_hi_1041 = {dataGroup_hi_hi_1041, dataGroup_hi_lo_1041};
  wire [7:0]    dataGroup_17_16 = dataGroup_lo_1041[831:824];
  wire [2047:0] dataGroup_lo_1042 = {dataGroup_lo_hi_1042, dataGroup_lo_lo_1042};
  wire [2047:0] dataGroup_hi_1042 = {dataGroup_hi_hi_1042, dataGroup_hi_lo_1042};
  wire [7:0]    dataGroup_18_16 = dataGroup_lo_1042[879:872];
  wire [2047:0] dataGroup_lo_1043 = {dataGroup_lo_hi_1043, dataGroup_lo_lo_1043};
  wire [2047:0] dataGroup_hi_1043 = {dataGroup_hi_hi_1043, dataGroup_hi_lo_1043};
  wire [7:0]    dataGroup_19_16 = dataGroup_lo_1043[927:920];
  wire [2047:0] dataGroup_lo_1044 = {dataGroup_lo_hi_1044, dataGroup_lo_lo_1044};
  wire [2047:0] dataGroup_hi_1044 = {dataGroup_hi_hi_1044, dataGroup_hi_lo_1044};
  wire [7:0]    dataGroup_20_16 = dataGroup_lo_1044[975:968];
  wire [2047:0] dataGroup_lo_1045 = {dataGroup_lo_hi_1045, dataGroup_lo_lo_1045};
  wire [2047:0] dataGroup_hi_1045 = {dataGroup_hi_hi_1045, dataGroup_hi_lo_1045};
  wire [7:0]    dataGroup_21_16 = dataGroup_lo_1045[1023:1016];
  wire [2047:0] dataGroup_lo_1046 = {dataGroup_lo_hi_1046, dataGroup_lo_lo_1046};
  wire [2047:0] dataGroup_hi_1046 = {dataGroup_hi_hi_1046, dataGroup_hi_lo_1046};
  wire [7:0]    dataGroup_22_16 = dataGroup_lo_1046[1071:1064];
  wire [2047:0] dataGroup_lo_1047 = {dataGroup_lo_hi_1047, dataGroup_lo_lo_1047};
  wire [2047:0] dataGroup_hi_1047 = {dataGroup_hi_hi_1047, dataGroup_hi_lo_1047};
  wire [7:0]    dataGroup_23_16 = dataGroup_lo_1047[1119:1112];
  wire [2047:0] dataGroup_lo_1048 = {dataGroup_lo_hi_1048, dataGroup_lo_lo_1048};
  wire [2047:0] dataGroup_hi_1048 = {dataGroup_hi_hi_1048, dataGroup_hi_lo_1048};
  wire [7:0]    dataGroup_24_16 = dataGroup_lo_1048[1167:1160];
  wire [2047:0] dataGroup_lo_1049 = {dataGroup_lo_hi_1049, dataGroup_lo_lo_1049};
  wire [2047:0] dataGroup_hi_1049 = {dataGroup_hi_hi_1049, dataGroup_hi_lo_1049};
  wire [7:0]    dataGroup_25_16 = dataGroup_lo_1049[1215:1208];
  wire [2047:0] dataGroup_lo_1050 = {dataGroup_lo_hi_1050, dataGroup_lo_lo_1050};
  wire [2047:0] dataGroup_hi_1050 = {dataGroup_hi_hi_1050, dataGroup_hi_lo_1050};
  wire [7:0]    dataGroup_26_16 = dataGroup_lo_1050[1263:1256];
  wire [2047:0] dataGroup_lo_1051 = {dataGroup_lo_hi_1051, dataGroup_lo_lo_1051};
  wire [2047:0] dataGroup_hi_1051 = {dataGroup_hi_hi_1051, dataGroup_hi_lo_1051};
  wire [7:0]    dataGroup_27_16 = dataGroup_lo_1051[1311:1304];
  wire [2047:0] dataGroup_lo_1052 = {dataGroup_lo_hi_1052, dataGroup_lo_lo_1052};
  wire [2047:0] dataGroup_hi_1052 = {dataGroup_hi_hi_1052, dataGroup_hi_lo_1052};
  wire [7:0]    dataGroup_28_16 = dataGroup_lo_1052[1359:1352];
  wire [2047:0] dataGroup_lo_1053 = {dataGroup_lo_hi_1053, dataGroup_lo_lo_1053};
  wire [2047:0] dataGroup_hi_1053 = {dataGroup_hi_hi_1053, dataGroup_hi_lo_1053};
  wire [7:0]    dataGroup_29_16 = dataGroup_lo_1053[1407:1400];
  wire [2047:0] dataGroup_lo_1054 = {dataGroup_lo_hi_1054, dataGroup_lo_lo_1054};
  wire [2047:0] dataGroup_hi_1054 = {dataGroup_hi_hi_1054, dataGroup_hi_lo_1054};
  wire [7:0]    dataGroup_30_16 = dataGroup_lo_1054[1455:1448];
  wire [2047:0] dataGroup_lo_1055 = {dataGroup_lo_hi_1055, dataGroup_lo_lo_1055};
  wire [2047:0] dataGroup_hi_1055 = {dataGroup_hi_hi_1055, dataGroup_hi_lo_1055};
  wire [7:0]    dataGroup_31_16 = dataGroup_lo_1055[1503:1496];
  wire [2047:0] dataGroup_lo_1056 = {dataGroup_lo_hi_1056, dataGroup_lo_lo_1056};
  wire [2047:0] dataGroup_hi_1056 = {dataGroup_hi_hi_1056, dataGroup_hi_lo_1056};
  wire [7:0]    dataGroup_32_16 = dataGroup_lo_1056[1551:1544];
  wire [2047:0] dataGroup_lo_1057 = {dataGroup_lo_hi_1057, dataGroup_lo_lo_1057};
  wire [2047:0] dataGroup_hi_1057 = {dataGroup_hi_hi_1057, dataGroup_hi_lo_1057};
  wire [7:0]    dataGroup_33_16 = dataGroup_lo_1057[1599:1592];
  wire [2047:0] dataGroup_lo_1058 = {dataGroup_lo_hi_1058, dataGroup_lo_lo_1058};
  wire [2047:0] dataGroup_hi_1058 = {dataGroup_hi_hi_1058, dataGroup_hi_lo_1058};
  wire [7:0]    dataGroup_34_16 = dataGroup_lo_1058[1647:1640];
  wire [2047:0] dataGroup_lo_1059 = {dataGroup_lo_hi_1059, dataGroup_lo_lo_1059};
  wire [2047:0] dataGroup_hi_1059 = {dataGroup_hi_hi_1059, dataGroup_hi_lo_1059};
  wire [7:0]    dataGroup_35_16 = dataGroup_lo_1059[1695:1688];
  wire [2047:0] dataGroup_lo_1060 = {dataGroup_lo_hi_1060, dataGroup_lo_lo_1060};
  wire [2047:0] dataGroup_hi_1060 = {dataGroup_hi_hi_1060, dataGroup_hi_lo_1060};
  wire [7:0]    dataGroup_36_16 = dataGroup_lo_1060[1743:1736];
  wire [2047:0] dataGroup_lo_1061 = {dataGroup_lo_hi_1061, dataGroup_lo_lo_1061};
  wire [2047:0] dataGroup_hi_1061 = {dataGroup_hi_hi_1061, dataGroup_hi_lo_1061};
  wire [7:0]    dataGroup_37_16 = dataGroup_lo_1061[1791:1784];
  wire [2047:0] dataGroup_lo_1062 = {dataGroup_lo_hi_1062, dataGroup_lo_lo_1062};
  wire [2047:0] dataGroup_hi_1062 = {dataGroup_hi_hi_1062, dataGroup_hi_lo_1062};
  wire [7:0]    dataGroup_38_16 = dataGroup_lo_1062[1839:1832];
  wire [2047:0] dataGroup_lo_1063 = {dataGroup_lo_hi_1063, dataGroup_lo_lo_1063};
  wire [2047:0] dataGroup_hi_1063 = {dataGroup_hi_hi_1063, dataGroup_hi_lo_1063};
  wire [7:0]    dataGroup_39_16 = dataGroup_lo_1063[1887:1880];
  wire [2047:0] dataGroup_lo_1064 = {dataGroup_lo_hi_1064, dataGroup_lo_lo_1064};
  wire [2047:0] dataGroup_hi_1064 = {dataGroup_hi_hi_1064, dataGroup_hi_lo_1064};
  wire [7:0]    dataGroup_40_16 = dataGroup_lo_1064[1935:1928];
  wire [2047:0] dataGroup_lo_1065 = {dataGroup_lo_hi_1065, dataGroup_lo_lo_1065};
  wire [2047:0] dataGroup_hi_1065 = {dataGroup_hi_hi_1065, dataGroup_hi_lo_1065};
  wire [7:0]    dataGroup_41_16 = dataGroup_lo_1065[1983:1976];
  wire [2047:0] dataGroup_lo_1066 = {dataGroup_lo_hi_1066, dataGroup_lo_lo_1066};
  wire [2047:0] dataGroup_hi_1066 = {dataGroup_hi_hi_1066, dataGroup_hi_lo_1066};
  wire [7:0]    dataGroup_42_16 = dataGroup_lo_1066[2031:2024];
  wire [2047:0] dataGroup_lo_1067 = {dataGroup_lo_hi_1067, dataGroup_lo_lo_1067};
  wire [2047:0] dataGroup_hi_1067 = {dataGroup_hi_hi_1067, dataGroup_hi_lo_1067};
  wire [7:0]    dataGroup_43_16 = dataGroup_hi_1067[31:24];
  wire [2047:0] dataGroup_lo_1068 = {dataGroup_lo_hi_1068, dataGroup_lo_lo_1068};
  wire [2047:0] dataGroup_hi_1068 = {dataGroup_hi_hi_1068, dataGroup_hi_lo_1068};
  wire [7:0]    dataGroup_44_16 = dataGroup_hi_1068[79:72];
  wire [2047:0] dataGroup_lo_1069 = {dataGroup_lo_hi_1069, dataGroup_lo_lo_1069};
  wire [2047:0] dataGroup_hi_1069 = {dataGroup_hi_hi_1069, dataGroup_hi_lo_1069};
  wire [7:0]    dataGroup_45_16 = dataGroup_hi_1069[127:120];
  wire [2047:0] dataGroup_lo_1070 = {dataGroup_lo_hi_1070, dataGroup_lo_lo_1070};
  wire [2047:0] dataGroup_hi_1070 = {dataGroup_hi_hi_1070, dataGroup_hi_lo_1070};
  wire [7:0]    dataGroup_46_16 = dataGroup_hi_1070[175:168];
  wire [2047:0] dataGroup_lo_1071 = {dataGroup_lo_hi_1071, dataGroup_lo_lo_1071};
  wire [2047:0] dataGroup_hi_1071 = {dataGroup_hi_hi_1071, dataGroup_hi_lo_1071};
  wire [7:0]    dataGroup_47_16 = dataGroup_hi_1071[223:216];
  wire [2047:0] dataGroup_lo_1072 = {dataGroup_lo_hi_1072, dataGroup_lo_lo_1072};
  wire [2047:0] dataGroup_hi_1072 = {dataGroup_hi_hi_1072, dataGroup_hi_lo_1072};
  wire [7:0]    dataGroup_48_16 = dataGroup_hi_1072[271:264];
  wire [2047:0] dataGroup_lo_1073 = {dataGroup_lo_hi_1073, dataGroup_lo_lo_1073};
  wire [2047:0] dataGroup_hi_1073 = {dataGroup_hi_hi_1073, dataGroup_hi_lo_1073};
  wire [7:0]    dataGroup_49_16 = dataGroup_hi_1073[319:312];
  wire [2047:0] dataGroup_lo_1074 = {dataGroup_lo_hi_1074, dataGroup_lo_lo_1074};
  wire [2047:0] dataGroup_hi_1074 = {dataGroup_hi_hi_1074, dataGroup_hi_lo_1074};
  wire [7:0]    dataGroup_50_16 = dataGroup_hi_1074[367:360];
  wire [2047:0] dataGroup_lo_1075 = {dataGroup_lo_hi_1075, dataGroup_lo_lo_1075};
  wire [2047:0] dataGroup_hi_1075 = {dataGroup_hi_hi_1075, dataGroup_hi_lo_1075};
  wire [7:0]    dataGroup_51_16 = dataGroup_hi_1075[415:408];
  wire [2047:0] dataGroup_lo_1076 = {dataGroup_lo_hi_1076, dataGroup_lo_lo_1076};
  wire [2047:0] dataGroup_hi_1076 = {dataGroup_hi_hi_1076, dataGroup_hi_lo_1076};
  wire [7:0]    dataGroup_52_16 = dataGroup_hi_1076[463:456];
  wire [2047:0] dataGroup_lo_1077 = {dataGroup_lo_hi_1077, dataGroup_lo_lo_1077};
  wire [2047:0] dataGroup_hi_1077 = {dataGroup_hi_hi_1077, dataGroup_hi_lo_1077};
  wire [7:0]    dataGroup_53_16 = dataGroup_hi_1077[511:504];
  wire [2047:0] dataGroup_lo_1078 = {dataGroup_lo_hi_1078, dataGroup_lo_lo_1078};
  wire [2047:0] dataGroup_hi_1078 = {dataGroup_hi_hi_1078, dataGroup_hi_lo_1078};
  wire [7:0]    dataGroup_54_16 = dataGroup_hi_1078[559:552];
  wire [2047:0] dataGroup_lo_1079 = {dataGroup_lo_hi_1079, dataGroup_lo_lo_1079};
  wire [2047:0] dataGroup_hi_1079 = {dataGroup_hi_hi_1079, dataGroup_hi_lo_1079};
  wire [7:0]    dataGroup_55_16 = dataGroup_hi_1079[607:600];
  wire [2047:0] dataGroup_lo_1080 = {dataGroup_lo_hi_1080, dataGroup_lo_lo_1080};
  wire [2047:0] dataGroup_hi_1080 = {dataGroup_hi_hi_1080, dataGroup_hi_lo_1080};
  wire [7:0]    dataGroup_56_16 = dataGroup_hi_1080[655:648];
  wire [2047:0] dataGroup_lo_1081 = {dataGroup_lo_hi_1081, dataGroup_lo_lo_1081};
  wire [2047:0] dataGroup_hi_1081 = {dataGroup_hi_hi_1081, dataGroup_hi_lo_1081};
  wire [7:0]    dataGroup_57_16 = dataGroup_hi_1081[703:696];
  wire [2047:0] dataGroup_lo_1082 = {dataGroup_lo_hi_1082, dataGroup_lo_lo_1082};
  wire [2047:0] dataGroup_hi_1082 = {dataGroup_hi_hi_1082, dataGroup_hi_lo_1082};
  wire [7:0]    dataGroup_58_16 = dataGroup_hi_1082[751:744];
  wire [2047:0] dataGroup_lo_1083 = {dataGroup_lo_hi_1083, dataGroup_lo_lo_1083};
  wire [2047:0] dataGroup_hi_1083 = {dataGroup_hi_hi_1083, dataGroup_hi_lo_1083};
  wire [7:0]    dataGroup_59_16 = dataGroup_hi_1083[799:792];
  wire [2047:0] dataGroup_lo_1084 = {dataGroup_lo_hi_1084, dataGroup_lo_lo_1084};
  wire [2047:0] dataGroup_hi_1084 = {dataGroup_hi_hi_1084, dataGroup_hi_lo_1084};
  wire [7:0]    dataGroup_60_16 = dataGroup_hi_1084[847:840];
  wire [2047:0] dataGroup_lo_1085 = {dataGroup_lo_hi_1085, dataGroup_lo_lo_1085};
  wire [2047:0] dataGroup_hi_1085 = {dataGroup_hi_hi_1085, dataGroup_hi_lo_1085};
  wire [7:0]    dataGroup_61_16 = dataGroup_hi_1085[895:888];
  wire [2047:0] dataGroup_lo_1086 = {dataGroup_lo_hi_1086, dataGroup_lo_lo_1086};
  wire [2047:0] dataGroup_hi_1086 = {dataGroup_hi_hi_1086, dataGroup_hi_lo_1086};
  wire [7:0]    dataGroup_62_16 = dataGroup_hi_1086[943:936];
  wire [2047:0] dataGroup_lo_1087 = {dataGroup_lo_hi_1087, dataGroup_lo_lo_1087};
  wire [2047:0] dataGroup_hi_1087 = {dataGroup_hi_hi_1087, dataGroup_hi_lo_1087};
  wire [7:0]    dataGroup_63_16 = dataGroup_hi_1087[991:984];
  wire [15:0]   res_lo_lo_lo_lo_lo_16 = {dataGroup_1_16, dataGroup_0_16};
  wire [15:0]   res_lo_lo_lo_lo_hi_16 = {dataGroup_3_16, dataGroup_2_16};
  wire [31:0]   res_lo_lo_lo_lo_16 = {res_lo_lo_lo_lo_hi_16, res_lo_lo_lo_lo_lo_16};
  wire [15:0]   res_lo_lo_lo_hi_lo_16 = {dataGroup_5_16, dataGroup_4_16};
  wire [15:0]   res_lo_lo_lo_hi_hi_16 = {dataGroup_7_16, dataGroup_6_16};
  wire [31:0]   res_lo_lo_lo_hi_16 = {res_lo_lo_lo_hi_hi_16, res_lo_lo_lo_hi_lo_16};
  wire [63:0]   res_lo_lo_lo_16 = {res_lo_lo_lo_hi_16, res_lo_lo_lo_lo_16};
  wire [15:0]   res_lo_lo_hi_lo_lo_16 = {dataGroup_9_16, dataGroup_8_16};
  wire [15:0]   res_lo_lo_hi_lo_hi_16 = {dataGroup_11_16, dataGroup_10_16};
  wire [31:0]   res_lo_lo_hi_lo_16 = {res_lo_lo_hi_lo_hi_16, res_lo_lo_hi_lo_lo_16};
  wire [15:0]   res_lo_lo_hi_hi_lo_16 = {dataGroup_13_16, dataGroup_12_16};
  wire [15:0]   res_lo_lo_hi_hi_hi_16 = {dataGroup_15_16, dataGroup_14_16};
  wire [31:0]   res_lo_lo_hi_hi_16 = {res_lo_lo_hi_hi_hi_16, res_lo_lo_hi_hi_lo_16};
  wire [63:0]   res_lo_lo_hi_16 = {res_lo_lo_hi_hi_16, res_lo_lo_hi_lo_16};
  wire [127:0]  res_lo_lo_16 = {res_lo_lo_hi_16, res_lo_lo_lo_16};
  wire [15:0]   res_lo_hi_lo_lo_lo_16 = {dataGroup_17_16, dataGroup_16_16};
  wire [15:0]   res_lo_hi_lo_lo_hi_16 = {dataGroup_19_16, dataGroup_18_16};
  wire [31:0]   res_lo_hi_lo_lo_16 = {res_lo_hi_lo_lo_hi_16, res_lo_hi_lo_lo_lo_16};
  wire [15:0]   res_lo_hi_lo_hi_lo_16 = {dataGroup_21_16, dataGroup_20_16};
  wire [15:0]   res_lo_hi_lo_hi_hi_16 = {dataGroup_23_16, dataGroup_22_16};
  wire [31:0]   res_lo_hi_lo_hi_16 = {res_lo_hi_lo_hi_hi_16, res_lo_hi_lo_hi_lo_16};
  wire [63:0]   res_lo_hi_lo_16 = {res_lo_hi_lo_hi_16, res_lo_hi_lo_lo_16};
  wire [15:0]   res_lo_hi_hi_lo_lo_16 = {dataGroup_25_16, dataGroup_24_16};
  wire [15:0]   res_lo_hi_hi_lo_hi_16 = {dataGroup_27_16, dataGroup_26_16};
  wire [31:0]   res_lo_hi_hi_lo_16 = {res_lo_hi_hi_lo_hi_16, res_lo_hi_hi_lo_lo_16};
  wire [15:0]   res_lo_hi_hi_hi_lo_16 = {dataGroup_29_16, dataGroup_28_16};
  wire [15:0]   res_lo_hi_hi_hi_hi_16 = {dataGroup_31_16, dataGroup_30_16};
  wire [31:0]   res_lo_hi_hi_hi_16 = {res_lo_hi_hi_hi_hi_16, res_lo_hi_hi_hi_lo_16};
  wire [63:0]   res_lo_hi_hi_16 = {res_lo_hi_hi_hi_16, res_lo_hi_hi_lo_16};
  wire [127:0]  res_lo_hi_16 = {res_lo_hi_hi_16, res_lo_hi_lo_16};
  wire [255:0]  res_lo_16 = {res_lo_hi_16, res_lo_lo_16};
  wire [15:0]   res_hi_lo_lo_lo_lo_16 = {dataGroup_33_16, dataGroup_32_16};
  wire [15:0]   res_hi_lo_lo_lo_hi_16 = {dataGroup_35_16, dataGroup_34_16};
  wire [31:0]   res_hi_lo_lo_lo_16 = {res_hi_lo_lo_lo_hi_16, res_hi_lo_lo_lo_lo_16};
  wire [15:0]   res_hi_lo_lo_hi_lo_16 = {dataGroup_37_16, dataGroup_36_16};
  wire [15:0]   res_hi_lo_lo_hi_hi_16 = {dataGroup_39_16, dataGroup_38_16};
  wire [31:0]   res_hi_lo_lo_hi_16 = {res_hi_lo_lo_hi_hi_16, res_hi_lo_lo_hi_lo_16};
  wire [63:0]   res_hi_lo_lo_16 = {res_hi_lo_lo_hi_16, res_hi_lo_lo_lo_16};
  wire [15:0]   res_hi_lo_hi_lo_lo_16 = {dataGroup_41_16, dataGroup_40_16};
  wire [15:0]   res_hi_lo_hi_lo_hi_16 = {dataGroup_43_16, dataGroup_42_16};
  wire [31:0]   res_hi_lo_hi_lo_16 = {res_hi_lo_hi_lo_hi_16, res_hi_lo_hi_lo_lo_16};
  wire [15:0]   res_hi_lo_hi_hi_lo_16 = {dataGroup_45_16, dataGroup_44_16};
  wire [15:0]   res_hi_lo_hi_hi_hi_16 = {dataGroup_47_16, dataGroup_46_16};
  wire [31:0]   res_hi_lo_hi_hi_16 = {res_hi_lo_hi_hi_hi_16, res_hi_lo_hi_hi_lo_16};
  wire [63:0]   res_hi_lo_hi_16 = {res_hi_lo_hi_hi_16, res_hi_lo_hi_lo_16};
  wire [127:0]  res_hi_lo_16 = {res_hi_lo_hi_16, res_hi_lo_lo_16};
  wire [15:0]   res_hi_hi_lo_lo_lo_16 = {dataGroup_49_16, dataGroup_48_16};
  wire [15:0]   res_hi_hi_lo_lo_hi_16 = {dataGroup_51_16, dataGroup_50_16};
  wire [31:0]   res_hi_hi_lo_lo_16 = {res_hi_hi_lo_lo_hi_16, res_hi_hi_lo_lo_lo_16};
  wire [15:0]   res_hi_hi_lo_hi_lo_16 = {dataGroup_53_16, dataGroup_52_16};
  wire [15:0]   res_hi_hi_lo_hi_hi_16 = {dataGroup_55_16, dataGroup_54_16};
  wire [31:0]   res_hi_hi_lo_hi_16 = {res_hi_hi_lo_hi_hi_16, res_hi_hi_lo_hi_lo_16};
  wire [63:0]   res_hi_hi_lo_16 = {res_hi_hi_lo_hi_16, res_hi_hi_lo_lo_16};
  wire [15:0]   res_hi_hi_hi_lo_lo_16 = {dataGroup_57_16, dataGroup_56_16};
  wire [15:0]   res_hi_hi_hi_lo_hi_16 = {dataGroup_59_16, dataGroup_58_16};
  wire [31:0]   res_hi_hi_hi_lo_16 = {res_hi_hi_hi_lo_hi_16, res_hi_hi_hi_lo_lo_16};
  wire [15:0]   res_hi_hi_hi_hi_lo_16 = {dataGroup_61_16, dataGroup_60_16};
  wire [15:0]   res_hi_hi_hi_hi_hi_16 = {dataGroup_63_16, dataGroup_62_16};
  wire [31:0]   res_hi_hi_hi_hi_16 = {res_hi_hi_hi_hi_hi_16, res_hi_hi_hi_hi_lo_16};
  wire [63:0]   res_hi_hi_hi_16 = {res_hi_hi_hi_hi_16, res_hi_hi_hi_lo_16};
  wire [127:0]  res_hi_hi_16 = {res_hi_hi_hi_16, res_hi_hi_lo_16};
  wire [255:0]  res_hi_16 = {res_hi_hi_16, res_hi_lo_16};
  wire [511:0]  res_41 = {res_hi_16, res_lo_16};
  wire [2047:0] dataGroup_lo_1088 = {dataGroup_lo_hi_1088, dataGroup_lo_lo_1088};
  wire [2047:0] dataGroup_hi_1088 = {dataGroup_hi_hi_1088, dataGroup_hi_lo_1088};
  wire [7:0]    dataGroup_0_17 = dataGroup_lo_1088[23:16];
  wire [2047:0] dataGroup_lo_1089 = {dataGroup_lo_hi_1089, dataGroup_lo_lo_1089};
  wire [2047:0] dataGroup_hi_1089 = {dataGroup_hi_hi_1089, dataGroup_hi_lo_1089};
  wire [7:0]    dataGroup_1_17 = dataGroup_lo_1089[71:64];
  wire [2047:0] dataGroup_lo_1090 = {dataGroup_lo_hi_1090, dataGroup_lo_lo_1090};
  wire [2047:0] dataGroup_hi_1090 = {dataGroup_hi_hi_1090, dataGroup_hi_lo_1090};
  wire [7:0]    dataGroup_2_17 = dataGroup_lo_1090[119:112];
  wire [2047:0] dataGroup_lo_1091 = {dataGroup_lo_hi_1091, dataGroup_lo_lo_1091};
  wire [2047:0] dataGroup_hi_1091 = {dataGroup_hi_hi_1091, dataGroup_hi_lo_1091};
  wire [7:0]    dataGroup_3_17 = dataGroup_lo_1091[167:160];
  wire [2047:0] dataGroup_lo_1092 = {dataGroup_lo_hi_1092, dataGroup_lo_lo_1092};
  wire [2047:0] dataGroup_hi_1092 = {dataGroup_hi_hi_1092, dataGroup_hi_lo_1092};
  wire [7:0]    dataGroup_4_17 = dataGroup_lo_1092[215:208];
  wire [2047:0] dataGroup_lo_1093 = {dataGroup_lo_hi_1093, dataGroup_lo_lo_1093};
  wire [2047:0] dataGroup_hi_1093 = {dataGroup_hi_hi_1093, dataGroup_hi_lo_1093};
  wire [7:0]    dataGroup_5_17 = dataGroup_lo_1093[263:256];
  wire [2047:0] dataGroup_lo_1094 = {dataGroup_lo_hi_1094, dataGroup_lo_lo_1094};
  wire [2047:0] dataGroup_hi_1094 = {dataGroup_hi_hi_1094, dataGroup_hi_lo_1094};
  wire [7:0]    dataGroup_6_17 = dataGroup_lo_1094[311:304];
  wire [2047:0] dataGroup_lo_1095 = {dataGroup_lo_hi_1095, dataGroup_lo_lo_1095};
  wire [2047:0] dataGroup_hi_1095 = {dataGroup_hi_hi_1095, dataGroup_hi_lo_1095};
  wire [7:0]    dataGroup_7_17 = dataGroup_lo_1095[359:352];
  wire [2047:0] dataGroup_lo_1096 = {dataGroup_lo_hi_1096, dataGroup_lo_lo_1096};
  wire [2047:0] dataGroup_hi_1096 = {dataGroup_hi_hi_1096, dataGroup_hi_lo_1096};
  wire [7:0]    dataGroup_8_17 = dataGroup_lo_1096[407:400];
  wire [2047:0] dataGroup_lo_1097 = {dataGroup_lo_hi_1097, dataGroup_lo_lo_1097};
  wire [2047:0] dataGroup_hi_1097 = {dataGroup_hi_hi_1097, dataGroup_hi_lo_1097};
  wire [7:0]    dataGroup_9_17 = dataGroup_lo_1097[455:448];
  wire [2047:0] dataGroup_lo_1098 = {dataGroup_lo_hi_1098, dataGroup_lo_lo_1098};
  wire [2047:0] dataGroup_hi_1098 = {dataGroup_hi_hi_1098, dataGroup_hi_lo_1098};
  wire [7:0]    dataGroup_10_17 = dataGroup_lo_1098[503:496];
  wire [2047:0] dataGroup_lo_1099 = {dataGroup_lo_hi_1099, dataGroup_lo_lo_1099};
  wire [2047:0] dataGroup_hi_1099 = {dataGroup_hi_hi_1099, dataGroup_hi_lo_1099};
  wire [7:0]    dataGroup_11_17 = dataGroup_lo_1099[551:544];
  wire [2047:0] dataGroup_lo_1100 = {dataGroup_lo_hi_1100, dataGroup_lo_lo_1100};
  wire [2047:0] dataGroup_hi_1100 = {dataGroup_hi_hi_1100, dataGroup_hi_lo_1100};
  wire [7:0]    dataGroup_12_17 = dataGroup_lo_1100[599:592];
  wire [2047:0] dataGroup_lo_1101 = {dataGroup_lo_hi_1101, dataGroup_lo_lo_1101};
  wire [2047:0] dataGroup_hi_1101 = {dataGroup_hi_hi_1101, dataGroup_hi_lo_1101};
  wire [7:0]    dataGroup_13_17 = dataGroup_lo_1101[647:640];
  wire [2047:0] dataGroup_lo_1102 = {dataGroup_lo_hi_1102, dataGroup_lo_lo_1102};
  wire [2047:0] dataGroup_hi_1102 = {dataGroup_hi_hi_1102, dataGroup_hi_lo_1102};
  wire [7:0]    dataGroup_14_17 = dataGroup_lo_1102[695:688];
  wire [2047:0] dataGroup_lo_1103 = {dataGroup_lo_hi_1103, dataGroup_lo_lo_1103};
  wire [2047:0] dataGroup_hi_1103 = {dataGroup_hi_hi_1103, dataGroup_hi_lo_1103};
  wire [7:0]    dataGroup_15_17 = dataGroup_lo_1103[743:736];
  wire [2047:0] dataGroup_lo_1104 = {dataGroup_lo_hi_1104, dataGroup_lo_lo_1104};
  wire [2047:0] dataGroup_hi_1104 = {dataGroup_hi_hi_1104, dataGroup_hi_lo_1104};
  wire [7:0]    dataGroup_16_17 = dataGroup_lo_1104[791:784];
  wire [2047:0] dataGroup_lo_1105 = {dataGroup_lo_hi_1105, dataGroup_lo_lo_1105};
  wire [2047:0] dataGroup_hi_1105 = {dataGroup_hi_hi_1105, dataGroup_hi_lo_1105};
  wire [7:0]    dataGroup_17_17 = dataGroup_lo_1105[839:832];
  wire [2047:0] dataGroup_lo_1106 = {dataGroup_lo_hi_1106, dataGroup_lo_lo_1106};
  wire [2047:0] dataGroup_hi_1106 = {dataGroup_hi_hi_1106, dataGroup_hi_lo_1106};
  wire [7:0]    dataGroup_18_17 = dataGroup_lo_1106[887:880];
  wire [2047:0] dataGroup_lo_1107 = {dataGroup_lo_hi_1107, dataGroup_lo_lo_1107};
  wire [2047:0] dataGroup_hi_1107 = {dataGroup_hi_hi_1107, dataGroup_hi_lo_1107};
  wire [7:0]    dataGroup_19_17 = dataGroup_lo_1107[935:928];
  wire [2047:0] dataGroup_lo_1108 = {dataGroup_lo_hi_1108, dataGroup_lo_lo_1108};
  wire [2047:0] dataGroup_hi_1108 = {dataGroup_hi_hi_1108, dataGroup_hi_lo_1108};
  wire [7:0]    dataGroup_20_17 = dataGroup_lo_1108[983:976];
  wire [2047:0] dataGroup_lo_1109 = {dataGroup_lo_hi_1109, dataGroup_lo_lo_1109};
  wire [2047:0] dataGroup_hi_1109 = {dataGroup_hi_hi_1109, dataGroup_hi_lo_1109};
  wire [7:0]    dataGroup_21_17 = dataGroup_lo_1109[1031:1024];
  wire [2047:0] dataGroup_lo_1110 = {dataGroup_lo_hi_1110, dataGroup_lo_lo_1110};
  wire [2047:0] dataGroup_hi_1110 = {dataGroup_hi_hi_1110, dataGroup_hi_lo_1110};
  wire [7:0]    dataGroup_22_17 = dataGroup_lo_1110[1079:1072];
  wire [2047:0] dataGroup_lo_1111 = {dataGroup_lo_hi_1111, dataGroup_lo_lo_1111};
  wire [2047:0] dataGroup_hi_1111 = {dataGroup_hi_hi_1111, dataGroup_hi_lo_1111};
  wire [7:0]    dataGroup_23_17 = dataGroup_lo_1111[1127:1120];
  wire [2047:0] dataGroup_lo_1112 = {dataGroup_lo_hi_1112, dataGroup_lo_lo_1112};
  wire [2047:0] dataGroup_hi_1112 = {dataGroup_hi_hi_1112, dataGroup_hi_lo_1112};
  wire [7:0]    dataGroup_24_17 = dataGroup_lo_1112[1175:1168];
  wire [2047:0] dataGroup_lo_1113 = {dataGroup_lo_hi_1113, dataGroup_lo_lo_1113};
  wire [2047:0] dataGroup_hi_1113 = {dataGroup_hi_hi_1113, dataGroup_hi_lo_1113};
  wire [7:0]    dataGroup_25_17 = dataGroup_lo_1113[1223:1216];
  wire [2047:0] dataGroup_lo_1114 = {dataGroup_lo_hi_1114, dataGroup_lo_lo_1114};
  wire [2047:0] dataGroup_hi_1114 = {dataGroup_hi_hi_1114, dataGroup_hi_lo_1114};
  wire [7:0]    dataGroup_26_17 = dataGroup_lo_1114[1271:1264];
  wire [2047:0] dataGroup_lo_1115 = {dataGroup_lo_hi_1115, dataGroup_lo_lo_1115};
  wire [2047:0] dataGroup_hi_1115 = {dataGroup_hi_hi_1115, dataGroup_hi_lo_1115};
  wire [7:0]    dataGroup_27_17 = dataGroup_lo_1115[1319:1312];
  wire [2047:0] dataGroup_lo_1116 = {dataGroup_lo_hi_1116, dataGroup_lo_lo_1116};
  wire [2047:0] dataGroup_hi_1116 = {dataGroup_hi_hi_1116, dataGroup_hi_lo_1116};
  wire [7:0]    dataGroup_28_17 = dataGroup_lo_1116[1367:1360];
  wire [2047:0] dataGroup_lo_1117 = {dataGroup_lo_hi_1117, dataGroup_lo_lo_1117};
  wire [2047:0] dataGroup_hi_1117 = {dataGroup_hi_hi_1117, dataGroup_hi_lo_1117};
  wire [7:0]    dataGroup_29_17 = dataGroup_lo_1117[1415:1408];
  wire [2047:0] dataGroup_lo_1118 = {dataGroup_lo_hi_1118, dataGroup_lo_lo_1118};
  wire [2047:0] dataGroup_hi_1118 = {dataGroup_hi_hi_1118, dataGroup_hi_lo_1118};
  wire [7:0]    dataGroup_30_17 = dataGroup_lo_1118[1463:1456];
  wire [2047:0] dataGroup_lo_1119 = {dataGroup_lo_hi_1119, dataGroup_lo_lo_1119};
  wire [2047:0] dataGroup_hi_1119 = {dataGroup_hi_hi_1119, dataGroup_hi_lo_1119};
  wire [7:0]    dataGroup_31_17 = dataGroup_lo_1119[1511:1504];
  wire [2047:0] dataGroup_lo_1120 = {dataGroup_lo_hi_1120, dataGroup_lo_lo_1120};
  wire [2047:0] dataGroup_hi_1120 = {dataGroup_hi_hi_1120, dataGroup_hi_lo_1120};
  wire [7:0]    dataGroup_32_17 = dataGroup_lo_1120[1559:1552];
  wire [2047:0] dataGroup_lo_1121 = {dataGroup_lo_hi_1121, dataGroup_lo_lo_1121};
  wire [2047:0] dataGroup_hi_1121 = {dataGroup_hi_hi_1121, dataGroup_hi_lo_1121};
  wire [7:0]    dataGroup_33_17 = dataGroup_lo_1121[1607:1600];
  wire [2047:0] dataGroup_lo_1122 = {dataGroup_lo_hi_1122, dataGroup_lo_lo_1122};
  wire [2047:0] dataGroup_hi_1122 = {dataGroup_hi_hi_1122, dataGroup_hi_lo_1122};
  wire [7:0]    dataGroup_34_17 = dataGroup_lo_1122[1655:1648];
  wire [2047:0] dataGroup_lo_1123 = {dataGroup_lo_hi_1123, dataGroup_lo_lo_1123};
  wire [2047:0] dataGroup_hi_1123 = {dataGroup_hi_hi_1123, dataGroup_hi_lo_1123};
  wire [7:0]    dataGroup_35_17 = dataGroup_lo_1123[1703:1696];
  wire [2047:0] dataGroup_lo_1124 = {dataGroup_lo_hi_1124, dataGroup_lo_lo_1124};
  wire [2047:0] dataGroup_hi_1124 = {dataGroup_hi_hi_1124, dataGroup_hi_lo_1124};
  wire [7:0]    dataGroup_36_17 = dataGroup_lo_1124[1751:1744];
  wire [2047:0] dataGroup_lo_1125 = {dataGroup_lo_hi_1125, dataGroup_lo_lo_1125};
  wire [2047:0] dataGroup_hi_1125 = {dataGroup_hi_hi_1125, dataGroup_hi_lo_1125};
  wire [7:0]    dataGroup_37_17 = dataGroup_lo_1125[1799:1792];
  wire [2047:0] dataGroup_lo_1126 = {dataGroup_lo_hi_1126, dataGroup_lo_lo_1126};
  wire [2047:0] dataGroup_hi_1126 = {dataGroup_hi_hi_1126, dataGroup_hi_lo_1126};
  wire [7:0]    dataGroup_38_17 = dataGroup_lo_1126[1847:1840];
  wire [2047:0] dataGroup_lo_1127 = {dataGroup_lo_hi_1127, dataGroup_lo_lo_1127};
  wire [2047:0] dataGroup_hi_1127 = {dataGroup_hi_hi_1127, dataGroup_hi_lo_1127};
  wire [7:0]    dataGroup_39_17 = dataGroup_lo_1127[1895:1888];
  wire [2047:0] dataGroup_lo_1128 = {dataGroup_lo_hi_1128, dataGroup_lo_lo_1128};
  wire [2047:0] dataGroup_hi_1128 = {dataGroup_hi_hi_1128, dataGroup_hi_lo_1128};
  wire [7:0]    dataGroup_40_17 = dataGroup_lo_1128[1943:1936];
  wire [2047:0] dataGroup_lo_1129 = {dataGroup_lo_hi_1129, dataGroup_lo_lo_1129};
  wire [2047:0] dataGroup_hi_1129 = {dataGroup_hi_hi_1129, dataGroup_hi_lo_1129};
  wire [7:0]    dataGroup_41_17 = dataGroup_lo_1129[1991:1984];
  wire [2047:0] dataGroup_lo_1130 = {dataGroup_lo_hi_1130, dataGroup_lo_lo_1130};
  wire [2047:0] dataGroup_hi_1130 = {dataGroup_hi_hi_1130, dataGroup_hi_lo_1130};
  wire [7:0]    dataGroup_42_17 = dataGroup_lo_1130[2039:2032];
  wire [2047:0] dataGroup_lo_1131 = {dataGroup_lo_hi_1131, dataGroup_lo_lo_1131};
  wire [2047:0] dataGroup_hi_1131 = {dataGroup_hi_hi_1131, dataGroup_hi_lo_1131};
  wire [7:0]    dataGroup_43_17 = dataGroup_hi_1131[39:32];
  wire [2047:0] dataGroup_lo_1132 = {dataGroup_lo_hi_1132, dataGroup_lo_lo_1132};
  wire [2047:0] dataGroup_hi_1132 = {dataGroup_hi_hi_1132, dataGroup_hi_lo_1132};
  wire [7:0]    dataGroup_44_17 = dataGroup_hi_1132[87:80];
  wire [2047:0] dataGroup_lo_1133 = {dataGroup_lo_hi_1133, dataGroup_lo_lo_1133};
  wire [2047:0] dataGroup_hi_1133 = {dataGroup_hi_hi_1133, dataGroup_hi_lo_1133};
  wire [7:0]    dataGroup_45_17 = dataGroup_hi_1133[135:128];
  wire [2047:0] dataGroup_lo_1134 = {dataGroup_lo_hi_1134, dataGroup_lo_lo_1134};
  wire [2047:0] dataGroup_hi_1134 = {dataGroup_hi_hi_1134, dataGroup_hi_lo_1134};
  wire [7:0]    dataGroup_46_17 = dataGroup_hi_1134[183:176];
  wire [2047:0] dataGroup_lo_1135 = {dataGroup_lo_hi_1135, dataGroup_lo_lo_1135};
  wire [2047:0] dataGroup_hi_1135 = {dataGroup_hi_hi_1135, dataGroup_hi_lo_1135};
  wire [7:0]    dataGroup_47_17 = dataGroup_hi_1135[231:224];
  wire [2047:0] dataGroup_lo_1136 = {dataGroup_lo_hi_1136, dataGroup_lo_lo_1136};
  wire [2047:0] dataGroup_hi_1136 = {dataGroup_hi_hi_1136, dataGroup_hi_lo_1136};
  wire [7:0]    dataGroup_48_17 = dataGroup_hi_1136[279:272];
  wire [2047:0] dataGroup_lo_1137 = {dataGroup_lo_hi_1137, dataGroup_lo_lo_1137};
  wire [2047:0] dataGroup_hi_1137 = {dataGroup_hi_hi_1137, dataGroup_hi_lo_1137};
  wire [7:0]    dataGroup_49_17 = dataGroup_hi_1137[327:320];
  wire [2047:0] dataGroup_lo_1138 = {dataGroup_lo_hi_1138, dataGroup_lo_lo_1138};
  wire [2047:0] dataGroup_hi_1138 = {dataGroup_hi_hi_1138, dataGroup_hi_lo_1138};
  wire [7:0]    dataGroup_50_17 = dataGroup_hi_1138[375:368];
  wire [2047:0] dataGroup_lo_1139 = {dataGroup_lo_hi_1139, dataGroup_lo_lo_1139};
  wire [2047:0] dataGroup_hi_1139 = {dataGroup_hi_hi_1139, dataGroup_hi_lo_1139};
  wire [7:0]    dataGroup_51_17 = dataGroup_hi_1139[423:416];
  wire [2047:0] dataGroup_lo_1140 = {dataGroup_lo_hi_1140, dataGroup_lo_lo_1140};
  wire [2047:0] dataGroup_hi_1140 = {dataGroup_hi_hi_1140, dataGroup_hi_lo_1140};
  wire [7:0]    dataGroup_52_17 = dataGroup_hi_1140[471:464];
  wire [2047:0] dataGroup_lo_1141 = {dataGroup_lo_hi_1141, dataGroup_lo_lo_1141};
  wire [2047:0] dataGroup_hi_1141 = {dataGroup_hi_hi_1141, dataGroup_hi_lo_1141};
  wire [7:0]    dataGroup_53_17 = dataGroup_hi_1141[519:512];
  wire [2047:0] dataGroup_lo_1142 = {dataGroup_lo_hi_1142, dataGroup_lo_lo_1142};
  wire [2047:0] dataGroup_hi_1142 = {dataGroup_hi_hi_1142, dataGroup_hi_lo_1142};
  wire [7:0]    dataGroup_54_17 = dataGroup_hi_1142[567:560];
  wire [2047:0] dataGroup_lo_1143 = {dataGroup_lo_hi_1143, dataGroup_lo_lo_1143};
  wire [2047:0] dataGroup_hi_1143 = {dataGroup_hi_hi_1143, dataGroup_hi_lo_1143};
  wire [7:0]    dataGroup_55_17 = dataGroup_hi_1143[615:608];
  wire [2047:0] dataGroup_lo_1144 = {dataGroup_lo_hi_1144, dataGroup_lo_lo_1144};
  wire [2047:0] dataGroup_hi_1144 = {dataGroup_hi_hi_1144, dataGroup_hi_lo_1144};
  wire [7:0]    dataGroup_56_17 = dataGroup_hi_1144[663:656];
  wire [2047:0] dataGroup_lo_1145 = {dataGroup_lo_hi_1145, dataGroup_lo_lo_1145};
  wire [2047:0] dataGroup_hi_1145 = {dataGroup_hi_hi_1145, dataGroup_hi_lo_1145};
  wire [7:0]    dataGroup_57_17 = dataGroup_hi_1145[711:704];
  wire [2047:0] dataGroup_lo_1146 = {dataGroup_lo_hi_1146, dataGroup_lo_lo_1146};
  wire [2047:0] dataGroup_hi_1146 = {dataGroup_hi_hi_1146, dataGroup_hi_lo_1146};
  wire [7:0]    dataGroup_58_17 = dataGroup_hi_1146[759:752];
  wire [2047:0] dataGroup_lo_1147 = {dataGroup_lo_hi_1147, dataGroup_lo_lo_1147};
  wire [2047:0] dataGroup_hi_1147 = {dataGroup_hi_hi_1147, dataGroup_hi_lo_1147};
  wire [7:0]    dataGroup_59_17 = dataGroup_hi_1147[807:800];
  wire [2047:0] dataGroup_lo_1148 = {dataGroup_lo_hi_1148, dataGroup_lo_lo_1148};
  wire [2047:0] dataGroup_hi_1148 = {dataGroup_hi_hi_1148, dataGroup_hi_lo_1148};
  wire [7:0]    dataGroup_60_17 = dataGroup_hi_1148[855:848];
  wire [2047:0] dataGroup_lo_1149 = {dataGroup_lo_hi_1149, dataGroup_lo_lo_1149};
  wire [2047:0] dataGroup_hi_1149 = {dataGroup_hi_hi_1149, dataGroup_hi_lo_1149};
  wire [7:0]    dataGroup_61_17 = dataGroup_hi_1149[903:896];
  wire [2047:0] dataGroup_lo_1150 = {dataGroup_lo_hi_1150, dataGroup_lo_lo_1150};
  wire [2047:0] dataGroup_hi_1150 = {dataGroup_hi_hi_1150, dataGroup_hi_lo_1150};
  wire [7:0]    dataGroup_62_17 = dataGroup_hi_1150[951:944];
  wire [2047:0] dataGroup_lo_1151 = {dataGroup_lo_hi_1151, dataGroup_lo_lo_1151};
  wire [2047:0] dataGroup_hi_1151 = {dataGroup_hi_hi_1151, dataGroup_hi_lo_1151};
  wire [7:0]    dataGroup_63_17 = dataGroup_hi_1151[999:992];
  wire [15:0]   res_lo_lo_lo_lo_lo_17 = {dataGroup_1_17, dataGroup_0_17};
  wire [15:0]   res_lo_lo_lo_lo_hi_17 = {dataGroup_3_17, dataGroup_2_17};
  wire [31:0]   res_lo_lo_lo_lo_17 = {res_lo_lo_lo_lo_hi_17, res_lo_lo_lo_lo_lo_17};
  wire [15:0]   res_lo_lo_lo_hi_lo_17 = {dataGroup_5_17, dataGroup_4_17};
  wire [15:0]   res_lo_lo_lo_hi_hi_17 = {dataGroup_7_17, dataGroup_6_17};
  wire [31:0]   res_lo_lo_lo_hi_17 = {res_lo_lo_lo_hi_hi_17, res_lo_lo_lo_hi_lo_17};
  wire [63:0]   res_lo_lo_lo_17 = {res_lo_lo_lo_hi_17, res_lo_lo_lo_lo_17};
  wire [15:0]   res_lo_lo_hi_lo_lo_17 = {dataGroup_9_17, dataGroup_8_17};
  wire [15:0]   res_lo_lo_hi_lo_hi_17 = {dataGroup_11_17, dataGroup_10_17};
  wire [31:0]   res_lo_lo_hi_lo_17 = {res_lo_lo_hi_lo_hi_17, res_lo_lo_hi_lo_lo_17};
  wire [15:0]   res_lo_lo_hi_hi_lo_17 = {dataGroup_13_17, dataGroup_12_17};
  wire [15:0]   res_lo_lo_hi_hi_hi_17 = {dataGroup_15_17, dataGroup_14_17};
  wire [31:0]   res_lo_lo_hi_hi_17 = {res_lo_lo_hi_hi_hi_17, res_lo_lo_hi_hi_lo_17};
  wire [63:0]   res_lo_lo_hi_17 = {res_lo_lo_hi_hi_17, res_lo_lo_hi_lo_17};
  wire [127:0]  res_lo_lo_17 = {res_lo_lo_hi_17, res_lo_lo_lo_17};
  wire [15:0]   res_lo_hi_lo_lo_lo_17 = {dataGroup_17_17, dataGroup_16_17};
  wire [15:0]   res_lo_hi_lo_lo_hi_17 = {dataGroup_19_17, dataGroup_18_17};
  wire [31:0]   res_lo_hi_lo_lo_17 = {res_lo_hi_lo_lo_hi_17, res_lo_hi_lo_lo_lo_17};
  wire [15:0]   res_lo_hi_lo_hi_lo_17 = {dataGroup_21_17, dataGroup_20_17};
  wire [15:0]   res_lo_hi_lo_hi_hi_17 = {dataGroup_23_17, dataGroup_22_17};
  wire [31:0]   res_lo_hi_lo_hi_17 = {res_lo_hi_lo_hi_hi_17, res_lo_hi_lo_hi_lo_17};
  wire [63:0]   res_lo_hi_lo_17 = {res_lo_hi_lo_hi_17, res_lo_hi_lo_lo_17};
  wire [15:0]   res_lo_hi_hi_lo_lo_17 = {dataGroup_25_17, dataGroup_24_17};
  wire [15:0]   res_lo_hi_hi_lo_hi_17 = {dataGroup_27_17, dataGroup_26_17};
  wire [31:0]   res_lo_hi_hi_lo_17 = {res_lo_hi_hi_lo_hi_17, res_lo_hi_hi_lo_lo_17};
  wire [15:0]   res_lo_hi_hi_hi_lo_17 = {dataGroup_29_17, dataGroup_28_17};
  wire [15:0]   res_lo_hi_hi_hi_hi_17 = {dataGroup_31_17, dataGroup_30_17};
  wire [31:0]   res_lo_hi_hi_hi_17 = {res_lo_hi_hi_hi_hi_17, res_lo_hi_hi_hi_lo_17};
  wire [63:0]   res_lo_hi_hi_17 = {res_lo_hi_hi_hi_17, res_lo_hi_hi_lo_17};
  wire [127:0]  res_lo_hi_17 = {res_lo_hi_hi_17, res_lo_hi_lo_17};
  wire [255:0]  res_lo_17 = {res_lo_hi_17, res_lo_lo_17};
  wire [15:0]   res_hi_lo_lo_lo_lo_17 = {dataGroup_33_17, dataGroup_32_17};
  wire [15:0]   res_hi_lo_lo_lo_hi_17 = {dataGroup_35_17, dataGroup_34_17};
  wire [31:0]   res_hi_lo_lo_lo_17 = {res_hi_lo_lo_lo_hi_17, res_hi_lo_lo_lo_lo_17};
  wire [15:0]   res_hi_lo_lo_hi_lo_17 = {dataGroup_37_17, dataGroup_36_17};
  wire [15:0]   res_hi_lo_lo_hi_hi_17 = {dataGroup_39_17, dataGroup_38_17};
  wire [31:0]   res_hi_lo_lo_hi_17 = {res_hi_lo_lo_hi_hi_17, res_hi_lo_lo_hi_lo_17};
  wire [63:0]   res_hi_lo_lo_17 = {res_hi_lo_lo_hi_17, res_hi_lo_lo_lo_17};
  wire [15:0]   res_hi_lo_hi_lo_lo_17 = {dataGroup_41_17, dataGroup_40_17};
  wire [15:0]   res_hi_lo_hi_lo_hi_17 = {dataGroup_43_17, dataGroup_42_17};
  wire [31:0]   res_hi_lo_hi_lo_17 = {res_hi_lo_hi_lo_hi_17, res_hi_lo_hi_lo_lo_17};
  wire [15:0]   res_hi_lo_hi_hi_lo_17 = {dataGroup_45_17, dataGroup_44_17};
  wire [15:0]   res_hi_lo_hi_hi_hi_17 = {dataGroup_47_17, dataGroup_46_17};
  wire [31:0]   res_hi_lo_hi_hi_17 = {res_hi_lo_hi_hi_hi_17, res_hi_lo_hi_hi_lo_17};
  wire [63:0]   res_hi_lo_hi_17 = {res_hi_lo_hi_hi_17, res_hi_lo_hi_lo_17};
  wire [127:0]  res_hi_lo_17 = {res_hi_lo_hi_17, res_hi_lo_lo_17};
  wire [15:0]   res_hi_hi_lo_lo_lo_17 = {dataGroup_49_17, dataGroup_48_17};
  wire [15:0]   res_hi_hi_lo_lo_hi_17 = {dataGroup_51_17, dataGroup_50_17};
  wire [31:0]   res_hi_hi_lo_lo_17 = {res_hi_hi_lo_lo_hi_17, res_hi_hi_lo_lo_lo_17};
  wire [15:0]   res_hi_hi_lo_hi_lo_17 = {dataGroup_53_17, dataGroup_52_17};
  wire [15:0]   res_hi_hi_lo_hi_hi_17 = {dataGroup_55_17, dataGroup_54_17};
  wire [31:0]   res_hi_hi_lo_hi_17 = {res_hi_hi_lo_hi_hi_17, res_hi_hi_lo_hi_lo_17};
  wire [63:0]   res_hi_hi_lo_17 = {res_hi_hi_lo_hi_17, res_hi_hi_lo_lo_17};
  wire [15:0]   res_hi_hi_hi_lo_lo_17 = {dataGroup_57_17, dataGroup_56_17};
  wire [15:0]   res_hi_hi_hi_lo_hi_17 = {dataGroup_59_17, dataGroup_58_17};
  wire [31:0]   res_hi_hi_hi_lo_17 = {res_hi_hi_hi_lo_hi_17, res_hi_hi_hi_lo_lo_17};
  wire [15:0]   res_hi_hi_hi_hi_lo_17 = {dataGroup_61_17, dataGroup_60_17};
  wire [15:0]   res_hi_hi_hi_hi_hi_17 = {dataGroup_63_17, dataGroup_62_17};
  wire [31:0]   res_hi_hi_hi_hi_17 = {res_hi_hi_hi_hi_hi_17, res_hi_hi_hi_hi_lo_17};
  wire [63:0]   res_hi_hi_hi_17 = {res_hi_hi_hi_hi_17, res_hi_hi_hi_lo_17};
  wire [127:0]  res_hi_hi_17 = {res_hi_hi_hi_17, res_hi_hi_lo_17};
  wire [255:0]  res_hi_17 = {res_hi_hi_17, res_hi_lo_17};
  wire [511:0]  res_42 = {res_hi_17, res_lo_17};
  wire [2047:0] dataGroup_lo_1152 = {dataGroup_lo_hi_1152, dataGroup_lo_lo_1152};
  wire [2047:0] dataGroup_hi_1152 = {dataGroup_hi_hi_1152, dataGroup_hi_lo_1152};
  wire [7:0]    dataGroup_0_18 = dataGroup_lo_1152[31:24];
  wire [2047:0] dataGroup_lo_1153 = {dataGroup_lo_hi_1153, dataGroup_lo_lo_1153};
  wire [2047:0] dataGroup_hi_1153 = {dataGroup_hi_hi_1153, dataGroup_hi_lo_1153};
  wire [7:0]    dataGroup_1_18 = dataGroup_lo_1153[79:72];
  wire [2047:0] dataGroup_lo_1154 = {dataGroup_lo_hi_1154, dataGroup_lo_lo_1154};
  wire [2047:0] dataGroup_hi_1154 = {dataGroup_hi_hi_1154, dataGroup_hi_lo_1154};
  wire [7:0]    dataGroup_2_18 = dataGroup_lo_1154[127:120];
  wire [2047:0] dataGroup_lo_1155 = {dataGroup_lo_hi_1155, dataGroup_lo_lo_1155};
  wire [2047:0] dataGroup_hi_1155 = {dataGroup_hi_hi_1155, dataGroup_hi_lo_1155};
  wire [7:0]    dataGroup_3_18 = dataGroup_lo_1155[175:168];
  wire [2047:0] dataGroup_lo_1156 = {dataGroup_lo_hi_1156, dataGroup_lo_lo_1156};
  wire [2047:0] dataGroup_hi_1156 = {dataGroup_hi_hi_1156, dataGroup_hi_lo_1156};
  wire [7:0]    dataGroup_4_18 = dataGroup_lo_1156[223:216];
  wire [2047:0] dataGroup_lo_1157 = {dataGroup_lo_hi_1157, dataGroup_lo_lo_1157};
  wire [2047:0] dataGroup_hi_1157 = {dataGroup_hi_hi_1157, dataGroup_hi_lo_1157};
  wire [7:0]    dataGroup_5_18 = dataGroup_lo_1157[271:264];
  wire [2047:0] dataGroup_lo_1158 = {dataGroup_lo_hi_1158, dataGroup_lo_lo_1158};
  wire [2047:0] dataGroup_hi_1158 = {dataGroup_hi_hi_1158, dataGroup_hi_lo_1158};
  wire [7:0]    dataGroup_6_18 = dataGroup_lo_1158[319:312];
  wire [2047:0] dataGroup_lo_1159 = {dataGroup_lo_hi_1159, dataGroup_lo_lo_1159};
  wire [2047:0] dataGroup_hi_1159 = {dataGroup_hi_hi_1159, dataGroup_hi_lo_1159};
  wire [7:0]    dataGroup_7_18 = dataGroup_lo_1159[367:360];
  wire [2047:0] dataGroup_lo_1160 = {dataGroup_lo_hi_1160, dataGroup_lo_lo_1160};
  wire [2047:0] dataGroup_hi_1160 = {dataGroup_hi_hi_1160, dataGroup_hi_lo_1160};
  wire [7:0]    dataGroup_8_18 = dataGroup_lo_1160[415:408];
  wire [2047:0] dataGroup_lo_1161 = {dataGroup_lo_hi_1161, dataGroup_lo_lo_1161};
  wire [2047:0] dataGroup_hi_1161 = {dataGroup_hi_hi_1161, dataGroup_hi_lo_1161};
  wire [7:0]    dataGroup_9_18 = dataGroup_lo_1161[463:456];
  wire [2047:0] dataGroup_lo_1162 = {dataGroup_lo_hi_1162, dataGroup_lo_lo_1162};
  wire [2047:0] dataGroup_hi_1162 = {dataGroup_hi_hi_1162, dataGroup_hi_lo_1162};
  wire [7:0]    dataGroup_10_18 = dataGroup_lo_1162[511:504];
  wire [2047:0] dataGroup_lo_1163 = {dataGroup_lo_hi_1163, dataGroup_lo_lo_1163};
  wire [2047:0] dataGroup_hi_1163 = {dataGroup_hi_hi_1163, dataGroup_hi_lo_1163};
  wire [7:0]    dataGroup_11_18 = dataGroup_lo_1163[559:552];
  wire [2047:0] dataGroup_lo_1164 = {dataGroup_lo_hi_1164, dataGroup_lo_lo_1164};
  wire [2047:0] dataGroup_hi_1164 = {dataGroup_hi_hi_1164, dataGroup_hi_lo_1164};
  wire [7:0]    dataGroup_12_18 = dataGroup_lo_1164[607:600];
  wire [2047:0] dataGroup_lo_1165 = {dataGroup_lo_hi_1165, dataGroup_lo_lo_1165};
  wire [2047:0] dataGroup_hi_1165 = {dataGroup_hi_hi_1165, dataGroup_hi_lo_1165};
  wire [7:0]    dataGroup_13_18 = dataGroup_lo_1165[655:648];
  wire [2047:0] dataGroup_lo_1166 = {dataGroup_lo_hi_1166, dataGroup_lo_lo_1166};
  wire [2047:0] dataGroup_hi_1166 = {dataGroup_hi_hi_1166, dataGroup_hi_lo_1166};
  wire [7:0]    dataGroup_14_18 = dataGroup_lo_1166[703:696];
  wire [2047:0] dataGroup_lo_1167 = {dataGroup_lo_hi_1167, dataGroup_lo_lo_1167};
  wire [2047:0] dataGroup_hi_1167 = {dataGroup_hi_hi_1167, dataGroup_hi_lo_1167};
  wire [7:0]    dataGroup_15_18 = dataGroup_lo_1167[751:744];
  wire [2047:0] dataGroup_lo_1168 = {dataGroup_lo_hi_1168, dataGroup_lo_lo_1168};
  wire [2047:0] dataGroup_hi_1168 = {dataGroup_hi_hi_1168, dataGroup_hi_lo_1168};
  wire [7:0]    dataGroup_16_18 = dataGroup_lo_1168[799:792];
  wire [2047:0] dataGroup_lo_1169 = {dataGroup_lo_hi_1169, dataGroup_lo_lo_1169};
  wire [2047:0] dataGroup_hi_1169 = {dataGroup_hi_hi_1169, dataGroup_hi_lo_1169};
  wire [7:0]    dataGroup_17_18 = dataGroup_lo_1169[847:840];
  wire [2047:0] dataGroup_lo_1170 = {dataGroup_lo_hi_1170, dataGroup_lo_lo_1170};
  wire [2047:0] dataGroup_hi_1170 = {dataGroup_hi_hi_1170, dataGroup_hi_lo_1170};
  wire [7:0]    dataGroup_18_18 = dataGroup_lo_1170[895:888];
  wire [2047:0] dataGroup_lo_1171 = {dataGroup_lo_hi_1171, dataGroup_lo_lo_1171};
  wire [2047:0] dataGroup_hi_1171 = {dataGroup_hi_hi_1171, dataGroup_hi_lo_1171};
  wire [7:0]    dataGroup_19_18 = dataGroup_lo_1171[943:936];
  wire [2047:0] dataGroup_lo_1172 = {dataGroup_lo_hi_1172, dataGroup_lo_lo_1172};
  wire [2047:0] dataGroup_hi_1172 = {dataGroup_hi_hi_1172, dataGroup_hi_lo_1172};
  wire [7:0]    dataGroup_20_18 = dataGroup_lo_1172[991:984];
  wire [2047:0] dataGroup_lo_1173 = {dataGroup_lo_hi_1173, dataGroup_lo_lo_1173};
  wire [2047:0] dataGroup_hi_1173 = {dataGroup_hi_hi_1173, dataGroup_hi_lo_1173};
  wire [7:0]    dataGroup_21_18 = dataGroup_lo_1173[1039:1032];
  wire [2047:0] dataGroup_lo_1174 = {dataGroup_lo_hi_1174, dataGroup_lo_lo_1174};
  wire [2047:0] dataGroup_hi_1174 = {dataGroup_hi_hi_1174, dataGroup_hi_lo_1174};
  wire [7:0]    dataGroup_22_18 = dataGroup_lo_1174[1087:1080];
  wire [2047:0] dataGroup_lo_1175 = {dataGroup_lo_hi_1175, dataGroup_lo_lo_1175};
  wire [2047:0] dataGroup_hi_1175 = {dataGroup_hi_hi_1175, dataGroup_hi_lo_1175};
  wire [7:0]    dataGroup_23_18 = dataGroup_lo_1175[1135:1128];
  wire [2047:0] dataGroup_lo_1176 = {dataGroup_lo_hi_1176, dataGroup_lo_lo_1176};
  wire [2047:0] dataGroup_hi_1176 = {dataGroup_hi_hi_1176, dataGroup_hi_lo_1176};
  wire [7:0]    dataGroup_24_18 = dataGroup_lo_1176[1183:1176];
  wire [2047:0] dataGroup_lo_1177 = {dataGroup_lo_hi_1177, dataGroup_lo_lo_1177};
  wire [2047:0] dataGroup_hi_1177 = {dataGroup_hi_hi_1177, dataGroup_hi_lo_1177};
  wire [7:0]    dataGroup_25_18 = dataGroup_lo_1177[1231:1224];
  wire [2047:0] dataGroup_lo_1178 = {dataGroup_lo_hi_1178, dataGroup_lo_lo_1178};
  wire [2047:0] dataGroup_hi_1178 = {dataGroup_hi_hi_1178, dataGroup_hi_lo_1178};
  wire [7:0]    dataGroup_26_18 = dataGroup_lo_1178[1279:1272];
  wire [2047:0] dataGroup_lo_1179 = {dataGroup_lo_hi_1179, dataGroup_lo_lo_1179};
  wire [2047:0] dataGroup_hi_1179 = {dataGroup_hi_hi_1179, dataGroup_hi_lo_1179};
  wire [7:0]    dataGroup_27_18 = dataGroup_lo_1179[1327:1320];
  wire [2047:0] dataGroup_lo_1180 = {dataGroup_lo_hi_1180, dataGroup_lo_lo_1180};
  wire [2047:0] dataGroup_hi_1180 = {dataGroup_hi_hi_1180, dataGroup_hi_lo_1180};
  wire [7:0]    dataGroup_28_18 = dataGroup_lo_1180[1375:1368];
  wire [2047:0] dataGroup_lo_1181 = {dataGroup_lo_hi_1181, dataGroup_lo_lo_1181};
  wire [2047:0] dataGroup_hi_1181 = {dataGroup_hi_hi_1181, dataGroup_hi_lo_1181};
  wire [7:0]    dataGroup_29_18 = dataGroup_lo_1181[1423:1416];
  wire [2047:0] dataGroup_lo_1182 = {dataGroup_lo_hi_1182, dataGroup_lo_lo_1182};
  wire [2047:0] dataGroup_hi_1182 = {dataGroup_hi_hi_1182, dataGroup_hi_lo_1182};
  wire [7:0]    dataGroup_30_18 = dataGroup_lo_1182[1471:1464];
  wire [2047:0] dataGroup_lo_1183 = {dataGroup_lo_hi_1183, dataGroup_lo_lo_1183};
  wire [2047:0] dataGroup_hi_1183 = {dataGroup_hi_hi_1183, dataGroup_hi_lo_1183};
  wire [7:0]    dataGroup_31_18 = dataGroup_lo_1183[1519:1512];
  wire [2047:0] dataGroup_lo_1184 = {dataGroup_lo_hi_1184, dataGroup_lo_lo_1184};
  wire [2047:0] dataGroup_hi_1184 = {dataGroup_hi_hi_1184, dataGroup_hi_lo_1184};
  wire [7:0]    dataGroup_32_18 = dataGroup_lo_1184[1567:1560];
  wire [2047:0] dataGroup_lo_1185 = {dataGroup_lo_hi_1185, dataGroup_lo_lo_1185};
  wire [2047:0] dataGroup_hi_1185 = {dataGroup_hi_hi_1185, dataGroup_hi_lo_1185};
  wire [7:0]    dataGroup_33_18 = dataGroup_lo_1185[1615:1608];
  wire [2047:0] dataGroup_lo_1186 = {dataGroup_lo_hi_1186, dataGroup_lo_lo_1186};
  wire [2047:0] dataGroup_hi_1186 = {dataGroup_hi_hi_1186, dataGroup_hi_lo_1186};
  wire [7:0]    dataGroup_34_18 = dataGroup_lo_1186[1663:1656];
  wire [2047:0] dataGroup_lo_1187 = {dataGroup_lo_hi_1187, dataGroup_lo_lo_1187};
  wire [2047:0] dataGroup_hi_1187 = {dataGroup_hi_hi_1187, dataGroup_hi_lo_1187};
  wire [7:0]    dataGroup_35_18 = dataGroup_lo_1187[1711:1704];
  wire [2047:0] dataGroup_lo_1188 = {dataGroup_lo_hi_1188, dataGroup_lo_lo_1188};
  wire [2047:0] dataGroup_hi_1188 = {dataGroup_hi_hi_1188, dataGroup_hi_lo_1188};
  wire [7:0]    dataGroup_36_18 = dataGroup_lo_1188[1759:1752];
  wire [2047:0] dataGroup_lo_1189 = {dataGroup_lo_hi_1189, dataGroup_lo_lo_1189};
  wire [2047:0] dataGroup_hi_1189 = {dataGroup_hi_hi_1189, dataGroup_hi_lo_1189};
  wire [7:0]    dataGroup_37_18 = dataGroup_lo_1189[1807:1800];
  wire [2047:0] dataGroup_lo_1190 = {dataGroup_lo_hi_1190, dataGroup_lo_lo_1190};
  wire [2047:0] dataGroup_hi_1190 = {dataGroup_hi_hi_1190, dataGroup_hi_lo_1190};
  wire [7:0]    dataGroup_38_18 = dataGroup_lo_1190[1855:1848];
  wire [2047:0] dataGroup_lo_1191 = {dataGroup_lo_hi_1191, dataGroup_lo_lo_1191};
  wire [2047:0] dataGroup_hi_1191 = {dataGroup_hi_hi_1191, dataGroup_hi_lo_1191};
  wire [7:0]    dataGroup_39_18 = dataGroup_lo_1191[1903:1896];
  wire [2047:0] dataGroup_lo_1192 = {dataGroup_lo_hi_1192, dataGroup_lo_lo_1192};
  wire [2047:0] dataGroup_hi_1192 = {dataGroup_hi_hi_1192, dataGroup_hi_lo_1192};
  wire [7:0]    dataGroup_40_18 = dataGroup_lo_1192[1951:1944];
  wire [2047:0] dataGroup_lo_1193 = {dataGroup_lo_hi_1193, dataGroup_lo_lo_1193};
  wire [2047:0] dataGroup_hi_1193 = {dataGroup_hi_hi_1193, dataGroup_hi_lo_1193};
  wire [7:0]    dataGroup_41_18 = dataGroup_lo_1193[1999:1992];
  wire [2047:0] dataGroup_lo_1194 = {dataGroup_lo_hi_1194, dataGroup_lo_lo_1194};
  wire [2047:0] dataGroup_hi_1194 = {dataGroup_hi_hi_1194, dataGroup_hi_lo_1194};
  wire [7:0]    dataGroup_42_18 = dataGroup_lo_1194[2047:2040];
  wire [2047:0] dataGroup_lo_1195 = {dataGroup_lo_hi_1195, dataGroup_lo_lo_1195};
  wire [2047:0] dataGroup_hi_1195 = {dataGroup_hi_hi_1195, dataGroup_hi_lo_1195};
  wire [7:0]    dataGroup_43_18 = dataGroup_hi_1195[47:40];
  wire [2047:0] dataGroup_lo_1196 = {dataGroup_lo_hi_1196, dataGroup_lo_lo_1196};
  wire [2047:0] dataGroup_hi_1196 = {dataGroup_hi_hi_1196, dataGroup_hi_lo_1196};
  wire [7:0]    dataGroup_44_18 = dataGroup_hi_1196[95:88];
  wire [2047:0] dataGroup_lo_1197 = {dataGroup_lo_hi_1197, dataGroup_lo_lo_1197};
  wire [2047:0] dataGroup_hi_1197 = {dataGroup_hi_hi_1197, dataGroup_hi_lo_1197};
  wire [7:0]    dataGroup_45_18 = dataGroup_hi_1197[143:136];
  wire [2047:0] dataGroup_lo_1198 = {dataGroup_lo_hi_1198, dataGroup_lo_lo_1198};
  wire [2047:0] dataGroup_hi_1198 = {dataGroup_hi_hi_1198, dataGroup_hi_lo_1198};
  wire [7:0]    dataGroup_46_18 = dataGroup_hi_1198[191:184];
  wire [2047:0] dataGroup_lo_1199 = {dataGroup_lo_hi_1199, dataGroup_lo_lo_1199};
  wire [2047:0] dataGroup_hi_1199 = {dataGroup_hi_hi_1199, dataGroup_hi_lo_1199};
  wire [7:0]    dataGroup_47_18 = dataGroup_hi_1199[239:232];
  wire [2047:0] dataGroup_lo_1200 = {dataGroup_lo_hi_1200, dataGroup_lo_lo_1200};
  wire [2047:0] dataGroup_hi_1200 = {dataGroup_hi_hi_1200, dataGroup_hi_lo_1200};
  wire [7:0]    dataGroup_48_18 = dataGroup_hi_1200[287:280];
  wire [2047:0] dataGroup_lo_1201 = {dataGroup_lo_hi_1201, dataGroup_lo_lo_1201};
  wire [2047:0] dataGroup_hi_1201 = {dataGroup_hi_hi_1201, dataGroup_hi_lo_1201};
  wire [7:0]    dataGroup_49_18 = dataGroup_hi_1201[335:328];
  wire [2047:0] dataGroup_lo_1202 = {dataGroup_lo_hi_1202, dataGroup_lo_lo_1202};
  wire [2047:0] dataGroup_hi_1202 = {dataGroup_hi_hi_1202, dataGroup_hi_lo_1202};
  wire [7:0]    dataGroup_50_18 = dataGroup_hi_1202[383:376];
  wire [2047:0] dataGroup_lo_1203 = {dataGroup_lo_hi_1203, dataGroup_lo_lo_1203};
  wire [2047:0] dataGroup_hi_1203 = {dataGroup_hi_hi_1203, dataGroup_hi_lo_1203};
  wire [7:0]    dataGroup_51_18 = dataGroup_hi_1203[431:424];
  wire [2047:0] dataGroup_lo_1204 = {dataGroup_lo_hi_1204, dataGroup_lo_lo_1204};
  wire [2047:0] dataGroup_hi_1204 = {dataGroup_hi_hi_1204, dataGroup_hi_lo_1204};
  wire [7:0]    dataGroup_52_18 = dataGroup_hi_1204[479:472];
  wire [2047:0] dataGroup_lo_1205 = {dataGroup_lo_hi_1205, dataGroup_lo_lo_1205};
  wire [2047:0] dataGroup_hi_1205 = {dataGroup_hi_hi_1205, dataGroup_hi_lo_1205};
  wire [7:0]    dataGroup_53_18 = dataGroup_hi_1205[527:520];
  wire [2047:0] dataGroup_lo_1206 = {dataGroup_lo_hi_1206, dataGroup_lo_lo_1206};
  wire [2047:0] dataGroup_hi_1206 = {dataGroup_hi_hi_1206, dataGroup_hi_lo_1206};
  wire [7:0]    dataGroup_54_18 = dataGroup_hi_1206[575:568];
  wire [2047:0] dataGroup_lo_1207 = {dataGroup_lo_hi_1207, dataGroup_lo_lo_1207};
  wire [2047:0] dataGroup_hi_1207 = {dataGroup_hi_hi_1207, dataGroup_hi_lo_1207};
  wire [7:0]    dataGroup_55_18 = dataGroup_hi_1207[623:616];
  wire [2047:0] dataGroup_lo_1208 = {dataGroup_lo_hi_1208, dataGroup_lo_lo_1208};
  wire [2047:0] dataGroup_hi_1208 = {dataGroup_hi_hi_1208, dataGroup_hi_lo_1208};
  wire [7:0]    dataGroup_56_18 = dataGroup_hi_1208[671:664];
  wire [2047:0] dataGroup_lo_1209 = {dataGroup_lo_hi_1209, dataGroup_lo_lo_1209};
  wire [2047:0] dataGroup_hi_1209 = {dataGroup_hi_hi_1209, dataGroup_hi_lo_1209};
  wire [7:0]    dataGroup_57_18 = dataGroup_hi_1209[719:712];
  wire [2047:0] dataGroup_lo_1210 = {dataGroup_lo_hi_1210, dataGroup_lo_lo_1210};
  wire [2047:0] dataGroup_hi_1210 = {dataGroup_hi_hi_1210, dataGroup_hi_lo_1210};
  wire [7:0]    dataGroup_58_18 = dataGroup_hi_1210[767:760];
  wire [2047:0] dataGroup_lo_1211 = {dataGroup_lo_hi_1211, dataGroup_lo_lo_1211};
  wire [2047:0] dataGroup_hi_1211 = {dataGroup_hi_hi_1211, dataGroup_hi_lo_1211};
  wire [7:0]    dataGroup_59_18 = dataGroup_hi_1211[815:808];
  wire [2047:0] dataGroup_lo_1212 = {dataGroup_lo_hi_1212, dataGroup_lo_lo_1212};
  wire [2047:0] dataGroup_hi_1212 = {dataGroup_hi_hi_1212, dataGroup_hi_lo_1212};
  wire [7:0]    dataGroup_60_18 = dataGroup_hi_1212[863:856];
  wire [2047:0] dataGroup_lo_1213 = {dataGroup_lo_hi_1213, dataGroup_lo_lo_1213};
  wire [2047:0] dataGroup_hi_1213 = {dataGroup_hi_hi_1213, dataGroup_hi_lo_1213};
  wire [7:0]    dataGroup_61_18 = dataGroup_hi_1213[911:904];
  wire [2047:0] dataGroup_lo_1214 = {dataGroup_lo_hi_1214, dataGroup_lo_lo_1214};
  wire [2047:0] dataGroup_hi_1214 = {dataGroup_hi_hi_1214, dataGroup_hi_lo_1214};
  wire [7:0]    dataGroup_62_18 = dataGroup_hi_1214[959:952];
  wire [2047:0] dataGroup_lo_1215 = {dataGroup_lo_hi_1215, dataGroup_lo_lo_1215};
  wire [2047:0] dataGroup_hi_1215 = {dataGroup_hi_hi_1215, dataGroup_hi_lo_1215};
  wire [7:0]    dataGroup_63_18 = dataGroup_hi_1215[1007:1000];
  wire [15:0]   res_lo_lo_lo_lo_lo_18 = {dataGroup_1_18, dataGroup_0_18};
  wire [15:0]   res_lo_lo_lo_lo_hi_18 = {dataGroup_3_18, dataGroup_2_18};
  wire [31:0]   res_lo_lo_lo_lo_18 = {res_lo_lo_lo_lo_hi_18, res_lo_lo_lo_lo_lo_18};
  wire [15:0]   res_lo_lo_lo_hi_lo_18 = {dataGroup_5_18, dataGroup_4_18};
  wire [15:0]   res_lo_lo_lo_hi_hi_18 = {dataGroup_7_18, dataGroup_6_18};
  wire [31:0]   res_lo_lo_lo_hi_18 = {res_lo_lo_lo_hi_hi_18, res_lo_lo_lo_hi_lo_18};
  wire [63:0]   res_lo_lo_lo_18 = {res_lo_lo_lo_hi_18, res_lo_lo_lo_lo_18};
  wire [15:0]   res_lo_lo_hi_lo_lo_18 = {dataGroup_9_18, dataGroup_8_18};
  wire [15:0]   res_lo_lo_hi_lo_hi_18 = {dataGroup_11_18, dataGroup_10_18};
  wire [31:0]   res_lo_lo_hi_lo_18 = {res_lo_lo_hi_lo_hi_18, res_lo_lo_hi_lo_lo_18};
  wire [15:0]   res_lo_lo_hi_hi_lo_18 = {dataGroup_13_18, dataGroup_12_18};
  wire [15:0]   res_lo_lo_hi_hi_hi_18 = {dataGroup_15_18, dataGroup_14_18};
  wire [31:0]   res_lo_lo_hi_hi_18 = {res_lo_lo_hi_hi_hi_18, res_lo_lo_hi_hi_lo_18};
  wire [63:0]   res_lo_lo_hi_18 = {res_lo_lo_hi_hi_18, res_lo_lo_hi_lo_18};
  wire [127:0]  res_lo_lo_18 = {res_lo_lo_hi_18, res_lo_lo_lo_18};
  wire [15:0]   res_lo_hi_lo_lo_lo_18 = {dataGroup_17_18, dataGroup_16_18};
  wire [15:0]   res_lo_hi_lo_lo_hi_18 = {dataGroup_19_18, dataGroup_18_18};
  wire [31:0]   res_lo_hi_lo_lo_18 = {res_lo_hi_lo_lo_hi_18, res_lo_hi_lo_lo_lo_18};
  wire [15:0]   res_lo_hi_lo_hi_lo_18 = {dataGroup_21_18, dataGroup_20_18};
  wire [15:0]   res_lo_hi_lo_hi_hi_18 = {dataGroup_23_18, dataGroup_22_18};
  wire [31:0]   res_lo_hi_lo_hi_18 = {res_lo_hi_lo_hi_hi_18, res_lo_hi_lo_hi_lo_18};
  wire [63:0]   res_lo_hi_lo_18 = {res_lo_hi_lo_hi_18, res_lo_hi_lo_lo_18};
  wire [15:0]   res_lo_hi_hi_lo_lo_18 = {dataGroup_25_18, dataGroup_24_18};
  wire [15:0]   res_lo_hi_hi_lo_hi_18 = {dataGroup_27_18, dataGroup_26_18};
  wire [31:0]   res_lo_hi_hi_lo_18 = {res_lo_hi_hi_lo_hi_18, res_lo_hi_hi_lo_lo_18};
  wire [15:0]   res_lo_hi_hi_hi_lo_18 = {dataGroup_29_18, dataGroup_28_18};
  wire [15:0]   res_lo_hi_hi_hi_hi_18 = {dataGroup_31_18, dataGroup_30_18};
  wire [31:0]   res_lo_hi_hi_hi_18 = {res_lo_hi_hi_hi_hi_18, res_lo_hi_hi_hi_lo_18};
  wire [63:0]   res_lo_hi_hi_18 = {res_lo_hi_hi_hi_18, res_lo_hi_hi_lo_18};
  wire [127:0]  res_lo_hi_18 = {res_lo_hi_hi_18, res_lo_hi_lo_18};
  wire [255:0]  res_lo_18 = {res_lo_hi_18, res_lo_lo_18};
  wire [15:0]   res_hi_lo_lo_lo_lo_18 = {dataGroup_33_18, dataGroup_32_18};
  wire [15:0]   res_hi_lo_lo_lo_hi_18 = {dataGroup_35_18, dataGroup_34_18};
  wire [31:0]   res_hi_lo_lo_lo_18 = {res_hi_lo_lo_lo_hi_18, res_hi_lo_lo_lo_lo_18};
  wire [15:0]   res_hi_lo_lo_hi_lo_18 = {dataGroup_37_18, dataGroup_36_18};
  wire [15:0]   res_hi_lo_lo_hi_hi_18 = {dataGroup_39_18, dataGroup_38_18};
  wire [31:0]   res_hi_lo_lo_hi_18 = {res_hi_lo_lo_hi_hi_18, res_hi_lo_lo_hi_lo_18};
  wire [63:0]   res_hi_lo_lo_18 = {res_hi_lo_lo_hi_18, res_hi_lo_lo_lo_18};
  wire [15:0]   res_hi_lo_hi_lo_lo_18 = {dataGroup_41_18, dataGroup_40_18};
  wire [15:0]   res_hi_lo_hi_lo_hi_18 = {dataGroup_43_18, dataGroup_42_18};
  wire [31:0]   res_hi_lo_hi_lo_18 = {res_hi_lo_hi_lo_hi_18, res_hi_lo_hi_lo_lo_18};
  wire [15:0]   res_hi_lo_hi_hi_lo_18 = {dataGroup_45_18, dataGroup_44_18};
  wire [15:0]   res_hi_lo_hi_hi_hi_18 = {dataGroup_47_18, dataGroup_46_18};
  wire [31:0]   res_hi_lo_hi_hi_18 = {res_hi_lo_hi_hi_hi_18, res_hi_lo_hi_hi_lo_18};
  wire [63:0]   res_hi_lo_hi_18 = {res_hi_lo_hi_hi_18, res_hi_lo_hi_lo_18};
  wire [127:0]  res_hi_lo_18 = {res_hi_lo_hi_18, res_hi_lo_lo_18};
  wire [15:0]   res_hi_hi_lo_lo_lo_18 = {dataGroup_49_18, dataGroup_48_18};
  wire [15:0]   res_hi_hi_lo_lo_hi_18 = {dataGroup_51_18, dataGroup_50_18};
  wire [31:0]   res_hi_hi_lo_lo_18 = {res_hi_hi_lo_lo_hi_18, res_hi_hi_lo_lo_lo_18};
  wire [15:0]   res_hi_hi_lo_hi_lo_18 = {dataGroup_53_18, dataGroup_52_18};
  wire [15:0]   res_hi_hi_lo_hi_hi_18 = {dataGroup_55_18, dataGroup_54_18};
  wire [31:0]   res_hi_hi_lo_hi_18 = {res_hi_hi_lo_hi_hi_18, res_hi_hi_lo_hi_lo_18};
  wire [63:0]   res_hi_hi_lo_18 = {res_hi_hi_lo_hi_18, res_hi_hi_lo_lo_18};
  wire [15:0]   res_hi_hi_hi_lo_lo_18 = {dataGroup_57_18, dataGroup_56_18};
  wire [15:0]   res_hi_hi_hi_lo_hi_18 = {dataGroup_59_18, dataGroup_58_18};
  wire [31:0]   res_hi_hi_hi_lo_18 = {res_hi_hi_hi_lo_hi_18, res_hi_hi_hi_lo_lo_18};
  wire [15:0]   res_hi_hi_hi_hi_lo_18 = {dataGroup_61_18, dataGroup_60_18};
  wire [15:0]   res_hi_hi_hi_hi_hi_18 = {dataGroup_63_18, dataGroup_62_18};
  wire [31:0]   res_hi_hi_hi_hi_18 = {res_hi_hi_hi_hi_hi_18, res_hi_hi_hi_hi_lo_18};
  wire [63:0]   res_hi_hi_hi_18 = {res_hi_hi_hi_hi_18, res_hi_hi_hi_lo_18};
  wire [127:0]  res_hi_hi_18 = {res_hi_hi_hi_18, res_hi_hi_lo_18};
  wire [255:0]  res_hi_18 = {res_hi_hi_18, res_hi_lo_18};
  wire [511:0]  res_43 = {res_hi_18, res_lo_18};
  wire [2047:0] dataGroup_lo_1216 = {dataGroup_lo_hi_1216, dataGroup_lo_lo_1216};
  wire [2047:0] dataGroup_hi_1216 = {dataGroup_hi_hi_1216, dataGroup_hi_lo_1216};
  wire [7:0]    dataGroup_0_19 = dataGroup_lo_1216[39:32];
  wire [2047:0] dataGroup_lo_1217 = {dataGroup_lo_hi_1217, dataGroup_lo_lo_1217};
  wire [2047:0] dataGroup_hi_1217 = {dataGroup_hi_hi_1217, dataGroup_hi_lo_1217};
  wire [7:0]    dataGroup_1_19 = dataGroup_lo_1217[87:80];
  wire [2047:0] dataGroup_lo_1218 = {dataGroup_lo_hi_1218, dataGroup_lo_lo_1218};
  wire [2047:0] dataGroup_hi_1218 = {dataGroup_hi_hi_1218, dataGroup_hi_lo_1218};
  wire [7:0]    dataGroup_2_19 = dataGroup_lo_1218[135:128];
  wire [2047:0] dataGroup_lo_1219 = {dataGroup_lo_hi_1219, dataGroup_lo_lo_1219};
  wire [2047:0] dataGroup_hi_1219 = {dataGroup_hi_hi_1219, dataGroup_hi_lo_1219};
  wire [7:0]    dataGroup_3_19 = dataGroup_lo_1219[183:176];
  wire [2047:0] dataGroup_lo_1220 = {dataGroup_lo_hi_1220, dataGroup_lo_lo_1220};
  wire [2047:0] dataGroup_hi_1220 = {dataGroup_hi_hi_1220, dataGroup_hi_lo_1220};
  wire [7:0]    dataGroup_4_19 = dataGroup_lo_1220[231:224];
  wire [2047:0] dataGroup_lo_1221 = {dataGroup_lo_hi_1221, dataGroup_lo_lo_1221};
  wire [2047:0] dataGroup_hi_1221 = {dataGroup_hi_hi_1221, dataGroup_hi_lo_1221};
  wire [7:0]    dataGroup_5_19 = dataGroup_lo_1221[279:272];
  wire [2047:0] dataGroup_lo_1222 = {dataGroup_lo_hi_1222, dataGroup_lo_lo_1222};
  wire [2047:0] dataGroup_hi_1222 = {dataGroup_hi_hi_1222, dataGroup_hi_lo_1222};
  wire [7:0]    dataGroup_6_19 = dataGroup_lo_1222[327:320];
  wire [2047:0] dataGroup_lo_1223 = {dataGroup_lo_hi_1223, dataGroup_lo_lo_1223};
  wire [2047:0] dataGroup_hi_1223 = {dataGroup_hi_hi_1223, dataGroup_hi_lo_1223};
  wire [7:0]    dataGroup_7_19 = dataGroup_lo_1223[375:368];
  wire [2047:0] dataGroup_lo_1224 = {dataGroup_lo_hi_1224, dataGroup_lo_lo_1224};
  wire [2047:0] dataGroup_hi_1224 = {dataGroup_hi_hi_1224, dataGroup_hi_lo_1224};
  wire [7:0]    dataGroup_8_19 = dataGroup_lo_1224[423:416];
  wire [2047:0] dataGroup_lo_1225 = {dataGroup_lo_hi_1225, dataGroup_lo_lo_1225};
  wire [2047:0] dataGroup_hi_1225 = {dataGroup_hi_hi_1225, dataGroup_hi_lo_1225};
  wire [7:0]    dataGroup_9_19 = dataGroup_lo_1225[471:464];
  wire [2047:0] dataGroup_lo_1226 = {dataGroup_lo_hi_1226, dataGroup_lo_lo_1226};
  wire [2047:0] dataGroup_hi_1226 = {dataGroup_hi_hi_1226, dataGroup_hi_lo_1226};
  wire [7:0]    dataGroup_10_19 = dataGroup_lo_1226[519:512];
  wire [2047:0] dataGroup_lo_1227 = {dataGroup_lo_hi_1227, dataGroup_lo_lo_1227};
  wire [2047:0] dataGroup_hi_1227 = {dataGroup_hi_hi_1227, dataGroup_hi_lo_1227};
  wire [7:0]    dataGroup_11_19 = dataGroup_lo_1227[567:560];
  wire [2047:0] dataGroup_lo_1228 = {dataGroup_lo_hi_1228, dataGroup_lo_lo_1228};
  wire [2047:0] dataGroup_hi_1228 = {dataGroup_hi_hi_1228, dataGroup_hi_lo_1228};
  wire [7:0]    dataGroup_12_19 = dataGroup_lo_1228[615:608];
  wire [2047:0] dataGroup_lo_1229 = {dataGroup_lo_hi_1229, dataGroup_lo_lo_1229};
  wire [2047:0] dataGroup_hi_1229 = {dataGroup_hi_hi_1229, dataGroup_hi_lo_1229};
  wire [7:0]    dataGroup_13_19 = dataGroup_lo_1229[663:656];
  wire [2047:0] dataGroup_lo_1230 = {dataGroup_lo_hi_1230, dataGroup_lo_lo_1230};
  wire [2047:0] dataGroup_hi_1230 = {dataGroup_hi_hi_1230, dataGroup_hi_lo_1230};
  wire [7:0]    dataGroup_14_19 = dataGroup_lo_1230[711:704];
  wire [2047:0] dataGroup_lo_1231 = {dataGroup_lo_hi_1231, dataGroup_lo_lo_1231};
  wire [2047:0] dataGroup_hi_1231 = {dataGroup_hi_hi_1231, dataGroup_hi_lo_1231};
  wire [7:0]    dataGroup_15_19 = dataGroup_lo_1231[759:752];
  wire [2047:0] dataGroup_lo_1232 = {dataGroup_lo_hi_1232, dataGroup_lo_lo_1232};
  wire [2047:0] dataGroup_hi_1232 = {dataGroup_hi_hi_1232, dataGroup_hi_lo_1232};
  wire [7:0]    dataGroup_16_19 = dataGroup_lo_1232[807:800];
  wire [2047:0] dataGroup_lo_1233 = {dataGroup_lo_hi_1233, dataGroup_lo_lo_1233};
  wire [2047:0] dataGroup_hi_1233 = {dataGroup_hi_hi_1233, dataGroup_hi_lo_1233};
  wire [7:0]    dataGroup_17_19 = dataGroup_lo_1233[855:848];
  wire [2047:0] dataGroup_lo_1234 = {dataGroup_lo_hi_1234, dataGroup_lo_lo_1234};
  wire [2047:0] dataGroup_hi_1234 = {dataGroup_hi_hi_1234, dataGroup_hi_lo_1234};
  wire [7:0]    dataGroup_18_19 = dataGroup_lo_1234[903:896];
  wire [2047:0] dataGroup_lo_1235 = {dataGroup_lo_hi_1235, dataGroup_lo_lo_1235};
  wire [2047:0] dataGroup_hi_1235 = {dataGroup_hi_hi_1235, dataGroup_hi_lo_1235};
  wire [7:0]    dataGroup_19_19 = dataGroup_lo_1235[951:944];
  wire [2047:0] dataGroup_lo_1236 = {dataGroup_lo_hi_1236, dataGroup_lo_lo_1236};
  wire [2047:0] dataGroup_hi_1236 = {dataGroup_hi_hi_1236, dataGroup_hi_lo_1236};
  wire [7:0]    dataGroup_20_19 = dataGroup_lo_1236[999:992];
  wire [2047:0] dataGroup_lo_1237 = {dataGroup_lo_hi_1237, dataGroup_lo_lo_1237};
  wire [2047:0] dataGroup_hi_1237 = {dataGroup_hi_hi_1237, dataGroup_hi_lo_1237};
  wire [7:0]    dataGroup_21_19 = dataGroup_lo_1237[1047:1040];
  wire [2047:0] dataGroup_lo_1238 = {dataGroup_lo_hi_1238, dataGroup_lo_lo_1238};
  wire [2047:0] dataGroup_hi_1238 = {dataGroup_hi_hi_1238, dataGroup_hi_lo_1238};
  wire [7:0]    dataGroup_22_19 = dataGroup_lo_1238[1095:1088];
  wire [2047:0] dataGroup_lo_1239 = {dataGroup_lo_hi_1239, dataGroup_lo_lo_1239};
  wire [2047:0] dataGroup_hi_1239 = {dataGroup_hi_hi_1239, dataGroup_hi_lo_1239};
  wire [7:0]    dataGroup_23_19 = dataGroup_lo_1239[1143:1136];
  wire [2047:0] dataGroup_lo_1240 = {dataGroup_lo_hi_1240, dataGroup_lo_lo_1240};
  wire [2047:0] dataGroup_hi_1240 = {dataGroup_hi_hi_1240, dataGroup_hi_lo_1240};
  wire [7:0]    dataGroup_24_19 = dataGroup_lo_1240[1191:1184];
  wire [2047:0] dataGroup_lo_1241 = {dataGroup_lo_hi_1241, dataGroup_lo_lo_1241};
  wire [2047:0] dataGroup_hi_1241 = {dataGroup_hi_hi_1241, dataGroup_hi_lo_1241};
  wire [7:0]    dataGroup_25_19 = dataGroup_lo_1241[1239:1232];
  wire [2047:0] dataGroup_lo_1242 = {dataGroup_lo_hi_1242, dataGroup_lo_lo_1242};
  wire [2047:0] dataGroup_hi_1242 = {dataGroup_hi_hi_1242, dataGroup_hi_lo_1242};
  wire [7:0]    dataGroup_26_19 = dataGroup_lo_1242[1287:1280];
  wire [2047:0] dataGroup_lo_1243 = {dataGroup_lo_hi_1243, dataGroup_lo_lo_1243};
  wire [2047:0] dataGroup_hi_1243 = {dataGroup_hi_hi_1243, dataGroup_hi_lo_1243};
  wire [7:0]    dataGroup_27_19 = dataGroup_lo_1243[1335:1328];
  wire [2047:0] dataGroup_lo_1244 = {dataGroup_lo_hi_1244, dataGroup_lo_lo_1244};
  wire [2047:0] dataGroup_hi_1244 = {dataGroup_hi_hi_1244, dataGroup_hi_lo_1244};
  wire [7:0]    dataGroup_28_19 = dataGroup_lo_1244[1383:1376];
  wire [2047:0] dataGroup_lo_1245 = {dataGroup_lo_hi_1245, dataGroup_lo_lo_1245};
  wire [2047:0] dataGroup_hi_1245 = {dataGroup_hi_hi_1245, dataGroup_hi_lo_1245};
  wire [7:0]    dataGroup_29_19 = dataGroup_lo_1245[1431:1424];
  wire [2047:0] dataGroup_lo_1246 = {dataGroup_lo_hi_1246, dataGroup_lo_lo_1246};
  wire [2047:0] dataGroup_hi_1246 = {dataGroup_hi_hi_1246, dataGroup_hi_lo_1246};
  wire [7:0]    dataGroup_30_19 = dataGroup_lo_1246[1479:1472];
  wire [2047:0] dataGroup_lo_1247 = {dataGroup_lo_hi_1247, dataGroup_lo_lo_1247};
  wire [2047:0] dataGroup_hi_1247 = {dataGroup_hi_hi_1247, dataGroup_hi_lo_1247};
  wire [7:0]    dataGroup_31_19 = dataGroup_lo_1247[1527:1520];
  wire [2047:0] dataGroup_lo_1248 = {dataGroup_lo_hi_1248, dataGroup_lo_lo_1248};
  wire [2047:0] dataGroup_hi_1248 = {dataGroup_hi_hi_1248, dataGroup_hi_lo_1248};
  wire [7:0]    dataGroup_32_19 = dataGroup_lo_1248[1575:1568];
  wire [2047:0] dataGroup_lo_1249 = {dataGroup_lo_hi_1249, dataGroup_lo_lo_1249};
  wire [2047:0] dataGroup_hi_1249 = {dataGroup_hi_hi_1249, dataGroup_hi_lo_1249};
  wire [7:0]    dataGroup_33_19 = dataGroup_lo_1249[1623:1616];
  wire [2047:0] dataGroup_lo_1250 = {dataGroup_lo_hi_1250, dataGroup_lo_lo_1250};
  wire [2047:0] dataGroup_hi_1250 = {dataGroup_hi_hi_1250, dataGroup_hi_lo_1250};
  wire [7:0]    dataGroup_34_19 = dataGroup_lo_1250[1671:1664];
  wire [2047:0] dataGroup_lo_1251 = {dataGroup_lo_hi_1251, dataGroup_lo_lo_1251};
  wire [2047:0] dataGroup_hi_1251 = {dataGroup_hi_hi_1251, dataGroup_hi_lo_1251};
  wire [7:0]    dataGroup_35_19 = dataGroup_lo_1251[1719:1712];
  wire [2047:0] dataGroup_lo_1252 = {dataGroup_lo_hi_1252, dataGroup_lo_lo_1252};
  wire [2047:0] dataGroup_hi_1252 = {dataGroup_hi_hi_1252, dataGroup_hi_lo_1252};
  wire [7:0]    dataGroup_36_19 = dataGroup_lo_1252[1767:1760];
  wire [2047:0] dataGroup_lo_1253 = {dataGroup_lo_hi_1253, dataGroup_lo_lo_1253};
  wire [2047:0] dataGroup_hi_1253 = {dataGroup_hi_hi_1253, dataGroup_hi_lo_1253};
  wire [7:0]    dataGroup_37_19 = dataGroup_lo_1253[1815:1808];
  wire [2047:0] dataGroup_lo_1254 = {dataGroup_lo_hi_1254, dataGroup_lo_lo_1254};
  wire [2047:0] dataGroup_hi_1254 = {dataGroup_hi_hi_1254, dataGroup_hi_lo_1254};
  wire [7:0]    dataGroup_38_19 = dataGroup_lo_1254[1863:1856];
  wire [2047:0] dataGroup_lo_1255 = {dataGroup_lo_hi_1255, dataGroup_lo_lo_1255};
  wire [2047:0] dataGroup_hi_1255 = {dataGroup_hi_hi_1255, dataGroup_hi_lo_1255};
  wire [7:0]    dataGroup_39_19 = dataGroup_lo_1255[1911:1904];
  wire [2047:0] dataGroup_lo_1256 = {dataGroup_lo_hi_1256, dataGroup_lo_lo_1256};
  wire [2047:0] dataGroup_hi_1256 = {dataGroup_hi_hi_1256, dataGroup_hi_lo_1256};
  wire [7:0]    dataGroup_40_19 = dataGroup_lo_1256[1959:1952];
  wire [2047:0] dataGroup_lo_1257 = {dataGroup_lo_hi_1257, dataGroup_lo_lo_1257};
  wire [2047:0] dataGroup_hi_1257 = {dataGroup_hi_hi_1257, dataGroup_hi_lo_1257};
  wire [7:0]    dataGroup_41_19 = dataGroup_lo_1257[2007:2000];
  wire [2047:0] dataGroup_lo_1258 = {dataGroup_lo_hi_1258, dataGroup_lo_lo_1258};
  wire [2047:0] dataGroup_hi_1258 = {dataGroup_hi_hi_1258, dataGroup_hi_lo_1258};
  wire [7:0]    dataGroup_42_19 = dataGroup_hi_1258[7:0];
  wire [2047:0] dataGroup_lo_1259 = {dataGroup_lo_hi_1259, dataGroup_lo_lo_1259};
  wire [2047:0] dataGroup_hi_1259 = {dataGroup_hi_hi_1259, dataGroup_hi_lo_1259};
  wire [7:0]    dataGroup_43_19 = dataGroup_hi_1259[55:48];
  wire [2047:0] dataGroup_lo_1260 = {dataGroup_lo_hi_1260, dataGroup_lo_lo_1260};
  wire [2047:0] dataGroup_hi_1260 = {dataGroup_hi_hi_1260, dataGroup_hi_lo_1260};
  wire [7:0]    dataGroup_44_19 = dataGroup_hi_1260[103:96];
  wire [2047:0] dataGroup_lo_1261 = {dataGroup_lo_hi_1261, dataGroup_lo_lo_1261};
  wire [2047:0] dataGroup_hi_1261 = {dataGroup_hi_hi_1261, dataGroup_hi_lo_1261};
  wire [7:0]    dataGroup_45_19 = dataGroup_hi_1261[151:144];
  wire [2047:0] dataGroup_lo_1262 = {dataGroup_lo_hi_1262, dataGroup_lo_lo_1262};
  wire [2047:0] dataGroup_hi_1262 = {dataGroup_hi_hi_1262, dataGroup_hi_lo_1262};
  wire [7:0]    dataGroup_46_19 = dataGroup_hi_1262[199:192];
  wire [2047:0] dataGroup_lo_1263 = {dataGroup_lo_hi_1263, dataGroup_lo_lo_1263};
  wire [2047:0] dataGroup_hi_1263 = {dataGroup_hi_hi_1263, dataGroup_hi_lo_1263};
  wire [7:0]    dataGroup_47_19 = dataGroup_hi_1263[247:240];
  wire [2047:0] dataGroup_lo_1264 = {dataGroup_lo_hi_1264, dataGroup_lo_lo_1264};
  wire [2047:0] dataGroup_hi_1264 = {dataGroup_hi_hi_1264, dataGroup_hi_lo_1264};
  wire [7:0]    dataGroup_48_19 = dataGroup_hi_1264[295:288];
  wire [2047:0] dataGroup_lo_1265 = {dataGroup_lo_hi_1265, dataGroup_lo_lo_1265};
  wire [2047:0] dataGroup_hi_1265 = {dataGroup_hi_hi_1265, dataGroup_hi_lo_1265};
  wire [7:0]    dataGroup_49_19 = dataGroup_hi_1265[343:336];
  wire [2047:0] dataGroup_lo_1266 = {dataGroup_lo_hi_1266, dataGroup_lo_lo_1266};
  wire [2047:0] dataGroup_hi_1266 = {dataGroup_hi_hi_1266, dataGroup_hi_lo_1266};
  wire [7:0]    dataGroup_50_19 = dataGroup_hi_1266[391:384];
  wire [2047:0] dataGroup_lo_1267 = {dataGroup_lo_hi_1267, dataGroup_lo_lo_1267};
  wire [2047:0] dataGroup_hi_1267 = {dataGroup_hi_hi_1267, dataGroup_hi_lo_1267};
  wire [7:0]    dataGroup_51_19 = dataGroup_hi_1267[439:432];
  wire [2047:0] dataGroup_lo_1268 = {dataGroup_lo_hi_1268, dataGroup_lo_lo_1268};
  wire [2047:0] dataGroup_hi_1268 = {dataGroup_hi_hi_1268, dataGroup_hi_lo_1268};
  wire [7:0]    dataGroup_52_19 = dataGroup_hi_1268[487:480];
  wire [2047:0] dataGroup_lo_1269 = {dataGroup_lo_hi_1269, dataGroup_lo_lo_1269};
  wire [2047:0] dataGroup_hi_1269 = {dataGroup_hi_hi_1269, dataGroup_hi_lo_1269};
  wire [7:0]    dataGroup_53_19 = dataGroup_hi_1269[535:528];
  wire [2047:0] dataGroup_lo_1270 = {dataGroup_lo_hi_1270, dataGroup_lo_lo_1270};
  wire [2047:0] dataGroup_hi_1270 = {dataGroup_hi_hi_1270, dataGroup_hi_lo_1270};
  wire [7:0]    dataGroup_54_19 = dataGroup_hi_1270[583:576];
  wire [2047:0] dataGroup_lo_1271 = {dataGroup_lo_hi_1271, dataGroup_lo_lo_1271};
  wire [2047:0] dataGroup_hi_1271 = {dataGroup_hi_hi_1271, dataGroup_hi_lo_1271};
  wire [7:0]    dataGroup_55_19 = dataGroup_hi_1271[631:624];
  wire [2047:0] dataGroup_lo_1272 = {dataGroup_lo_hi_1272, dataGroup_lo_lo_1272};
  wire [2047:0] dataGroup_hi_1272 = {dataGroup_hi_hi_1272, dataGroup_hi_lo_1272};
  wire [7:0]    dataGroup_56_19 = dataGroup_hi_1272[679:672];
  wire [2047:0] dataGroup_lo_1273 = {dataGroup_lo_hi_1273, dataGroup_lo_lo_1273};
  wire [2047:0] dataGroup_hi_1273 = {dataGroup_hi_hi_1273, dataGroup_hi_lo_1273};
  wire [7:0]    dataGroup_57_19 = dataGroup_hi_1273[727:720];
  wire [2047:0] dataGroup_lo_1274 = {dataGroup_lo_hi_1274, dataGroup_lo_lo_1274};
  wire [2047:0] dataGroup_hi_1274 = {dataGroup_hi_hi_1274, dataGroup_hi_lo_1274};
  wire [7:0]    dataGroup_58_19 = dataGroup_hi_1274[775:768];
  wire [2047:0] dataGroup_lo_1275 = {dataGroup_lo_hi_1275, dataGroup_lo_lo_1275};
  wire [2047:0] dataGroup_hi_1275 = {dataGroup_hi_hi_1275, dataGroup_hi_lo_1275};
  wire [7:0]    dataGroup_59_19 = dataGroup_hi_1275[823:816];
  wire [2047:0] dataGroup_lo_1276 = {dataGroup_lo_hi_1276, dataGroup_lo_lo_1276};
  wire [2047:0] dataGroup_hi_1276 = {dataGroup_hi_hi_1276, dataGroup_hi_lo_1276};
  wire [7:0]    dataGroup_60_19 = dataGroup_hi_1276[871:864];
  wire [2047:0] dataGroup_lo_1277 = {dataGroup_lo_hi_1277, dataGroup_lo_lo_1277};
  wire [2047:0] dataGroup_hi_1277 = {dataGroup_hi_hi_1277, dataGroup_hi_lo_1277};
  wire [7:0]    dataGroup_61_19 = dataGroup_hi_1277[919:912];
  wire [2047:0] dataGroup_lo_1278 = {dataGroup_lo_hi_1278, dataGroup_lo_lo_1278};
  wire [2047:0] dataGroup_hi_1278 = {dataGroup_hi_hi_1278, dataGroup_hi_lo_1278};
  wire [7:0]    dataGroup_62_19 = dataGroup_hi_1278[967:960];
  wire [2047:0] dataGroup_lo_1279 = {dataGroup_lo_hi_1279, dataGroup_lo_lo_1279};
  wire [2047:0] dataGroup_hi_1279 = {dataGroup_hi_hi_1279, dataGroup_hi_lo_1279};
  wire [7:0]    dataGroup_63_19 = dataGroup_hi_1279[1015:1008];
  wire [15:0]   res_lo_lo_lo_lo_lo_19 = {dataGroup_1_19, dataGroup_0_19};
  wire [15:0]   res_lo_lo_lo_lo_hi_19 = {dataGroup_3_19, dataGroup_2_19};
  wire [31:0]   res_lo_lo_lo_lo_19 = {res_lo_lo_lo_lo_hi_19, res_lo_lo_lo_lo_lo_19};
  wire [15:0]   res_lo_lo_lo_hi_lo_19 = {dataGroup_5_19, dataGroup_4_19};
  wire [15:0]   res_lo_lo_lo_hi_hi_19 = {dataGroup_7_19, dataGroup_6_19};
  wire [31:0]   res_lo_lo_lo_hi_19 = {res_lo_lo_lo_hi_hi_19, res_lo_lo_lo_hi_lo_19};
  wire [63:0]   res_lo_lo_lo_19 = {res_lo_lo_lo_hi_19, res_lo_lo_lo_lo_19};
  wire [15:0]   res_lo_lo_hi_lo_lo_19 = {dataGroup_9_19, dataGroup_8_19};
  wire [15:0]   res_lo_lo_hi_lo_hi_19 = {dataGroup_11_19, dataGroup_10_19};
  wire [31:0]   res_lo_lo_hi_lo_19 = {res_lo_lo_hi_lo_hi_19, res_lo_lo_hi_lo_lo_19};
  wire [15:0]   res_lo_lo_hi_hi_lo_19 = {dataGroup_13_19, dataGroup_12_19};
  wire [15:0]   res_lo_lo_hi_hi_hi_19 = {dataGroup_15_19, dataGroup_14_19};
  wire [31:0]   res_lo_lo_hi_hi_19 = {res_lo_lo_hi_hi_hi_19, res_lo_lo_hi_hi_lo_19};
  wire [63:0]   res_lo_lo_hi_19 = {res_lo_lo_hi_hi_19, res_lo_lo_hi_lo_19};
  wire [127:0]  res_lo_lo_19 = {res_lo_lo_hi_19, res_lo_lo_lo_19};
  wire [15:0]   res_lo_hi_lo_lo_lo_19 = {dataGroup_17_19, dataGroup_16_19};
  wire [15:0]   res_lo_hi_lo_lo_hi_19 = {dataGroup_19_19, dataGroup_18_19};
  wire [31:0]   res_lo_hi_lo_lo_19 = {res_lo_hi_lo_lo_hi_19, res_lo_hi_lo_lo_lo_19};
  wire [15:0]   res_lo_hi_lo_hi_lo_19 = {dataGroup_21_19, dataGroup_20_19};
  wire [15:0]   res_lo_hi_lo_hi_hi_19 = {dataGroup_23_19, dataGroup_22_19};
  wire [31:0]   res_lo_hi_lo_hi_19 = {res_lo_hi_lo_hi_hi_19, res_lo_hi_lo_hi_lo_19};
  wire [63:0]   res_lo_hi_lo_19 = {res_lo_hi_lo_hi_19, res_lo_hi_lo_lo_19};
  wire [15:0]   res_lo_hi_hi_lo_lo_19 = {dataGroup_25_19, dataGroup_24_19};
  wire [15:0]   res_lo_hi_hi_lo_hi_19 = {dataGroup_27_19, dataGroup_26_19};
  wire [31:0]   res_lo_hi_hi_lo_19 = {res_lo_hi_hi_lo_hi_19, res_lo_hi_hi_lo_lo_19};
  wire [15:0]   res_lo_hi_hi_hi_lo_19 = {dataGroup_29_19, dataGroup_28_19};
  wire [15:0]   res_lo_hi_hi_hi_hi_19 = {dataGroup_31_19, dataGroup_30_19};
  wire [31:0]   res_lo_hi_hi_hi_19 = {res_lo_hi_hi_hi_hi_19, res_lo_hi_hi_hi_lo_19};
  wire [63:0]   res_lo_hi_hi_19 = {res_lo_hi_hi_hi_19, res_lo_hi_hi_lo_19};
  wire [127:0]  res_lo_hi_19 = {res_lo_hi_hi_19, res_lo_hi_lo_19};
  wire [255:0]  res_lo_19 = {res_lo_hi_19, res_lo_lo_19};
  wire [15:0]   res_hi_lo_lo_lo_lo_19 = {dataGroup_33_19, dataGroup_32_19};
  wire [15:0]   res_hi_lo_lo_lo_hi_19 = {dataGroup_35_19, dataGroup_34_19};
  wire [31:0]   res_hi_lo_lo_lo_19 = {res_hi_lo_lo_lo_hi_19, res_hi_lo_lo_lo_lo_19};
  wire [15:0]   res_hi_lo_lo_hi_lo_19 = {dataGroup_37_19, dataGroup_36_19};
  wire [15:0]   res_hi_lo_lo_hi_hi_19 = {dataGroup_39_19, dataGroup_38_19};
  wire [31:0]   res_hi_lo_lo_hi_19 = {res_hi_lo_lo_hi_hi_19, res_hi_lo_lo_hi_lo_19};
  wire [63:0]   res_hi_lo_lo_19 = {res_hi_lo_lo_hi_19, res_hi_lo_lo_lo_19};
  wire [15:0]   res_hi_lo_hi_lo_lo_19 = {dataGroup_41_19, dataGroup_40_19};
  wire [15:0]   res_hi_lo_hi_lo_hi_19 = {dataGroup_43_19, dataGroup_42_19};
  wire [31:0]   res_hi_lo_hi_lo_19 = {res_hi_lo_hi_lo_hi_19, res_hi_lo_hi_lo_lo_19};
  wire [15:0]   res_hi_lo_hi_hi_lo_19 = {dataGroup_45_19, dataGroup_44_19};
  wire [15:0]   res_hi_lo_hi_hi_hi_19 = {dataGroup_47_19, dataGroup_46_19};
  wire [31:0]   res_hi_lo_hi_hi_19 = {res_hi_lo_hi_hi_hi_19, res_hi_lo_hi_hi_lo_19};
  wire [63:0]   res_hi_lo_hi_19 = {res_hi_lo_hi_hi_19, res_hi_lo_hi_lo_19};
  wire [127:0]  res_hi_lo_19 = {res_hi_lo_hi_19, res_hi_lo_lo_19};
  wire [15:0]   res_hi_hi_lo_lo_lo_19 = {dataGroup_49_19, dataGroup_48_19};
  wire [15:0]   res_hi_hi_lo_lo_hi_19 = {dataGroup_51_19, dataGroup_50_19};
  wire [31:0]   res_hi_hi_lo_lo_19 = {res_hi_hi_lo_lo_hi_19, res_hi_hi_lo_lo_lo_19};
  wire [15:0]   res_hi_hi_lo_hi_lo_19 = {dataGroup_53_19, dataGroup_52_19};
  wire [15:0]   res_hi_hi_lo_hi_hi_19 = {dataGroup_55_19, dataGroup_54_19};
  wire [31:0]   res_hi_hi_lo_hi_19 = {res_hi_hi_lo_hi_hi_19, res_hi_hi_lo_hi_lo_19};
  wire [63:0]   res_hi_hi_lo_19 = {res_hi_hi_lo_hi_19, res_hi_hi_lo_lo_19};
  wire [15:0]   res_hi_hi_hi_lo_lo_19 = {dataGroup_57_19, dataGroup_56_19};
  wire [15:0]   res_hi_hi_hi_lo_hi_19 = {dataGroup_59_19, dataGroup_58_19};
  wire [31:0]   res_hi_hi_hi_lo_19 = {res_hi_hi_hi_lo_hi_19, res_hi_hi_hi_lo_lo_19};
  wire [15:0]   res_hi_hi_hi_hi_lo_19 = {dataGroup_61_19, dataGroup_60_19};
  wire [15:0]   res_hi_hi_hi_hi_hi_19 = {dataGroup_63_19, dataGroup_62_19};
  wire [31:0]   res_hi_hi_hi_hi_19 = {res_hi_hi_hi_hi_hi_19, res_hi_hi_hi_hi_lo_19};
  wire [63:0]   res_hi_hi_hi_19 = {res_hi_hi_hi_hi_19, res_hi_hi_hi_lo_19};
  wire [127:0]  res_hi_hi_19 = {res_hi_hi_hi_19, res_hi_hi_lo_19};
  wire [255:0]  res_hi_19 = {res_hi_hi_19, res_hi_lo_19};
  wire [511:0]  res_44 = {res_hi_19, res_lo_19};
  wire [2047:0] dataGroup_lo_1280 = {dataGroup_lo_hi_1280, dataGroup_lo_lo_1280};
  wire [2047:0] dataGroup_hi_1280 = {dataGroup_hi_hi_1280, dataGroup_hi_lo_1280};
  wire [7:0]    dataGroup_0_20 = dataGroup_lo_1280[47:40];
  wire [2047:0] dataGroup_lo_1281 = {dataGroup_lo_hi_1281, dataGroup_lo_lo_1281};
  wire [2047:0] dataGroup_hi_1281 = {dataGroup_hi_hi_1281, dataGroup_hi_lo_1281};
  wire [7:0]    dataGroup_1_20 = dataGroup_lo_1281[95:88];
  wire [2047:0] dataGroup_lo_1282 = {dataGroup_lo_hi_1282, dataGroup_lo_lo_1282};
  wire [2047:0] dataGroup_hi_1282 = {dataGroup_hi_hi_1282, dataGroup_hi_lo_1282};
  wire [7:0]    dataGroup_2_20 = dataGroup_lo_1282[143:136];
  wire [2047:0] dataGroup_lo_1283 = {dataGroup_lo_hi_1283, dataGroup_lo_lo_1283};
  wire [2047:0] dataGroup_hi_1283 = {dataGroup_hi_hi_1283, dataGroup_hi_lo_1283};
  wire [7:0]    dataGroup_3_20 = dataGroup_lo_1283[191:184];
  wire [2047:0] dataGroup_lo_1284 = {dataGroup_lo_hi_1284, dataGroup_lo_lo_1284};
  wire [2047:0] dataGroup_hi_1284 = {dataGroup_hi_hi_1284, dataGroup_hi_lo_1284};
  wire [7:0]    dataGroup_4_20 = dataGroup_lo_1284[239:232];
  wire [2047:0] dataGroup_lo_1285 = {dataGroup_lo_hi_1285, dataGroup_lo_lo_1285};
  wire [2047:0] dataGroup_hi_1285 = {dataGroup_hi_hi_1285, dataGroup_hi_lo_1285};
  wire [7:0]    dataGroup_5_20 = dataGroup_lo_1285[287:280];
  wire [2047:0] dataGroup_lo_1286 = {dataGroup_lo_hi_1286, dataGroup_lo_lo_1286};
  wire [2047:0] dataGroup_hi_1286 = {dataGroup_hi_hi_1286, dataGroup_hi_lo_1286};
  wire [7:0]    dataGroup_6_20 = dataGroup_lo_1286[335:328];
  wire [2047:0] dataGroup_lo_1287 = {dataGroup_lo_hi_1287, dataGroup_lo_lo_1287};
  wire [2047:0] dataGroup_hi_1287 = {dataGroup_hi_hi_1287, dataGroup_hi_lo_1287};
  wire [7:0]    dataGroup_7_20 = dataGroup_lo_1287[383:376];
  wire [2047:0] dataGroup_lo_1288 = {dataGroup_lo_hi_1288, dataGroup_lo_lo_1288};
  wire [2047:0] dataGroup_hi_1288 = {dataGroup_hi_hi_1288, dataGroup_hi_lo_1288};
  wire [7:0]    dataGroup_8_20 = dataGroup_lo_1288[431:424];
  wire [2047:0] dataGroup_lo_1289 = {dataGroup_lo_hi_1289, dataGroup_lo_lo_1289};
  wire [2047:0] dataGroup_hi_1289 = {dataGroup_hi_hi_1289, dataGroup_hi_lo_1289};
  wire [7:0]    dataGroup_9_20 = dataGroup_lo_1289[479:472];
  wire [2047:0] dataGroup_lo_1290 = {dataGroup_lo_hi_1290, dataGroup_lo_lo_1290};
  wire [2047:0] dataGroup_hi_1290 = {dataGroup_hi_hi_1290, dataGroup_hi_lo_1290};
  wire [7:0]    dataGroup_10_20 = dataGroup_lo_1290[527:520];
  wire [2047:0] dataGroup_lo_1291 = {dataGroup_lo_hi_1291, dataGroup_lo_lo_1291};
  wire [2047:0] dataGroup_hi_1291 = {dataGroup_hi_hi_1291, dataGroup_hi_lo_1291};
  wire [7:0]    dataGroup_11_20 = dataGroup_lo_1291[575:568];
  wire [2047:0] dataGroup_lo_1292 = {dataGroup_lo_hi_1292, dataGroup_lo_lo_1292};
  wire [2047:0] dataGroup_hi_1292 = {dataGroup_hi_hi_1292, dataGroup_hi_lo_1292};
  wire [7:0]    dataGroup_12_20 = dataGroup_lo_1292[623:616];
  wire [2047:0] dataGroup_lo_1293 = {dataGroup_lo_hi_1293, dataGroup_lo_lo_1293};
  wire [2047:0] dataGroup_hi_1293 = {dataGroup_hi_hi_1293, dataGroup_hi_lo_1293};
  wire [7:0]    dataGroup_13_20 = dataGroup_lo_1293[671:664];
  wire [2047:0] dataGroup_lo_1294 = {dataGroup_lo_hi_1294, dataGroup_lo_lo_1294};
  wire [2047:0] dataGroup_hi_1294 = {dataGroup_hi_hi_1294, dataGroup_hi_lo_1294};
  wire [7:0]    dataGroup_14_20 = dataGroup_lo_1294[719:712];
  wire [2047:0] dataGroup_lo_1295 = {dataGroup_lo_hi_1295, dataGroup_lo_lo_1295};
  wire [2047:0] dataGroup_hi_1295 = {dataGroup_hi_hi_1295, dataGroup_hi_lo_1295};
  wire [7:0]    dataGroup_15_20 = dataGroup_lo_1295[767:760];
  wire [2047:0] dataGroup_lo_1296 = {dataGroup_lo_hi_1296, dataGroup_lo_lo_1296};
  wire [2047:0] dataGroup_hi_1296 = {dataGroup_hi_hi_1296, dataGroup_hi_lo_1296};
  wire [7:0]    dataGroup_16_20 = dataGroup_lo_1296[815:808];
  wire [2047:0] dataGroup_lo_1297 = {dataGroup_lo_hi_1297, dataGroup_lo_lo_1297};
  wire [2047:0] dataGroup_hi_1297 = {dataGroup_hi_hi_1297, dataGroup_hi_lo_1297};
  wire [7:0]    dataGroup_17_20 = dataGroup_lo_1297[863:856];
  wire [2047:0] dataGroup_lo_1298 = {dataGroup_lo_hi_1298, dataGroup_lo_lo_1298};
  wire [2047:0] dataGroup_hi_1298 = {dataGroup_hi_hi_1298, dataGroup_hi_lo_1298};
  wire [7:0]    dataGroup_18_20 = dataGroup_lo_1298[911:904];
  wire [2047:0] dataGroup_lo_1299 = {dataGroup_lo_hi_1299, dataGroup_lo_lo_1299};
  wire [2047:0] dataGroup_hi_1299 = {dataGroup_hi_hi_1299, dataGroup_hi_lo_1299};
  wire [7:0]    dataGroup_19_20 = dataGroup_lo_1299[959:952];
  wire [2047:0] dataGroup_lo_1300 = {dataGroup_lo_hi_1300, dataGroup_lo_lo_1300};
  wire [2047:0] dataGroup_hi_1300 = {dataGroup_hi_hi_1300, dataGroup_hi_lo_1300};
  wire [7:0]    dataGroup_20_20 = dataGroup_lo_1300[1007:1000];
  wire [2047:0] dataGroup_lo_1301 = {dataGroup_lo_hi_1301, dataGroup_lo_lo_1301};
  wire [2047:0] dataGroup_hi_1301 = {dataGroup_hi_hi_1301, dataGroup_hi_lo_1301};
  wire [7:0]    dataGroup_21_20 = dataGroup_lo_1301[1055:1048];
  wire [2047:0] dataGroup_lo_1302 = {dataGroup_lo_hi_1302, dataGroup_lo_lo_1302};
  wire [2047:0] dataGroup_hi_1302 = {dataGroup_hi_hi_1302, dataGroup_hi_lo_1302};
  wire [7:0]    dataGroup_22_20 = dataGroup_lo_1302[1103:1096];
  wire [2047:0] dataGroup_lo_1303 = {dataGroup_lo_hi_1303, dataGroup_lo_lo_1303};
  wire [2047:0] dataGroup_hi_1303 = {dataGroup_hi_hi_1303, dataGroup_hi_lo_1303};
  wire [7:0]    dataGroup_23_20 = dataGroup_lo_1303[1151:1144];
  wire [2047:0] dataGroup_lo_1304 = {dataGroup_lo_hi_1304, dataGroup_lo_lo_1304};
  wire [2047:0] dataGroup_hi_1304 = {dataGroup_hi_hi_1304, dataGroup_hi_lo_1304};
  wire [7:0]    dataGroup_24_20 = dataGroup_lo_1304[1199:1192];
  wire [2047:0] dataGroup_lo_1305 = {dataGroup_lo_hi_1305, dataGroup_lo_lo_1305};
  wire [2047:0] dataGroup_hi_1305 = {dataGroup_hi_hi_1305, dataGroup_hi_lo_1305};
  wire [7:0]    dataGroup_25_20 = dataGroup_lo_1305[1247:1240];
  wire [2047:0] dataGroup_lo_1306 = {dataGroup_lo_hi_1306, dataGroup_lo_lo_1306};
  wire [2047:0] dataGroup_hi_1306 = {dataGroup_hi_hi_1306, dataGroup_hi_lo_1306};
  wire [7:0]    dataGroup_26_20 = dataGroup_lo_1306[1295:1288];
  wire [2047:0] dataGroup_lo_1307 = {dataGroup_lo_hi_1307, dataGroup_lo_lo_1307};
  wire [2047:0] dataGroup_hi_1307 = {dataGroup_hi_hi_1307, dataGroup_hi_lo_1307};
  wire [7:0]    dataGroup_27_20 = dataGroup_lo_1307[1343:1336];
  wire [2047:0] dataGroup_lo_1308 = {dataGroup_lo_hi_1308, dataGroup_lo_lo_1308};
  wire [2047:0] dataGroup_hi_1308 = {dataGroup_hi_hi_1308, dataGroup_hi_lo_1308};
  wire [7:0]    dataGroup_28_20 = dataGroup_lo_1308[1391:1384];
  wire [2047:0] dataGroup_lo_1309 = {dataGroup_lo_hi_1309, dataGroup_lo_lo_1309};
  wire [2047:0] dataGroup_hi_1309 = {dataGroup_hi_hi_1309, dataGroup_hi_lo_1309};
  wire [7:0]    dataGroup_29_20 = dataGroup_lo_1309[1439:1432];
  wire [2047:0] dataGroup_lo_1310 = {dataGroup_lo_hi_1310, dataGroup_lo_lo_1310};
  wire [2047:0] dataGroup_hi_1310 = {dataGroup_hi_hi_1310, dataGroup_hi_lo_1310};
  wire [7:0]    dataGroup_30_20 = dataGroup_lo_1310[1487:1480];
  wire [2047:0] dataGroup_lo_1311 = {dataGroup_lo_hi_1311, dataGroup_lo_lo_1311};
  wire [2047:0] dataGroup_hi_1311 = {dataGroup_hi_hi_1311, dataGroup_hi_lo_1311};
  wire [7:0]    dataGroup_31_20 = dataGroup_lo_1311[1535:1528];
  wire [2047:0] dataGroup_lo_1312 = {dataGroup_lo_hi_1312, dataGroup_lo_lo_1312};
  wire [2047:0] dataGroup_hi_1312 = {dataGroup_hi_hi_1312, dataGroup_hi_lo_1312};
  wire [7:0]    dataGroup_32_20 = dataGroup_lo_1312[1583:1576];
  wire [2047:0] dataGroup_lo_1313 = {dataGroup_lo_hi_1313, dataGroup_lo_lo_1313};
  wire [2047:0] dataGroup_hi_1313 = {dataGroup_hi_hi_1313, dataGroup_hi_lo_1313};
  wire [7:0]    dataGroup_33_20 = dataGroup_lo_1313[1631:1624];
  wire [2047:0] dataGroup_lo_1314 = {dataGroup_lo_hi_1314, dataGroup_lo_lo_1314};
  wire [2047:0] dataGroup_hi_1314 = {dataGroup_hi_hi_1314, dataGroup_hi_lo_1314};
  wire [7:0]    dataGroup_34_20 = dataGroup_lo_1314[1679:1672];
  wire [2047:0] dataGroup_lo_1315 = {dataGroup_lo_hi_1315, dataGroup_lo_lo_1315};
  wire [2047:0] dataGroup_hi_1315 = {dataGroup_hi_hi_1315, dataGroup_hi_lo_1315};
  wire [7:0]    dataGroup_35_20 = dataGroup_lo_1315[1727:1720];
  wire [2047:0] dataGroup_lo_1316 = {dataGroup_lo_hi_1316, dataGroup_lo_lo_1316};
  wire [2047:0] dataGroup_hi_1316 = {dataGroup_hi_hi_1316, dataGroup_hi_lo_1316};
  wire [7:0]    dataGroup_36_20 = dataGroup_lo_1316[1775:1768];
  wire [2047:0] dataGroup_lo_1317 = {dataGroup_lo_hi_1317, dataGroup_lo_lo_1317};
  wire [2047:0] dataGroup_hi_1317 = {dataGroup_hi_hi_1317, dataGroup_hi_lo_1317};
  wire [7:0]    dataGroup_37_20 = dataGroup_lo_1317[1823:1816];
  wire [2047:0] dataGroup_lo_1318 = {dataGroup_lo_hi_1318, dataGroup_lo_lo_1318};
  wire [2047:0] dataGroup_hi_1318 = {dataGroup_hi_hi_1318, dataGroup_hi_lo_1318};
  wire [7:0]    dataGroup_38_20 = dataGroup_lo_1318[1871:1864];
  wire [2047:0] dataGroup_lo_1319 = {dataGroup_lo_hi_1319, dataGroup_lo_lo_1319};
  wire [2047:0] dataGroup_hi_1319 = {dataGroup_hi_hi_1319, dataGroup_hi_lo_1319};
  wire [7:0]    dataGroup_39_20 = dataGroup_lo_1319[1919:1912];
  wire [2047:0] dataGroup_lo_1320 = {dataGroup_lo_hi_1320, dataGroup_lo_lo_1320};
  wire [2047:0] dataGroup_hi_1320 = {dataGroup_hi_hi_1320, dataGroup_hi_lo_1320};
  wire [7:0]    dataGroup_40_20 = dataGroup_lo_1320[1967:1960];
  wire [2047:0] dataGroup_lo_1321 = {dataGroup_lo_hi_1321, dataGroup_lo_lo_1321};
  wire [2047:0] dataGroup_hi_1321 = {dataGroup_hi_hi_1321, dataGroup_hi_lo_1321};
  wire [7:0]    dataGroup_41_20 = dataGroup_lo_1321[2015:2008];
  wire [2047:0] dataGroup_lo_1322 = {dataGroup_lo_hi_1322, dataGroup_lo_lo_1322};
  wire [2047:0] dataGroup_hi_1322 = {dataGroup_hi_hi_1322, dataGroup_hi_lo_1322};
  wire [7:0]    dataGroup_42_20 = dataGroup_hi_1322[15:8];
  wire [2047:0] dataGroup_lo_1323 = {dataGroup_lo_hi_1323, dataGroup_lo_lo_1323};
  wire [2047:0] dataGroup_hi_1323 = {dataGroup_hi_hi_1323, dataGroup_hi_lo_1323};
  wire [7:0]    dataGroup_43_20 = dataGroup_hi_1323[63:56];
  wire [2047:0] dataGroup_lo_1324 = {dataGroup_lo_hi_1324, dataGroup_lo_lo_1324};
  wire [2047:0] dataGroup_hi_1324 = {dataGroup_hi_hi_1324, dataGroup_hi_lo_1324};
  wire [7:0]    dataGroup_44_20 = dataGroup_hi_1324[111:104];
  wire [2047:0] dataGroup_lo_1325 = {dataGroup_lo_hi_1325, dataGroup_lo_lo_1325};
  wire [2047:0] dataGroup_hi_1325 = {dataGroup_hi_hi_1325, dataGroup_hi_lo_1325};
  wire [7:0]    dataGroup_45_20 = dataGroup_hi_1325[159:152];
  wire [2047:0] dataGroup_lo_1326 = {dataGroup_lo_hi_1326, dataGroup_lo_lo_1326};
  wire [2047:0] dataGroup_hi_1326 = {dataGroup_hi_hi_1326, dataGroup_hi_lo_1326};
  wire [7:0]    dataGroup_46_20 = dataGroup_hi_1326[207:200];
  wire [2047:0] dataGroup_lo_1327 = {dataGroup_lo_hi_1327, dataGroup_lo_lo_1327};
  wire [2047:0] dataGroup_hi_1327 = {dataGroup_hi_hi_1327, dataGroup_hi_lo_1327};
  wire [7:0]    dataGroup_47_20 = dataGroup_hi_1327[255:248];
  wire [2047:0] dataGroup_lo_1328 = {dataGroup_lo_hi_1328, dataGroup_lo_lo_1328};
  wire [2047:0] dataGroup_hi_1328 = {dataGroup_hi_hi_1328, dataGroup_hi_lo_1328};
  wire [7:0]    dataGroup_48_20 = dataGroup_hi_1328[303:296];
  wire [2047:0] dataGroup_lo_1329 = {dataGroup_lo_hi_1329, dataGroup_lo_lo_1329};
  wire [2047:0] dataGroup_hi_1329 = {dataGroup_hi_hi_1329, dataGroup_hi_lo_1329};
  wire [7:0]    dataGroup_49_20 = dataGroup_hi_1329[351:344];
  wire [2047:0] dataGroup_lo_1330 = {dataGroup_lo_hi_1330, dataGroup_lo_lo_1330};
  wire [2047:0] dataGroup_hi_1330 = {dataGroup_hi_hi_1330, dataGroup_hi_lo_1330};
  wire [7:0]    dataGroup_50_20 = dataGroup_hi_1330[399:392];
  wire [2047:0] dataGroup_lo_1331 = {dataGroup_lo_hi_1331, dataGroup_lo_lo_1331};
  wire [2047:0] dataGroup_hi_1331 = {dataGroup_hi_hi_1331, dataGroup_hi_lo_1331};
  wire [7:0]    dataGroup_51_20 = dataGroup_hi_1331[447:440];
  wire [2047:0] dataGroup_lo_1332 = {dataGroup_lo_hi_1332, dataGroup_lo_lo_1332};
  wire [2047:0] dataGroup_hi_1332 = {dataGroup_hi_hi_1332, dataGroup_hi_lo_1332};
  wire [7:0]    dataGroup_52_20 = dataGroup_hi_1332[495:488];
  wire [2047:0] dataGroup_lo_1333 = {dataGroup_lo_hi_1333, dataGroup_lo_lo_1333};
  wire [2047:0] dataGroup_hi_1333 = {dataGroup_hi_hi_1333, dataGroup_hi_lo_1333};
  wire [7:0]    dataGroup_53_20 = dataGroup_hi_1333[543:536];
  wire [2047:0] dataGroup_lo_1334 = {dataGroup_lo_hi_1334, dataGroup_lo_lo_1334};
  wire [2047:0] dataGroup_hi_1334 = {dataGroup_hi_hi_1334, dataGroup_hi_lo_1334};
  wire [7:0]    dataGroup_54_20 = dataGroup_hi_1334[591:584];
  wire [2047:0] dataGroup_lo_1335 = {dataGroup_lo_hi_1335, dataGroup_lo_lo_1335};
  wire [2047:0] dataGroup_hi_1335 = {dataGroup_hi_hi_1335, dataGroup_hi_lo_1335};
  wire [7:0]    dataGroup_55_20 = dataGroup_hi_1335[639:632];
  wire [2047:0] dataGroup_lo_1336 = {dataGroup_lo_hi_1336, dataGroup_lo_lo_1336};
  wire [2047:0] dataGroup_hi_1336 = {dataGroup_hi_hi_1336, dataGroup_hi_lo_1336};
  wire [7:0]    dataGroup_56_20 = dataGroup_hi_1336[687:680];
  wire [2047:0] dataGroup_lo_1337 = {dataGroup_lo_hi_1337, dataGroup_lo_lo_1337};
  wire [2047:0] dataGroup_hi_1337 = {dataGroup_hi_hi_1337, dataGroup_hi_lo_1337};
  wire [7:0]    dataGroup_57_20 = dataGroup_hi_1337[735:728];
  wire [2047:0] dataGroup_lo_1338 = {dataGroup_lo_hi_1338, dataGroup_lo_lo_1338};
  wire [2047:0] dataGroup_hi_1338 = {dataGroup_hi_hi_1338, dataGroup_hi_lo_1338};
  wire [7:0]    dataGroup_58_20 = dataGroup_hi_1338[783:776];
  wire [2047:0] dataGroup_lo_1339 = {dataGroup_lo_hi_1339, dataGroup_lo_lo_1339};
  wire [2047:0] dataGroup_hi_1339 = {dataGroup_hi_hi_1339, dataGroup_hi_lo_1339};
  wire [7:0]    dataGroup_59_20 = dataGroup_hi_1339[831:824];
  wire [2047:0] dataGroup_lo_1340 = {dataGroup_lo_hi_1340, dataGroup_lo_lo_1340};
  wire [2047:0] dataGroup_hi_1340 = {dataGroup_hi_hi_1340, dataGroup_hi_lo_1340};
  wire [7:0]    dataGroup_60_20 = dataGroup_hi_1340[879:872];
  wire [2047:0] dataGroup_lo_1341 = {dataGroup_lo_hi_1341, dataGroup_lo_lo_1341};
  wire [2047:0] dataGroup_hi_1341 = {dataGroup_hi_hi_1341, dataGroup_hi_lo_1341};
  wire [7:0]    dataGroup_61_20 = dataGroup_hi_1341[927:920];
  wire [2047:0] dataGroup_lo_1342 = {dataGroup_lo_hi_1342, dataGroup_lo_lo_1342};
  wire [2047:0] dataGroup_hi_1342 = {dataGroup_hi_hi_1342, dataGroup_hi_lo_1342};
  wire [7:0]    dataGroup_62_20 = dataGroup_hi_1342[975:968];
  wire [2047:0] dataGroup_lo_1343 = {dataGroup_lo_hi_1343, dataGroup_lo_lo_1343};
  wire [2047:0] dataGroup_hi_1343 = {dataGroup_hi_hi_1343, dataGroup_hi_lo_1343};
  wire [7:0]    dataGroup_63_20 = dataGroup_hi_1343[1023:1016];
  wire [15:0]   res_lo_lo_lo_lo_lo_20 = {dataGroup_1_20, dataGroup_0_20};
  wire [15:0]   res_lo_lo_lo_lo_hi_20 = {dataGroup_3_20, dataGroup_2_20};
  wire [31:0]   res_lo_lo_lo_lo_20 = {res_lo_lo_lo_lo_hi_20, res_lo_lo_lo_lo_lo_20};
  wire [15:0]   res_lo_lo_lo_hi_lo_20 = {dataGroup_5_20, dataGroup_4_20};
  wire [15:0]   res_lo_lo_lo_hi_hi_20 = {dataGroup_7_20, dataGroup_6_20};
  wire [31:0]   res_lo_lo_lo_hi_20 = {res_lo_lo_lo_hi_hi_20, res_lo_lo_lo_hi_lo_20};
  wire [63:0]   res_lo_lo_lo_20 = {res_lo_lo_lo_hi_20, res_lo_lo_lo_lo_20};
  wire [15:0]   res_lo_lo_hi_lo_lo_20 = {dataGroup_9_20, dataGroup_8_20};
  wire [15:0]   res_lo_lo_hi_lo_hi_20 = {dataGroup_11_20, dataGroup_10_20};
  wire [31:0]   res_lo_lo_hi_lo_20 = {res_lo_lo_hi_lo_hi_20, res_lo_lo_hi_lo_lo_20};
  wire [15:0]   res_lo_lo_hi_hi_lo_20 = {dataGroup_13_20, dataGroup_12_20};
  wire [15:0]   res_lo_lo_hi_hi_hi_20 = {dataGroup_15_20, dataGroup_14_20};
  wire [31:0]   res_lo_lo_hi_hi_20 = {res_lo_lo_hi_hi_hi_20, res_lo_lo_hi_hi_lo_20};
  wire [63:0]   res_lo_lo_hi_20 = {res_lo_lo_hi_hi_20, res_lo_lo_hi_lo_20};
  wire [127:0]  res_lo_lo_20 = {res_lo_lo_hi_20, res_lo_lo_lo_20};
  wire [15:0]   res_lo_hi_lo_lo_lo_20 = {dataGroup_17_20, dataGroup_16_20};
  wire [15:0]   res_lo_hi_lo_lo_hi_20 = {dataGroup_19_20, dataGroup_18_20};
  wire [31:0]   res_lo_hi_lo_lo_20 = {res_lo_hi_lo_lo_hi_20, res_lo_hi_lo_lo_lo_20};
  wire [15:0]   res_lo_hi_lo_hi_lo_20 = {dataGroup_21_20, dataGroup_20_20};
  wire [15:0]   res_lo_hi_lo_hi_hi_20 = {dataGroup_23_20, dataGroup_22_20};
  wire [31:0]   res_lo_hi_lo_hi_20 = {res_lo_hi_lo_hi_hi_20, res_lo_hi_lo_hi_lo_20};
  wire [63:0]   res_lo_hi_lo_20 = {res_lo_hi_lo_hi_20, res_lo_hi_lo_lo_20};
  wire [15:0]   res_lo_hi_hi_lo_lo_20 = {dataGroup_25_20, dataGroup_24_20};
  wire [15:0]   res_lo_hi_hi_lo_hi_20 = {dataGroup_27_20, dataGroup_26_20};
  wire [31:0]   res_lo_hi_hi_lo_20 = {res_lo_hi_hi_lo_hi_20, res_lo_hi_hi_lo_lo_20};
  wire [15:0]   res_lo_hi_hi_hi_lo_20 = {dataGroup_29_20, dataGroup_28_20};
  wire [15:0]   res_lo_hi_hi_hi_hi_20 = {dataGroup_31_20, dataGroup_30_20};
  wire [31:0]   res_lo_hi_hi_hi_20 = {res_lo_hi_hi_hi_hi_20, res_lo_hi_hi_hi_lo_20};
  wire [63:0]   res_lo_hi_hi_20 = {res_lo_hi_hi_hi_20, res_lo_hi_hi_lo_20};
  wire [127:0]  res_lo_hi_20 = {res_lo_hi_hi_20, res_lo_hi_lo_20};
  wire [255:0]  res_lo_20 = {res_lo_hi_20, res_lo_lo_20};
  wire [15:0]   res_hi_lo_lo_lo_lo_20 = {dataGroup_33_20, dataGroup_32_20};
  wire [15:0]   res_hi_lo_lo_lo_hi_20 = {dataGroup_35_20, dataGroup_34_20};
  wire [31:0]   res_hi_lo_lo_lo_20 = {res_hi_lo_lo_lo_hi_20, res_hi_lo_lo_lo_lo_20};
  wire [15:0]   res_hi_lo_lo_hi_lo_20 = {dataGroup_37_20, dataGroup_36_20};
  wire [15:0]   res_hi_lo_lo_hi_hi_20 = {dataGroup_39_20, dataGroup_38_20};
  wire [31:0]   res_hi_lo_lo_hi_20 = {res_hi_lo_lo_hi_hi_20, res_hi_lo_lo_hi_lo_20};
  wire [63:0]   res_hi_lo_lo_20 = {res_hi_lo_lo_hi_20, res_hi_lo_lo_lo_20};
  wire [15:0]   res_hi_lo_hi_lo_lo_20 = {dataGroup_41_20, dataGroup_40_20};
  wire [15:0]   res_hi_lo_hi_lo_hi_20 = {dataGroup_43_20, dataGroup_42_20};
  wire [31:0]   res_hi_lo_hi_lo_20 = {res_hi_lo_hi_lo_hi_20, res_hi_lo_hi_lo_lo_20};
  wire [15:0]   res_hi_lo_hi_hi_lo_20 = {dataGroup_45_20, dataGroup_44_20};
  wire [15:0]   res_hi_lo_hi_hi_hi_20 = {dataGroup_47_20, dataGroup_46_20};
  wire [31:0]   res_hi_lo_hi_hi_20 = {res_hi_lo_hi_hi_hi_20, res_hi_lo_hi_hi_lo_20};
  wire [63:0]   res_hi_lo_hi_20 = {res_hi_lo_hi_hi_20, res_hi_lo_hi_lo_20};
  wire [127:0]  res_hi_lo_20 = {res_hi_lo_hi_20, res_hi_lo_lo_20};
  wire [15:0]   res_hi_hi_lo_lo_lo_20 = {dataGroup_49_20, dataGroup_48_20};
  wire [15:0]   res_hi_hi_lo_lo_hi_20 = {dataGroup_51_20, dataGroup_50_20};
  wire [31:0]   res_hi_hi_lo_lo_20 = {res_hi_hi_lo_lo_hi_20, res_hi_hi_lo_lo_lo_20};
  wire [15:0]   res_hi_hi_lo_hi_lo_20 = {dataGroup_53_20, dataGroup_52_20};
  wire [15:0]   res_hi_hi_lo_hi_hi_20 = {dataGroup_55_20, dataGroup_54_20};
  wire [31:0]   res_hi_hi_lo_hi_20 = {res_hi_hi_lo_hi_hi_20, res_hi_hi_lo_hi_lo_20};
  wire [63:0]   res_hi_hi_lo_20 = {res_hi_hi_lo_hi_20, res_hi_hi_lo_lo_20};
  wire [15:0]   res_hi_hi_hi_lo_lo_20 = {dataGroup_57_20, dataGroup_56_20};
  wire [15:0]   res_hi_hi_hi_lo_hi_20 = {dataGroup_59_20, dataGroup_58_20};
  wire [31:0]   res_hi_hi_hi_lo_20 = {res_hi_hi_hi_lo_hi_20, res_hi_hi_hi_lo_lo_20};
  wire [15:0]   res_hi_hi_hi_hi_lo_20 = {dataGroup_61_20, dataGroup_60_20};
  wire [15:0]   res_hi_hi_hi_hi_hi_20 = {dataGroup_63_20, dataGroup_62_20};
  wire [31:0]   res_hi_hi_hi_hi_20 = {res_hi_hi_hi_hi_hi_20, res_hi_hi_hi_hi_lo_20};
  wire [63:0]   res_hi_hi_hi_20 = {res_hi_hi_hi_hi_20, res_hi_hi_hi_lo_20};
  wire [127:0]  res_hi_hi_20 = {res_hi_hi_hi_20, res_hi_hi_lo_20};
  wire [255:0]  res_hi_20 = {res_hi_hi_20, res_hi_lo_20};
  wire [511:0]  res_45 = {res_hi_20, res_lo_20};
  wire [1023:0] lo_lo_5 = {res_41, res_40};
  wire [1023:0] lo_hi_5 = {res_43, res_42};
  wire [2047:0] lo_5 = {lo_hi_5, lo_lo_5};
  wire [1023:0] hi_lo_5 = {res_45, res_44};
  wire [2047:0] hi_5 = {1024'h0, hi_lo_5};
  wire [4095:0] regroupLoadData_0_5 = {hi_5, lo_5};
  wire [2047:0] dataGroup_lo_1344 = {dataGroup_lo_hi_1344, dataGroup_lo_lo_1344};
  wire [2047:0] dataGroup_hi_1344 = {dataGroup_hi_hi_1344, dataGroup_hi_lo_1344};
  wire [7:0]    dataGroup_0_21 = dataGroup_lo_1344[7:0];
  wire [2047:0] dataGroup_lo_1345 = {dataGroup_lo_hi_1345, dataGroup_lo_lo_1345};
  wire [2047:0] dataGroup_hi_1345 = {dataGroup_hi_hi_1345, dataGroup_hi_lo_1345};
  wire [7:0]    dataGroup_1_21 = dataGroup_lo_1345[63:56];
  wire [2047:0] dataGroup_lo_1346 = {dataGroup_lo_hi_1346, dataGroup_lo_lo_1346};
  wire [2047:0] dataGroup_hi_1346 = {dataGroup_hi_hi_1346, dataGroup_hi_lo_1346};
  wire [7:0]    dataGroup_2_21 = dataGroup_lo_1346[119:112];
  wire [2047:0] dataGroup_lo_1347 = {dataGroup_lo_hi_1347, dataGroup_lo_lo_1347};
  wire [2047:0] dataGroup_hi_1347 = {dataGroup_hi_hi_1347, dataGroup_hi_lo_1347};
  wire [7:0]    dataGroup_3_21 = dataGroup_lo_1347[175:168];
  wire [2047:0] dataGroup_lo_1348 = {dataGroup_lo_hi_1348, dataGroup_lo_lo_1348};
  wire [2047:0] dataGroup_hi_1348 = {dataGroup_hi_hi_1348, dataGroup_hi_lo_1348};
  wire [7:0]    dataGroup_4_21 = dataGroup_lo_1348[231:224];
  wire [2047:0] dataGroup_lo_1349 = {dataGroup_lo_hi_1349, dataGroup_lo_lo_1349};
  wire [2047:0] dataGroup_hi_1349 = {dataGroup_hi_hi_1349, dataGroup_hi_lo_1349};
  wire [7:0]    dataGroup_5_21 = dataGroup_lo_1349[287:280];
  wire [2047:0] dataGroup_lo_1350 = {dataGroup_lo_hi_1350, dataGroup_lo_lo_1350};
  wire [2047:0] dataGroup_hi_1350 = {dataGroup_hi_hi_1350, dataGroup_hi_lo_1350};
  wire [7:0]    dataGroup_6_21 = dataGroup_lo_1350[343:336];
  wire [2047:0] dataGroup_lo_1351 = {dataGroup_lo_hi_1351, dataGroup_lo_lo_1351};
  wire [2047:0] dataGroup_hi_1351 = {dataGroup_hi_hi_1351, dataGroup_hi_lo_1351};
  wire [7:0]    dataGroup_7_21 = dataGroup_lo_1351[399:392];
  wire [2047:0] dataGroup_lo_1352 = {dataGroup_lo_hi_1352, dataGroup_lo_lo_1352};
  wire [2047:0] dataGroup_hi_1352 = {dataGroup_hi_hi_1352, dataGroup_hi_lo_1352};
  wire [7:0]    dataGroup_8_21 = dataGroup_lo_1352[455:448];
  wire [2047:0] dataGroup_lo_1353 = {dataGroup_lo_hi_1353, dataGroup_lo_lo_1353};
  wire [2047:0] dataGroup_hi_1353 = {dataGroup_hi_hi_1353, dataGroup_hi_lo_1353};
  wire [7:0]    dataGroup_9_21 = dataGroup_lo_1353[511:504];
  wire [2047:0] dataGroup_lo_1354 = {dataGroup_lo_hi_1354, dataGroup_lo_lo_1354};
  wire [2047:0] dataGroup_hi_1354 = {dataGroup_hi_hi_1354, dataGroup_hi_lo_1354};
  wire [7:0]    dataGroup_10_21 = dataGroup_lo_1354[567:560];
  wire [2047:0] dataGroup_lo_1355 = {dataGroup_lo_hi_1355, dataGroup_lo_lo_1355};
  wire [2047:0] dataGroup_hi_1355 = {dataGroup_hi_hi_1355, dataGroup_hi_lo_1355};
  wire [7:0]    dataGroup_11_21 = dataGroup_lo_1355[623:616];
  wire [2047:0] dataGroup_lo_1356 = {dataGroup_lo_hi_1356, dataGroup_lo_lo_1356};
  wire [2047:0] dataGroup_hi_1356 = {dataGroup_hi_hi_1356, dataGroup_hi_lo_1356};
  wire [7:0]    dataGroup_12_21 = dataGroup_lo_1356[679:672];
  wire [2047:0] dataGroup_lo_1357 = {dataGroup_lo_hi_1357, dataGroup_lo_lo_1357};
  wire [2047:0] dataGroup_hi_1357 = {dataGroup_hi_hi_1357, dataGroup_hi_lo_1357};
  wire [7:0]    dataGroup_13_21 = dataGroup_lo_1357[735:728];
  wire [2047:0] dataGroup_lo_1358 = {dataGroup_lo_hi_1358, dataGroup_lo_lo_1358};
  wire [2047:0] dataGroup_hi_1358 = {dataGroup_hi_hi_1358, dataGroup_hi_lo_1358};
  wire [7:0]    dataGroup_14_21 = dataGroup_lo_1358[791:784];
  wire [2047:0] dataGroup_lo_1359 = {dataGroup_lo_hi_1359, dataGroup_lo_lo_1359};
  wire [2047:0] dataGroup_hi_1359 = {dataGroup_hi_hi_1359, dataGroup_hi_lo_1359};
  wire [7:0]    dataGroup_15_21 = dataGroup_lo_1359[847:840];
  wire [2047:0] dataGroup_lo_1360 = {dataGroup_lo_hi_1360, dataGroup_lo_lo_1360};
  wire [2047:0] dataGroup_hi_1360 = {dataGroup_hi_hi_1360, dataGroup_hi_lo_1360};
  wire [7:0]    dataGroup_16_21 = dataGroup_lo_1360[903:896];
  wire [2047:0] dataGroup_lo_1361 = {dataGroup_lo_hi_1361, dataGroup_lo_lo_1361};
  wire [2047:0] dataGroup_hi_1361 = {dataGroup_hi_hi_1361, dataGroup_hi_lo_1361};
  wire [7:0]    dataGroup_17_21 = dataGroup_lo_1361[959:952];
  wire [2047:0] dataGroup_lo_1362 = {dataGroup_lo_hi_1362, dataGroup_lo_lo_1362};
  wire [2047:0] dataGroup_hi_1362 = {dataGroup_hi_hi_1362, dataGroup_hi_lo_1362};
  wire [7:0]    dataGroup_18_21 = dataGroup_lo_1362[1015:1008];
  wire [2047:0] dataGroup_lo_1363 = {dataGroup_lo_hi_1363, dataGroup_lo_lo_1363};
  wire [2047:0] dataGroup_hi_1363 = {dataGroup_hi_hi_1363, dataGroup_hi_lo_1363};
  wire [7:0]    dataGroup_19_21 = dataGroup_lo_1363[1071:1064];
  wire [2047:0] dataGroup_lo_1364 = {dataGroup_lo_hi_1364, dataGroup_lo_lo_1364};
  wire [2047:0] dataGroup_hi_1364 = {dataGroup_hi_hi_1364, dataGroup_hi_lo_1364};
  wire [7:0]    dataGroup_20_21 = dataGroup_lo_1364[1127:1120];
  wire [2047:0] dataGroup_lo_1365 = {dataGroup_lo_hi_1365, dataGroup_lo_lo_1365};
  wire [2047:0] dataGroup_hi_1365 = {dataGroup_hi_hi_1365, dataGroup_hi_lo_1365};
  wire [7:0]    dataGroup_21_21 = dataGroup_lo_1365[1183:1176];
  wire [2047:0] dataGroup_lo_1366 = {dataGroup_lo_hi_1366, dataGroup_lo_lo_1366};
  wire [2047:0] dataGroup_hi_1366 = {dataGroup_hi_hi_1366, dataGroup_hi_lo_1366};
  wire [7:0]    dataGroup_22_21 = dataGroup_lo_1366[1239:1232];
  wire [2047:0] dataGroup_lo_1367 = {dataGroup_lo_hi_1367, dataGroup_lo_lo_1367};
  wire [2047:0] dataGroup_hi_1367 = {dataGroup_hi_hi_1367, dataGroup_hi_lo_1367};
  wire [7:0]    dataGroup_23_21 = dataGroup_lo_1367[1295:1288];
  wire [2047:0] dataGroup_lo_1368 = {dataGroup_lo_hi_1368, dataGroup_lo_lo_1368};
  wire [2047:0] dataGroup_hi_1368 = {dataGroup_hi_hi_1368, dataGroup_hi_lo_1368};
  wire [7:0]    dataGroup_24_21 = dataGroup_lo_1368[1351:1344];
  wire [2047:0] dataGroup_lo_1369 = {dataGroup_lo_hi_1369, dataGroup_lo_lo_1369};
  wire [2047:0] dataGroup_hi_1369 = {dataGroup_hi_hi_1369, dataGroup_hi_lo_1369};
  wire [7:0]    dataGroup_25_21 = dataGroup_lo_1369[1407:1400];
  wire [2047:0] dataGroup_lo_1370 = {dataGroup_lo_hi_1370, dataGroup_lo_lo_1370};
  wire [2047:0] dataGroup_hi_1370 = {dataGroup_hi_hi_1370, dataGroup_hi_lo_1370};
  wire [7:0]    dataGroup_26_21 = dataGroup_lo_1370[1463:1456];
  wire [2047:0] dataGroup_lo_1371 = {dataGroup_lo_hi_1371, dataGroup_lo_lo_1371};
  wire [2047:0] dataGroup_hi_1371 = {dataGroup_hi_hi_1371, dataGroup_hi_lo_1371};
  wire [7:0]    dataGroup_27_21 = dataGroup_lo_1371[1519:1512];
  wire [2047:0] dataGroup_lo_1372 = {dataGroup_lo_hi_1372, dataGroup_lo_lo_1372};
  wire [2047:0] dataGroup_hi_1372 = {dataGroup_hi_hi_1372, dataGroup_hi_lo_1372};
  wire [7:0]    dataGroup_28_21 = dataGroup_lo_1372[1575:1568];
  wire [2047:0] dataGroup_lo_1373 = {dataGroup_lo_hi_1373, dataGroup_lo_lo_1373};
  wire [2047:0] dataGroup_hi_1373 = {dataGroup_hi_hi_1373, dataGroup_hi_lo_1373};
  wire [7:0]    dataGroup_29_21 = dataGroup_lo_1373[1631:1624];
  wire [2047:0] dataGroup_lo_1374 = {dataGroup_lo_hi_1374, dataGroup_lo_lo_1374};
  wire [2047:0] dataGroup_hi_1374 = {dataGroup_hi_hi_1374, dataGroup_hi_lo_1374};
  wire [7:0]    dataGroup_30_21 = dataGroup_lo_1374[1687:1680];
  wire [2047:0] dataGroup_lo_1375 = {dataGroup_lo_hi_1375, dataGroup_lo_lo_1375};
  wire [2047:0] dataGroup_hi_1375 = {dataGroup_hi_hi_1375, dataGroup_hi_lo_1375};
  wire [7:0]    dataGroup_31_21 = dataGroup_lo_1375[1743:1736];
  wire [2047:0] dataGroup_lo_1376 = {dataGroup_lo_hi_1376, dataGroup_lo_lo_1376};
  wire [2047:0] dataGroup_hi_1376 = {dataGroup_hi_hi_1376, dataGroup_hi_lo_1376};
  wire [7:0]    dataGroup_32_21 = dataGroup_lo_1376[1799:1792];
  wire [2047:0] dataGroup_lo_1377 = {dataGroup_lo_hi_1377, dataGroup_lo_lo_1377};
  wire [2047:0] dataGroup_hi_1377 = {dataGroup_hi_hi_1377, dataGroup_hi_lo_1377};
  wire [7:0]    dataGroup_33_21 = dataGroup_lo_1377[1855:1848];
  wire [2047:0] dataGroup_lo_1378 = {dataGroup_lo_hi_1378, dataGroup_lo_lo_1378};
  wire [2047:0] dataGroup_hi_1378 = {dataGroup_hi_hi_1378, dataGroup_hi_lo_1378};
  wire [7:0]    dataGroup_34_21 = dataGroup_lo_1378[1911:1904];
  wire [2047:0] dataGroup_lo_1379 = {dataGroup_lo_hi_1379, dataGroup_lo_lo_1379};
  wire [2047:0] dataGroup_hi_1379 = {dataGroup_hi_hi_1379, dataGroup_hi_lo_1379};
  wire [7:0]    dataGroup_35_21 = dataGroup_lo_1379[1967:1960];
  wire [2047:0] dataGroup_lo_1380 = {dataGroup_lo_hi_1380, dataGroup_lo_lo_1380};
  wire [2047:0] dataGroup_hi_1380 = {dataGroup_hi_hi_1380, dataGroup_hi_lo_1380};
  wire [7:0]    dataGroup_36_21 = dataGroup_lo_1380[2023:2016];
  wire [2047:0] dataGroup_lo_1381 = {dataGroup_lo_hi_1381, dataGroup_lo_lo_1381};
  wire [2047:0] dataGroup_hi_1381 = {dataGroup_hi_hi_1381, dataGroup_hi_lo_1381};
  wire [7:0]    dataGroup_37_21 = dataGroup_hi_1381[31:24];
  wire [2047:0] dataGroup_lo_1382 = {dataGroup_lo_hi_1382, dataGroup_lo_lo_1382};
  wire [2047:0] dataGroup_hi_1382 = {dataGroup_hi_hi_1382, dataGroup_hi_lo_1382};
  wire [7:0]    dataGroup_38_21 = dataGroup_hi_1382[87:80];
  wire [2047:0] dataGroup_lo_1383 = {dataGroup_lo_hi_1383, dataGroup_lo_lo_1383};
  wire [2047:0] dataGroup_hi_1383 = {dataGroup_hi_hi_1383, dataGroup_hi_lo_1383};
  wire [7:0]    dataGroup_39_21 = dataGroup_hi_1383[143:136];
  wire [2047:0] dataGroup_lo_1384 = {dataGroup_lo_hi_1384, dataGroup_lo_lo_1384};
  wire [2047:0] dataGroup_hi_1384 = {dataGroup_hi_hi_1384, dataGroup_hi_lo_1384};
  wire [7:0]    dataGroup_40_21 = dataGroup_hi_1384[199:192];
  wire [2047:0] dataGroup_lo_1385 = {dataGroup_lo_hi_1385, dataGroup_lo_lo_1385};
  wire [2047:0] dataGroup_hi_1385 = {dataGroup_hi_hi_1385, dataGroup_hi_lo_1385};
  wire [7:0]    dataGroup_41_21 = dataGroup_hi_1385[255:248];
  wire [2047:0] dataGroup_lo_1386 = {dataGroup_lo_hi_1386, dataGroup_lo_lo_1386};
  wire [2047:0] dataGroup_hi_1386 = {dataGroup_hi_hi_1386, dataGroup_hi_lo_1386};
  wire [7:0]    dataGroup_42_21 = dataGroup_hi_1386[311:304];
  wire [2047:0] dataGroup_lo_1387 = {dataGroup_lo_hi_1387, dataGroup_lo_lo_1387};
  wire [2047:0] dataGroup_hi_1387 = {dataGroup_hi_hi_1387, dataGroup_hi_lo_1387};
  wire [7:0]    dataGroup_43_21 = dataGroup_hi_1387[367:360];
  wire [2047:0] dataGroup_lo_1388 = {dataGroup_lo_hi_1388, dataGroup_lo_lo_1388};
  wire [2047:0] dataGroup_hi_1388 = {dataGroup_hi_hi_1388, dataGroup_hi_lo_1388};
  wire [7:0]    dataGroup_44_21 = dataGroup_hi_1388[423:416];
  wire [2047:0] dataGroup_lo_1389 = {dataGroup_lo_hi_1389, dataGroup_lo_lo_1389};
  wire [2047:0] dataGroup_hi_1389 = {dataGroup_hi_hi_1389, dataGroup_hi_lo_1389};
  wire [7:0]    dataGroup_45_21 = dataGroup_hi_1389[479:472];
  wire [2047:0] dataGroup_lo_1390 = {dataGroup_lo_hi_1390, dataGroup_lo_lo_1390};
  wire [2047:0] dataGroup_hi_1390 = {dataGroup_hi_hi_1390, dataGroup_hi_lo_1390};
  wire [7:0]    dataGroup_46_21 = dataGroup_hi_1390[535:528];
  wire [2047:0] dataGroup_lo_1391 = {dataGroup_lo_hi_1391, dataGroup_lo_lo_1391};
  wire [2047:0] dataGroup_hi_1391 = {dataGroup_hi_hi_1391, dataGroup_hi_lo_1391};
  wire [7:0]    dataGroup_47_21 = dataGroup_hi_1391[591:584];
  wire [2047:0] dataGroup_lo_1392 = {dataGroup_lo_hi_1392, dataGroup_lo_lo_1392};
  wire [2047:0] dataGroup_hi_1392 = {dataGroup_hi_hi_1392, dataGroup_hi_lo_1392};
  wire [7:0]    dataGroup_48_21 = dataGroup_hi_1392[647:640];
  wire [2047:0] dataGroup_lo_1393 = {dataGroup_lo_hi_1393, dataGroup_lo_lo_1393};
  wire [2047:0] dataGroup_hi_1393 = {dataGroup_hi_hi_1393, dataGroup_hi_lo_1393};
  wire [7:0]    dataGroup_49_21 = dataGroup_hi_1393[703:696];
  wire [2047:0] dataGroup_lo_1394 = {dataGroup_lo_hi_1394, dataGroup_lo_lo_1394};
  wire [2047:0] dataGroup_hi_1394 = {dataGroup_hi_hi_1394, dataGroup_hi_lo_1394};
  wire [7:0]    dataGroup_50_21 = dataGroup_hi_1394[759:752];
  wire [2047:0] dataGroup_lo_1395 = {dataGroup_lo_hi_1395, dataGroup_lo_lo_1395};
  wire [2047:0] dataGroup_hi_1395 = {dataGroup_hi_hi_1395, dataGroup_hi_lo_1395};
  wire [7:0]    dataGroup_51_21 = dataGroup_hi_1395[815:808];
  wire [2047:0] dataGroup_lo_1396 = {dataGroup_lo_hi_1396, dataGroup_lo_lo_1396};
  wire [2047:0] dataGroup_hi_1396 = {dataGroup_hi_hi_1396, dataGroup_hi_lo_1396};
  wire [7:0]    dataGroup_52_21 = dataGroup_hi_1396[871:864];
  wire [2047:0] dataGroup_lo_1397 = {dataGroup_lo_hi_1397, dataGroup_lo_lo_1397};
  wire [2047:0] dataGroup_hi_1397 = {dataGroup_hi_hi_1397, dataGroup_hi_lo_1397};
  wire [7:0]    dataGroup_53_21 = dataGroup_hi_1397[927:920];
  wire [2047:0] dataGroup_lo_1398 = {dataGroup_lo_hi_1398, dataGroup_lo_lo_1398};
  wire [2047:0] dataGroup_hi_1398 = {dataGroup_hi_hi_1398, dataGroup_hi_lo_1398};
  wire [7:0]    dataGroup_54_21 = dataGroup_hi_1398[983:976];
  wire [2047:0] dataGroup_lo_1399 = {dataGroup_lo_hi_1399, dataGroup_lo_lo_1399};
  wire [2047:0] dataGroup_hi_1399 = {dataGroup_hi_hi_1399, dataGroup_hi_lo_1399};
  wire [7:0]    dataGroup_55_21 = dataGroup_hi_1399[1039:1032];
  wire [2047:0] dataGroup_lo_1400 = {dataGroup_lo_hi_1400, dataGroup_lo_lo_1400};
  wire [2047:0] dataGroup_hi_1400 = {dataGroup_hi_hi_1400, dataGroup_hi_lo_1400};
  wire [7:0]    dataGroup_56_21 = dataGroup_hi_1400[1095:1088];
  wire [2047:0] dataGroup_lo_1401 = {dataGroup_lo_hi_1401, dataGroup_lo_lo_1401};
  wire [2047:0] dataGroup_hi_1401 = {dataGroup_hi_hi_1401, dataGroup_hi_lo_1401};
  wire [7:0]    dataGroup_57_21 = dataGroup_hi_1401[1151:1144];
  wire [2047:0] dataGroup_lo_1402 = {dataGroup_lo_hi_1402, dataGroup_lo_lo_1402};
  wire [2047:0] dataGroup_hi_1402 = {dataGroup_hi_hi_1402, dataGroup_hi_lo_1402};
  wire [7:0]    dataGroup_58_21 = dataGroup_hi_1402[1207:1200];
  wire [2047:0] dataGroup_lo_1403 = {dataGroup_lo_hi_1403, dataGroup_lo_lo_1403};
  wire [2047:0] dataGroup_hi_1403 = {dataGroup_hi_hi_1403, dataGroup_hi_lo_1403};
  wire [7:0]    dataGroup_59_21 = dataGroup_hi_1403[1263:1256];
  wire [2047:0] dataGroup_lo_1404 = {dataGroup_lo_hi_1404, dataGroup_lo_lo_1404};
  wire [2047:0] dataGroup_hi_1404 = {dataGroup_hi_hi_1404, dataGroup_hi_lo_1404};
  wire [7:0]    dataGroup_60_21 = dataGroup_hi_1404[1319:1312];
  wire [2047:0] dataGroup_lo_1405 = {dataGroup_lo_hi_1405, dataGroup_lo_lo_1405};
  wire [2047:0] dataGroup_hi_1405 = {dataGroup_hi_hi_1405, dataGroup_hi_lo_1405};
  wire [7:0]    dataGroup_61_21 = dataGroup_hi_1405[1375:1368];
  wire [2047:0] dataGroup_lo_1406 = {dataGroup_lo_hi_1406, dataGroup_lo_lo_1406};
  wire [2047:0] dataGroup_hi_1406 = {dataGroup_hi_hi_1406, dataGroup_hi_lo_1406};
  wire [7:0]    dataGroup_62_21 = dataGroup_hi_1406[1431:1424];
  wire [2047:0] dataGroup_lo_1407 = {dataGroup_lo_hi_1407, dataGroup_lo_lo_1407};
  wire [2047:0] dataGroup_hi_1407 = {dataGroup_hi_hi_1407, dataGroup_hi_lo_1407};
  wire [7:0]    dataGroup_63_21 = dataGroup_hi_1407[1487:1480];
  wire [15:0]   res_lo_lo_lo_lo_lo_21 = {dataGroup_1_21, dataGroup_0_21};
  wire [15:0]   res_lo_lo_lo_lo_hi_21 = {dataGroup_3_21, dataGroup_2_21};
  wire [31:0]   res_lo_lo_lo_lo_21 = {res_lo_lo_lo_lo_hi_21, res_lo_lo_lo_lo_lo_21};
  wire [15:0]   res_lo_lo_lo_hi_lo_21 = {dataGroup_5_21, dataGroup_4_21};
  wire [15:0]   res_lo_lo_lo_hi_hi_21 = {dataGroup_7_21, dataGroup_6_21};
  wire [31:0]   res_lo_lo_lo_hi_21 = {res_lo_lo_lo_hi_hi_21, res_lo_lo_lo_hi_lo_21};
  wire [63:0]   res_lo_lo_lo_21 = {res_lo_lo_lo_hi_21, res_lo_lo_lo_lo_21};
  wire [15:0]   res_lo_lo_hi_lo_lo_21 = {dataGroup_9_21, dataGroup_8_21};
  wire [15:0]   res_lo_lo_hi_lo_hi_21 = {dataGroup_11_21, dataGroup_10_21};
  wire [31:0]   res_lo_lo_hi_lo_21 = {res_lo_lo_hi_lo_hi_21, res_lo_lo_hi_lo_lo_21};
  wire [15:0]   res_lo_lo_hi_hi_lo_21 = {dataGroup_13_21, dataGroup_12_21};
  wire [15:0]   res_lo_lo_hi_hi_hi_21 = {dataGroup_15_21, dataGroup_14_21};
  wire [31:0]   res_lo_lo_hi_hi_21 = {res_lo_lo_hi_hi_hi_21, res_lo_lo_hi_hi_lo_21};
  wire [63:0]   res_lo_lo_hi_21 = {res_lo_lo_hi_hi_21, res_lo_lo_hi_lo_21};
  wire [127:0]  res_lo_lo_21 = {res_lo_lo_hi_21, res_lo_lo_lo_21};
  wire [15:0]   res_lo_hi_lo_lo_lo_21 = {dataGroup_17_21, dataGroup_16_21};
  wire [15:0]   res_lo_hi_lo_lo_hi_21 = {dataGroup_19_21, dataGroup_18_21};
  wire [31:0]   res_lo_hi_lo_lo_21 = {res_lo_hi_lo_lo_hi_21, res_lo_hi_lo_lo_lo_21};
  wire [15:0]   res_lo_hi_lo_hi_lo_21 = {dataGroup_21_21, dataGroup_20_21};
  wire [15:0]   res_lo_hi_lo_hi_hi_21 = {dataGroup_23_21, dataGroup_22_21};
  wire [31:0]   res_lo_hi_lo_hi_21 = {res_lo_hi_lo_hi_hi_21, res_lo_hi_lo_hi_lo_21};
  wire [63:0]   res_lo_hi_lo_21 = {res_lo_hi_lo_hi_21, res_lo_hi_lo_lo_21};
  wire [15:0]   res_lo_hi_hi_lo_lo_21 = {dataGroup_25_21, dataGroup_24_21};
  wire [15:0]   res_lo_hi_hi_lo_hi_21 = {dataGroup_27_21, dataGroup_26_21};
  wire [31:0]   res_lo_hi_hi_lo_21 = {res_lo_hi_hi_lo_hi_21, res_lo_hi_hi_lo_lo_21};
  wire [15:0]   res_lo_hi_hi_hi_lo_21 = {dataGroup_29_21, dataGroup_28_21};
  wire [15:0]   res_lo_hi_hi_hi_hi_21 = {dataGroup_31_21, dataGroup_30_21};
  wire [31:0]   res_lo_hi_hi_hi_21 = {res_lo_hi_hi_hi_hi_21, res_lo_hi_hi_hi_lo_21};
  wire [63:0]   res_lo_hi_hi_21 = {res_lo_hi_hi_hi_21, res_lo_hi_hi_lo_21};
  wire [127:0]  res_lo_hi_21 = {res_lo_hi_hi_21, res_lo_hi_lo_21};
  wire [255:0]  res_lo_21 = {res_lo_hi_21, res_lo_lo_21};
  wire [15:0]   res_hi_lo_lo_lo_lo_21 = {dataGroup_33_21, dataGroup_32_21};
  wire [15:0]   res_hi_lo_lo_lo_hi_21 = {dataGroup_35_21, dataGroup_34_21};
  wire [31:0]   res_hi_lo_lo_lo_21 = {res_hi_lo_lo_lo_hi_21, res_hi_lo_lo_lo_lo_21};
  wire [15:0]   res_hi_lo_lo_hi_lo_21 = {dataGroup_37_21, dataGroup_36_21};
  wire [15:0]   res_hi_lo_lo_hi_hi_21 = {dataGroup_39_21, dataGroup_38_21};
  wire [31:0]   res_hi_lo_lo_hi_21 = {res_hi_lo_lo_hi_hi_21, res_hi_lo_lo_hi_lo_21};
  wire [63:0]   res_hi_lo_lo_21 = {res_hi_lo_lo_hi_21, res_hi_lo_lo_lo_21};
  wire [15:0]   res_hi_lo_hi_lo_lo_21 = {dataGroup_41_21, dataGroup_40_21};
  wire [15:0]   res_hi_lo_hi_lo_hi_21 = {dataGroup_43_21, dataGroup_42_21};
  wire [31:0]   res_hi_lo_hi_lo_21 = {res_hi_lo_hi_lo_hi_21, res_hi_lo_hi_lo_lo_21};
  wire [15:0]   res_hi_lo_hi_hi_lo_21 = {dataGroup_45_21, dataGroup_44_21};
  wire [15:0]   res_hi_lo_hi_hi_hi_21 = {dataGroup_47_21, dataGroup_46_21};
  wire [31:0]   res_hi_lo_hi_hi_21 = {res_hi_lo_hi_hi_hi_21, res_hi_lo_hi_hi_lo_21};
  wire [63:0]   res_hi_lo_hi_21 = {res_hi_lo_hi_hi_21, res_hi_lo_hi_lo_21};
  wire [127:0]  res_hi_lo_21 = {res_hi_lo_hi_21, res_hi_lo_lo_21};
  wire [15:0]   res_hi_hi_lo_lo_lo_21 = {dataGroup_49_21, dataGroup_48_21};
  wire [15:0]   res_hi_hi_lo_lo_hi_21 = {dataGroup_51_21, dataGroup_50_21};
  wire [31:0]   res_hi_hi_lo_lo_21 = {res_hi_hi_lo_lo_hi_21, res_hi_hi_lo_lo_lo_21};
  wire [15:0]   res_hi_hi_lo_hi_lo_21 = {dataGroup_53_21, dataGroup_52_21};
  wire [15:0]   res_hi_hi_lo_hi_hi_21 = {dataGroup_55_21, dataGroup_54_21};
  wire [31:0]   res_hi_hi_lo_hi_21 = {res_hi_hi_lo_hi_hi_21, res_hi_hi_lo_hi_lo_21};
  wire [63:0]   res_hi_hi_lo_21 = {res_hi_hi_lo_hi_21, res_hi_hi_lo_lo_21};
  wire [15:0]   res_hi_hi_hi_lo_lo_21 = {dataGroup_57_21, dataGroup_56_21};
  wire [15:0]   res_hi_hi_hi_lo_hi_21 = {dataGroup_59_21, dataGroup_58_21};
  wire [31:0]   res_hi_hi_hi_lo_21 = {res_hi_hi_hi_lo_hi_21, res_hi_hi_hi_lo_lo_21};
  wire [15:0]   res_hi_hi_hi_hi_lo_21 = {dataGroup_61_21, dataGroup_60_21};
  wire [15:0]   res_hi_hi_hi_hi_hi_21 = {dataGroup_63_21, dataGroup_62_21};
  wire [31:0]   res_hi_hi_hi_hi_21 = {res_hi_hi_hi_hi_hi_21, res_hi_hi_hi_hi_lo_21};
  wire [63:0]   res_hi_hi_hi_21 = {res_hi_hi_hi_hi_21, res_hi_hi_hi_lo_21};
  wire [127:0]  res_hi_hi_21 = {res_hi_hi_hi_21, res_hi_hi_lo_21};
  wire [255:0]  res_hi_21 = {res_hi_hi_21, res_hi_lo_21};
  wire [511:0]  res_48 = {res_hi_21, res_lo_21};
  wire [2047:0] dataGroup_lo_1408 = {dataGroup_lo_hi_1408, dataGroup_lo_lo_1408};
  wire [2047:0] dataGroup_hi_1408 = {dataGroup_hi_hi_1408, dataGroup_hi_lo_1408};
  wire [7:0]    dataGroup_0_22 = dataGroup_lo_1408[15:8];
  wire [2047:0] dataGroup_lo_1409 = {dataGroup_lo_hi_1409, dataGroup_lo_lo_1409};
  wire [2047:0] dataGroup_hi_1409 = {dataGroup_hi_hi_1409, dataGroup_hi_lo_1409};
  wire [7:0]    dataGroup_1_22 = dataGroup_lo_1409[71:64];
  wire [2047:0] dataGroup_lo_1410 = {dataGroup_lo_hi_1410, dataGroup_lo_lo_1410};
  wire [2047:0] dataGroup_hi_1410 = {dataGroup_hi_hi_1410, dataGroup_hi_lo_1410};
  wire [7:0]    dataGroup_2_22 = dataGroup_lo_1410[127:120];
  wire [2047:0] dataGroup_lo_1411 = {dataGroup_lo_hi_1411, dataGroup_lo_lo_1411};
  wire [2047:0] dataGroup_hi_1411 = {dataGroup_hi_hi_1411, dataGroup_hi_lo_1411};
  wire [7:0]    dataGroup_3_22 = dataGroup_lo_1411[183:176];
  wire [2047:0] dataGroup_lo_1412 = {dataGroup_lo_hi_1412, dataGroup_lo_lo_1412};
  wire [2047:0] dataGroup_hi_1412 = {dataGroup_hi_hi_1412, dataGroup_hi_lo_1412};
  wire [7:0]    dataGroup_4_22 = dataGroup_lo_1412[239:232];
  wire [2047:0] dataGroup_lo_1413 = {dataGroup_lo_hi_1413, dataGroup_lo_lo_1413};
  wire [2047:0] dataGroup_hi_1413 = {dataGroup_hi_hi_1413, dataGroup_hi_lo_1413};
  wire [7:0]    dataGroup_5_22 = dataGroup_lo_1413[295:288];
  wire [2047:0] dataGroup_lo_1414 = {dataGroup_lo_hi_1414, dataGroup_lo_lo_1414};
  wire [2047:0] dataGroup_hi_1414 = {dataGroup_hi_hi_1414, dataGroup_hi_lo_1414};
  wire [7:0]    dataGroup_6_22 = dataGroup_lo_1414[351:344];
  wire [2047:0] dataGroup_lo_1415 = {dataGroup_lo_hi_1415, dataGroup_lo_lo_1415};
  wire [2047:0] dataGroup_hi_1415 = {dataGroup_hi_hi_1415, dataGroup_hi_lo_1415};
  wire [7:0]    dataGroup_7_22 = dataGroup_lo_1415[407:400];
  wire [2047:0] dataGroup_lo_1416 = {dataGroup_lo_hi_1416, dataGroup_lo_lo_1416};
  wire [2047:0] dataGroup_hi_1416 = {dataGroup_hi_hi_1416, dataGroup_hi_lo_1416};
  wire [7:0]    dataGroup_8_22 = dataGroup_lo_1416[463:456];
  wire [2047:0] dataGroup_lo_1417 = {dataGroup_lo_hi_1417, dataGroup_lo_lo_1417};
  wire [2047:0] dataGroup_hi_1417 = {dataGroup_hi_hi_1417, dataGroup_hi_lo_1417};
  wire [7:0]    dataGroup_9_22 = dataGroup_lo_1417[519:512];
  wire [2047:0] dataGroup_lo_1418 = {dataGroup_lo_hi_1418, dataGroup_lo_lo_1418};
  wire [2047:0] dataGroup_hi_1418 = {dataGroup_hi_hi_1418, dataGroup_hi_lo_1418};
  wire [7:0]    dataGroup_10_22 = dataGroup_lo_1418[575:568];
  wire [2047:0] dataGroup_lo_1419 = {dataGroup_lo_hi_1419, dataGroup_lo_lo_1419};
  wire [2047:0] dataGroup_hi_1419 = {dataGroup_hi_hi_1419, dataGroup_hi_lo_1419};
  wire [7:0]    dataGroup_11_22 = dataGroup_lo_1419[631:624];
  wire [2047:0] dataGroup_lo_1420 = {dataGroup_lo_hi_1420, dataGroup_lo_lo_1420};
  wire [2047:0] dataGroup_hi_1420 = {dataGroup_hi_hi_1420, dataGroup_hi_lo_1420};
  wire [7:0]    dataGroup_12_22 = dataGroup_lo_1420[687:680];
  wire [2047:0] dataGroup_lo_1421 = {dataGroup_lo_hi_1421, dataGroup_lo_lo_1421};
  wire [2047:0] dataGroup_hi_1421 = {dataGroup_hi_hi_1421, dataGroup_hi_lo_1421};
  wire [7:0]    dataGroup_13_22 = dataGroup_lo_1421[743:736];
  wire [2047:0] dataGroup_lo_1422 = {dataGroup_lo_hi_1422, dataGroup_lo_lo_1422};
  wire [2047:0] dataGroup_hi_1422 = {dataGroup_hi_hi_1422, dataGroup_hi_lo_1422};
  wire [7:0]    dataGroup_14_22 = dataGroup_lo_1422[799:792];
  wire [2047:0] dataGroup_lo_1423 = {dataGroup_lo_hi_1423, dataGroup_lo_lo_1423};
  wire [2047:0] dataGroup_hi_1423 = {dataGroup_hi_hi_1423, dataGroup_hi_lo_1423};
  wire [7:0]    dataGroup_15_22 = dataGroup_lo_1423[855:848];
  wire [2047:0] dataGroup_lo_1424 = {dataGroup_lo_hi_1424, dataGroup_lo_lo_1424};
  wire [2047:0] dataGroup_hi_1424 = {dataGroup_hi_hi_1424, dataGroup_hi_lo_1424};
  wire [7:0]    dataGroup_16_22 = dataGroup_lo_1424[911:904];
  wire [2047:0] dataGroup_lo_1425 = {dataGroup_lo_hi_1425, dataGroup_lo_lo_1425};
  wire [2047:0] dataGroup_hi_1425 = {dataGroup_hi_hi_1425, dataGroup_hi_lo_1425};
  wire [7:0]    dataGroup_17_22 = dataGroup_lo_1425[967:960];
  wire [2047:0] dataGroup_lo_1426 = {dataGroup_lo_hi_1426, dataGroup_lo_lo_1426};
  wire [2047:0] dataGroup_hi_1426 = {dataGroup_hi_hi_1426, dataGroup_hi_lo_1426};
  wire [7:0]    dataGroup_18_22 = dataGroup_lo_1426[1023:1016];
  wire [2047:0] dataGroup_lo_1427 = {dataGroup_lo_hi_1427, dataGroup_lo_lo_1427};
  wire [2047:0] dataGroup_hi_1427 = {dataGroup_hi_hi_1427, dataGroup_hi_lo_1427};
  wire [7:0]    dataGroup_19_22 = dataGroup_lo_1427[1079:1072];
  wire [2047:0] dataGroup_lo_1428 = {dataGroup_lo_hi_1428, dataGroup_lo_lo_1428};
  wire [2047:0] dataGroup_hi_1428 = {dataGroup_hi_hi_1428, dataGroup_hi_lo_1428};
  wire [7:0]    dataGroup_20_22 = dataGroup_lo_1428[1135:1128];
  wire [2047:0] dataGroup_lo_1429 = {dataGroup_lo_hi_1429, dataGroup_lo_lo_1429};
  wire [2047:0] dataGroup_hi_1429 = {dataGroup_hi_hi_1429, dataGroup_hi_lo_1429};
  wire [7:0]    dataGroup_21_22 = dataGroup_lo_1429[1191:1184];
  wire [2047:0] dataGroup_lo_1430 = {dataGroup_lo_hi_1430, dataGroup_lo_lo_1430};
  wire [2047:0] dataGroup_hi_1430 = {dataGroup_hi_hi_1430, dataGroup_hi_lo_1430};
  wire [7:0]    dataGroup_22_22 = dataGroup_lo_1430[1247:1240];
  wire [2047:0] dataGroup_lo_1431 = {dataGroup_lo_hi_1431, dataGroup_lo_lo_1431};
  wire [2047:0] dataGroup_hi_1431 = {dataGroup_hi_hi_1431, dataGroup_hi_lo_1431};
  wire [7:0]    dataGroup_23_22 = dataGroup_lo_1431[1303:1296];
  wire [2047:0] dataGroup_lo_1432 = {dataGroup_lo_hi_1432, dataGroup_lo_lo_1432};
  wire [2047:0] dataGroup_hi_1432 = {dataGroup_hi_hi_1432, dataGroup_hi_lo_1432};
  wire [7:0]    dataGroup_24_22 = dataGroup_lo_1432[1359:1352];
  wire [2047:0] dataGroup_lo_1433 = {dataGroup_lo_hi_1433, dataGroup_lo_lo_1433};
  wire [2047:0] dataGroup_hi_1433 = {dataGroup_hi_hi_1433, dataGroup_hi_lo_1433};
  wire [7:0]    dataGroup_25_22 = dataGroup_lo_1433[1415:1408];
  wire [2047:0] dataGroup_lo_1434 = {dataGroup_lo_hi_1434, dataGroup_lo_lo_1434};
  wire [2047:0] dataGroup_hi_1434 = {dataGroup_hi_hi_1434, dataGroup_hi_lo_1434};
  wire [7:0]    dataGroup_26_22 = dataGroup_lo_1434[1471:1464];
  wire [2047:0] dataGroup_lo_1435 = {dataGroup_lo_hi_1435, dataGroup_lo_lo_1435};
  wire [2047:0] dataGroup_hi_1435 = {dataGroup_hi_hi_1435, dataGroup_hi_lo_1435};
  wire [7:0]    dataGroup_27_22 = dataGroup_lo_1435[1527:1520];
  wire [2047:0] dataGroup_lo_1436 = {dataGroup_lo_hi_1436, dataGroup_lo_lo_1436};
  wire [2047:0] dataGroup_hi_1436 = {dataGroup_hi_hi_1436, dataGroup_hi_lo_1436};
  wire [7:0]    dataGroup_28_22 = dataGroup_lo_1436[1583:1576];
  wire [2047:0] dataGroup_lo_1437 = {dataGroup_lo_hi_1437, dataGroup_lo_lo_1437};
  wire [2047:0] dataGroup_hi_1437 = {dataGroup_hi_hi_1437, dataGroup_hi_lo_1437};
  wire [7:0]    dataGroup_29_22 = dataGroup_lo_1437[1639:1632];
  wire [2047:0] dataGroup_lo_1438 = {dataGroup_lo_hi_1438, dataGroup_lo_lo_1438};
  wire [2047:0] dataGroup_hi_1438 = {dataGroup_hi_hi_1438, dataGroup_hi_lo_1438};
  wire [7:0]    dataGroup_30_22 = dataGroup_lo_1438[1695:1688];
  wire [2047:0] dataGroup_lo_1439 = {dataGroup_lo_hi_1439, dataGroup_lo_lo_1439};
  wire [2047:0] dataGroup_hi_1439 = {dataGroup_hi_hi_1439, dataGroup_hi_lo_1439};
  wire [7:0]    dataGroup_31_22 = dataGroup_lo_1439[1751:1744];
  wire [2047:0] dataGroup_lo_1440 = {dataGroup_lo_hi_1440, dataGroup_lo_lo_1440};
  wire [2047:0] dataGroup_hi_1440 = {dataGroup_hi_hi_1440, dataGroup_hi_lo_1440};
  wire [7:0]    dataGroup_32_22 = dataGroup_lo_1440[1807:1800];
  wire [2047:0] dataGroup_lo_1441 = {dataGroup_lo_hi_1441, dataGroup_lo_lo_1441};
  wire [2047:0] dataGroup_hi_1441 = {dataGroup_hi_hi_1441, dataGroup_hi_lo_1441};
  wire [7:0]    dataGroup_33_22 = dataGroup_lo_1441[1863:1856];
  wire [2047:0] dataGroup_lo_1442 = {dataGroup_lo_hi_1442, dataGroup_lo_lo_1442};
  wire [2047:0] dataGroup_hi_1442 = {dataGroup_hi_hi_1442, dataGroup_hi_lo_1442};
  wire [7:0]    dataGroup_34_22 = dataGroup_lo_1442[1919:1912];
  wire [2047:0] dataGroup_lo_1443 = {dataGroup_lo_hi_1443, dataGroup_lo_lo_1443};
  wire [2047:0] dataGroup_hi_1443 = {dataGroup_hi_hi_1443, dataGroup_hi_lo_1443};
  wire [7:0]    dataGroup_35_22 = dataGroup_lo_1443[1975:1968];
  wire [2047:0] dataGroup_lo_1444 = {dataGroup_lo_hi_1444, dataGroup_lo_lo_1444};
  wire [2047:0] dataGroup_hi_1444 = {dataGroup_hi_hi_1444, dataGroup_hi_lo_1444};
  wire [7:0]    dataGroup_36_22 = dataGroup_lo_1444[2031:2024];
  wire [2047:0] dataGroup_lo_1445 = {dataGroup_lo_hi_1445, dataGroup_lo_lo_1445};
  wire [2047:0] dataGroup_hi_1445 = {dataGroup_hi_hi_1445, dataGroup_hi_lo_1445};
  wire [7:0]    dataGroup_37_22 = dataGroup_hi_1445[39:32];
  wire [2047:0] dataGroup_lo_1446 = {dataGroup_lo_hi_1446, dataGroup_lo_lo_1446};
  wire [2047:0] dataGroup_hi_1446 = {dataGroup_hi_hi_1446, dataGroup_hi_lo_1446};
  wire [7:0]    dataGroup_38_22 = dataGroup_hi_1446[95:88];
  wire [2047:0] dataGroup_lo_1447 = {dataGroup_lo_hi_1447, dataGroup_lo_lo_1447};
  wire [2047:0] dataGroup_hi_1447 = {dataGroup_hi_hi_1447, dataGroup_hi_lo_1447};
  wire [7:0]    dataGroup_39_22 = dataGroup_hi_1447[151:144];
  wire [2047:0] dataGroup_lo_1448 = {dataGroup_lo_hi_1448, dataGroup_lo_lo_1448};
  wire [2047:0] dataGroup_hi_1448 = {dataGroup_hi_hi_1448, dataGroup_hi_lo_1448};
  wire [7:0]    dataGroup_40_22 = dataGroup_hi_1448[207:200];
  wire [2047:0] dataGroup_lo_1449 = {dataGroup_lo_hi_1449, dataGroup_lo_lo_1449};
  wire [2047:0] dataGroup_hi_1449 = {dataGroup_hi_hi_1449, dataGroup_hi_lo_1449};
  wire [7:0]    dataGroup_41_22 = dataGroup_hi_1449[263:256];
  wire [2047:0] dataGroup_lo_1450 = {dataGroup_lo_hi_1450, dataGroup_lo_lo_1450};
  wire [2047:0] dataGroup_hi_1450 = {dataGroup_hi_hi_1450, dataGroup_hi_lo_1450};
  wire [7:0]    dataGroup_42_22 = dataGroup_hi_1450[319:312];
  wire [2047:0] dataGroup_lo_1451 = {dataGroup_lo_hi_1451, dataGroup_lo_lo_1451};
  wire [2047:0] dataGroup_hi_1451 = {dataGroup_hi_hi_1451, dataGroup_hi_lo_1451};
  wire [7:0]    dataGroup_43_22 = dataGroup_hi_1451[375:368];
  wire [2047:0] dataGroup_lo_1452 = {dataGroup_lo_hi_1452, dataGroup_lo_lo_1452};
  wire [2047:0] dataGroup_hi_1452 = {dataGroup_hi_hi_1452, dataGroup_hi_lo_1452};
  wire [7:0]    dataGroup_44_22 = dataGroup_hi_1452[431:424];
  wire [2047:0] dataGroup_lo_1453 = {dataGroup_lo_hi_1453, dataGroup_lo_lo_1453};
  wire [2047:0] dataGroup_hi_1453 = {dataGroup_hi_hi_1453, dataGroup_hi_lo_1453};
  wire [7:0]    dataGroup_45_22 = dataGroup_hi_1453[487:480];
  wire [2047:0] dataGroup_lo_1454 = {dataGroup_lo_hi_1454, dataGroup_lo_lo_1454};
  wire [2047:0] dataGroup_hi_1454 = {dataGroup_hi_hi_1454, dataGroup_hi_lo_1454};
  wire [7:0]    dataGroup_46_22 = dataGroup_hi_1454[543:536];
  wire [2047:0] dataGroup_lo_1455 = {dataGroup_lo_hi_1455, dataGroup_lo_lo_1455};
  wire [2047:0] dataGroup_hi_1455 = {dataGroup_hi_hi_1455, dataGroup_hi_lo_1455};
  wire [7:0]    dataGroup_47_22 = dataGroup_hi_1455[599:592];
  wire [2047:0] dataGroup_lo_1456 = {dataGroup_lo_hi_1456, dataGroup_lo_lo_1456};
  wire [2047:0] dataGroup_hi_1456 = {dataGroup_hi_hi_1456, dataGroup_hi_lo_1456};
  wire [7:0]    dataGroup_48_22 = dataGroup_hi_1456[655:648];
  wire [2047:0] dataGroup_lo_1457 = {dataGroup_lo_hi_1457, dataGroup_lo_lo_1457};
  wire [2047:0] dataGroup_hi_1457 = {dataGroup_hi_hi_1457, dataGroup_hi_lo_1457};
  wire [7:0]    dataGroup_49_22 = dataGroup_hi_1457[711:704];
  wire [2047:0] dataGroup_lo_1458 = {dataGroup_lo_hi_1458, dataGroup_lo_lo_1458};
  wire [2047:0] dataGroup_hi_1458 = {dataGroup_hi_hi_1458, dataGroup_hi_lo_1458};
  wire [7:0]    dataGroup_50_22 = dataGroup_hi_1458[767:760];
  wire [2047:0] dataGroup_lo_1459 = {dataGroup_lo_hi_1459, dataGroup_lo_lo_1459};
  wire [2047:0] dataGroup_hi_1459 = {dataGroup_hi_hi_1459, dataGroup_hi_lo_1459};
  wire [7:0]    dataGroup_51_22 = dataGroup_hi_1459[823:816];
  wire [2047:0] dataGroup_lo_1460 = {dataGroup_lo_hi_1460, dataGroup_lo_lo_1460};
  wire [2047:0] dataGroup_hi_1460 = {dataGroup_hi_hi_1460, dataGroup_hi_lo_1460};
  wire [7:0]    dataGroup_52_22 = dataGroup_hi_1460[879:872];
  wire [2047:0] dataGroup_lo_1461 = {dataGroup_lo_hi_1461, dataGroup_lo_lo_1461};
  wire [2047:0] dataGroup_hi_1461 = {dataGroup_hi_hi_1461, dataGroup_hi_lo_1461};
  wire [7:0]    dataGroup_53_22 = dataGroup_hi_1461[935:928];
  wire [2047:0] dataGroup_lo_1462 = {dataGroup_lo_hi_1462, dataGroup_lo_lo_1462};
  wire [2047:0] dataGroup_hi_1462 = {dataGroup_hi_hi_1462, dataGroup_hi_lo_1462};
  wire [7:0]    dataGroup_54_22 = dataGroup_hi_1462[991:984];
  wire [2047:0] dataGroup_lo_1463 = {dataGroup_lo_hi_1463, dataGroup_lo_lo_1463};
  wire [2047:0] dataGroup_hi_1463 = {dataGroup_hi_hi_1463, dataGroup_hi_lo_1463};
  wire [7:0]    dataGroup_55_22 = dataGroup_hi_1463[1047:1040];
  wire [2047:0] dataGroup_lo_1464 = {dataGroup_lo_hi_1464, dataGroup_lo_lo_1464};
  wire [2047:0] dataGroup_hi_1464 = {dataGroup_hi_hi_1464, dataGroup_hi_lo_1464};
  wire [7:0]    dataGroup_56_22 = dataGroup_hi_1464[1103:1096];
  wire [2047:0] dataGroup_lo_1465 = {dataGroup_lo_hi_1465, dataGroup_lo_lo_1465};
  wire [2047:0] dataGroup_hi_1465 = {dataGroup_hi_hi_1465, dataGroup_hi_lo_1465};
  wire [7:0]    dataGroup_57_22 = dataGroup_hi_1465[1159:1152];
  wire [2047:0] dataGroup_lo_1466 = {dataGroup_lo_hi_1466, dataGroup_lo_lo_1466};
  wire [2047:0] dataGroup_hi_1466 = {dataGroup_hi_hi_1466, dataGroup_hi_lo_1466};
  wire [7:0]    dataGroup_58_22 = dataGroup_hi_1466[1215:1208];
  wire [2047:0] dataGroup_lo_1467 = {dataGroup_lo_hi_1467, dataGroup_lo_lo_1467};
  wire [2047:0] dataGroup_hi_1467 = {dataGroup_hi_hi_1467, dataGroup_hi_lo_1467};
  wire [7:0]    dataGroup_59_22 = dataGroup_hi_1467[1271:1264];
  wire [2047:0] dataGroup_lo_1468 = {dataGroup_lo_hi_1468, dataGroup_lo_lo_1468};
  wire [2047:0] dataGroup_hi_1468 = {dataGroup_hi_hi_1468, dataGroup_hi_lo_1468};
  wire [7:0]    dataGroup_60_22 = dataGroup_hi_1468[1327:1320];
  wire [2047:0] dataGroup_lo_1469 = {dataGroup_lo_hi_1469, dataGroup_lo_lo_1469};
  wire [2047:0] dataGroup_hi_1469 = {dataGroup_hi_hi_1469, dataGroup_hi_lo_1469};
  wire [7:0]    dataGroup_61_22 = dataGroup_hi_1469[1383:1376];
  wire [2047:0] dataGroup_lo_1470 = {dataGroup_lo_hi_1470, dataGroup_lo_lo_1470};
  wire [2047:0] dataGroup_hi_1470 = {dataGroup_hi_hi_1470, dataGroup_hi_lo_1470};
  wire [7:0]    dataGroup_62_22 = dataGroup_hi_1470[1439:1432];
  wire [2047:0] dataGroup_lo_1471 = {dataGroup_lo_hi_1471, dataGroup_lo_lo_1471};
  wire [2047:0] dataGroup_hi_1471 = {dataGroup_hi_hi_1471, dataGroup_hi_lo_1471};
  wire [7:0]    dataGroup_63_22 = dataGroup_hi_1471[1495:1488];
  wire [15:0]   res_lo_lo_lo_lo_lo_22 = {dataGroup_1_22, dataGroup_0_22};
  wire [15:0]   res_lo_lo_lo_lo_hi_22 = {dataGroup_3_22, dataGroup_2_22};
  wire [31:0]   res_lo_lo_lo_lo_22 = {res_lo_lo_lo_lo_hi_22, res_lo_lo_lo_lo_lo_22};
  wire [15:0]   res_lo_lo_lo_hi_lo_22 = {dataGroup_5_22, dataGroup_4_22};
  wire [15:0]   res_lo_lo_lo_hi_hi_22 = {dataGroup_7_22, dataGroup_6_22};
  wire [31:0]   res_lo_lo_lo_hi_22 = {res_lo_lo_lo_hi_hi_22, res_lo_lo_lo_hi_lo_22};
  wire [63:0]   res_lo_lo_lo_22 = {res_lo_lo_lo_hi_22, res_lo_lo_lo_lo_22};
  wire [15:0]   res_lo_lo_hi_lo_lo_22 = {dataGroup_9_22, dataGroup_8_22};
  wire [15:0]   res_lo_lo_hi_lo_hi_22 = {dataGroup_11_22, dataGroup_10_22};
  wire [31:0]   res_lo_lo_hi_lo_22 = {res_lo_lo_hi_lo_hi_22, res_lo_lo_hi_lo_lo_22};
  wire [15:0]   res_lo_lo_hi_hi_lo_22 = {dataGroup_13_22, dataGroup_12_22};
  wire [15:0]   res_lo_lo_hi_hi_hi_22 = {dataGroup_15_22, dataGroup_14_22};
  wire [31:0]   res_lo_lo_hi_hi_22 = {res_lo_lo_hi_hi_hi_22, res_lo_lo_hi_hi_lo_22};
  wire [63:0]   res_lo_lo_hi_22 = {res_lo_lo_hi_hi_22, res_lo_lo_hi_lo_22};
  wire [127:0]  res_lo_lo_22 = {res_lo_lo_hi_22, res_lo_lo_lo_22};
  wire [15:0]   res_lo_hi_lo_lo_lo_22 = {dataGroup_17_22, dataGroup_16_22};
  wire [15:0]   res_lo_hi_lo_lo_hi_22 = {dataGroup_19_22, dataGroup_18_22};
  wire [31:0]   res_lo_hi_lo_lo_22 = {res_lo_hi_lo_lo_hi_22, res_lo_hi_lo_lo_lo_22};
  wire [15:0]   res_lo_hi_lo_hi_lo_22 = {dataGroup_21_22, dataGroup_20_22};
  wire [15:0]   res_lo_hi_lo_hi_hi_22 = {dataGroup_23_22, dataGroup_22_22};
  wire [31:0]   res_lo_hi_lo_hi_22 = {res_lo_hi_lo_hi_hi_22, res_lo_hi_lo_hi_lo_22};
  wire [63:0]   res_lo_hi_lo_22 = {res_lo_hi_lo_hi_22, res_lo_hi_lo_lo_22};
  wire [15:0]   res_lo_hi_hi_lo_lo_22 = {dataGroup_25_22, dataGroup_24_22};
  wire [15:0]   res_lo_hi_hi_lo_hi_22 = {dataGroup_27_22, dataGroup_26_22};
  wire [31:0]   res_lo_hi_hi_lo_22 = {res_lo_hi_hi_lo_hi_22, res_lo_hi_hi_lo_lo_22};
  wire [15:0]   res_lo_hi_hi_hi_lo_22 = {dataGroup_29_22, dataGroup_28_22};
  wire [15:0]   res_lo_hi_hi_hi_hi_22 = {dataGroup_31_22, dataGroup_30_22};
  wire [31:0]   res_lo_hi_hi_hi_22 = {res_lo_hi_hi_hi_hi_22, res_lo_hi_hi_hi_lo_22};
  wire [63:0]   res_lo_hi_hi_22 = {res_lo_hi_hi_hi_22, res_lo_hi_hi_lo_22};
  wire [127:0]  res_lo_hi_22 = {res_lo_hi_hi_22, res_lo_hi_lo_22};
  wire [255:0]  res_lo_22 = {res_lo_hi_22, res_lo_lo_22};
  wire [15:0]   res_hi_lo_lo_lo_lo_22 = {dataGroup_33_22, dataGroup_32_22};
  wire [15:0]   res_hi_lo_lo_lo_hi_22 = {dataGroup_35_22, dataGroup_34_22};
  wire [31:0]   res_hi_lo_lo_lo_22 = {res_hi_lo_lo_lo_hi_22, res_hi_lo_lo_lo_lo_22};
  wire [15:0]   res_hi_lo_lo_hi_lo_22 = {dataGroup_37_22, dataGroup_36_22};
  wire [15:0]   res_hi_lo_lo_hi_hi_22 = {dataGroup_39_22, dataGroup_38_22};
  wire [31:0]   res_hi_lo_lo_hi_22 = {res_hi_lo_lo_hi_hi_22, res_hi_lo_lo_hi_lo_22};
  wire [63:0]   res_hi_lo_lo_22 = {res_hi_lo_lo_hi_22, res_hi_lo_lo_lo_22};
  wire [15:0]   res_hi_lo_hi_lo_lo_22 = {dataGroup_41_22, dataGroup_40_22};
  wire [15:0]   res_hi_lo_hi_lo_hi_22 = {dataGroup_43_22, dataGroup_42_22};
  wire [31:0]   res_hi_lo_hi_lo_22 = {res_hi_lo_hi_lo_hi_22, res_hi_lo_hi_lo_lo_22};
  wire [15:0]   res_hi_lo_hi_hi_lo_22 = {dataGroup_45_22, dataGroup_44_22};
  wire [15:0]   res_hi_lo_hi_hi_hi_22 = {dataGroup_47_22, dataGroup_46_22};
  wire [31:0]   res_hi_lo_hi_hi_22 = {res_hi_lo_hi_hi_hi_22, res_hi_lo_hi_hi_lo_22};
  wire [63:0]   res_hi_lo_hi_22 = {res_hi_lo_hi_hi_22, res_hi_lo_hi_lo_22};
  wire [127:0]  res_hi_lo_22 = {res_hi_lo_hi_22, res_hi_lo_lo_22};
  wire [15:0]   res_hi_hi_lo_lo_lo_22 = {dataGroup_49_22, dataGroup_48_22};
  wire [15:0]   res_hi_hi_lo_lo_hi_22 = {dataGroup_51_22, dataGroup_50_22};
  wire [31:0]   res_hi_hi_lo_lo_22 = {res_hi_hi_lo_lo_hi_22, res_hi_hi_lo_lo_lo_22};
  wire [15:0]   res_hi_hi_lo_hi_lo_22 = {dataGroup_53_22, dataGroup_52_22};
  wire [15:0]   res_hi_hi_lo_hi_hi_22 = {dataGroup_55_22, dataGroup_54_22};
  wire [31:0]   res_hi_hi_lo_hi_22 = {res_hi_hi_lo_hi_hi_22, res_hi_hi_lo_hi_lo_22};
  wire [63:0]   res_hi_hi_lo_22 = {res_hi_hi_lo_hi_22, res_hi_hi_lo_lo_22};
  wire [15:0]   res_hi_hi_hi_lo_lo_22 = {dataGroup_57_22, dataGroup_56_22};
  wire [15:0]   res_hi_hi_hi_lo_hi_22 = {dataGroup_59_22, dataGroup_58_22};
  wire [31:0]   res_hi_hi_hi_lo_22 = {res_hi_hi_hi_lo_hi_22, res_hi_hi_hi_lo_lo_22};
  wire [15:0]   res_hi_hi_hi_hi_lo_22 = {dataGroup_61_22, dataGroup_60_22};
  wire [15:0]   res_hi_hi_hi_hi_hi_22 = {dataGroup_63_22, dataGroup_62_22};
  wire [31:0]   res_hi_hi_hi_hi_22 = {res_hi_hi_hi_hi_hi_22, res_hi_hi_hi_hi_lo_22};
  wire [63:0]   res_hi_hi_hi_22 = {res_hi_hi_hi_hi_22, res_hi_hi_hi_lo_22};
  wire [127:0]  res_hi_hi_22 = {res_hi_hi_hi_22, res_hi_hi_lo_22};
  wire [255:0]  res_hi_22 = {res_hi_hi_22, res_hi_lo_22};
  wire [511:0]  res_49 = {res_hi_22, res_lo_22};
  wire [2047:0] dataGroup_lo_1472 = {dataGroup_lo_hi_1472, dataGroup_lo_lo_1472};
  wire [2047:0] dataGroup_hi_1472 = {dataGroup_hi_hi_1472, dataGroup_hi_lo_1472};
  wire [7:0]    dataGroup_0_23 = dataGroup_lo_1472[23:16];
  wire [2047:0] dataGroup_lo_1473 = {dataGroup_lo_hi_1473, dataGroup_lo_lo_1473};
  wire [2047:0] dataGroup_hi_1473 = {dataGroup_hi_hi_1473, dataGroup_hi_lo_1473};
  wire [7:0]    dataGroup_1_23 = dataGroup_lo_1473[79:72];
  wire [2047:0] dataGroup_lo_1474 = {dataGroup_lo_hi_1474, dataGroup_lo_lo_1474};
  wire [2047:0] dataGroup_hi_1474 = {dataGroup_hi_hi_1474, dataGroup_hi_lo_1474};
  wire [7:0]    dataGroup_2_23 = dataGroup_lo_1474[135:128];
  wire [2047:0] dataGroup_lo_1475 = {dataGroup_lo_hi_1475, dataGroup_lo_lo_1475};
  wire [2047:0] dataGroup_hi_1475 = {dataGroup_hi_hi_1475, dataGroup_hi_lo_1475};
  wire [7:0]    dataGroup_3_23 = dataGroup_lo_1475[191:184];
  wire [2047:0] dataGroup_lo_1476 = {dataGroup_lo_hi_1476, dataGroup_lo_lo_1476};
  wire [2047:0] dataGroup_hi_1476 = {dataGroup_hi_hi_1476, dataGroup_hi_lo_1476};
  wire [7:0]    dataGroup_4_23 = dataGroup_lo_1476[247:240];
  wire [2047:0] dataGroup_lo_1477 = {dataGroup_lo_hi_1477, dataGroup_lo_lo_1477};
  wire [2047:0] dataGroup_hi_1477 = {dataGroup_hi_hi_1477, dataGroup_hi_lo_1477};
  wire [7:0]    dataGroup_5_23 = dataGroup_lo_1477[303:296];
  wire [2047:0] dataGroup_lo_1478 = {dataGroup_lo_hi_1478, dataGroup_lo_lo_1478};
  wire [2047:0] dataGroup_hi_1478 = {dataGroup_hi_hi_1478, dataGroup_hi_lo_1478};
  wire [7:0]    dataGroup_6_23 = dataGroup_lo_1478[359:352];
  wire [2047:0] dataGroup_lo_1479 = {dataGroup_lo_hi_1479, dataGroup_lo_lo_1479};
  wire [2047:0] dataGroup_hi_1479 = {dataGroup_hi_hi_1479, dataGroup_hi_lo_1479};
  wire [7:0]    dataGroup_7_23 = dataGroup_lo_1479[415:408];
  wire [2047:0] dataGroup_lo_1480 = {dataGroup_lo_hi_1480, dataGroup_lo_lo_1480};
  wire [2047:0] dataGroup_hi_1480 = {dataGroup_hi_hi_1480, dataGroup_hi_lo_1480};
  wire [7:0]    dataGroup_8_23 = dataGroup_lo_1480[471:464];
  wire [2047:0] dataGroup_lo_1481 = {dataGroup_lo_hi_1481, dataGroup_lo_lo_1481};
  wire [2047:0] dataGroup_hi_1481 = {dataGroup_hi_hi_1481, dataGroup_hi_lo_1481};
  wire [7:0]    dataGroup_9_23 = dataGroup_lo_1481[527:520];
  wire [2047:0] dataGroup_lo_1482 = {dataGroup_lo_hi_1482, dataGroup_lo_lo_1482};
  wire [2047:0] dataGroup_hi_1482 = {dataGroup_hi_hi_1482, dataGroup_hi_lo_1482};
  wire [7:0]    dataGroup_10_23 = dataGroup_lo_1482[583:576];
  wire [2047:0] dataGroup_lo_1483 = {dataGroup_lo_hi_1483, dataGroup_lo_lo_1483};
  wire [2047:0] dataGroup_hi_1483 = {dataGroup_hi_hi_1483, dataGroup_hi_lo_1483};
  wire [7:0]    dataGroup_11_23 = dataGroup_lo_1483[639:632];
  wire [2047:0] dataGroup_lo_1484 = {dataGroup_lo_hi_1484, dataGroup_lo_lo_1484};
  wire [2047:0] dataGroup_hi_1484 = {dataGroup_hi_hi_1484, dataGroup_hi_lo_1484};
  wire [7:0]    dataGroup_12_23 = dataGroup_lo_1484[695:688];
  wire [2047:0] dataGroup_lo_1485 = {dataGroup_lo_hi_1485, dataGroup_lo_lo_1485};
  wire [2047:0] dataGroup_hi_1485 = {dataGroup_hi_hi_1485, dataGroup_hi_lo_1485};
  wire [7:0]    dataGroup_13_23 = dataGroup_lo_1485[751:744];
  wire [2047:0] dataGroup_lo_1486 = {dataGroup_lo_hi_1486, dataGroup_lo_lo_1486};
  wire [2047:0] dataGroup_hi_1486 = {dataGroup_hi_hi_1486, dataGroup_hi_lo_1486};
  wire [7:0]    dataGroup_14_23 = dataGroup_lo_1486[807:800];
  wire [2047:0] dataGroup_lo_1487 = {dataGroup_lo_hi_1487, dataGroup_lo_lo_1487};
  wire [2047:0] dataGroup_hi_1487 = {dataGroup_hi_hi_1487, dataGroup_hi_lo_1487};
  wire [7:0]    dataGroup_15_23 = dataGroup_lo_1487[863:856];
  wire [2047:0] dataGroup_lo_1488 = {dataGroup_lo_hi_1488, dataGroup_lo_lo_1488};
  wire [2047:0] dataGroup_hi_1488 = {dataGroup_hi_hi_1488, dataGroup_hi_lo_1488};
  wire [7:0]    dataGroup_16_23 = dataGroup_lo_1488[919:912];
  wire [2047:0] dataGroup_lo_1489 = {dataGroup_lo_hi_1489, dataGroup_lo_lo_1489};
  wire [2047:0] dataGroup_hi_1489 = {dataGroup_hi_hi_1489, dataGroup_hi_lo_1489};
  wire [7:0]    dataGroup_17_23 = dataGroup_lo_1489[975:968];
  wire [2047:0] dataGroup_lo_1490 = {dataGroup_lo_hi_1490, dataGroup_lo_lo_1490};
  wire [2047:0] dataGroup_hi_1490 = {dataGroup_hi_hi_1490, dataGroup_hi_lo_1490};
  wire [7:0]    dataGroup_18_23 = dataGroup_lo_1490[1031:1024];
  wire [2047:0] dataGroup_lo_1491 = {dataGroup_lo_hi_1491, dataGroup_lo_lo_1491};
  wire [2047:0] dataGroup_hi_1491 = {dataGroup_hi_hi_1491, dataGroup_hi_lo_1491};
  wire [7:0]    dataGroup_19_23 = dataGroup_lo_1491[1087:1080];
  wire [2047:0] dataGroup_lo_1492 = {dataGroup_lo_hi_1492, dataGroup_lo_lo_1492};
  wire [2047:0] dataGroup_hi_1492 = {dataGroup_hi_hi_1492, dataGroup_hi_lo_1492};
  wire [7:0]    dataGroup_20_23 = dataGroup_lo_1492[1143:1136];
  wire [2047:0] dataGroup_lo_1493 = {dataGroup_lo_hi_1493, dataGroup_lo_lo_1493};
  wire [2047:0] dataGroup_hi_1493 = {dataGroup_hi_hi_1493, dataGroup_hi_lo_1493};
  wire [7:0]    dataGroup_21_23 = dataGroup_lo_1493[1199:1192];
  wire [2047:0] dataGroup_lo_1494 = {dataGroup_lo_hi_1494, dataGroup_lo_lo_1494};
  wire [2047:0] dataGroup_hi_1494 = {dataGroup_hi_hi_1494, dataGroup_hi_lo_1494};
  wire [7:0]    dataGroup_22_23 = dataGroup_lo_1494[1255:1248];
  wire [2047:0] dataGroup_lo_1495 = {dataGroup_lo_hi_1495, dataGroup_lo_lo_1495};
  wire [2047:0] dataGroup_hi_1495 = {dataGroup_hi_hi_1495, dataGroup_hi_lo_1495};
  wire [7:0]    dataGroup_23_23 = dataGroup_lo_1495[1311:1304];
  wire [2047:0] dataGroup_lo_1496 = {dataGroup_lo_hi_1496, dataGroup_lo_lo_1496};
  wire [2047:0] dataGroup_hi_1496 = {dataGroup_hi_hi_1496, dataGroup_hi_lo_1496};
  wire [7:0]    dataGroup_24_23 = dataGroup_lo_1496[1367:1360];
  wire [2047:0] dataGroup_lo_1497 = {dataGroup_lo_hi_1497, dataGroup_lo_lo_1497};
  wire [2047:0] dataGroup_hi_1497 = {dataGroup_hi_hi_1497, dataGroup_hi_lo_1497};
  wire [7:0]    dataGroup_25_23 = dataGroup_lo_1497[1423:1416];
  wire [2047:0] dataGroup_lo_1498 = {dataGroup_lo_hi_1498, dataGroup_lo_lo_1498};
  wire [2047:0] dataGroup_hi_1498 = {dataGroup_hi_hi_1498, dataGroup_hi_lo_1498};
  wire [7:0]    dataGroup_26_23 = dataGroup_lo_1498[1479:1472];
  wire [2047:0] dataGroup_lo_1499 = {dataGroup_lo_hi_1499, dataGroup_lo_lo_1499};
  wire [2047:0] dataGroup_hi_1499 = {dataGroup_hi_hi_1499, dataGroup_hi_lo_1499};
  wire [7:0]    dataGroup_27_23 = dataGroup_lo_1499[1535:1528];
  wire [2047:0] dataGroup_lo_1500 = {dataGroup_lo_hi_1500, dataGroup_lo_lo_1500};
  wire [2047:0] dataGroup_hi_1500 = {dataGroup_hi_hi_1500, dataGroup_hi_lo_1500};
  wire [7:0]    dataGroup_28_23 = dataGroup_lo_1500[1591:1584];
  wire [2047:0] dataGroup_lo_1501 = {dataGroup_lo_hi_1501, dataGroup_lo_lo_1501};
  wire [2047:0] dataGroup_hi_1501 = {dataGroup_hi_hi_1501, dataGroup_hi_lo_1501};
  wire [7:0]    dataGroup_29_23 = dataGroup_lo_1501[1647:1640];
  wire [2047:0] dataGroup_lo_1502 = {dataGroup_lo_hi_1502, dataGroup_lo_lo_1502};
  wire [2047:0] dataGroup_hi_1502 = {dataGroup_hi_hi_1502, dataGroup_hi_lo_1502};
  wire [7:0]    dataGroup_30_23 = dataGroup_lo_1502[1703:1696];
  wire [2047:0] dataGroup_lo_1503 = {dataGroup_lo_hi_1503, dataGroup_lo_lo_1503};
  wire [2047:0] dataGroup_hi_1503 = {dataGroup_hi_hi_1503, dataGroup_hi_lo_1503};
  wire [7:0]    dataGroup_31_23 = dataGroup_lo_1503[1759:1752];
  wire [2047:0] dataGroup_lo_1504 = {dataGroup_lo_hi_1504, dataGroup_lo_lo_1504};
  wire [2047:0] dataGroup_hi_1504 = {dataGroup_hi_hi_1504, dataGroup_hi_lo_1504};
  wire [7:0]    dataGroup_32_23 = dataGroup_lo_1504[1815:1808];
  wire [2047:0] dataGroup_lo_1505 = {dataGroup_lo_hi_1505, dataGroup_lo_lo_1505};
  wire [2047:0] dataGroup_hi_1505 = {dataGroup_hi_hi_1505, dataGroup_hi_lo_1505};
  wire [7:0]    dataGroup_33_23 = dataGroup_lo_1505[1871:1864];
  wire [2047:0] dataGroup_lo_1506 = {dataGroup_lo_hi_1506, dataGroup_lo_lo_1506};
  wire [2047:0] dataGroup_hi_1506 = {dataGroup_hi_hi_1506, dataGroup_hi_lo_1506};
  wire [7:0]    dataGroup_34_23 = dataGroup_lo_1506[1927:1920];
  wire [2047:0] dataGroup_lo_1507 = {dataGroup_lo_hi_1507, dataGroup_lo_lo_1507};
  wire [2047:0] dataGroup_hi_1507 = {dataGroup_hi_hi_1507, dataGroup_hi_lo_1507};
  wire [7:0]    dataGroup_35_23 = dataGroup_lo_1507[1983:1976];
  wire [2047:0] dataGroup_lo_1508 = {dataGroup_lo_hi_1508, dataGroup_lo_lo_1508};
  wire [2047:0] dataGroup_hi_1508 = {dataGroup_hi_hi_1508, dataGroup_hi_lo_1508};
  wire [7:0]    dataGroup_36_23 = dataGroup_lo_1508[2039:2032];
  wire [2047:0] dataGroup_lo_1509 = {dataGroup_lo_hi_1509, dataGroup_lo_lo_1509};
  wire [2047:0] dataGroup_hi_1509 = {dataGroup_hi_hi_1509, dataGroup_hi_lo_1509};
  wire [7:0]    dataGroup_37_23 = dataGroup_hi_1509[47:40];
  wire [2047:0] dataGroup_lo_1510 = {dataGroup_lo_hi_1510, dataGroup_lo_lo_1510};
  wire [2047:0] dataGroup_hi_1510 = {dataGroup_hi_hi_1510, dataGroup_hi_lo_1510};
  wire [7:0]    dataGroup_38_23 = dataGroup_hi_1510[103:96];
  wire [2047:0] dataGroup_lo_1511 = {dataGroup_lo_hi_1511, dataGroup_lo_lo_1511};
  wire [2047:0] dataGroup_hi_1511 = {dataGroup_hi_hi_1511, dataGroup_hi_lo_1511};
  wire [7:0]    dataGroup_39_23 = dataGroup_hi_1511[159:152];
  wire [2047:0] dataGroup_lo_1512 = {dataGroup_lo_hi_1512, dataGroup_lo_lo_1512};
  wire [2047:0] dataGroup_hi_1512 = {dataGroup_hi_hi_1512, dataGroup_hi_lo_1512};
  wire [7:0]    dataGroup_40_23 = dataGroup_hi_1512[215:208];
  wire [2047:0] dataGroup_lo_1513 = {dataGroup_lo_hi_1513, dataGroup_lo_lo_1513};
  wire [2047:0] dataGroup_hi_1513 = {dataGroup_hi_hi_1513, dataGroup_hi_lo_1513};
  wire [7:0]    dataGroup_41_23 = dataGroup_hi_1513[271:264];
  wire [2047:0] dataGroup_lo_1514 = {dataGroup_lo_hi_1514, dataGroup_lo_lo_1514};
  wire [2047:0] dataGroup_hi_1514 = {dataGroup_hi_hi_1514, dataGroup_hi_lo_1514};
  wire [7:0]    dataGroup_42_23 = dataGroup_hi_1514[327:320];
  wire [2047:0] dataGroup_lo_1515 = {dataGroup_lo_hi_1515, dataGroup_lo_lo_1515};
  wire [2047:0] dataGroup_hi_1515 = {dataGroup_hi_hi_1515, dataGroup_hi_lo_1515};
  wire [7:0]    dataGroup_43_23 = dataGroup_hi_1515[383:376];
  wire [2047:0] dataGroup_lo_1516 = {dataGroup_lo_hi_1516, dataGroup_lo_lo_1516};
  wire [2047:0] dataGroup_hi_1516 = {dataGroup_hi_hi_1516, dataGroup_hi_lo_1516};
  wire [7:0]    dataGroup_44_23 = dataGroup_hi_1516[439:432];
  wire [2047:0] dataGroup_lo_1517 = {dataGroup_lo_hi_1517, dataGroup_lo_lo_1517};
  wire [2047:0] dataGroup_hi_1517 = {dataGroup_hi_hi_1517, dataGroup_hi_lo_1517};
  wire [7:0]    dataGroup_45_23 = dataGroup_hi_1517[495:488];
  wire [2047:0] dataGroup_lo_1518 = {dataGroup_lo_hi_1518, dataGroup_lo_lo_1518};
  wire [2047:0] dataGroup_hi_1518 = {dataGroup_hi_hi_1518, dataGroup_hi_lo_1518};
  wire [7:0]    dataGroup_46_23 = dataGroup_hi_1518[551:544];
  wire [2047:0] dataGroup_lo_1519 = {dataGroup_lo_hi_1519, dataGroup_lo_lo_1519};
  wire [2047:0] dataGroup_hi_1519 = {dataGroup_hi_hi_1519, dataGroup_hi_lo_1519};
  wire [7:0]    dataGroup_47_23 = dataGroup_hi_1519[607:600];
  wire [2047:0] dataGroup_lo_1520 = {dataGroup_lo_hi_1520, dataGroup_lo_lo_1520};
  wire [2047:0] dataGroup_hi_1520 = {dataGroup_hi_hi_1520, dataGroup_hi_lo_1520};
  wire [7:0]    dataGroup_48_23 = dataGroup_hi_1520[663:656];
  wire [2047:0] dataGroup_lo_1521 = {dataGroup_lo_hi_1521, dataGroup_lo_lo_1521};
  wire [2047:0] dataGroup_hi_1521 = {dataGroup_hi_hi_1521, dataGroup_hi_lo_1521};
  wire [7:0]    dataGroup_49_23 = dataGroup_hi_1521[719:712];
  wire [2047:0] dataGroup_lo_1522 = {dataGroup_lo_hi_1522, dataGroup_lo_lo_1522};
  wire [2047:0] dataGroup_hi_1522 = {dataGroup_hi_hi_1522, dataGroup_hi_lo_1522};
  wire [7:0]    dataGroup_50_23 = dataGroup_hi_1522[775:768];
  wire [2047:0] dataGroup_lo_1523 = {dataGroup_lo_hi_1523, dataGroup_lo_lo_1523};
  wire [2047:0] dataGroup_hi_1523 = {dataGroup_hi_hi_1523, dataGroup_hi_lo_1523};
  wire [7:0]    dataGroup_51_23 = dataGroup_hi_1523[831:824];
  wire [2047:0] dataGroup_lo_1524 = {dataGroup_lo_hi_1524, dataGroup_lo_lo_1524};
  wire [2047:0] dataGroup_hi_1524 = {dataGroup_hi_hi_1524, dataGroup_hi_lo_1524};
  wire [7:0]    dataGroup_52_23 = dataGroup_hi_1524[887:880];
  wire [2047:0] dataGroup_lo_1525 = {dataGroup_lo_hi_1525, dataGroup_lo_lo_1525};
  wire [2047:0] dataGroup_hi_1525 = {dataGroup_hi_hi_1525, dataGroup_hi_lo_1525};
  wire [7:0]    dataGroup_53_23 = dataGroup_hi_1525[943:936];
  wire [2047:0] dataGroup_lo_1526 = {dataGroup_lo_hi_1526, dataGroup_lo_lo_1526};
  wire [2047:0] dataGroup_hi_1526 = {dataGroup_hi_hi_1526, dataGroup_hi_lo_1526};
  wire [7:0]    dataGroup_54_23 = dataGroup_hi_1526[999:992];
  wire [2047:0] dataGroup_lo_1527 = {dataGroup_lo_hi_1527, dataGroup_lo_lo_1527};
  wire [2047:0] dataGroup_hi_1527 = {dataGroup_hi_hi_1527, dataGroup_hi_lo_1527};
  wire [7:0]    dataGroup_55_23 = dataGroup_hi_1527[1055:1048];
  wire [2047:0] dataGroup_lo_1528 = {dataGroup_lo_hi_1528, dataGroup_lo_lo_1528};
  wire [2047:0] dataGroup_hi_1528 = {dataGroup_hi_hi_1528, dataGroup_hi_lo_1528};
  wire [7:0]    dataGroup_56_23 = dataGroup_hi_1528[1111:1104];
  wire [2047:0] dataGroup_lo_1529 = {dataGroup_lo_hi_1529, dataGroup_lo_lo_1529};
  wire [2047:0] dataGroup_hi_1529 = {dataGroup_hi_hi_1529, dataGroup_hi_lo_1529};
  wire [7:0]    dataGroup_57_23 = dataGroup_hi_1529[1167:1160];
  wire [2047:0] dataGroup_lo_1530 = {dataGroup_lo_hi_1530, dataGroup_lo_lo_1530};
  wire [2047:0] dataGroup_hi_1530 = {dataGroup_hi_hi_1530, dataGroup_hi_lo_1530};
  wire [7:0]    dataGroup_58_23 = dataGroup_hi_1530[1223:1216];
  wire [2047:0] dataGroup_lo_1531 = {dataGroup_lo_hi_1531, dataGroup_lo_lo_1531};
  wire [2047:0] dataGroup_hi_1531 = {dataGroup_hi_hi_1531, dataGroup_hi_lo_1531};
  wire [7:0]    dataGroup_59_23 = dataGroup_hi_1531[1279:1272];
  wire [2047:0] dataGroup_lo_1532 = {dataGroup_lo_hi_1532, dataGroup_lo_lo_1532};
  wire [2047:0] dataGroup_hi_1532 = {dataGroup_hi_hi_1532, dataGroup_hi_lo_1532};
  wire [7:0]    dataGroup_60_23 = dataGroup_hi_1532[1335:1328];
  wire [2047:0] dataGroup_lo_1533 = {dataGroup_lo_hi_1533, dataGroup_lo_lo_1533};
  wire [2047:0] dataGroup_hi_1533 = {dataGroup_hi_hi_1533, dataGroup_hi_lo_1533};
  wire [7:0]    dataGroup_61_23 = dataGroup_hi_1533[1391:1384];
  wire [2047:0] dataGroup_lo_1534 = {dataGroup_lo_hi_1534, dataGroup_lo_lo_1534};
  wire [2047:0] dataGroup_hi_1534 = {dataGroup_hi_hi_1534, dataGroup_hi_lo_1534};
  wire [7:0]    dataGroup_62_23 = dataGroup_hi_1534[1447:1440];
  wire [2047:0] dataGroup_lo_1535 = {dataGroup_lo_hi_1535, dataGroup_lo_lo_1535};
  wire [2047:0] dataGroup_hi_1535 = {dataGroup_hi_hi_1535, dataGroup_hi_lo_1535};
  wire [7:0]    dataGroup_63_23 = dataGroup_hi_1535[1503:1496];
  wire [15:0]   res_lo_lo_lo_lo_lo_23 = {dataGroup_1_23, dataGroup_0_23};
  wire [15:0]   res_lo_lo_lo_lo_hi_23 = {dataGroup_3_23, dataGroup_2_23};
  wire [31:0]   res_lo_lo_lo_lo_23 = {res_lo_lo_lo_lo_hi_23, res_lo_lo_lo_lo_lo_23};
  wire [15:0]   res_lo_lo_lo_hi_lo_23 = {dataGroup_5_23, dataGroup_4_23};
  wire [15:0]   res_lo_lo_lo_hi_hi_23 = {dataGroup_7_23, dataGroup_6_23};
  wire [31:0]   res_lo_lo_lo_hi_23 = {res_lo_lo_lo_hi_hi_23, res_lo_lo_lo_hi_lo_23};
  wire [63:0]   res_lo_lo_lo_23 = {res_lo_lo_lo_hi_23, res_lo_lo_lo_lo_23};
  wire [15:0]   res_lo_lo_hi_lo_lo_23 = {dataGroup_9_23, dataGroup_8_23};
  wire [15:0]   res_lo_lo_hi_lo_hi_23 = {dataGroup_11_23, dataGroup_10_23};
  wire [31:0]   res_lo_lo_hi_lo_23 = {res_lo_lo_hi_lo_hi_23, res_lo_lo_hi_lo_lo_23};
  wire [15:0]   res_lo_lo_hi_hi_lo_23 = {dataGroup_13_23, dataGroup_12_23};
  wire [15:0]   res_lo_lo_hi_hi_hi_23 = {dataGroup_15_23, dataGroup_14_23};
  wire [31:0]   res_lo_lo_hi_hi_23 = {res_lo_lo_hi_hi_hi_23, res_lo_lo_hi_hi_lo_23};
  wire [63:0]   res_lo_lo_hi_23 = {res_lo_lo_hi_hi_23, res_lo_lo_hi_lo_23};
  wire [127:0]  res_lo_lo_23 = {res_lo_lo_hi_23, res_lo_lo_lo_23};
  wire [15:0]   res_lo_hi_lo_lo_lo_23 = {dataGroup_17_23, dataGroup_16_23};
  wire [15:0]   res_lo_hi_lo_lo_hi_23 = {dataGroup_19_23, dataGroup_18_23};
  wire [31:0]   res_lo_hi_lo_lo_23 = {res_lo_hi_lo_lo_hi_23, res_lo_hi_lo_lo_lo_23};
  wire [15:0]   res_lo_hi_lo_hi_lo_23 = {dataGroup_21_23, dataGroup_20_23};
  wire [15:0]   res_lo_hi_lo_hi_hi_23 = {dataGroup_23_23, dataGroup_22_23};
  wire [31:0]   res_lo_hi_lo_hi_23 = {res_lo_hi_lo_hi_hi_23, res_lo_hi_lo_hi_lo_23};
  wire [63:0]   res_lo_hi_lo_23 = {res_lo_hi_lo_hi_23, res_lo_hi_lo_lo_23};
  wire [15:0]   res_lo_hi_hi_lo_lo_23 = {dataGroup_25_23, dataGroup_24_23};
  wire [15:0]   res_lo_hi_hi_lo_hi_23 = {dataGroup_27_23, dataGroup_26_23};
  wire [31:0]   res_lo_hi_hi_lo_23 = {res_lo_hi_hi_lo_hi_23, res_lo_hi_hi_lo_lo_23};
  wire [15:0]   res_lo_hi_hi_hi_lo_23 = {dataGroup_29_23, dataGroup_28_23};
  wire [15:0]   res_lo_hi_hi_hi_hi_23 = {dataGroup_31_23, dataGroup_30_23};
  wire [31:0]   res_lo_hi_hi_hi_23 = {res_lo_hi_hi_hi_hi_23, res_lo_hi_hi_hi_lo_23};
  wire [63:0]   res_lo_hi_hi_23 = {res_lo_hi_hi_hi_23, res_lo_hi_hi_lo_23};
  wire [127:0]  res_lo_hi_23 = {res_lo_hi_hi_23, res_lo_hi_lo_23};
  wire [255:0]  res_lo_23 = {res_lo_hi_23, res_lo_lo_23};
  wire [15:0]   res_hi_lo_lo_lo_lo_23 = {dataGroup_33_23, dataGroup_32_23};
  wire [15:0]   res_hi_lo_lo_lo_hi_23 = {dataGroup_35_23, dataGroup_34_23};
  wire [31:0]   res_hi_lo_lo_lo_23 = {res_hi_lo_lo_lo_hi_23, res_hi_lo_lo_lo_lo_23};
  wire [15:0]   res_hi_lo_lo_hi_lo_23 = {dataGroup_37_23, dataGroup_36_23};
  wire [15:0]   res_hi_lo_lo_hi_hi_23 = {dataGroup_39_23, dataGroup_38_23};
  wire [31:0]   res_hi_lo_lo_hi_23 = {res_hi_lo_lo_hi_hi_23, res_hi_lo_lo_hi_lo_23};
  wire [63:0]   res_hi_lo_lo_23 = {res_hi_lo_lo_hi_23, res_hi_lo_lo_lo_23};
  wire [15:0]   res_hi_lo_hi_lo_lo_23 = {dataGroup_41_23, dataGroup_40_23};
  wire [15:0]   res_hi_lo_hi_lo_hi_23 = {dataGroup_43_23, dataGroup_42_23};
  wire [31:0]   res_hi_lo_hi_lo_23 = {res_hi_lo_hi_lo_hi_23, res_hi_lo_hi_lo_lo_23};
  wire [15:0]   res_hi_lo_hi_hi_lo_23 = {dataGroup_45_23, dataGroup_44_23};
  wire [15:0]   res_hi_lo_hi_hi_hi_23 = {dataGroup_47_23, dataGroup_46_23};
  wire [31:0]   res_hi_lo_hi_hi_23 = {res_hi_lo_hi_hi_hi_23, res_hi_lo_hi_hi_lo_23};
  wire [63:0]   res_hi_lo_hi_23 = {res_hi_lo_hi_hi_23, res_hi_lo_hi_lo_23};
  wire [127:0]  res_hi_lo_23 = {res_hi_lo_hi_23, res_hi_lo_lo_23};
  wire [15:0]   res_hi_hi_lo_lo_lo_23 = {dataGroup_49_23, dataGroup_48_23};
  wire [15:0]   res_hi_hi_lo_lo_hi_23 = {dataGroup_51_23, dataGroup_50_23};
  wire [31:0]   res_hi_hi_lo_lo_23 = {res_hi_hi_lo_lo_hi_23, res_hi_hi_lo_lo_lo_23};
  wire [15:0]   res_hi_hi_lo_hi_lo_23 = {dataGroup_53_23, dataGroup_52_23};
  wire [15:0]   res_hi_hi_lo_hi_hi_23 = {dataGroup_55_23, dataGroup_54_23};
  wire [31:0]   res_hi_hi_lo_hi_23 = {res_hi_hi_lo_hi_hi_23, res_hi_hi_lo_hi_lo_23};
  wire [63:0]   res_hi_hi_lo_23 = {res_hi_hi_lo_hi_23, res_hi_hi_lo_lo_23};
  wire [15:0]   res_hi_hi_hi_lo_lo_23 = {dataGroup_57_23, dataGroup_56_23};
  wire [15:0]   res_hi_hi_hi_lo_hi_23 = {dataGroup_59_23, dataGroup_58_23};
  wire [31:0]   res_hi_hi_hi_lo_23 = {res_hi_hi_hi_lo_hi_23, res_hi_hi_hi_lo_lo_23};
  wire [15:0]   res_hi_hi_hi_hi_lo_23 = {dataGroup_61_23, dataGroup_60_23};
  wire [15:0]   res_hi_hi_hi_hi_hi_23 = {dataGroup_63_23, dataGroup_62_23};
  wire [31:0]   res_hi_hi_hi_hi_23 = {res_hi_hi_hi_hi_hi_23, res_hi_hi_hi_hi_lo_23};
  wire [63:0]   res_hi_hi_hi_23 = {res_hi_hi_hi_hi_23, res_hi_hi_hi_lo_23};
  wire [127:0]  res_hi_hi_23 = {res_hi_hi_hi_23, res_hi_hi_lo_23};
  wire [255:0]  res_hi_23 = {res_hi_hi_23, res_hi_lo_23};
  wire [511:0]  res_50 = {res_hi_23, res_lo_23};
  wire [2047:0] dataGroup_lo_1536 = {dataGroup_lo_hi_1536, dataGroup_lo_lo_1536};
  wire [2047:0] dataGroup_hi_1536 = {dataGroup_hi_hi_1536, dataGroup_hi_lo_1536};
  wire [7:0]    dataGroup_0_24 = dataGroup_lo_1536[31:24];
  wire [2047:0] dataGroup_lo_1537 = {dataGroup_lo_hi_1537, dataGroup_lo_lo_1537};
  wire [2047:0] dataGroup_hi_1537 = {dataGroup_hi_hi_1537, dataGroup_hi_lo_1537};
  wire [7:0]    dataGroup_1_24 = dataGroup_lo_1537[87:80];
  wire [2047:0] dataGroup_lo_1538 = {dataGroup_lo_hi_1538, dataGroup_lo_lo_1538};
  wire [2047:0] dataGroup_hi_1538 = {dataGroup_hi_hi_1538, dataGroup_hi_lo_1538};
  wire [7:0]    dataGroup_2_24 = dataGroup_lo_1538[143:136];
  wire [2047:0] dataGroup_lo_1539 = {dataGroup_lo_hi_1539, dataGroup_lo_lo_1539};
  wire [2047:0] dataGroup_hi_1539 = {dataGroup_hi_hi_1539, dataGroup_hi_lo_1539};
  wire [7:0]    dataGroup_3_24 = dataGroup_lo_1539[199:192];
  wire [2047:0] dataGroup_lo_1540 = {dataGroup_lo_hi_1540, dataGroup_lo_lo_1540};
  wire [2047:0] dataGroup_hi_1540 = {dataGroup_hi_hi_1540, dataGroup_hi_lo_1540};
  wire [7:0]    dataGroup_4_24 = dataGroup_lo_1540[255:248];
  wire [2047:0] dataGroup_lo_1541 = {dataGroup_lo_hi_1541, dataGroup_lo_lo_1541};
  wire [2047:0] dataGroup_hi_1541 = {dataGroup_hi_hi_1541, dataGroup_hi_lo_1541};
  wire [7:0]    dataGroup_5_24 = dataGroup_lo_1541[311:304];
  wire [2047:0] dataGroup_lo_1542 = {dataGroup_lo_hi_1542, dataGroup_lo_lo_1542};
  wire [2047:0] dataGroup_hi_1542 = {dataGroup_hi_hi_1542, dataGroup_hi_lo_1542};
  wire [7:0]    dataGroup_6_24 = dataGroup_lo_1542[367:360];
  wire [2047:0] dataGroup_lo_1543 = {dataGroup_lo_hi_1543, dataGroup_lo_lo_1543};
  wire [2047:0] dataGroup_hi_1543 = {dataGroup_hi_hi_1543, dataGroup_hi_lo_1543};
  wire [7:0]    dataGroup_7_24 = dataGroup_lo_1543[423:416];
  wire [2047:0] dataGroup_lo_1544 = {dataGroup_lo_hi_1544, dataGroup_lo_lo_1544};
  wire [2047:0] dataGroup_hi_1544 = {dataGroup_hi_hi_1544, dataGroup_hi_lo_1544};
  wire [7:0]    dataGroup_8_24 = dataGroup_lo_1544[479:472];
  wire [2047:0] dataGroup_lo_1545 = {dataGroup_lo_hi_1545, dataGroup_lo_lo_1545};
  wire [2047:0] dataGroup_hi_1545 = {dataGroup_hi_hi_1545, dataGroup_hi_lo_1545};
  wire [7:0]    dataGroup_9_24 = dataGroup_lo_1545[535:528];
  wire [2047:0] dataGroup_lo_1546 = {dataGroup_lo_hi_1546, dataGroup_lo_lo_1546};
  wire [2047:0] dataGroup_hi_1546 = {dataGroup_hi_hi_1546, dataGroup_hi_lo_1546};
  wire [7:0]    dataGroup_10_24 = dataGroup_lo_1546[591:584];
  wire [2047:0] dataGroup_lo_1547 = {dataGroup_lo_hi_1547, dataGroup_lo_lo_1547};
  wire [2047:0] dataGroup_hi_1547 = {dataGroup_hi_hi_1547, dataGroup_hi_lo_1547};
  wire [7:0]    dataGroup_11_24 = dataGroup_lo_1547[647:640];
  wire [2047:0] dataGroup_lo_1548 = {dataGroup_lo_hi_1548, dataGroup_lo_lo_1548};
  wire [2047:0] dataGroup_hi_1548 = {dataGroup_hi_hi_1548, dataGroup_hi_lo_1548};
  wire [7:0]    dataGroup_12_24 = dataGroup_lo_1548[703:696];
  wire [2047:0] dataGroup_lo_1549 = {dataGroup_lo_hi_1549, dataGroup_lo_lo_1549};
  wire [2047:0] dataGroup_hi_1549 = {dataGroup_hi_hi_1549, dataGroup_hi_lo_1549};
  wire [7:0]    dataGroup_13_24 = dataGroup_lo_1549[759:752];
  wire [2047:0] dataGroup_lo_1550 = {dataGroup_lo_hi_1550, dataGroup_lo_lo_1550};
  wire [2047:0] dataGroup_hi_1550 = {dataGroup_hi_hi_1550, dataGroup_hi_lo_1550};
  wire [7:0]    dataGroup_14_24 = dataGroup_lo_1550[815:808];
  wire [2047:0] dataGroup_lo_1551 = {dataGroup_lo_hi_1551, dataGroup_lo_lo_1551};
  wire [2047:0] dataGroup_hi_1551 = {dataGroup_hi_hi_1551, dataGroup_hi_lo_1551};
  wire [7:0]    dataGroup_15_24 = dataGroup_lo_1551[871:864];
  wire [2047:0] dataGroup_lo_1552 = {dataGroup_lo_hi_1552, dataGroup_lo_lo_1552};
  wire [2047:0] dataGroup_hi_1552 = {dataGroup_hi_hi_1552, dataGroup_hi_lo_1552};
  wire [7:0]    dataGroup_16_24 = dataGroup_lo_1552[927:920];
  wire [2047:0] dataGroup_lo_1553 = {dataGroup_lo_hi_1553, dataGroup_lo_lo_1553};
  wire [2047:0] dataGroup_hi_1553 = {dataGroup_hi_hi_1553, dataGroup_hi_lo_1553};
  wire [7:0]    dataGroup_17_24 = dataGroup_lo_1553[983:976];
  wire [2047:0] dataGroup_lo_1554 = {dataGroup_lo_hi_1554, dataGroup_lo_lo_1554};
  wire [2047:0] dataGroup_hi_1554 = {dataGroup_hi_hi_1554, dataGroup_hi_lo_1554};
  wire [7:0]    dataGroup_18_24 = dataGroup_lo_1554[1039:1032];
  wire [2047:0] dataGroup_lo_1555 = {dataGroup_lo_hi_1555, dataGroup_lo_lo_1555};
  wire [2047:0] dataGroup_hi_1555 = {dataGroup_hi_hi_1555, dataGroup_hi_lo_1555};
  wire [7:0]    dataGroup_19_24 = dataGroup_lo_1555[1095:1088];
  wire [2047:0] dataGroup_lo_1556 = {dataGroup_lo_hi_1556, dataGroup_lo_lo_1556};
  wire [2047:0] dataGroup_hi_1556 = {dataGroup_hi_hi_1556, dataGroup_hi_lo_1556};
  wire [7:0]    dataGroup_20_24 = dataGroup_lo_1556[1151:1144];
  wire [2047:0] dataGroup_lo_1557 = {dataGroup_lo_hi_1557, dataGroup_lo_lo_1557};
  wire [2047:0] dataGroup_hi_1557 = {dataGroup_hi_hi_1557, dataGroup_hi_lo_1557};
  wire [7:0]    dataGroup_21_24 = dataGroup_lo_1557[1207:1200];
  wire [2047:0] dataGroup_lo_1558 = {dataGroup_lo_hi_1558, dataGroup_lo_lo_1558};
  wire [2047:0] dataGroup_hi_1558 = {dataGroup_hi_hi_1558, dataGroup_hi_lo_1558};
  wire [7:0]    dataGroup_22_24 = dataGroup_lo_1558[1263:1256];
  wire [2047:0] dataGroup_lo_1559 = {dataGroup_lo_hi_1559, dataGroup_lo_lo_1559};
  wire [2047:0] dataGroup_hi_1559 = {dataGroup_hi_hi_1559, dataGroup_hi_lo_1559};
  wire [7:0]    dataGroup_23_24 = dataGroup_lo_1559[1319:1312];
  wire [2047:0] dataGroup_lo_1560 = {dataGroup_lo_hi_1560, dataGroup_lo_lo_1560};
  wire [2047:0] dataGroup_hi_1560 = {dataGroup_hi_hi_1560, dataGroup_hi_lo_1560};
  wire [7:0]    dataGroup_24_24 = dataGroup_lo_1560[1375:1368];
  wire [2047:0] dataGroup_lo_1561 = {dataGroup_lo_hi_1561, dataGroup_lo_lo_1561};
  wire [2047:0] dataGroup_hi_1561 = {dataGroup_hi_hi_1561, dataGroup_hi_lo_1561};
  wire [7:0]    dataGroup_25_24 = dataGroup_lo_1561[1431:1424];
  wire [2047:0] dataGroup_lo_1562 = {dataGroup_lo_hi_1562, dataGroup_lo_lo_1562};
  wire [2047:0] dataGroup_hi_1562 = {dataGroup_hi_hi_1562, dataGroup_hi_lo_1562};
  wire [7:0]    dataGroup_26_24 = dataGroup_lo_1562[1487:1480];
  wire [2047:0] dataGroup_lo_1563 = {dataGroup_lo_hi_1563, dataGroup_lo_lo_1563};
  wire [2047:0] dataGroup_hi_1563 = {dataGroup_hi_hi_1563, dataGroup_hi_lo_1563};
  wire [7:0]    dataGroup_27_24 = dataGroup_lo_1563[1543:1536];
  wire [2047:0] dataGroup_lo_1564 = {dataGroup_lo_hi_1564, dataGroup_lo_lo_1564};
  wire [2047:0] dataGroup_hi_1564 = {dataGroup_hi_hi_1564, dataGroup_hi_lo_1564};
  wire [7:0]    dataGroup_28_24 = dataGroup_lo_1564[1599:1592];
  wire [2047:0] dataGroup_lo_1565 = {dataGroup_lo_hi_1565, dataGroup_lo_lo_1565};
  wire [2047:0] dataGroup_hi_1565 = {dataGroup_hi_hi_1565, dataGroup_hi_lo_1565};
  wire [7:0]    dataGroup_29_24 = dataGroup_lo_1565[1655:1648];
  wire [2047:0] dataGroup_lo_1566 = {dataGroup_lo_hi_1566, dataGroup_lo_lo_1566};
  wire [2047:0] dataGroup_hi_1566 = {dataGroup_hi_hi_1566, dataGroup_hi_lo_1566};
  wire [7:0]    dataGroup_30_24 = dataGroup_lo_1566[1711:1704];
  wire [2047:0] dataGroup_lo_1567 = {dataGroup_lo_hi_1567, dataGroup_lo_lo_1567};
  wire [2047:0] dataGroup_hi_1567 = {dataGroup_hi_hi_1567, dataGroup_hi_lo_1567};
  wire [7:0]    dataGroup_31_24 = dataGroup_lo_1567[1767:1760];
  wire [2047:0] dataGroup_lo_1568 = {dataGroup_lo_hi_1568, dataGroup_lo_lo_1568};
  wire [2047:0] dataGroup_hi_1568 = {dataGroup_hi_hi_1568, dataGroup_hi_lo_1568};
  wire [7:0]    dataGroup_32_24 = dataGroup_lo_1568[1823:1816];
  wire [2047:0] dataGroup_lo_1569 = {dataGroup_lo_hi_1569, dataGroup_lo_lo_1569};
  wire [2047:0] dataGroup_hi_1569 = {dataGroup_hi_hi_1569, dataGroup_hi_lo_1569};
  wire [7:0]    dataGroup_33_24 = dataGroup_lo_1569[1879:1872];
  wire [2047:0] dataGroup_lo_1570 = {dataGroup_lo_hi_1570, dataGroup_lo_lo_1570};
  wire [2047:0] dataGroup_hi_1570 = {dataGroup_hi_hi_1570, dataGroup_hi_lo_1570};
  wire [7:0]    dataGroup_34_24 = dataGroup_lo_1570[1935:1928];
  wire [2047:0] dataGroup_lo_1571 = {dataGroup_lo_hi_1571, dataGroup_lo_lo_1571};
  wire [2047:0] dataGroup_hi_1571 = {dataGroup_hi_hi_1571, dataGroup_hi_lo_1571};
  wire [7:0]    dataGroup_35_24 = dataGroup_lo_1571[1991:1984];
  wire [2047:0] dataGroup_lo_1572 = {dataGroup_lo_hi_1572, dataGroup_lo_lo_1572};
  wire [2047:0] dataGroup_hi_1572 = {dataGroup_hi_hi_1572, dataGroup_hi_lo_1572};
  wire [7:0]    dataGroup_36_24 = dataGroup_lo_1572[2047:2040];
  wire [2047:0] dataGroup_lo_1573 = {dataGroup_lo_hi_1573, dataGroup_lo_lo_1573};
  wire [2047:0] dataGroup_hi_1573 = {dataGroup_hi_hi_1573, dataGroup_hi_lo_1573};
  wire [7:0]    dataGroup_37_24 = dataGroup_hi_1573[55:48];
  wire [2047:0] dataGroup_lo_1574 = {dataGroup_lo_hi_1574, dataGroup_lo_lo_1574};
  wire [2047:0] dataGroup_hi_1574 = {dataGroup_hi_hi_1574, dataGroup_hi_lo_1574};
  wire [7:0]    dataGroup_38_24 = dataGroup_hi_1574[111:104];
  wire [2047:0] dataGroup_lo_1575 = {dataGroup_lo_hi_1575, dataGroup_lo_lo_1575};
  wire [2047:0] dataGroup_hi_1575 = {dataGroup_hi_hi_1575, dataGroup_hi_lo_1575};
  wire [7:0]    dataGroup_39_24 = dataGroup_hi_1575[167:160];
  wire [2047:0] dataGroup_lo_1576 = {dataGroup_lo_hi_1576, dataGroup_lo_lo_1576};
  wire [2047:0] dataGroup_hi_1576 = {dataGroup_hi_hi_1576, dataGroup_hi_lo_1576};
  wire [7:0]    dataGroup_40_24 = dataGroup_hi_1576[223:216];
  wire [2047:0] dataGroup_lo_1577 = {dataGroup_lo_hi_1577, dataGroup_lo_lo_1577};
  wire [2047:0] dataGroup_hi_1577 = {dataGroup_hi_hi_1577, dataGroup_hi_lo_1577};
  wire [7:0]    dataGroup_41_24 = dataGroup_hi_1577[279:272];
  wire [2047:0] dataGroup_lo_1578 = {dataGroup_lo_hi_1578, dataGroup_lo_lo_1578};
  wire [2047:0] dataGroup_hi_1578 = {dataGroup_hi_hi_1578, dataGroup_hi_lo_1578};
  wire [7:0]    dataGroup_42_24 = dataGroup_hi_1578[335:328];
  wire [2047:0] dataGroup_lo_1579 = {dataGroup_lo_hi_1579, dataGroup_lo_lo_1579};
  wire [2047:0] dataGroup_hi_1579 = {dataGroup_hi_hi_1579, dataGroup_hi_lo_1579};
  wire [7:0]    dataGroup_43_24 = dataGroup_hi_1579[391:384];
  wire [2047:0] dataGroup_lo_1580 = {dataGroup_lo_hi_1580, dataGroup_lo_lo_1580};
  wire [2047:0] dataGroup_hi_1580 = {dataGroup_hi_hi_1580, dataGroup_hi_lo_1580};
  wire [7:0]    dataGroup_44_24 = dataGroup_hi_1580[447:440];
  wire [2047:0] dataGroup_lo_1581 = {dataGroup_lo_hi_1581, dataGroup_lo_lo_1581};
  wire [2047:0] dataGroup_hi_1581 = {dataGroup_hi_hi_1581, dataGroup_hi_lo_1581};
  wire [7:0]    dataGroup_45_24 = dataGroup_hi_1581[503:496];
  wire [2047:0] dataGroup_lo_1582 = {dataGroup_lo_hi_1582, dataGroup_lo_lo_1582};
  wire [2047:0] dataGroup_hi_1582 = {dataGroup_hi_hi_1582, dataGroup_hi_lo_1582};
  wire [7:0]    dataGroup_46_24 = dataGroup_hi_1582[559:552];
  wire [2047:0] dataGroup_lo_1583 = {dataGroup_lo_hi_1583, dataGroup_lo_lo_1583};
  wire [2047:0] dataGroup_hi_1583 = {dataGroup_hi_hi_1583, dataGroup_hi_lo_1583};
  wire [7:0]    dataGroup_47_24 = dataGroup_hi_1583[615:608];
  wire [2047:0] dataGroup_lo_1584 = {dataGroup_lo_hi_1584, dataGroup_lo_lo_1584};
  wire [2047:0] dataGroup_hi_1584 = {dataGroup_hi_hi_1584, dataGroup_hi_lo_1584};
  wire [7:0]    dataGroup_48_24 = dataGroup_hi_1584[671:664];
  wire [2047:0] dataGroup_lo_1585 = {dataGroup_lo_hi_1585, dataGroup_lo_lo_1585};
  wire [2047:0] dataGroup_hi_1585 = {dataGroup_hi_hi_1585, dataGroup_hi_lo_1585};
  wire [7:0]    dataGroup_49_24 = dataGroup_hi_1585[727:720];
  wire [2047:0] dataGroup_lo_1586 = {dataGroup_lo_hi_1586, dataGroup_lo_lo_1586};
  wire [2047:0] dataGroup_hi_1586 = {dataGroup_hi_hi_1586, dataGroup_hi_lo_1586};
  wire [7:0]    dataGroup_50_24 = dataGroup_hi_1586[783:776];
  wire [2047:0] dataGroup_lo_1587 = {dataGroup_lo_hi_1587, dataGroup_lo_lo_1587};
  wire [2047:0] dataGroup_hi_1587 = {dataGroup_hi_hi_1587, dataGroup_hi_lo_1587};
  wire [7:0]    dataGroup_51_24 = dataGroup_hi_1587[839:832];
  wire [2047:0] dataGroup_lo_1588 = {dataGroup_lo_hi_1588, dataGroup_lo_lo_1588};
  wire [2047:0] dataGroup_hi_1588 = {dataGroup_hi_hi_1588, dataGroup_hi_lo_1588};
  wire [7:0]    dataGroup_52_24 = dataGroup_hi_1588[895:888];
  wire [2047:0] dataGroup_lo_1589 = {dataGroup_lo_hi_1589, dataGroup_lo_lo_1589};
  wire [2047:0] dataGroup_hi_1589 = {dataGroup_hi_hi_1589, dataGroup_hi_lo_1589};
  wire [7:0]    dataGroup_53_24 = dataGroup_hi_1589[951:944];
  wire [2047:0] dataGroup_lo_1590 = {dataGroup_lo_hi_1590, dataGroup_lo_lo_1590};
  wire [2047:0] dataGroup_hi_1590 = {dataGroup_hi_hi_1590, dataGroup_hi_lo_1590};
  wire [7:0]    dataGroup_54_24 = dataGroup_hi_1590[1007:1000];
  wire [2047:0] dataGroup_lo_1591 = {dataGroup_lo_hi_1591, dataGroup_lo_lo_1591};
  wire [2047:0] dataGroup_hi_1591 = {dataGroup_hi_hi_1591, dataGroup_hi_lo_1591};
  wire [7:0]    dataGroup_55_24 = dataGroup_hi_1591[1063:1056];
  wire [2047:0] dataGroup_lo_1592 = {dataGroup_lo_hi_1592, dataGroup_lo_lo_1592};
  wire [2047:0] dataGroup_hi_1592 = {dataGroup_hi_hi_1592, dataGroup_hi_lo_1592};
  wire [7:0]    dataGroup_56_24 = dataGroup_hi_1592[1119:1112];
  wire [2047:0] dataGroup_lo_1593 = {dataGroup_lo_hi_1593, dataGroup_lo_lo_1593};
  wire [2047:0] dataGroup_hi_1593 = {dataGroup_hi_hi_1593, dataGroup_hi_lo_1593};
  wire [7:0]    dataGroup_57_24 = dataGroup_hi_1593[1175:1168];
  wire [2047:0] dataGroup_lo_1594 = {dataGroup_lo_hi_1594, dataGroup_lo_lo_1594};
  wire [2047:0] dataGroup_hi_1594 = {dataGroup_hi_hi_1594, dataGroup_hi_lo_1594};
  wire [7:0]    dataGroup_58_24 = dataGroup_hi_1594[1231:1224];
  wire [2047:0] dataGroup_lo_1595 = {dataGroup_lo_hi_1595, dataGroup_lo_lo_1595};
  wire [2047:0] dataGroup_hi_1595 = {dataGroup_hi_hi_1595, dataGroup_hi_lo_1595};
  wire [7:0]    dataGroup_59_24 = dataGroup_hi_1595[1287:1280];
  wire [2047:0] dataGroup_lo_1596 = {dataGroup_lo_hi_1596, dataGroup_lo_lo_1596};
  wire [2047:0] dataGroup_hi_1596 = {dataGroup_hi_hi_1596, dataGroup_hi_lo_1596};
  wire [7:0]    dataGroup_60_24 = dataGroup_hi_1596[1343:1336];
  wire [2047:0] dataGroup_lo_1597 = {dataGroup_lo_hi_1597, dataGroup_lo_lo_1597};
  wire [2047:0] dataGroup_hi_1597 = {dataGroup_hi_hi_1597, dataGroup_hi_lo_1597};
  wire [7:0]    dataGroup_61_24 = dataGroup_hi_1597[1399:1392];
  wire [2047:0] dataGroup_lo_1598 = {dataGroup_lo_hi_1598, dataGroup_lo_lo_1598};
  wire [2047:0] dataGroup_hi_1598 = {dataGroup_hi_hi_1598, dataGroup_hi_lo_1598};
  wire [7:0]    dataGroup_62_24 = dataGroup_hi_1598[1455:1448];
  wire [2047:0] dataGroup_lo_1599 = {dataGroup_lo_hi_1599, dataGroup_lo_lo_1599};
  wire [2047:0] dataGroup_hi_1599 = {dataGroup_hi_hi_1599, dataGroup_hi_lo_1599};
  wire [7:0]    dataGroup_63_24 = dataGroup_hi_1599[1511:1504];
  wire [15:0]   res_lo_lo_lo_lo_lo_24 = {dataGroup_1_24, dataGroup_0_24};
  wire [15:0]   res_lo_lo_lo_lo_hi_24 = {dataGroup_3_24, dataGroup_2_24};
  wire [31:0]   res_lo_lo_lo_lo_24 = {res_lo_lo_lo_lo_hi_24, res_lo_lo_lo_lo_lo_24};
  wire [15:0]   res_lo_lo_lo_hi_lo_24 = {dataGroup_5_24, dataGroup_4_24};
  wire [15:0]   res_lo_lo_lo_hi_hi_24 = {dataGroup_7_24, dataGroup_6_24};
  wire [31:0]   res_lo_lo_lo_hi_24 = {res_lo_lo_lo_hi_hi_24, res_lo_lo_lo_hi_lo_24};
  wire [63:0]   res_lo_lo_lo_24 = {res_lo_lo_lo_hi_24, res_lo_lo_lo_lo_24};
  wire [15:0]   res_lo_lo_hi_lo_lo_24 = {dataGroup_9_24, dataGroup_8_24};
  wire [15:0]   res_lo_lo_hi_lo_hi_24 = {dataGroup_11_24, dataGroup_10_24};
  wire [31:0]   res_lo_lo_hi_lo_24 = {res_lo_lo_hi_lo_hi_24, res_lo_lo_hi_lo_lo_24};
  wire [15:0]   res_lo_lo_hi_hi_lo_24 = {dataGroup_13_24, dataGroup_12_24};
  wire [15:0]   res_lo_lo_hi_hi_hi_24 = {dataGroup_15_24, dataGroup_14_24};
  wire [31:0]   res_lo_lo_hi_hi_24 = {res_lo_lo_hi_hi_hi_24, res_lo_lo_hi_hi_lo_24};
  wire [63:0]   res_lo_lo_hi_24 = {res_lo_lo_hi_hi_24, res_lo_lo_hi_lo_24};
  wire [127:0]  res_lo_lo_24 = {res_lo_lo_hi_24, res_lo_lo_lo_24};
  wire [15:0]   res_lo_hi_lo_lo_lo_24 = {dataGroup_17_24, dataGroup_16_24};
  wire [15:0]   res_lo_hi_lo_lo_hi_24 = {dataGroup_19_24, dataGroup_18_24};
  wire [31:0]   res_lo_hi_lo_lo_24 = {res_lo_hi_lo_lo_hi_24, res_lo_hi_lo_lo_lo_24};
  wire [15:0]   res_lo_hi_lo_hi_lo_24 = {dataGroup_21_24, dataGroup_20_24};
  wire [15:0]   res_lo_hi_lo_hi_hi_24 = {dataGroup_23_24, dataGroup_22_24};
  wire [31:0]   res_lo_hi_lo_hi_24 = {res_lo_hi_lo_hi_hi_24, res_lo_hi_lo_hi_lo_24};
  wire [63:0]   res_lo_hi_lo_24 = {res_lo_hi_lo_hi_24, res_lo_hi_lo_lo_24};
  wire [15:0]   res_lo_hi_hi_lo_lo_24 = {dataGroup_25_24, dataGroup_24_24};
  wire [15:0]   res_lo_hi_hi_lo_hi_24 = {dataGroup_27_24, dataGroup_26_24};
  wire [31:0]   res_lo_hi_hi_lo_24 = {res_lo_hi_hi_lo_hi_24, res_lo_hi_hi_lo_lo_24};
  wire [15:0]   res_lo_hi_hi_hi_lo_24 = {dataGroup_29_24, dataGroup_28_24};
  wire [15:0]   res_lo_hi_hi_hi_hi_24 = {dataGroup_31_24, dataGroup_30_24};
  wire [31:0]   res_lo_hi_hi_hi_24 = {res_lo_hi_hi_hi_hi_24, res_lo_hi_hi_hi_lo_24};
  wire [63:0]   res_lo_hi_hi_24 = {res_lo_hi_hi_hi_24, res_lo_hi_hi_lo_24};
  wire [127:0]  res_lo_hi_24 = {res_lo_hi_hi_24, res_lo_hi_lo_24};
  wire [255:0]  res_lo_24 = {res_lo_hi_24, res_lo_lo_24};
  wire [15:0]   res_hi_lo_lo_lo_lo_24 = {dataGroup_33_24, dataGroup_32_24};
  wire [15:0]   res_hi_lo_lo_lo_hi_24 = {dataGroup_35_24, dataGroup_34_24};
  wire [31:0]   res_hi_lo_lo_lo_24 = {res_hi_lo_lo_lo_hi_24, res_hi_lo_lo_lo_lo_24};
  wire [15:0]   res_hi_lo_lo_hi_lo_24 = {dataGroup_37_24, dataGroup_36_24};
  wire [15:0]   res_hi_lo_lo_hi_hi_24 = {dataGroup_39_24, dataGroup_38_24};
  wire [31:0]   res_hi_lo_lo_hi_24 = {res_hi_lo_lo_hi_hi_24, res_hi_lo_lo_hi_lo_24};
  wire [63:0]   res_hi_lo_lo_24 = {res_hi_lo_lo_hi_24, res_hi_lo_lo_lo_24};
  wire [15:0]   res_hi_lo_hi_lo_lo_24 = {dataGroup_41_24, dataGroup_40_24};
  wire [15:0]   res_hi_lo_hi_lo_hi_24 = {dataGroup_43_24, dataGroup_42_24};
  wire [31:0]   res_hi_lo_hi_lo_24 = {res_hi_lo_hi_lo_hi_24, res_hi_lo_hi_lo_lo_24};
  wire [15:0]   res_hi_lo_hi_hi_lo_24 = {dataGroup_45_24, dataGroup_44_24};
  wire [15:0]   res_hi_lo_hi_hi_hi_24 = {dataGroup_47_24, dataGroup_46_24};
  wire [31:0]   res_hi_lo_hi_hi_24 = {res_hi_lo_hi_hi_hi_24, res_hi_lo_hi_hi_lo_24};
  wire [63:0]   res_hi_lo_hi_24 = {res_hi_lo_hi_hi_24, res_hi_lo_hi_lo_24};
  wire [127:0]  res_hi_lo_24 = {res_hi_lo_hi_24, res_hi_lo_lo_24};
  wire [15:0]   res_hi_hi_lo_lo_lo_24 = {dataGroup_49_24, dataGroup_48_24};
  wire [15:0]   res_hi_hi_lo_lo_hi_24 = {dataGroup_51_24, dataGroup_50_24};
  wire [31:0]   res_hi_hi_lo_lo_24 = {res_hi_hi_lo_lo_hi_24, res_hi_hi_lo_lo_lo_24};
  wire [15:0]   res_hi_hi_lo_hi_lo_24 = {dataGroup_53_24, dataGroup_52_24};
  wire [15:0]   res_hi_hi_lo_hi_hi_24 = {dataGroup_55_24, dataGroup_54_24};
  wire [31:0]   res_hi_hi_lo_hi_24 = {res_hi_hi_lo_hi_hi_24, res_hi_hi_lo_hi_lo_24};
  wire [63:0]   res_hi_hi_lo_24 = {res_hi_hi_lo_hi_24, res_hi_hi_lo_lo_24};
  wire [15:0]   res_hi_hi_hi_lo_lo_24 = {dataGroup_57_24, dataGroup_56_24};
  wire [15:0]   res_hi_hi_hi_lo_hi_24 = {dataGroup_59_24, dataGroup_58_24};
  wire [31:0]   res_hi_hi_hi_lo_24 = {res_hi_hi_hi_lo_hi_24, res_hi_hi_hi_lo_lo_24};
  wire [15:0]   res_hi_hi_hi_hi_lo_24 = {dataGroup_61_24, dataGroup_60_24};
  wire [15:0]   res_hi_hi_hi_hi_hi_24 = {dataGroup_63_24, dataGroup_62_24};
  wire [31:0]   res_hi_hi_hi_hi_24 = {res_hi_hi_hi_hi_hi_24, res_hi_hi_hi_hi_lo_24};
  wire [63:0]   res_hi_hi_hi_24 = {res_hi_hi_hi_hi_24, res_hi_hi_hi_lo_24};
  wire [127:0]  res_hi_hi_24 = {res_hi_hi_hi_24, res_hi_hi_lo_24};
  wire [255:0]  res_hi_24 = {res_hi_hi_24, res_hi_lo_24};
  wire [511:0]  res_51 = {res_hi_24, res_lo_24};
  wire [2047:0] dataGroup_lo_1600 = {dataGroup_lo_hi_1600, dataGroup_lo_lo_1600};
  wire [2047:0] dataGroup_hi_1600 = {dataGroup_hi_hi_1600, dataGroup_hi_lo_1600};
  wire [7:0]    dataGroup_0_25 = dataGroup_lo_1600[39:32];
  wire [2047:0] dataGroup_lo_1601 = {dataGroup_lo_hi_1601, dataGroup_lo_lo_1601};
  wire [2047:0] dataGroup_hi_1601 = {dataGroup_hi_hi_1601, dataGroup_hi_lo_1601};
  wire [7:0]    dataGroup_1_25 = dataGroup_lo_1601[95:88];
  wire [2047:0] dataGroup_lo_1602 = {dataGroup_lo_hi_1602, dataGroup_lo_lo_1602};
  wire [2047:0] dataGroup_hi_1602 = {dataGroup_hi_hi_1602, dataGroup_hi_lo_1602};
  wire [7:0]    dataGroup_2_25 = dataGroup_lo_1602[151:144];
  wire [2047:0] dataGroup_lo_1603 = {dataGroup_lo_hi_1603, dataGroup_lo_lo_1603};
  wire [2047:0] dataGroup_hi_1603 = {dataGroup_hi_hi_1603, dataGroup_hi_lo_1603};
  wire [7:0]    dataGroup_3_25 = dataGroup_lo_1603[207:200];
  wire [2047:0] dataGroup_lo_1604 = {dataGroup_lo_hi_1604, dataGroup_lo_lo_1604};
  wire [2047:0] dataGroup_hi_1604 = {dataGroup_hi_hi_1604, dataGroup_hi_lo_1604};
  wire [7:0]    dataGroup_4_25 = dataGroup_lo_1604[263:256];
  wire [2047:0] dataGroup_lo_1605 = {dataGroup_lo_hi_1605, dataGroup_lo_lo_1605};
  wire [2047:0] dataGroup_hi_1605 = {dataGroup_hi_hi_1605, dataGroup_hi_lo_1605};
  wire [7:0]    dataGroup_5_25 = dataGroup_lo_1605[319:312];
  wire [2047:0] dataGroup_lo_1606 = {dataGroup_lo_hi_1606, dataGroup_lo_lo_1606};
  wire [2047:0] dataGroup_hi_1606 = {dataGroup_hi_hi_1606, dataGroup_hi_lo_1606};
  wire [7:0]    dataGroup_6_25 = dataGroup_lo_1606[375:368];
  wire [2047:0] dataGroup_lo_1607 = {dataGroup_lo_hi_1607, dataGroup_lo_lo_1607};
  wire [2047:0] dataGroup_hi_1607 = {dataGroup_hi_hi_1607, dataGroup_hi_lo_1607};
  wire [7:0]    dataGroup_7_25 = dataGroup_lo_1607[431:424];
  wire [2047:0] dataGroup_lo_1608 = {dataGroup_lo_hi_1608, dataGroup_lo_lo_1608};
  wire [2047:0] dataGroup_hi_1608 = {dataGroup_hi_hi_1608, dataGroup_hi_lo_1608};
  wire [7:0]    dataGroup_8_25 = dataGroup_lo_1608[487:480];
  wire [2047:0] dataGroup_lo_1609 = {dataGroup_lo_hi_1609, dataGroup_lo_lo_1609};
  wire [2047:0] dataGroup_hi_1609 = {dataGroup_hi_hi_1609, dataGroup_hi_lo_1609};
  wire [7:0]    dataGroup_9_25 = dataGroup_lo_1609[543:536];
  wire [2047:0] dataGroup_lo_1610 = {dataGroup_lo_hi_1610, dataGroup_lo_lo_1610};
  wire [2047:0] dataGroup_hi_1610 = {dataGroup_hi_hi_1610, dataGroup_hi_lo_1610};
  wire [7:0]    dataGroup_10_25 = dataGroup_lo_1610[599:592];
  wire [2047:0] dataGroup_lo_1611 = {dataGroup_lo_hi_1611, dataGroup_lo_lo_1611};
  wire [2047:0] dataGroup_hi_1611 = {dataGroup_hi_hi_1611, dataGroup_hi_lo_1611};
  wire [7:0]    dataGroup_11_25 = dataGroup_lo_1611[655:648];
  wire [2047:0] dataGroup_lo_1612 = {dataGroup_lo_hi_1612, dataGroup_lo_lo_1612};
  wire [2047:0] dataGroup_hi_1612 = {dataGroup_hi_hi_1612, dataGroup_hi_lo_1612};
  wire [7:0]    dataGroup_12_25 = dataGroup_lo_1612[711:704];
  wire [2047:0] dataGroup_lo_1613 = {dataGroup_lo_hi_1613, dataGroup_lo_lo_1613};
  wire [2047:0] dataGroup_hi_1613 = {dataGroup_hi_hi_1613, dataGroup_hi_lo_1613};
  wire [7:0]    dataGroup_13_25 = dataGroup_lo_1613[767:760];
  wire [2047:0] dataGroup_lo_1614 = {dataGroup_lo_hi_1614, dataGroup_lo_lo_1614};
  wire [2047:0] dataGroup_hi_1614 = {dataGroup_hi_hi_1614, dataGroup_hi_lo_1614};
  wire [7:0]    dataGroup_14_25 = dataGroup_lo_1614[823:816];
  wire [2047:0] dataGroup_lo_1615 = {dataGroup_lo_hi_1615, dataGroup_lo_lo_1615};
  wire [2047:0] dataGroup_hi_1615 = {dataGroup_hi_hi_1615, dataGroup_hi_lo_1615};
  wire [7:0]    dataGroup_15_25 = dataGroup_lo_1615[879:872];
  wire [2047:0] dataGroup_lo_1616 = {dataGroup_lo_hi_1616, dataGroup_lo_lo_1616};
  wire [2047:0] dataGroup_hi_1616 = {dataGroup_hi_hi_1616, dataGroup_hi_lo_1616};
  wire [7:0]    dataGroup_16_25 = dataGroup_lo_1616[935:928];
  wire [2047:0] dataGroup_lo_1617 = {dataGroup_lo_hi_1617, dataGroup_lo_lo_1617};
  wire [2047:0] dataGroup_hi_1617 = {dataGroup_hi_hi_1617, dataGroup_hi_lo_1617};
  wire [7:0]    dataGroup_17_25 = dataGroup_lo_1617[991:984];
  wire [2047:0] dataGroup_lo_1618 = {dataGroup_lo_hi_1618, dataGroup_lo_lo_1618};
  wire [2047:0] dataGroup_hi_1618 = {dataGroup_hi_hi_1618, dataGroup_hi_lo_1618};
  wire [7:0]    dataGroup_18_25 = dataGroup_lo_1618[1047:1040];
  wire [2047:0] dataGroup_lo_1619 = {dataGroup_lo_hi_1619, dataGroup_lo_lo_1619};
  wire [2047:0] dataGroup_hi_1619 = {dataGroup_hi_hi_1619, dataGroup_hi_lo_1619};
  wire [7:0]    dataGroup_19_25 = dataGroup_lo_1619[1103:1096];
  wire [2047:0] dataGroup_lo_1620 = {dataGroup_lo_hi_1620, dataGroup_lo_lo_1620};
  wire [2047:0] dataGroup_hi_1620 = {dataGroup_hi_hi_1620, dataGroup_hi_lo_1620};
  wire [7:0]    dataGroup_20_25 = dataGroup_lo_1620[1159:1152];
  wire [2047:0] dataGroup_lo_1621 = {dataGroup_lo_hi_1621, dataGroup_lo_lo_1621};
  wire [2047:0] dataGroup_hi_1621 = {dataGroup_hi_hi_1621, dataGroup_hi_lo_1621};
  wire [7:0]    dataGroup_21_25 = dataGroup_lo_1621[1215:1208];
  wire [2047:0] dataGroup_lo_1622 = {dataGroup_lo_hi_1622, dataGroup_lo_lo_1622};
  wire [2047:0] dataGroup_hi_1622 = {dataGroup_hi_hi_1622, dataGroup_hi_lo_1622};
  wire [7:0]    dataGroup_22_25 = dataGroup_lo_1622[1271:1264];
  wire [2047:0] dataGroup_lo_1623 = {dataGroup_lo_hi_1623, dataGroup_lo_lo_1623};
  wire [2047:0] dataGroup_hi_1623 = {dataGroup_hi_hi_1623, dataGroup_hi_lo_1623};
  wire [7:0]    dataGroup_23_25 = dataGroup_lo_1623[1327:1320];
  wire [2047:0] dataGroup_lo_1624 = {dataGroup_lo_hi_1624, dataGroup_lo_lo_1624};
  wire [2047:0] dataGroup_hi_1624 = {dataGroup_hi_hi_1624, dataGroup_hi_lo_1624};
  wire [7:0]    dataGroup_24_25 = dataGroup_lo_1624[1383:1376];
  wire [2047:0] dataGroup_lo_1625 = {dataGroup_lo_hi_1625, dataGroup_lo_lo_1625};
  wire [2047:0] dataGroup_hi_1625 = {dataGroup_hi_hi_1625, dataGroup_hi_lo_1625};
  wire [7:0]    dataGroup_25_25 = dataGroup_lo_1625[1439:1432];
  wire [2047:0] dataGroup_lo_1626 = {dataGroup_lo_hi_1626, dataGroup_lo_lo_1626};
  wire [2047:0] dataGroup_hi_1626 = {dataGroup_hi_hi_1626, dataGroup_hi_lo_1626};
  wire [7:0]    dataGroup_26_25 = dataGroup_lo_1626[1495:1488];
  wire [2047:0] dataGroup_lo_1627 = {dataGroup_lo_hi_1627, dataGroup_lo_lo_1627};
  wire [2047:0] dataGroup_hi_1627 = {dataGroup_hi_hi_1627, dataGroup_hi_lo_1627};
  wire [7:0]    dataGroup_27_25 = dataGroup_lo_1627[1551:1544];
  wire [2047:0] dataGroup_lo_1628 = {dataGroup_lo_hi_1628, dataGroup_lo_lo_1628};
  wire [2047:0] dataGroup_hi_1628 = {dataGroup_hi_hi_1628, dataGroup_hi_lo_1628};
  wire [7:0]    dataGroup_28_25 = dataGroup_lo_1628[1607:1600];
  wire [2047:0] dataGroup_lo_1629 = {dataGroup_lo_hi_1629, dataGroup_lo_lo_1629};
  wire [2047:0] dataGroup_hi_1629 = {dataGroup_hi_hi_1629, dataGroup_hi_lo_1629};
  wire [7:0]    dataGroup_29_25 = dataGroup_lo_1629[1663:1656];
  wire [2047:0] dataGroup_lo_1630 = {dataGroup_lo_hi_1630, dataGroup_lo_lo_1630};
  wire [2047:0] dataGroup_hi_1630 = {dataGroup_hi_hi_1630, dataGroup_hi_lo_1630};
  wire [7:0]    dataGroup_30_25 = dataGroup_lo_1630[1719:1712];
  wire [2047:0] dataGroup_lo_1631 = {dataGroup_lo_hi_1631, dataGroup_lo_lo_1631};
  wire [2047:0] dataGroup_hi_1631 = {dataGroup_hi_hi_1631, dataGroup_hi_lo_1631};
  wire [7:0]    dataGroup_31_25 = dataGroup_lo_1631[1775:1768];
  wire [2047:0] dataGroup_lo_1632 = {dataGroup_lo_hi_1632, dataGroup_lo_lo_1632};
  wire [2047:0] dataGroup_hi_1632 = {dataGroup_hi_hi_1632, dataGroup_hi_lo_1632};
  wire [7:0]    dataGroup_32_25 = dataGroup_lo_1632[1831:1824];
  wire [2047:0] dataGroup_lo_1633 = {dataGroup_lo_hi_1633, dataGroup_lo_lo_1633};
  wire [2047:0] dataGroup_hi_1633 = {dataGroup_hi_hi_1633, dataGroup_hi_lo_1633};
  wire [7:0]    dataGroup_33_25 = dataGroup_lo_1633[1887:1880];
  wire [2047:0] dataGroup_lo_1634 = {dataGroup_lo_hi_1634, dataGroup_lo_lo_1634};
  wire [2047:0] dataGroup_hi_1634 = {dataGroup_hi_hi_1634, dataGroup_hi_lo_1634};
  wire [7:0]    dataGroup_34_25 = dataGroup_lo_1634[1943:1936];
  wire [2047:0] dataGroup_lo_1635 = {dataGroup_lo_hi_1635, dataGroup_lo_lo_1635};
  wire [2047:0] dataGroup_hi_1635 = {dataGroup_hi_hi_1635, dataGroup_hi_lo_1635};
  wire [7:0]    dataGroup_35_25 = dataGroup_lo_1635[1999:1992];
  wire [2047:0] dataGroup_lo_1636 = {dataGroup_lo_hi_1636, dataGroup_lo_lo_1636};
  wire [2047:0] dataGroup_hi_1636 = {dataGroup_hi_hi_1636, dataGroup_hi_lo_1636};
  wire [7:0]    dataGroup_36_25 = dataGroup_hi_1636[7:0];
  wire [2047:0] dataGroup_lo_1637 = {dataGroup_lo_hi_1637, dataGroup_lo_lo_1637};
  wire [2047:0] dataGroup_hi_1637 = {dataGroup_hi_hi_1637, dataGroup_hi_lo_1637};
  wire [7:0]    dataGroup_37_25 = dataGroup_hi_1637[63:56];
  wire [2047:0] dataGroup_lo_1638 = {dataGroup_lo_hi_1638, dataGroup_lo_lo_1638};
  wire [2047:0] dataGroup_hi_1638 = {dataGroup_hi_hi_1638, dataGroup_hi_lo_1638};
  wire [7:0]    dataGroup_38_25 = dataGroup_hi_1638[119:112];
  wire [2047:0] dataGroup_lo_1639 = {dataGroup_lo_hi_1639, dataGroup_lo_lo_1639};
  wire [2047:0] dataGroup_hi_1639 = {dataGroup_hi_hi_1639, dataGroup_hi_lo_1639};
  wire [7:0]    dataGroup_39_25 = dataGroup_hi_1639[175:168];
  wire [2047:0] dataGroup_lo_1640 = {dataGroup_lo_hi_1640, dataGroup_lo_lo_1640};
  wire [2047:0] dataGroup_hi_1640 = {dataGroup_hi_hi_1640, dataGroup_hi_lo_1640};
  wire [7:0]    dataGroup_40_25 = dataGroup_hi_1640[231:224];
  wire [2047:0] dataGroup_lo_1641 = {dataGroup_lo_hi_1641, dataGroup_lo_lo_1641};
  wire [2047:0] dataGroup_hi_1641 = {dataGroup_hi_hi_1641, dataGroup_hi_lo_1641};
  wire [7:0]    dataGroup_41_25 = dataGroup_hi_1641[287:280];
  wire [2047:0] dataGroup_lo_1642 = {dataGroup_lo_hi_1642, dataGroup_lo_lo_1642};
  wire [2047:0] dataGroup_hi_1642 = {dataGroup_hi_hi_1642, dataGroup_hi_lo_1642};
  wire [7:0]    dataGroup_42_25 = dataGroup_hi_1642[343:336];
  wire [2047:0] dataGroup_lo_1643 = {dataGroup_lo_hi_1643, dataGroup_lo_lo_1643};
  wire [2047:0] dataGroup_hi_1643 = {dataGroup_hi_hi_1643, dataGroup_hi_lo_1643};
  wire [7:0]    dataGroup_43_25 = dataGroup_hi_1643[399:392];
  wire [2047:0] dataGroup_lo_1644 = {dataGroup_lo_hi_1644, dataGroup_lo_lo_1644};
  wire [2047:0] dataGroup_hi_1644 = {dataGroup_hi_hi_1644, dataGroup_hi_lo_1644};
  wire [7:0]    dataGroup_44_25 = dataGroup_hi_1644[455:448];
  wire [2047:0] dataGroup_lo_1645 = {dataGroup_lo_hi_1645, dataGroup_lo_lo_1645};
  wire [2047:0] dataGroup_hi_1645 = {dataGroup_hi_hi_1645, dataGroup_hi_lo_1645};
  wire [7:0]    dataGroup_45_25 = dataGroup_hi_1645[511:504];
  wire [2047:0] dataGroup_lo_1646 = {dataGroup_lo_hi_1646, dataGroup_lo_lo_1646};
  wire [2047:0] dataGroup_hi_1646 = {dataGroup_hi_hi_1646, dataGroup_hi_lo_1646};
  wire [7:0]    dataGroup_46_25 = dataGroup_hi_1646[567:560];
  wire [2047:0] dataGroup_lo_1647 = {dataGroup_lo_hi_1647, dataGroup_lo_lo_1647};
  wire [2047:0] dataGroup_hi_1647 = {dataGroup_hi_hi_1647, dataGroup_hi_lo_1647};
  wire [7:0]    dataGroup_47_25 = dataGroup_hi_1647[623:616];
  wire [2047:0] dataGroup_lo_1648 = {dataGroup_lo_hi_1648, dataGroup_lo_lo_1648};
  wire [2047:0] dataGroup_hi_1648 = {dataGroup_hi_hi_1648, dataGroup_hi_lo_1648};
  wire [7:0]    dataGroup_48_25 = dataGroup_hi_1648[679:672];
  wire [2047:0] dataGroup_lo_1649 = {dataGroup_lo_hi_1649, dataGroup_lo_lo_1649};
  wire [2047:0] dataGroup_hi_1649 = {dataGroup_hi_hi_1649, dataGroup_hi_lo_1649};
  wire [7:0]    dataGroup_49_25 = dataGroup_hi_1649[735:728];
  wire [2047:0] dataGroup_lo_1650 = {dataGroup_lo_hi_1650, dataGroup_lo_lo_1650};
  wire [2047:0] dataGroup_hi_1650 = {dataGroup_hi_hi_1650, dataGroup_hi_lo_1650};
  wire [7:0]    dataGroup_50_25 = dataGroup_hi_1650[791:784];
  wire [2047:0] dataGroup_lo_1651 = {dataGroup_lo_hi_1651, dataGroup_lo_lo_1651};
  wire [2047:0] dataGroup_hi_1651 = {dataGroup_hi_hi_1651, dataGroup_hi_lo_1651};
  wire [7:0]    dataGroup_51_25 = dataGroup_hi_1651[847:840];
  wire [2047:0] dataGroup_lo_1652 = {dataGroup_lo_hi_1652, dataGroup_lo_lo_1652};
  wire [2047:0] dataGroup_hi_1652 = {dataGroup_hi_hi_1652, dataGroup_hi_lo_1652};
  wire [7:0]    dataGroup_52_25 = dataGroup_hi_1652[903:896];
  wire [2047:0] dataGroup_lo_1653 = {dataGroup_lo_hi_1653, dataGroup_lo_lo_1653};
  wire [2047:0] dataGroup_hi_1653 = {dataGroup_hi_hi_1653, dataGroup_hi_lo_1653};
  wire [7:0]    dataGroup_53_25 = dataGroup_hi_1653[959:952];
  wire [2047:0] dataGroup_lo_1654 = {dataGroup_lo_hi_1654, dataGroup_lo_lo_1654};
  wire [2047:0] dataGroup_hi_1654 = {dataGroup_hi_hi_1654, dataGroup_hi_lo_1654};
  wire [7:0]    dataGroup_54_25 = dataGroup_hi_1654[1015:1008];
  wire [2047:0] dataGroup_lo_1655 = {dataGroup_lo_hi_1655, dataGroup_lo_lo_1655};
  wire [2047:0] dataGroup_hi_1655 = {dataGroup_hi_hi_1655, dataGroup_hi_lo_1655};
  wire [7:0]    dataGroup_55_25 = dataGroup_hi_1655[1071:1064];
  wire [2047:0] dataGroup_lo_1656 = {dataGroup_lo_hi_1656, dataGroup_lo_lo_1656};
  wire [2047:0] dataGroup_hi_1656 = {dataGroup_hi_hi_1656, dataGroup_hi_lo_1656};
  wire [7:0]    dataGroup_56_25 = dataGroup_hi_1656[1127:1120];
  wire [2047:0] dataGroup_lo_1657 = {dataGroup_lo_hi_1657, dataGroup_lo_lo_1657};
  wire [2047:0] dataGroup_hi_1657 = {dataGroup_hi_hi_1657, dataGroup_hi_lo_1657};
  wire [7:0]    dataGroup_57_25 = dataGroup_hi_1657[1183:1176];
  wire [2047:0] dataGroup_lo_1658 = {dataGroup_lo_hi_1658, dataGroup_lo_lo_1658};
  wire [2047:0] dataGroup_hi_1658 = {dataGroup_hi_hi_1658, dataGroup_hi_lo_1658};
  wire [7:0]    dataGroup_58_25 = dataGroup_hi_1658[1239:1232];
  wire [2047:0] dataGroup_lo_1659 = {dataGroup_lo_hi_1659, dataGroup_lo_lo_1659};
  wire [2047:0] dataGroup_hi_1659 = {dataGroup_hi_hi_1659, dataGroup_hi_lo_1659};
  wire [7:0]    dataGroup_59_25 = dataGroup_hi_1659[1295:1288];
  wire [2047:0] dataGroup_lo_1660 = {dataGroup_lo_hi_1660, dataGroup_lo_lo_1660};
  wire [2047:0] dataGroup_hi_1660 = {dataGroup_hi_hi_1660, dataGroup_hi_lo_1660};
  wire [7:0]    dataGroup_60_25 = dataGroup_hi_1660[1351:1344];
  wire [2047:0] dataGroup_lo_1661 = {dataGroup_lo_hi_1661, dataGroup_lo_lo_1661};
  wire [2047:0] dataGroup_hi_1661 = {dataGroup_hi_hi_1661, dataGroup_hi_lo_1661};
  wire [7:0]    dataGroup_61_25 = dataGroup_hi_1661[1407:1400];
  wire [2047:0] dataGroup_lo_1662 = {dataGroup_lo_hi_1662, dataGroup_lo_lo_1662};
  wire [2047:0] dataGroup_hi_1662 = {dataGroup_hi_hi_1662, dataGroup_hi_lo_1662};
  wire [7:0]    dataGroup_62_25 = dataGroup_hi_1662[1463:1456];
  wire [2047:0] dataGroup_lo_1663 = {dataGroup_lo_hi_1663, dataGroup_lo_lo_1663};
  wire [2047:0] dataGroup_hi_1663 = {dataGroup_hi_hi_1663, dataGroup_hi_lo_1663};
  wire [7:0]    dataGroup_63_25 = dataGroup_hi_1663[1519:1512];
  wire [15:0]   res_lo_lo_lo_lo_lo_25 = {dataGroup_1_25, dataGroup_0_25};
  wire [15:0]   res_lo_lo_lo_lo_hi_25 = {dataGroup_3_25, dataGroup_2_25};
  wire [31:0]   res_lo_lo_lo_lo_25 = {res_lo_lo_lo_lo_hi_25, res_lo_lo_lo_lo_lo_25};
  wire [15:0]   res_lo_lo_lo_hi_lo_25 = {dataGroup_5_25, dataGroup_4_25};
  wire [15:0]   res_lo_lo_lo_hi_hi_25 = {dataGroup_7_25, dataGroup_6_25};
  wire [31:0]   res_lo_lo_lo_hi_25 = {res_lo_lo_lo_hi_hi_25, res_lo_lo_lo_hi_lo_25};
  wire [63:0]   res_lo_lo_lo_25 = {res_lo_lo_lo_hi_25, res_lo_lo_lo_lo_25};
  wire [15:0]   res_lo_lo_hi_lo_lo_25 = {dataGroup_9_25, dataGroup_8_25};
  wire [15:0]   res_lo_lo_hi_lo_hi_25 = {dataGroup_11_25, dataGroup_10_25};
  wire [31:0]   res_lo_lo_hi_lo_25 = {res_lo_lo_hi_lo_hi_25, res_lo_lo_hi_lo_lo_25};
  wire [15:0]   res_lo_lo_hi_hi_lo_25 = {dataGroup_13_25, dataGroup_12_25};
  wire [15:0]   res_lo_lo_hi_hi_hi_25 = {dataGroup_15_25, dataGroup_14_25};
  wire [31:0]   res_lo_lo_hi_hi_25 = {res_lo_lo_hi_hi_hi_25, res_lo_lo_hi_hi_lo_25};
  wire [63:0]   res_lo_lo_hi_25 = {res_lo_lo_hi_hi_25, res_lo_lo_hi_lo_25};
  wire [127:0]  res_lo_lo_25 = {res_lo_lo_hi_25, res_lo_lo_lo_25};
  wire [15:0]   res_lo_hi_lo_lo_lo_25 = {dataGroup_17_25, dataGroup_16_25};
  wire [15:0]   res_lo_hi_lo_lo_hi_25 = {dataGroup_19_25, dataGroup_18_25};
  wire [31:0]   res_lo_hi_lo_lo_25 = {res_lo_hi_lo_lo_hi_25, res_lo_hi_lo_lo_lo_25};
  wire [15:0]   res_lo_hi_lo_hi_lo_25 = {dataGroup_21_25, dataGroup_20_25};
  wire [15:0]   res_lo_hi_lo_hi_hi_25 = {dataGroup_23_25, dataGroup_22_25};
  wire [31:0]   res_lo_hi_lo_hi_25 = {res_lo_hi_lo_hi_hi_25, res_lo_hi_lo_hi_lo_25};
  wire [63:0]   res_lo_hi_lo_25 = {res_lo_hi_lo_hi_25, res_lo_hi_lo_lo_25};
  wire [15:0]   res_lo_hi_hi_lo_lo_25 = {dataGroup_25_25, dataGroup_24_25};
  wire [15:0]   res_lo_hi_hi_lo_hi_25 = {dataGroup_27_25, dataGroup_26_25};
  wire [31:0]   res_lo_hi_hi_lo_25 = {res_lo_hi_hi_lo_hi_25, res_lo_hi_hi_lo_lo_25};
  wire [15:0]   res_lo_hi_hi_hi_lo_25 = {dataGroup_29_25, dataGroup_28_25};
  wire [15:0]   res_lo_hi_hi_hi_hi_25 = {dataGroup_31_25, dataGroup_30_25};
  wire [31:0]   res_lo_hi_hi_hi_25 = {res_lo_hi_hi_hi_hi_25, res_lo_hi_hi_hi_lo_25};
  wire [63:0]   res_lo_hi_hi_25 = {res_lo_hi_hi_hi_25, res_lo_hi_hi_lo_25};
  wire [127:0]  res_lo_hi_25 = {res_lo_hi_hi_25, res_lo_hi_lo_25};
  wire [255:0]  res_lo_25 = {res_lo_hi_25, res_lo_lo_25};
  wire [15:0]   res_hi_lo_lo_lo_lo_25 = {dataGroup_33_25, dataGroup_32_25};
  wire [15:0]   res_hi_lo_lo_lo_hi_25 = {dataGroup_35_25, dataGroup_34_25};
  wire [31:0]   res_hi_lo_lo_lo_25 = {res_hi_lo_lo_lo_hi_25, res_hi_lo_lo_lo_lo_25};
  wire [15:0]   res_hi_lo_lo_hi_lo_25 = {dataGroup_37_25, dataGroup_36_25};
  wire [15:0]   res_hi_lo_lo_hi_hi_25 = {dataGroup_39_25, dataGroup_38_25};
  wire [31:0]   res_hi_lo_lo_hi_25 = {res_hi_lo_lo_hi_hi_25, res_hi_lo_lo_hi_lo_25};
  wire [63:0]   res_hi_lo_lo_25 = {res_hi_lo_lo_hi_25, res_hi_lo_lo_lo_25};
  wire [15:0]   res_hi_lo_hi_lo_lo_25 = {dataGroup_41_25, dataGroup_40_25};
  wire [15:0]   res_hi_lo_hi_lo_hi_25 = {dataGroup_43_25, dataGroup_42_25};
  wire [31:0]   res_hi_lo_hi_lo_25 = {res_hi_lo_hi_lo_hi_25, res_hi_lo_hi_lo_lo_25};
  wire [15:0]   res_hi_lo_hi_hi_lo_25 = {dataGroup_45_25, dataGroup_44_25};
  wire [15:0]   res_hi_lo_hi_hi_hi_25 = {dataGroup_47_25, dataGroup_46_25};
  wire [31:0]   res_hi_lo_hi_hi_25 = {res_hi_lo_hi_hi_hi_25, res_hi_lo_hi_hi_lo_25};
  wire [63:0]   res_hi_lo_hi_25 = {res_hi_lo_hi_hi_25, res_hi_lo_hi_lo_25};
  wire [127:0]  res_hi_lo_25 = {res_hi_lo_hi_25, res_hi_lo_lo_25};
  wire [15:0]   res_hi_hi_lo_lo_lo_25 = {dataGroup_49_25, dataGroup_48_25};
  wire [15:0]   res_hi_hi_lo_lo_hi_25 = {dataGroup_51_25, dataGroup_50_25};
  wire [31:0]   res_hi_hi_lo_lo_25 = {res_hi_hi_lo_lo_hi_25, res_hi_hi_lo_lo_lo_25};
  wire [15:0]   res_hi_hi_lo_hi_lo_25 = {dataGroup_53_25, dataGroup_52_25};
  wire [15:0]   res_hi_hi_lo_hi_hi_25 = {dataGroup_55_25, dataGroup_54_25};
  wire [31:0]   res_hi_hi_lo_hi_25 = {res_hi_hi_lo_hi_hi_25, res_hi_hi_lo_hi_lo_25};
  wire [63:0]   res_hi_hi_lo_25 = {res_hi_hi_lo_hi_25, res_hi_hi_lo_lo_25};
  wire [15:0]   res_hi_hi_hi_lo_lo_25 = {dataGroup_57_25, dataGroup_56_25};
  wire [15:0]   res_hi_hi_hi_lo_hi_25 = {dataGroup_59_25, dataGroup_58_25};
  wire [31:0]   res_hi_hi_hi_lo_25 = {res_hi_hi_hi_lo_hi_25, res_hi_hi_hi_lo_lo_25};
  wire [15:0]   res_hi_hi_hi_hi_lo_25 = {dataGroup_61_25, dataGroup_60_25};
  wire [15:0]   res_hi_hi_hi_hi_hi_25 = {dataGroup_63_25, dataGroup_62_25};
  wire [31:0]   res_hi_hi_hi_hi_25 = {res_hi_hi_hi_hi_hi_25, res_hi_hi_hi_hi_lo_25};
  wire [63:0]   res_hi_hi_hi_25 = {res_hi_hi_hi_hi_25, res_hi_hi_hi_lo_25};
  wire [127:0]  res_hi_hi_25 = {res_hi_hi_hi_25, res_hi_hi_lo_25};
  wire [255:0]  res_hi_25 = {res_hi_hi_25, res_hi_lo_25};
  wire [511:0]  res_52 = {res_hi_25, res_lo_25};
  wire [2047:0] dataGroup_lo_1664 = {dataGroup_lo_hi_1664, dataGroup_lo_lo_1664};
  wire [2047:0] dataGroup_hi_1664 = {dataGroup_hi_hi_1664, dataGroup_hi_lo_1664};
  wire [7:0]    dataGroup_0_26 = dataGroup_lo_1664[47:40];
  wire [2047:0] dataGroup_lo_1665 = {dataGroup_lo_hi_1665, dataGroup_lo_lo_1665};
  wire [2047:0] dataGroup_hi_1665 = {dataGroup_hi_hi_1665, dataGroup_hi_lo_1665};
  wire [7:0]    dataGroup_1_26 = dataGroup_lo_1665[103:96];
  wire [2047:0] dataGroup_lo_1666 = {dataGroup_lo_hi_1666, dataGroup_lo_lo_1666};
  wire [2047:0] dataGroup_hi_1666 = {dataGroup_hi_hi_1666, dataGroup_hi_lo_1666};
  wire [7:0]    dataGroup_2_26 = dataGroup_lo_1666[159:152];
  wire [2047:0] dataGroup_lo_1667 = {dataGroup_lo_hi_1667, dataGroup_lo_lo_1667};
  wire [2047:0] dataGroup_hi_1667 = {dataGroup_hi_hi_1667, dataGroup_hi_lo_1667};
  wire [7:0]    dataGroup_3_26 = dataGroup_lo_1667[215:208];
  wire [2047:0] dataGroup_lo_1668 = {dataGroup_lo_hi_1668, dataGroup_lo_lo_1668};
  wire [2047:0] dataGroup_hi_1668 = {dataGroup_hi_hi_1668, dataGroup_hi_lo_1668};
  wire [7:0]    dataGroup_4_26 = dataGroup_lo_1668[271:264];
  wire [2047:0] dataGroup_lo_1669 = {dataGroup_lo_hi_1669, dataGroup_lo_lo_1669};
  wire [2047:0] dataGroup_hi_1669 = {dataGroup_hi_hi_1669, dataGroup_hi_lo_1669};
  wire [7:0]    dataGroup_5_26 = dataGroup_lo_1669[327:320];
  wire [2047:0] dataGroup_lo_1670 = {dataGroup_lo_hi_1670, dataGroup_lo_lo_1670};
  wire [2047:0] dataGroup_hi_1670 = {dataGroup_hi_hi_1670, dataGroup_hi_lo_1670};
  wire [7:0]    dataGroup_6_26 = dataGroup_lo_1670[383:376];
  wire [2047:0] dataGroup_lo_1671 = {dataGroup_lo_hi_1671, dataGroup_lo_lo_1671};
  wire [2047:0] dataGroup_hi_1671 = {dataGroup_hi_hi_1671, dataGroup_hi_lo_1671};
  wire [7:0]    dataGroup_7_26 = dataGroup_lo_1671[439:432];
  wire [2047:0] dataGroup_lo_1672 = {dataGroup_lo_hi_1672, dataGroup_lo_lo_1672};
  wire [2047:0] dataGroup_hi_1672 = {dataGroup_hi_hi_1672, dataGroup_hi_lo_1672};
  wire [7:0]    dataGroup_8_26 = dataGroup_lo_1672[495:488];
  wire [2047:0] dataGroup_lo_1673 = {dataGroup_lo_hi_1673, dataGroup_lo_lo_1673};
  wire [2047:0] dataGroup_hi_1673 = {dataGroup_hi_hi_1673, dataGroup_hi_lo_1673};
  wire [7:0]    dataGroup_9_26 = dataGroup_lo_1673[551:544];
  wire [2047:0] dataGroup_lo_1674 = {dataGroup_lo_hi_1674, dataGroup_lo_lo_1674};
  wire [2047:0] dataGroup_hi_1674 = {dataGroup_hi_hi_1674, dataGroup_hi_lo_1674};
  wire [7:0]    dataGroup_10_26 = dataGroup_lo_1674[607:600];
  wire [2047:0] dataGroup_lo_1675 = {dataGroup_lo_hi_1675, dataGroup_lo_lo_1675};
  wire [2047:0] dataGroup_hi_1675 = {dataGroup_hi_hi_1675, dataGroup_hi_lo_1675};
  wire [7:0]    dataGroup_11_26 = dataGroup_lo_1675[663:656];
  wire [2047:0] dataGroup_lo_1676 = {dataGroup_lo_hi_1676, dataGroup_lo_lo_1676};
  wire [2047:0] dataGroup_hi_1676 = {dataGroup_hi_hi_1676, dataGroup_hi_lo_1676};
  wire [7:0]    dataGroup_12_26 = dataGroup_lo_1676[719:712];
  wire [2047:0] dataGroup_lo_1677 = {dataGroup_lo_hi_1677, dataGroup_lo_lo_1677};
  wire [2047:0] dataGroup_hi_1677 = {dataGroup_hi_hi_1677, dataGroup_hi_lo_1677};
  wire [7:0]    dataGroup_13_26 = dataGroup_lo_1677[775:768];
  wire [2047:0] dataGroup_lo_1678 = {dataGroup_lo_hi_1678, dataGroup_lo_lo_1678};
  wire [2047:0] dataGroup_hi_1678 = {dataGroup_hi_hi_1678, dataGroup_hi_lo_1678};
  wire [7:0]    dataGroup_14_26 = dataGroup_lo_1678[831:824];
  wire [2047:0] dataGroup_lo_1679 = {dataGroup_lo_hi_1679, dataGroup_lo_lo_1679};
  wire [2047:0] dataGroup_hi_1679 = {dataGroup_hi_hi_1679, dataGroup_hi_lo_1679};
  wire [7:0]    dataGroup_15_26 = dataGroup_lo_1679[887:880];
  wire [2047:0] dataGroup_lo_1680 = {dataGroup_lo_hi_1680, dataGroup_lo_lo_1680};
  wire [2047:0] dataGroup_hi_1680 = {dataGroup_hi_hi_1680, dataGroup_hi_lo_1680};
  wire [7:0]    dataGroup_16_26 = dataGroup_lo_1680[943:936];
  wire [2047:0] dataGroup_lo_1681 = {dataGroup_lo_hi_1681, dataGroup_lo_lo_1681};
  wire [2047:0] dataGroup_hi_1681 = {dataGroup_hi_hi_1681, dataGroup_hi_lo_1681};
  wire [7:0]    dataGroup_17_26 = dataGroup_lo_1681[999:992];
  wire [2047:0] dataGroup_lo_1682 = {dataGroup_lo_hi_1682, dataGroup_lo_lo_1682};
  wire [2047:0] dataGroup_hi_1682 = {dataGroup_hi_hi_1682, dataGroup_hi_lo_1682};
  wire [7:0]    dataGroup_18_26 = dataGroup_lo_1682[1055:1048];
  wire [2047:0] dataGroup_lo_1683 = {dataGroup_lo_hi_1683, dataGroup_lo_lo_1683};
  wire [2047:0] dataGroup_hi_1683 = {dataGroup_hi_hi_1683, dataGroup_hi_lo_1683};
  wire [7:0]    dataGroup_19_26 = dataGroup_lo_1683[1111:1104];
  wire [2047:0] dataGroup_lo_1684 = {dataGroup_lo_hi_1684, dataGroup_lo_lo_1684};
  wire [2047:0] dataGroup_hi_1684 = {dataGroup_hi_hi_1684, dataGroup_hi_lo_1684};
  wire [7:0]    dataGroup_20_26 = dataGroup_lo_1684[1167:1160];
  wire [2047:0] dataGroup_lo_1685 = {dataGroup_lo_hi_1685, dataGroup_lo_lo_1685};
  wire [2047:0] dataGroup_hi_1685 = {dataGroup_hi_hi_1685, dataGroup_hi_lo_1685};
  wire [7:0]    dataGroup_21_26 = dataGroup_lo_1685[1223:1216];
  wire [2047:0] dataGroup_lo_1686 = {dataGroup_lo_hi_1686, dataGroup_lo_lo_1686};
  wire [2047:0] dataGroup_hi_1686 = {dataGroup_hi_hi_1686, dataGroup_hi_lo_1686};
  wire [7:0]    dataGroup_22_26 = dataGroup_lo_1686[1279:1272];
  wire [2047:0] dataGroup_lo_1687 = {dataGroup_lo_hi_1687, dataGroup_lo_lo_1687};
  wire [2047:0] dataGroup_hi_1687 = {dataGroup_hi_hi_1687, dataGroup_hi_lo_1687};
  wire [7:0]    dataGroup_23_26 = dataGroup_lo_1687[1335:1328];
  wire [2047:0] dataGroup_lo_1688 = {dataGroup_lo_hi_1688, dataGroup_lo_lo_1688};
  wire [2047:0] dataGroup_hi_1688 = {dataGroup_hi_hi_1688, dataGroup_hi_lo_1688};
  wire [7:0]    dataGroup_24_26 = dataGroup_lo_1688[1391:1384];
  wire [2047:0] dataGroup_lo_1689 = {dataGroup_lo_hi_1689, dataGroup_lo_lo_1689};
  wire [2047:0] dataGroup_hi_1689 = {dataGroup_hi_hi_1689, dataGroup_hi_lo_1689};
  wire [7:0]    dataGroup_25_26 = dataGroup_lo_1689[1447:1440];
  wire [2047:0] dataGroup_lo_1690 = {dataGroup_lo_hi_1690, dataGroup_lo_lo_1690};
  wire [2047:0] dataGroup_hi_1690 = {dataGroup_hi_hi_1690, dataGroup_hi_lo_1690};
  wire [7:0]    dataGroup_26_26 = dataGroup_lo_1690[1503:1496];
  wire [2047:0] dataGroup_lo_1691 = {dataGroup_lo_hi_1691, dataGroup_lo_lo_1691};
  wire [2047:0] dataGroup_hi_1691 = {dataGroup_hi_hi_1691, dataGroup_hi_lo_1691};
  wire [7:0]    dataGroup_27_26 = dataGroup_lo_1691[1559:1552];
  wire [2047:0] dataGroup_lo_1692 = {dataGroup_lo_hi_1692, dataGroup_lo_lo_1692};
  wire [2047:0] dataGroup_hi_1692 = {dataGroup_hi_hi_1692, dataGroup_hi_lo_1692};
  wire [7:0]    dataGroup_28_26 = dataGroup_lo_1692[1615:1608];
  wire [2047:0] dataGroup_lo_1693 = {dataGroup_lo_hi_1693, dataGroup_lo_lo_1693};
  wire [2047:0] dataGroup_hi_1693 = {dataGroup_hi_hi_1693, dataGroup_hi_lo_1693};
  wire [7:0]    dataGroup_29_26 = dataGroup_lo_1693[1671:1664];
  wire [2047:0] dataGroup_lo_1694 = {dataGroup_lo_hi_1694, dataGroup_lo_lo_1694};
  wire [2047:0] dataGroup_hi_1694 = {dataGroup_hi_hi_1694, dataGroup_hi_lo_1694};
  wire [7:0]    dataGroup_30_26 = dataGroup_lo_1694[1727:1720];
  wire [2047:0] dataGroup_lo_1695 = {dataGroup_lo_hi_1695, dataGroup_lo_lo_1695};
  wire [2047:0] dataGroup_hi_1695 = {dataGroup_hi_hi_1695, dataGroup_hi_lo_1695};
  wire [7:0]    dataGroup_31_26 = dataGroup_lo_1695[1783:1776];
  wire [2047:0] dataGroup_lo_1696 = {dataGroup_lo_hi_1696, dataGroup_lo_lo_1696};
  wire [2047:0] dataGroup_hi_1696 = {dataGroup_hi_hi_1696, dataGroup_hi_lo_1696};
  wire [7:0]    dataGroup_32_26 = dataGroup_lo_1696[1839:1832];
  wire [2047:0] dataGroup_lo_1697 = {dataGroup_lo_hi_1697, dataGroup_lo_lo_1697};
  wire [2047:0] dataGroup_hi_1697 = {dataGroup_hi_hi_1697, dataGroup_hi_lo_1697};
  wire [7:0]    dataGroup_33_26 = dataGroup_lo_1697[1895:1888];
  wire [2047:0] dataGroup_lo_1698 = {dataGroup_lo_hi_1698, dataGroup_lo_lo_1698};
  wire [2047:0] dataGroup_hi_1698 = {dataGroup_hi_hi_1698, dataGroup_hi_lo_1698};
  wire [7:0]    dataGroup_34_26 = dataGroup_lo_1698[1951:1944];
  wire [2047:0] dataGroup_lo_1699 = {dataGroup_lo_hi_1699, dataGroup_lo_lo_1699};
  wire [2047:0] dataGroup_hi_1699 = {dataGroup_hi_hi_1699, dataGroup_hi_lo_1699};
  wire [7:0]    dataGroup_35_26 = dataGroup_lo_1699[2007:2000];
  wire [2047:0] dataGroup_lo_1700 = {dataGroup_lo_hi_1700, dataGroup_lo_lo_1700};
  wire [2047:0] dataGroup_hi_1700 = {dataGroup_hi_hi_1700, dataGroup_hi_lo_1700};
  wire [7:0]    dataGroup_36_26 = dataGroup_hi_1700[15:8];
  wire [2047:0] dataGroup_lo_1701 = {dataGroup_lo_hi_1701, dataGroup_lo_lo_1701};
  wire [2047:0] dataGroup_hi_1701 = {dataGroup_hi_hi_1701, dataGroup_hi_lo_1701};
  wire [7:0]    dataGroup_37_26 = dataGroup_hi_1701[71:64];
  wire [2047:0] dataGroup_lo_1702 = {dataGroup_lo_hi_1702, dataGroup_lo_lo_1702};
  wire [2047:0] dataGroup_hi_1702 = {dataGroup_hi_hi_1702, dataGroup_hi_lo_1702};
  wire [7:0]    dataGroup_38_26 = dataGroup_hi_1702[127:120];
  wire [2047:0] dataGroup_lo_1703 = {dataGroup_lo_hi_1703, dataGroup_lo_lo_1703};
  wire [2047:0] dataGroup_hi_1703 = {dataGroup_hi_hi_1703, dataGroup_hi_lo_1703};
  wire [7:0]    dataGroup_39_26 = dataGroup_hi_1703[183:176];
  wire [2047:0] dataGroup_lo_1704 = {dataGroup_lo_hi_1704, dataGroup_lo_lo_1704};
  wire [2047:0] dataGroup_hi_1704 = {dataGroup_hi_hi_1704, dataGroup_hi_lo_1704};
  wire [7:0]    dataGroup_40_26 = dataGroup_hi_1704[239:232];
  wire [2047:0] dataGroup_lo_1705 = {dataGroup_lo_hi_1705, dataGroup_lo_lo_1705};
  wire [2047:0] dataGroup_hi_1705 = {dataGroup_hi_hi_1705, dataGroup_hi_lo_1705};
  wire [7:0]    dataGroup_41_26 = dataGroup_hi_1705[295:288];
  wire [2047:0] dataGroup_lo_1706 = {dataGroup_lo_hi_1706, dataGroup_lo_lo_1706};
  wire [2047:0] dataGroup_hi_1706 = {dataGroup_hi_hi_1706, dataGroup_hi_lo_1706};
  wire [7:0]    dataGroup_42_26 = dataGroup_hi_1706[351:344];
  wire [2047:0] dataGroup_lo_1707 = {dataGroup_lo_hi_1707, dataGroup_lo_lo_1707};
  wire [2047:0] dataGroup_hi_1707 = {dataGroup_hi_hi_1707, dataGroup_hi_lo_1707};
  wire [7:0]    dataGroup_43_26 = dataGroup_hi_1707[407:400];
  wire [2047:0] dataGroup_lo_1708 = {dataGroup_lo_hi_1708, dataGroup_lo_lo_1708};
  wire [2047:0] dataGroup_hi_1708 = {dataGroup_hi_hi_1708, dataGroup_hi_lo_1708};
  wire [7:0]    dataGroup_44_26 = dataGroup_hi_1708[463:456];
  wire [2047:0] dataGroup_lo_1709 = {dataGroup_lo_hi_1709, dataGroup_lo_lo_1709};
  wire [2047:0] dataGroup_hi_1709 = {dataGroup_hi_hi_1709, dataGroup_hi_lo_1709};
  wire [7:0]    dataGroup_45_26 = dataGroup_hi_1709[519:512];
  wire [2047:0] dataGroup_lo_1710 = {dataGroup_lo_hi_1710, dataGroup_lo_lo_1710};
  wire [2047:0] dataGroup_hi_1710 = {dataGroup_hi_hi_1710, dataGroup_hi_lo_1710};
  wire [7:0]    dataGroup_46_26 = dataGroup_hi_1710[575:568];
  wire [2047:0] dataGroup_lo_1711 = {dataGroup_lo_hi_1711, dataGroup_lo_lo_1711};
  wire [2047:0] dataGroup_hi_1711 = {dataGroup_hi_hi_1711, dataGroup_hi_lo_1711};
  wire [7:0]    dataGroup_47_26 = dataGroup_hi_1711[631:624];
  wire [2047:0] dataGroup_lo_1712 = {dataGroup_lo_hi_1712, dataGroup_lo_lo_1712};
  wire [2047:0] dataGroup_hi_1712 = {dataGroup_hi_hi_1712, dataGroup_hi_lo_1712};
  wire [7:0]    dataGroup_48_26 = dataGroup_hi_1712[687:680];
  wire [2047:0] dataGroup_lo_1713 = {dataGroup_lo_hi_1713, dataGroup_lo_lo_1713};
  wire [2047:0] dataGroup_hi_1713 = {dataGroup_hi_hi_1713, dataGroup_hi_lo_1713};
  wire [7:0]    dataGroup_49_26 = dataGroup_hi_1713[743:736];
  wire [2047:0] dataGroup_lo_1714 = {dataGroup_lo_hi_1714, dataGroup_lo_lo_1714};
  wire [2047:0] dataGroup_hi_1714 = {dataGroup_hi_hi_1714, dataGroup_hi_lo_1714};
  wire [7:0]    dataGroup_50_26 = dataGroup_hi_1714[799:792];
  wire [2047:0] dataGroup_lo_1715 = {dataGroup_lo_hi_1715, dataGroup_lo_lo_1715};
  wire [2047:0] dataGroup_hi_1715 = {dataGroup_hi_hi_1715, dataGroup_hi_lo_1715};
  wire [7:0]    dataGroup_51_26 = dataGroup_hi_1715[855:848];
  wire [2047:0] dataGroup_lo_1716 = {dataGroup_lo_hi_1716, dataGroup_lo_lo_1716};
  wire [2047:0] dataGroup_hi_1716 = {dataGroup_hi_hi_1716, dataGroup_hi_lo_1716};
  wire [7:0]    dataGroup_52_26 = dataGroup_hi_1716[911:904];
  wire [2047:0] dataGroup_lo_1717 = {dataGroup_lo_hi_1717, dataGroup_lo_lo_1717};
  wire [2047:0] dataGroup_hi_1717 = {dataGroup_hi_hi_1717, dataGroup_hi_lo_1717};
  wire [7:0]    dataGroup_53_26 = dataGroup_hi_1717[967:960];
  wire [2047:0] dataGroup_lo_1718 = {dataGroup_lo_hi_1718, dataGroup_lo_lo_1718};
  wire [2047:0] dataGroup_hi_1718 = {dataGroup_hi_hi_1718, dataGroup_hi_lo_1718};
  wire [7:0]    dataGroup_54_26 = dataGroup_hi_1718[1023:1016];
  wire [2047:0] dataGroup_lo_1719 = {dataGroup_lo_hi_1719, dataGroup_lo_lo_1719};
  wire [2047:0] dataGroup_hi_1719 = {dataGroup_hi_hi_1719, dataGroup_hi_lo_1719};
  wire [7:0]    dataGroup_55_26 = dataGroup_hi_1719[1079:1072];
  wire [2047:0] dataGroup_lo_1720 = {dataGroup_lo_hi_1720, dataGroup_lo_lo_1720};
  wire [2047:0] dataGroup_hi_1720 = {dataGroup_hi_hi_1720, dataGroup_hi_lo_1720};
  wire [7:0]    dataGroup_56_26 = dataGroup_hi_1720[1135:1128];
  wire [2047:0] dataGroup_lo_1721 = {dataGroup_lo_hi_1721, dataGroup_lo_lo_1721};
  wire [2047:0] dataGroup_hi_1721 = {dataGroup_hi_hi_1721, dataGroup_hi_lo_1721};
  wire [7:0]    dataGroup_57_26 = dataGroup_hi_1721[1191:1184];
  wire [2047:0] dataGroup_lo_1722 = {dataGroup_lo_hi_1722, dataGroup_lo_lo_1722};
  wire [2047:0] dataGroup_hi_1722 = {dataGroup_hi_hi_1722, dataGroup_hi_lo_1722};
  wire [7:0]    dataGroup_58_26 = dataGroup_hi_1722[1247:1240];
  wire [2047:0] dataGroup_lo_1723 = {dataGroup_lo_hi_1723, dataGroup_lo_lo_1723};
  wire [2047:0] dataGroup_hi_1723 = {dataGroup_hi_hi_1723, dataGroup_hi_lo_1723};
  wire [7:0]    dataGroup_59_26 = dataGroup_hi_1723[1303:1296];
  wire [2047:0] dataGroup_lo_1724 = {dataGroup_lo_hi_1724, dataGroup_lo_lo_1724};
  wire [2047:0] dataGroup_hi_1724 = {dataGroup_hi_hi_1724, dataGroup_hi_lo_1724};
  wire [7:0]    dataGroup_60_26 = dataGroup_hi_1724[1359:1352];
  wire [2047:0] dataGroup_lo_1725 = {dataGroup_lo_hi_1725, dataGroup_lo_lo_1725};
  wire [2047:0] dataGroup_hi_1725 = {dataGroup_hi_hi_1725, dataGroup_hi_lo_1725};
  wire [7:0]    dataGroup_61_26 = dataGroup_hi_1725[1415:1408];
  wire [2047:0] dataGroup_lo_1726 = {dataGroup_lo_hi_1726, dataGroup_lo_lo_1726};
  wire [2047:0] dataGroup_hi_1726 = {dataGroup_hi_hi_1726, dataGroup_hi_lo_1726};
  wire [7:0]    dataGroup_62_26 = dataGroup_hi_1726[1471:1464];
  wire [2047:0] dataGroup_lo_1727 = {dataGroup_lo_hi_1727, dataGroup_lo_lo_1727};
  wire [2047:0] dataGroup_hi_1727 = {dataGroup_hi_hi_1727, dataGroup_hi_lo_1727};
  wire [7:0]    dataGroup_63_26 = dataGroup_hi_1727[1527:1520];
  wire [15:0]   res_lo_lo_lo_lo_lo_26 = {dataGroup_1_26, dataGroup_0_26};
  wire [15:0]   res_lo_lo_lo_lo_hi_26 = {dataGroup_3_26, dataGroup_2_26};
  wire [31:0]   res_lo_lo_lo_lo_26 = {res_lo_lo_lo_lo_hi_26, res_lo_lo_lo_lo_lo_26};
  wire [15:0]   res_lo_lo_lo_hi_lo_26 = {dataGroup_5_26, dataGroup_4_26};
  wire [15:0]   res_lo_lo_lo_hi_hi_26 = {dataGroup_7_26, dataGroup_6_26};
  wire [31:0]   res_lo_lo_lo_hi_26 = {res_lo_lo_lo_hi_hi_26, res_lo_lo_lo_hi_lo_26};
  wire [63:0]   res_lo_lo_lo_26 = {res_lo_lo_lo_hi_26, res_lo_lo_lo_lo_26};
  wire [15:0]   res_lo_lo_hi_lo_lo_26 = {dataGroup_9_26, dataGroup_8_26};
  wire [15:0]   res_lo_lo_hi_lo_hi_26 = {dataGroup_11_26, dataGroup_10_26};
  wire [31:0]   res_lo_lo_hi_lo_26 = {res_lo_lo_hi_lo_hi_26, res_lo_lo_hi_lo_lo_26};
  wire [15:0]   res_lo_lo_hi_hi_lo_26 = {dataGroup_13_26, dataGroup_12_26};
  wire [15:0]   res_lo_lo_hi_hi_hi_26 = {dataGroup_15_26, dataGroup_14_26};
  wire [31:0]   res_lo_lo_hi_hi_26 = {res_lo_lo_hi_hi_hi_26, res_lo_lo_hi_hi_lo_26};
  wire [63:0]   res_lo_lo_hi_26 = {res_lo_lo_hi_hi_26, res_lo_lo_hi_lo_26};
  wire [127:0]  res_lo_lo_26 = {res_lo_lo_hi_26, res_lo_lo_lo_26};
  wire [15:0]   res_lo_hi_lo_lo_lo_26 = {dataGroup_17_26, dataGroup_16_26};
  wire [15:0]   res_lo_hi_lo_lo_hi_26 = {dataGroup_19_26, dataGroup_18_26};
  wire [31:0]   res_lo_hi_lo_lo_26 = {res_lo_hi_lo_lo_hi_26, res_lo_hi_lo_lo_lo_26};
  wire [15:0]   res_lo_hi_lo_hi_lo_26 = {dataGroup_21_26, dataGroup_20_26};
  wire [15:0]   res_lo_hi_lo_hi_hi_26 = {dataGroup_23_26, dataGroup_22_26};
  wire [31:0]   res_lo_hi_lo_hi_26 = {res_lo_hi_lo_hi_hi_26, res_lo_hi_lo_hi_lo_26};
  wire [63:0]   res_lo_hi_lo_26 = {res_lo_hi_lo_hi_26, res_lo_hi_lo_lo_26};
  wire [15:0]   res_lo_hi_hi_lo_lo_26 = {dataGroup_25_26, dataGroup_24_26};
  wire [15:0]   res_lo_hi_hi_lo_hi_26 = {dataGroup_27_26, dataGroup_26_26};
  wire [31:0]   res_lo_hi_hi_lo_26 = {res_lo_hi_hi_lo_hi_26, res_lo_hi_hi_lo_lo_26};
  wire [15:0]   res_lo_hi_hi_hi_lo_26 = {dataGroup_29_26, dataGroup_28_26};
  wire [15:0]   res_lo_hi_hi_hi_hi_26 = {dataGroup_31_26, dataGroup_30_26};
  wire [31:0]   res_lo_hi_hi_hi_26 = {res_lo_hi_hi_hi_hi_26, res_lo_hi_hi_hi_lo_26};
  wire [63:0]   res_lo_hi_hi_26 = {res_lo_hi_hi_hi_26, res_lo_hi_hi_lo_26};
  wire [127:0]  res_lo_hi_26 = {res_lo_hi_hi_26, res_lo_hi_lo_26};
  wire [255:0]  res_lo_26 = {res_lo_hi_26, res_lo_lo_26};
  wire [15:0]   res_hi_lo_lo_lo_lo_26 = {dataGroup_33_26, dataGroup_32_26};
  wire [15:0]   res_hi_lo_lo_lo_hi_26 = {dataGroup_35_26, dataGroup_34_26};
  wire [31:0]   res_hi_lo_lo_lo_26 = {res_hi_lo_lo_lo_hi_26, res_hi_lo_lo_lo_lo_26};
  wire [15:0]   res_hi_lo_lo_hi_lo_26 = {dataGroup_37_26, dataGroup_36_26};
  wire [15:0]   res_hi_lo_lo_hi_hi_26 = {dataGroup_39_26, dataGroup_38_26};
  wire [31:0]   res_hi_lo_lo_hi_26 = {res_hi_lo_lo_hi_hi_26, res_hi_lo_lo_hi_lo_26};
  wire [63:0]   res_hi_lo_lo_26 = {res_hi_lo_lo_hi_26, res_hi_lo_lo_lo_26};
  wire [15:0]   res_hi_lo_hi_lo_lo_26 = {dataGroup_41_26, dataGroup_40_26};
  wire [15:0]   res_hi_lo_hi_lo_hi_26 = {dataGroup_43_26, dataGroup_42_26};
  wire [31:0]   res_hi_lo_hi_lo_26 = {res_hi_lo_hi_lo_hi_26, res_hi_lo_hi_lo_lo_26};
  wire [15:0]   res_hi_lo_hi_hi_lo_26 = {dataGroup_45_26, dataGroup_44_26};
  wire [15:0]   res_hi_lo_hi_hi_hi_26 = {dataGroup_47_26, dataGroup_46_26};
  wire [31:0]   res_hi_lo_hi_hi_26 = {res_hi_lo_hi_hi_hi_26, res_hi_lo_hi_hi_lo_26};
  wire [63:0]   res_hi_lo_hi_26 = {res_hi_lo_hi_hi_26, res_hi_lo_hi_lo_26};
  wire [127:0]  res_hi_lo_26 = {res_hi_lo_hi_26, res_hi_lo_lo_26};
  wire [15:0]   res_hi_hi_lo_lo_lo_26 = {dataGroup_49_26, dataGroup_48_26};
  wire [15:0]   res_hi_hi_lo_lo_hi_26 = {dataGroup_51_26, dataGroup_50_26};
  wire [31:0]   res_hi_hi_lo_lo_26 = {res_hi_hi_lo_lo_hi_26, res_hi_hi_lo_lo_lo_26};
  wire [15:0]   res_hi_hi_lo_hi_lo_26 = {dataGroup_53_26, dataGroup_52_26};
  wire [15:0]   res_hi_hi_lo_hi_hi_26 = {dataGroup_55_26, dataGroup_54_26};
  wire [31:0]   res_hi_hi_lo_hi_26 = {res_hi_hi_lo_hi_hi_26, res_hi_hi_lo_hi_lo_26};
  wire [63:0]   res_hi_hi_lo_26 = {res_hi_hi_lo_hi_26, res_hi_hi_lo_lo_26};
  wire [15:0]   res_hi_hi_hi_lo_lo_26 = {dataGroup_57_26, dataGroup_56_26};
  wire [15:0]   res_hi_hi_hi_lo_hi_26 = {dataGroup_59_26, dataGroup_58_26};
  wire [31:0]   res_hi_hi_hi_lo_26 = {res_hi_hi_hi_lo_hi_26, res_hi_hi_hi_lo_lo_26};
  wire [15:0]   res_hi_hi_hi_hi_lo_26 = {dataGroup_61_26, dataGroup_60_26};
  wire [15:0]   res_hi_hi_hi_hi_hi_26 = {dataGroup_63_26, dataGroup_62_26};
  wire [31:0]   res_hi_hi_hi_hi_26 = {res_hi_hi_hi_hi_hi_26, res_hi_hi_hi_hi_lo_26};
  wire [63:0]   res_hi_hi_hi_26 = {res_hi_hi_hi_hi_26, res_hi_hi_hi_lo_26};
  wire [127:0]  res_hi_hi_26 = {res_hi_hi_hi_26, res_hi_hi_lo_26};
  wire [255:0]  res_hi_26 = {res_hi_hi_26, res_hi_lo_26};
  wire [511:0]  res_53 = {res_hi_26, res_lo_26};
  wire [2047:0] dataGroup_lo_1728 = {dataGroup_lo_hi_1728, dataGroup_lo_lo_1728};
  wire [2047:0] dataGroup_hi_1728 = {dataGroup_hi_hi_1728, dataGroup_hi_lo_1728};
  wire [7:0]    dataGroup_0_27 = dataGroup_lo_1728[55:48];
  wire [2047:0] dataGroup_lo_1729 = {dataGroup_lo_hi_1729, dataGroup_lo_lo_1729};
  wire [2047:0] dataGroup_hi_1729 = {dataGroup_hi_hi_1729, dataGroup_hi_lo_1729};
  wire [7:0]    dataGroup_1_27 = dataGroup_lo_1729[111:104];
  wire [2047:0] dataGroup_lo_1730 = {dataGroup_lo_hi_1730, dataGroup_lo_lo_1730};
  wire [2047:0] dataGroup_hi_1730 = {dataGroup_hi_hi_1730, dataGroup_hi_lo_1730};
  wire [7:0]    dataGroup_2_27 = dataGroup_lo_1730[167:160];
  wire [2047:0] dataGroup_lo_1731 = {dataGroup_lo_hi_1731, dataGroup_lo_lo_1731};
  wire [2047:0] dataGroup_hi_1731 = {dataGroup_hi_hi_1731, dataGroup_hi_lo_1731};
  wire [7:0]    dataGroup_3_27 = dataGroup_lo_1731[223:216];
  wire [2047:0] dataGroup_lo_1732 = {dataGroup_lo_hi_1732, dataGroup_lo_lo_1732};
  wire [2047:0] dataGroup_hi_1732 = {dataGroup_hi_hi_1732, dataGroup_hi_lo_1732};
  wire [7:0]    dataGroup_4_27 = dataGroup_lo_1732[279:272];
  wire [2047:0] dataGroup_lo_1733 = {dataGroup_lo_hi_1733, dataGroup_lo_lo_1733};
  wire [2047:0] dataGroup_hi_1733 = {dataGroup_hi_hi_1733, dataGroup_hi_lo_1733};
  wire [7:0]    dataGroup_5_27 = dataGroup_lo_1733[335:328];
  wire [2047:0] dataGroup_lo_1734 = {dataGroup_lo_hi_1734, dataGroup_lo_lo_1734};
  wire [2047:0] dataGroup_hi_1734 = {dataGroup_hi_hi_1734, dataGroup_hi_lo_1734};
  wire [7:0]    dataGroup_6_27 = dataGroup_lo_1734[391:384];
  wire [2047:0] dataGroup_lo_1735 = {dataGroup_lo_hi_1735, dataGroup_lo_lo_1735};
  wire [2047:0] dataGroup_hi_1735 = {dataGroup_hi_hi_1735, dataGroup_hi_lo_1735};
  wire [7:0]    dataGroup_7_27 = dataGroup_lo_1735[447:440];
  wire [2047:0] dataGroup_lo_1736 = {dataGroup_lo_hi_1736, dataGroup_lo_lo_1736};
  wire [2047:0] dataGroup_hi_1736 = {dataGroup_hi_hi_1736, dataGroup_hi_lo_1736};
  wire [7:0]    dataGroup_8_27 = dataGroup_lo_1736[503:496];
  wire [2047:0] dataGroup_lo_1737 = {dataGroup_lo_hi_1737, dataGroup_lo_lo_1737};
  wire [2047:0] dataGroup_hi_1737 = {dataGroup_hi_hi_1737, dataGroup_hi_lo_1737};
  wire [7:0]    dataGroup_9_27 = dataGroup_lo_1737[559:552];
  wire [2047:0] dataGroup_lo_1738 = {dataGroup_lo_hi_1738, dataGroup_lo_lo_1738};
  wire [2047:0] dataGroup_hi_1738 = {dataGroup_hi_hi_1738, dataGroup_hi_lo_1738};
  wire [7:0]    dataGroup_10_27 = dataGroup_lo_1738[615:608];
  wire [2047:0] dataGroup_lo_1739 = {dataGroup_lo_hi_1739, dataGroup_lo_lo_1739};
  wire [2047:0] dataGroup_hi_1739 = {dataGroup_hi_hi_1739, dataGroup_hi_lo_1739};
  wire [7:0]    dataGroup_11_27 = dataGroup_lo_1739[671:664];
  wire [2047:0] dataGroup_lo_1740 = {dataGroup_lo_hi_1740, dataGroup_lo_lo_1740};
  wire [2047:0] dataGroup_hi_1740 = {dataGroup_hi_hi_1740, dataGroup_hi_lo_1740};
  wire [7:0]    dataGroup_12_27 = dataGroup_lo_1740[727:720];
  wire [2047:0] dataGroup_lo_1741 = {dataGroup_lo_hi_1741, dataGroup_lo_lo_1741};
  wire [2047:0] dataGroup_hi_1741 = {dataGroup_hi_hi_1741, dataGroup_hi_lo_1741};
  wire [7:0]    dataGroup_13_27 = dataGroup_lo_1741[783:776];
  wire [2047:0] dataGroup_lo_1742 = {dataGroup_lo_hi_1742, dataGroup_lo_lo_1742};
  wire [2047:0] dataGroup_hi_1742 = {dataGroup_hi_hi_1742, dataGroup_hi_lo_1742};
  wire [7:0]    dataGroup_14_27 = dataGroup_lo_1742[839:832];
  wire [2047:0] dataGroup_lo_1743 = {dataGroup_lo_hi_1743, dataGroup_lo_lo_1743};
  wire [2047:0] dataGroup_hi_1743 = {dataGroup_hi_hi_1743, dataGroup_hi_lo_1743};
  wire [7:0]    dataGroup_15_27 = dataGroup_lo_1743[895:888];
  wire [2047:0] dataGroup_lo_1744 = {dataGroup_lo_hi_1744, dataGroup_lo_lo_1744};
  wire [2047:0] dataGroup_hi_1744 = {dataGroup_hi_hi_1744, dataGroup_hi_lo_1744};
  wire [7:0]    dataGroup_16_27 = dataGroup_lo_1744[951:944];
  wire [2047:0] dataGroup_lo_1745 = {dataGroup_lo_hi_1745, dataGroup_lo_lo_1745};
  wire [2047:0] dataGroup_hi_1745 = {dataGroup_hi_hi_1745, dataGroup_hi_lo_1745};
  wire [7:0]    dataGroup_17_27 = dataGroup_lo_1745[1007:1000];
  wire [2047:0] dataGroup_lo_1746 = {dataGroup_lo_hi_1746, dataGroup_lo_lo_1746};
  wire [2047:0] dataGroup_hi_1746 = {dataGroup_hi_hi_1746, dataGroup_hi_lo_1746};
  wire [7:0]    dataGroup_18_27 = dataGroup_lo_1746[1063:1056];
  wire [2047:0] dataGroup_lo_1747 = {dataGroup_lo_hi_1747, dataGroup_lo_lo_1747};
  wire [2047:0] dataGroup_hi_1747 = {dataGroup_hi_hi_1747, dataGroup_hi_lo_1747};
  wire [7:0]    dataGroup_19_27 = dataGroup_lo_1747[1119:1112];
  wire [2047:0] dataGroup_lo_1748 = {dataGroup_lo_hi_1748, dataGroup_lo_lo_1748};
  wire [2047:0] dataGroup_hi_1748 = {dataGroup_hi_hi_1748, dataGroup_hi_lo_1748};
  wire [7:0]    dataGroup_20_27 = dataGroup_lo_1748[1175:1168];
  wire [2047:0] dataGroup_lo_1749 = {dataGroup_lo_hi_1749, dataGroup_lo_lo_1749};
  wire [2047:0] dataGroup_hi_1749 = {dataGroup_hi_hi_1749, dataGroup_hi_lo_1749};
  wire [7:0]    dataGroup_21_27 = dataGroup_lo_1749[1231:1224];
  wire [2047:0] dataGroup_lo_1750 = {dataGroup_lo_hi_1750, dataGroup_lo_lo_1750};
  wire [2047:0] dataGroup_hi_1750 = {dataGroup_hi_hi_1750, dataGroup_hi_lo_1750};
  wire [7:0]    dataGroup_22_27 = dataGroup_lo_1750[1287:1280];
  wire [2047:0] dataGroup_lo_1751 = {dataGroup_lo_hi_1751, dataGroup_lo_lo_1751};
  wire [2047:0] dataGroup_hi_1751 = {dataGroup_hi_hi_1751, dataGroup_hi_lo_1751};
  wire [7:0]    dataGroup_23_27 = dataGroup_lo_1751[1343:1336];
  wire [2047:0] dataGroup_lo_1752 = {dataGroup_lo_hi_1752, dataGroup_lo_lo_1752};
  wire [2047:0] dataGroup_hi_1752 = {dataGroup_hi_hi_1752, dataGroup_hi_lo_1752};
  wire [7:0]    dataGroup_24_27 = dataGroup_lo_1752[1399:1392];
  wire [2047:0] dataGroup_lo_1753 = {dataGroup_lo_hi_1753, dataGroup_lo_lo_1753};
  wire [2047:0] dataGroup_hi_1753 = {dataGroup_hi_hi_1753, dataGroup_hi_lo_1753};
  wire [7:0]    dataGroup_25_27 = dataGroup_lo_1753[1455:1448];
  wire [2047:0] dataGroup_lo_1754 = {dataGroup_lo_hi_1754, dataGroup_lo_lo_1754};
  wire [2047:0] dataGroup_hi_1754 = {dataGroup_hi_hi_1754, dataGroup_hi_lo_1754};
  wire [7:0]    dataGroup_26_27 = dataGroup_lo_1754[1511:1504];
  wire [2047:0] dataGroup_lo_1755 = {dataGroup_lo_hi_1755, dataGroup_lo_lo_1755};
  wire [2047:0] dataGroup_hi_1755 = {dataGroup_hi_hi_1755, dataGroup_hi_lo_1755};
  wire [7:0]    dataGroup_27_27 = dataGroup_lo_1755[1567:1560];
  wire [2047:0] dataGroup_lo_1756 = {dataGroup_lo_hi_1756, dataGroup_lo_lo_1756};
  wire [2047:0] dataGroup_hi_1756 = {dataGroup_hi_hi_1756, dataGroup_hi_lo_1756};
  wire [7:0]    dataGroup_28_27 = dataGroup_lo_1756[1623:1616];
  wire [2047:0] dataGroup_lo_1757 = {dataGroup_lo_hi_1757, dataGroup_lo_lo_1757};
  wire [2047:0] dataGroup_hi_1757 = {dataGroup_hi_hi_1757, dataGroup_hi_lo_1757};
  wire [7:0]    dataGroup_29_27 = dataGroup_lo_1757[1679:1672];
  wire [2047:0] dataGroup_lo_1758 = {dataGroup_lo_hi_1758, dataGroup_lo_lo_1758};
  wire [2047:0] dataGroup_hi_1758 = {dataGroup_hi_hi_1758, dataGroup_hi_lo_1758};
  wire [7:0]    dataGroup_30_27 = dataGroup_lo_1758[1735:1728];
  wire [2047:0] dataGroup_lo_1759 = {dataGroup_lo_hi_1759, dataGroup_lo_lo_1759};
  wire [2047:0] dataGroup_hi_1759 = {dataGroup_hi_hi_1759, dataGroup_hi_lo_1759};
  wire [7:0]    dataGroup_31_27 = dataGroup_lo_1759[1791:1784];
  wire [2047:0] dataGroup_lo_1760 = {dataGroup_lo_hi_1760, dataGroup_lo_lo_1760};
  wire [2047:0] dataGroup_hi_1760 = {dataGroup_hi_hi_1760, dataGroup_hi_lo_1760};
  wire [7:0]    dataGroup_32_27 = dataGroup_lo_1760[1847:1840];
  wire [2047:0] dataGroup_lo_1761 = {dataGroup_lo_hi_1761, dataGroup_lo_lo_1761};
  wire [2047:0] dataGroup_hi_1761 = {dataGroup_hi_hi_1761, dataGroup_hi_lo_1761};
  wire [7:0]    dataGroup_33_27 = dataGroup_lo_1761[1903:1896];
  wire [2047:0] dataGroup_lo_1762 = {dataGroup_lo_hi_1762, dataGroup_lo_lo_1762};
  wire [2047:0] dataGroup_hi_1762 = {dataGroup_hi_hi_1762, dataGroup_hi_lo_1762};
  wire [7:0]    dataGroup_34_27 = dataGroup_lo_1762[1959:1952];
  wire [2047:0] dataGroup_lo_1763 = {dataGroup_lo_hi_1763, dataGroup_lo_lo_1763};
  wire [2047:0] dataGroup_hi_1763 = {dataGroup_hi_hi_1763, dataGroup_hi_lo_1763};
  wire [7:0]    dataGroup_35_27 = dataGroup_lo_1763[2015:2008];
  wire [2047:0] dataGroup_lo_1764 = {dataGroup_lo_hi_1764, dataGroup_lo_lo_1764};
  wire [2047:0] dataGroup_hi_1764 = {dataGroup_hi_hi_1764, dataGroup_hi_lo_1764};
  wire [7:0]    dataGroup_36_27 = dataGroup_hi_1764[23:16];
  wire [2047:0] dataGroup_lo_1765 = {dataGroup_lo_hi_1765, dataGroup_lo_lo_1765};
  wire [2047:0] dataGroup_hi_1765 = {dataGroup_hi_hi_1765, dataGroup_hi_lo_1765};
  wire [7:0]    dataGroup_37_27 = dataGroup_hi_1765[79:72];
  wire [2047:0] dataGroup_lo_1766 = {dataGroup_lo_hi_1766, dataGroup_lo_lo_1766};
  wire [2047:0] dataGroup_hi_1766 = {dataGroup_hi_hi_1766, dataGroup_hi_lo_1766};
  wire [7:0]    dataGroup_38_27 = dataGroup_hi_1766[135:128];
  wire [2047:0] dataGroup_lo_1767 = {dataGroup_lo_hi_1767, dataGroup_lo_lo_1767};
  wire [2047:0] dataGroup_hi_1767 = {dataGroup_hi_hi_1767, dataGroup_hi_lo_1767};
  wire [7:0]    dataGroup_39_27 = dataGroup_hi_1767[191:184];
  wire [2047:0] dataGroup_lo_1768 = {dataGroup_lo_hi_1768, dataGroup_lo_lo_1768};
  wire [2047:0] dataGroup_hi_1768 = {dataGroup_hi_hi_1768, dataGroup_hi_lo_1768};
  wire [7:0]    dataGroup_40_27 = dataGroup_hi_1768[247:240];
  wire [2047:0] dataGroup_lo_1769 = {dataGroup_lo_hi_1769, dataGroup_lo_lo_1769};
  wire [2047:0] dataGroup_hi_1769 = {dataGroup_hi_hi_1769, dataGroup_hi_lo_1769};
  wire [7:0]    dataGroup_41_27 = dataGroup_hi_1769[303:296];
  wire [2047:0] dataGroup_lo_1770 = {dataGroup_lo_hi_1770, dataGroup_lo_lo_1770};
  wire [2047:0] dataGroup_hi_1770 = {dataGroup_hi_hi_1770, dataGroup_hi_lo_1770};
  wire [7:0]    dataGroup_42_27 = dataGroup_hi_1770[359:352];
  wire [2047:0] dataGroup_lo_1771 = {dataGroup_lo_hi_1771, dataGroup_lo_lo_1771};
  wire [2047:0] dataGroup_hi_1771 = {dataGroup_hi_hi_1771, dataGroup_hi_lo_1771};
  wire [7:0]    dataGroup_43_27 = dataGroup_hi_1771[415:408];
  wire [2047:0] dataGroup_lo_1772 = {dataGroup_lo_hi_1772, dataGroup_lo_lo_1772};
  wire [2047:0] dataGroup_hi_1772 = {dataGroup_hi_hi_1772, dataGroup_hi_lo_1772};
  wire [7:0]    dataGroup_44_27 = dataGroup_hi_1772[471:464];
  wire [2047:0] dataGroup_lo_1773 = {dataGroup_lo_hi_1773, dataGroup_lo_lo_1773};
  wire [2047:0] dataGroup_hi_1773 = {dataGroup_hi_hi_1773, dataGroup_hi_lo_1773};
  wire [7:0]    dataGroup_45_27 = dataGroup_hi_1773[527:520];
  wire [2047:0] dataGroup_lo_1774 = {dataGroup_lo_hi_1774, dataGroup_lo_lo_1774};
  wire [2047:0] dataGroup_hi_1774 = {dataGroup_hi_hi_1774, dataGroup_hi_lo_1774};
  wire [7:0]    dataGroup_46_27 = dataGroup_hi_1774[583:576];
  wire [2047:0] dataGroup_lo_1775 = {dataGroup_lo_hi_1775, dataGroup_lo_lo_1775};
  wire [2047:0] dataGroup_hi_1775 = {dataGroup_hi_hi_1775, dataGroup_hi_lo_1775};
  wire [7:0]    dataGroup_47_27 = dataGroup_hi_1775[639:632];
  wire [2047:0] dataGroup_lo_1776 = {dataGroup_lo_hi_1776, dataGroup_lo_lo_1776};
  wire [2047:0] dataGroup_hi_1776 = {dataGroup_hi_hi_1776, dataGroup_hi_lo_1776};
  wire [7:0]    dataGroup_48_27 = dataGroup_hi_1776[695:688];
  wire [2047:0] dataGroup_lo_1777 = {dataGroup_lo_hi_1777, dataGroup_lo_lo_1777};
  wire [2047:0] dataGroup_hi_1777 = {dataGroup_hi_hi_1777, dataGroup_hi_lo_1777};
  wire [7:0]    dataGroup_49_27 = dataGroup_hi_1777[751:744];
  wire [2047:0] dataGroup_lo_1778 = {dataGroup_lo_hi_1778, dataGroup_lo_lo_1778};
  wire [2047:0] dataGroup_hi_1778 = {dataGroup_hi_hi_1778, dataGroup_hi_lo_1778};
  wire [7:0]    dataGroup_50_27 = dataGroup_hi_1778[807:800];
  wire [2047:0] dataGroup_lo_1779 = {dataGroup_lo_hi_1779, dataGroup_lo_lo_1779};
  wire [2047:0] dataGroup_hi_1779 = {dataGroup_hi_hi_1779, dataGroup_hi_lo_1779};
  wire [7:0]    dataGroup_51_27 = dataGroup_hi_1779[863:856];
  wire [2047:0] dataGroup_lo_1780 = {dataGroup_lo_hi_1780, dataGroup_lo_lo_1780};
  wire [2047:0] dataGroup_hi_1780 = {dataGroup_hi_hi_1780, dataGroup_hi_lo_1780};
  wire [7:0]    dataGroup_52_27 = dataGroup_hi_1780[919:912];
  wire [2047:0] dataGroup_lo_1781 = {dataGroup_lo_hi_1781, dataGroup_lo_lo_1781};
  wire [2047:0] dataGroup_hi_1781 = {dataGroup_hi_hi_1781, dataGroup_hi_lo_1781};
  wire [7:0]    dataGroup_53_27 = dataGroup_hi_1781[975:968];
  wire [2047:0] dataGroup_lo_1782 = {dataGroup_lo_hi_1782, dataGroup_lo_lo_1782};
  wire [2047:0] dataGroup_hi_1782 = {dataGroup_hi_hi_1782, dataGroup_hi_lo_1782};
  wire [7:0]    dataGroup_54_27 = dataGroup_hi_1782[1031:1024];
  wire [2047:0] dataGroup_lo_1783 = {dataGroup_lo_hi_1783, dataGroup_lo_lo_1783};
  wire [2047:0] dataGroup_hi_1783 = {dataGroup_hi_hi_1783, dataGroup_hi_lo_1783};
  wire [7:0]    dataGroup_55_27 = dataGroup_hi_1783[1087:1080];
  wire [2047:0] dataGroup_lo_1784 = {dataGroup_lo_hi_1784, dataGroup_lo_lo_1784};
  wire [2047:0] dataGroup_hi_1784 = {dataGroup_hi_hi_1784, dataGroup_hi_lo_1784};
  wire [7:0]    dataGroup_56_27 = dataGroup_hi_1784[1143:1136];
  wire [2047:0] dataGroup_lo_1785 = {dataGroup_lo_hi_1785, dataGroup_lo_lo_1785};
  wire [2047:0] dataGroup_hi_1785 = {dataGroup_hi_hi_1785, dataGroup_hi_lo_1785};
  wire [7:0]    dataGroup_57_27 = dataGroup_hi_1785[1199:1192];
  wire [2047:0] dataGroup_lo_1786 = {dataGroup_lo_hi_1786, dataGroup_lo_lo_1786};
  wire [2047:0] dataGroup_hi_1786 = {dataGroup_hi_hi_1786, dataGroup_hi_lo_1786};
  wire [7:0]    dataGroup_58_27 = dataGroup_hi_1786[1255:1248];
  wire [2047:0] dataGroup_lo_1787 = {dataGroup_lo_hi_1787, dataGroup_lo_lo_1787};
  wire [2047:0] dataGroup_hi_1787 = {dataGroup_hi_hi_1787, dataGroup_hi_lo_1787};
  wire [7:0]    dataGroup_59_27 = dataGroup_hi_1787[1311:1304];
  wire [2047:0] dataGroup_lo_1788 = {dataGroup_lo_hi_1788, dataGroup_lo_lo_1788};
  wire [2047:0] dataGroup_hi_1788 = {dataGroup_hi_hi_1788, dataGroup_hi_lo_1788};
  wire [7:0]    dataGroup_60_27 = dataGroup_hi_1788[1367:1360];
  wire [2047:0] dataGroup_lo_1789 = {dataGroup_lo_hi_1789, dataGroup_lo_lo_1789};
  wire [2047:0] dataGroup_hi_1789 = {dataGroup_hi_hi_1789, dataGroup_hi_lo_1789};
  wire [7:0]    dataGroup_61_27 = dataGroup_hi_1789[1423:1416];
  wire [2047:0] dataGroup_lo_1790 = {dataGroup_lo_hi_1790, dataGroup_lo_lo_1790};
  wire [2047:0] dataGroup_hi_1790 = {dataGroup_hi_hi_1790, dataGroup_hi_lo_1790};
  wire [7:0]    dataGroup_62_27 = dataGroup_hi_1790[1479:1472];
  wire [2047:0] dataGroup_lo_1791 = {dataGroup_lo_hi_1791, dataGroup_lo_lo_1791};
  wire [2047:0] dataGroup_hi_1791 = {dataGroup_hi_hi_1791, dataGroup_hi_lo_1791};
  wire [7:0]    dataGroup_63_27 = dataGroup_hi_1791[1535:1528];
  wire [15:0]   res_lo_lo_lo_lo_lo_27 = {dataGroup_1_27, dataGroup_0_27};
  wire [15:0]   res_lo_lo_lo_lo_hi_27 = {dataGroup_3_27, dataGroup_2_27};
  wire [31:0]   res_lo_lo_lo_lo_27 = {res_lo_lo_lo_lo_hi_27, res_lo_lo_lo_lo_lo_27};
  wire [15:0]   res_lo_lo_lo_hi_lo_27 = {dataGroup_5_27, dataGroup_4_27};
  wire [15:0]   res_lo_lo_lo_hi_hi_27 = {dataGroup_7_27, dataGroup_6_27};
  wire [31:0]   res_lo_lo_lo_hi_27 = {res_lo_lo_lo_hi_hi_27, res_lo_lo_lo_hi_lo_27};
  wire [63:0]   res_lo_lo_lo_27 = {res_lo_lo_lo_hi_27, res_lo_lo_lo_lo_27};
  wire [15:0]   res_lo_lo_hi_lo_lo_27 = {dataGroup_9_27, dataGroup_8_27};
  wire [15:0]   res_lo_lo_hi_lo_hi_27 = {dataGroup_11_27, dataGroup_10_27};
  wire [31:0]   res_lo_lo_hi_lo_27 = {res_lo_lo_hi_lo_hi_27, res_lo_lo_hi_lo_lo_27};
  wire [15:0]   res_lo_lo_hi_hi_lo_27 = {dataGroup_13_27, dataGroup_12_27};
  wire [15:0]   res_lo_lo_hi_hi_hi_27 = {dataGroup_15_27, dataGroup_14_27};
  wire [31:0]   res_lo_lo_hi_hi_27 = {res_lo_lo_hi_hi_hi_27, res_lo_lo_hi_hi_lo_27};
  wire [63:0]   res_lo_lo_hi_27 = {res_lo_lo_hi_hi_27, res_lo_lo_hi_lo_27};
  wire [127:0]  res_lo_lo_27 = {res_lo_lo_hi_27, res_lo_lo_lo_27};
  wire [15:0]   res_lo_hi_lo_lo_lo_27 = {dataGroup_17_27, dataGroup_16_27};
  wire [15:0]   res_lo_hi_lo_lo_hi_27 = {dataGroup_19_27, dataGroup_18_27};
  wire [31:0]   res_lo_hi_lo_lo_27 = {res_lo_hi_lo_lo_hi_27, res_lo_hi_lo_lo_lo_27};
  wire [15:0]   res_lo_hi_lo_hi_lo_27 = {dataGroup_21_27, dataGroup_20_27};
  wire [15:0]   res_lo_hi_lo_hi_hi_27 = {dataGroup_23_27, dataGroup_22_27};
  wire [31:0]   res_lo_hi_lo_hi_27 = {res_lo_hi_lo_hi_hi_27, res_lo_hi_lo_hi_lo_27};
  wire [63:0]   res_lo_hi_lo_27 = {res_lo_hi_lo_hi_27, res_lo_hi_lo_lo_27};
  wire [15:0]   res_lo_hi_hi_lo_lo_27 = {dataGroup_25_27, dataGroup_24_27};
  wire [15:0]   res_lo_hi_hi_lo_hi_27 = {dataGroup_27_27, dataGroup_26_27};
  wire [31:0]   res_lo_hi_hi_lo_27 = {res_lo_hi_hi_lo_hi_27, res_lo_hi_hi_lo_lo_27};
  wire [15:0]   res_lo_hi_hi_hi_lo_27 = {dataGroup_29_27, dataGroup_28_27};
  wire [15:0]   res_lo_hi_hi_hi_hi_27 = {dataGroup_31_27, dataGroup_30_27};
  wire [31:0]   res_lo_hi_hi_hi_27 = {res_lo_hi_hi_hi_hi_27, res_lo_hi_hi_hi_lo_27};
  wire [63:0]   res_lo_hi_hi_27 = {res_lo_hi_hi_hi_27, res_lo_hi_hi_lo_27};
  wire [127:0]  res_lo_hi_27 = {res_lo_hi_hi_27, res_lo_hi_lo_27};
  wire [255:0]  res_lo_27 = {res_lo_hi_27, res_lo_lo_27};
  wire [15:0]   res_hi_lo_lo_lo_lo_27 = {dataGroup_33_27, dataGroup_32_27};
  wire [15:0]   res_hi_lo_lo_lo_hi_27 = {dataGroup_35_27, dataGroup_34_27};
  wire [31:0]   res_hi_lo_lo_lo_27 = {res_hi_lo_lo_lo_hi_27, res_hi_lo_lo_lo_lo_27};
  wire [15:0]   res_hi_lo_lo_hi_lo_27 = {dataGroup_37_27, dataGroup_36_27};
  wire [15:0]   res_hi_lo_lo_hi_hi_27 = {dataGroup_39_27, dataGroup_38_27};
  wire [31:0]   res_hi_lo_lo_hi_27 = {res_hi_lo_lo_hi_hi_27, res_hi_lo_lo_hi_lo_27};
  wire [63:0]   res_hi_lo_lo_27 = {res_hi_lo_lo_hi_27, res_hi_lo_lo_lo_27};
  wire [15:0]   res_hi_lo_hi_lo_lo_27 = {dataGroup_41_27, dataGroup_40_27};
  wire [15:0]   res_hi_lo_hi_lo_hi_27 = {dataGroup_43_27, dataGroup_42_27};
  wire [31:0]   res_hi_lo_hi_lo_27 = {res_hi_lo_hi_lo_hi_27, res_hi_lo_hi_lo_lo_27};
  wire [15:0]   res_hi_lo_hi_hi_lo_27 = {dataGroup_45_27, dataGroup_44_27};
  wire [15:0]   res_hi_lo_hi_hi_hi_27 = {dataGroup_47_27, dataGroup_46_27};
  wire [31:0]   res_hi_lo_hi_hi_27 = {res_hi_lo_hi_hi_hi_27, res_hi_lo_hi_hi_lo_27};
  wire [63:0]   res_hi_lo_hi_27 = {res_hi_lo_hi_hi_27, res_hi_lo_hi_lo_27};
  wire [127:0]  res_hi_lo_27 = {res_hi_lo_hi_27, res_hi_lo_lo_27};
  wire [15:0]   res_hi_hi_lo_lo_lo_27 = {dataGroup_49_27, dataGroup_48_27};
  wire [15:0]   res_hi_hi_lo_lo_hi_27 = {dataGroup_51_27, dataGroup_50_27};
  wire [31:0]   res_hi_hi_lo_lo_27 = {res_hi_hi_lo_lo_hi_27, res_hi_hi_lo_lo_lo_27};
  wire [15:0]   res_hi_hi_lo_hi_lo_27 = {dataGroup_53_27, dataGroup_52_27};
  wire [15:0]   res_hi_hi_lo_hi_hi_27 = {dataGroup_55_27, dataGroup_54_27};
  wire [31:0]   res_hi_hi_lo_hi_27 = {res_hi_hi_lo_hi_hi_27, res_hi_hi_lo_hi_lo_27};
  wire [63:0]   res_hi_hi_lo_27 = {res_hi_hi_lo_hi_27, res_hi_hi_lo_lo_27};
  wire [15:0]   res_hi_hi_hi_lo_lo_27 = {dataGroup_57_27, dataGroup_56_27};
  wire [15:0]   res_hi_hi_hi_lo_hi_27 = {dataGroup_59_27, dataGroup_58_27};
  wire [31:0]   res_hi_hi_hi_lo_27 = {res_hi_hi_hi_lo_hi_27, res_hi_hi_hi_lo_lo_27};
  wire [15:0]   res_hi_hi_hi_hi_lo_27 = {dataGroup_61_27, dataGroup_60_27};
  wire [15:0]   res_hi_hi_hi_hi_hi_27 = {dataGroup_63_27, dataGroup_62_27};
  wire [31:0]   res_hi_hi_hi_hi_27 = {res_hi_hi_hi_hi_hi_27, res_hi_hi_hi_hi_lo_27};
  wire [63:0]   res_hi_hi_hi_27 = {res_hi_hi_hi_hi_27, res_hi_hi_hi_lo_27};
  wire [127:0]  res_hi_hi_27 = {res_hi_hi_hi_27, res_hi_hi_lo_27};
  wire [255:0]  res_hi_27 = {res_hi_hi_27, res_hi_lo_27};
  wire [511:0]  res_54 = {res_hi_27, res_lo_27};
  wire [1023:0] lo_lo_6 = {res_49, res_48};
  wire [1023:0] lo_hi_6 = {res_51, res_50};
  wire [2047:0] lo_6 = {lo_hi_6, lo_lo_6};
  wire [1023:0] hi_lo_6 = {res_53, res_52};
  wire [1023:0] hi_hi_6 = {512'h0, res_54};
  wire [2047:0] hi_6 = {hi_hi_6, hi_lo_6};
  wire [4095:0] regroupLoadData_0_6 = {hi_6, lo_6};
  wire [2047:0] dataGroup_lo_1792 = {dataGroup_lo_hi_1792, dataGroup_lo_lo_1792};
  wire [2047:0] dataGroup_hi_1792 = {dataGroup_hi_hi_1792, dataGroup_hi_lo_1792};
  wire [7:0]    dataGroup_0_28 = dataGroup_lo_1792[7:0];
  wire [2047:0] dataGroup_lo_1793 = {dataGroup_lo_hi_1793, dataGroup_lo_lo_1793};
  wire [2047:0] dataGroup_hi_1793 = {dataGroup_hi_hi_1793, dataGroup_hi_lo_1793};
  wire [7:0]    dataGroup_1_28 = dataGroup_lo_1793[71:64];
  wire [2047:0] dataGroup_lo_1794 = {dataGroup_lo_hi_1794, dataGroup_lo_lo_1794};
  wire [2047:0] dataGroup_hi_1794 = {dataGroup_hi_hi_1794, dataGroup_hi_lo_1794};
  wire [7:0]    dataGroup_2_28 = dataGroup_lo_1794[135:128];
  wire [2047:0] dataGroup_lo_1795 = {dataGroup_lo_hi_1795, dataGroup_lo_lo_1795};
  wire [2047:0] dataGroup_hi_1795 = {dataGroup_hi_hi_1795, dataGroup_hi_lo_1795};
  wire [7:0]    dataGroup_3_28 = dataGroup_lo_1795[199:192];
  wire [2047:0] dataGroup_lo_1796 = {dataGroup_lo_hi_1796, dataGroup_lo_lo_1796};
  wire [2047:0] dataGroup_hi_1796 = {dataGroup_hi_hi_1796, dataGroup_hi_lo_1796};
  wire [7:0]    dataGroup_4_28 = dataGroup_lo_1796[263:256];
  wire [2047:0] dataGroup_lo_1797 = {dataGroup_lo_hi_1797, dataGroup_lo_lo_1797};
  wire [2047:0] dataGroup_hi_1797 = {dataGroup_hi_hi_1797, dataGroup_hi_lo_1797};
  wire [7:0]    dataGroup_5_28 = dataGroup_lo_1797[327:320];
  wire [2047:0] dataGroup_lo_1798 = {dataGroup_lo_hi_1798, dataGroup_lo_lo_1798};
  wire [2047:0] dataGroup_hi_1798 = {dataGroup_hi_hi_1798, dataGroup_hi_lo_1798};
  wire [7:0]    dataGroup_6_28 = dataGroup_lo_1798[391:384];
  wire [2047:0] dataGroup_lo_1799 = {dataGroup_lo_hi_1799, dataGroup_lo_lo_1799};
  wire [2047:0] dataGroup_hi_1799 = {dataGroup_hi_hi_1799, dataGroup_hi_lo_1799};
  wire [7:0]    dataGroup_7_28 = dataGroup_lo_1799[455:448];
  wire [2047:0] dataGroup_lo_1800 = {dataGroup_lo_hi_1800, dataGroup_lo_lo_1800};
  wire [2047:0] dataGroup_hi_1800 = {dataGroup_hi_hi_1800, dataGroup_hi_lo_1800};
  wire [7:0]    dataGroup_8_28 = dataGroup_lo_1800[519:512];
  wire [2047:0] dataGroup_lo_1801 = {dataGroup_lo_hi_1801, dataGroup_lo_lo_1801};
  wire [2047:0] dataGroup_hi_1801 = {dataGroup_hi_hi_1801, dataGroup_hi_lo_1801};
  wire [7:0]    dataGroup_9_28 = dataGroup_lo_1801[583:576];
  wire [2047:0] dataGroup_lo_1802 = {dataGroup_lo_hi_1802, dataGroup_lo_lo_1802};
  wire [2047:0] dataGroup_hi_1802 = {dataGroup_hi_hi_1802, dataGroup_hi_lo_1802};
  wire [7:0]    dataGroup_10_28 = dataGroup_lo_1802[647:640];
  wire [2047:0] dataGroup_lo_1803 = {dataGroup_lo_hi_1803, dataGroup_lo_lo_1803};
  wire [2047:0] dataGroup_hi_1803 = {dataGroup_hi_hi_1803, dataGroup_hi_lo_1803};
  wire [7:0]    dataGroup_11_28 = dataGroup_lo_1803[711:704];
  wire [2047:0] dataGroup_lo_1804 = {dataGroup_lo_hi_1804, dataGroup_lo_lo_1804};
  wire [2047:0] dataGroup_hi_1804 = {dataGroup_hi_hi_1804, dataGroup_hi_lo_1804};
  wire [7:0]    dataGroup_12_28 = dataGroup_lo_1804[775:768];
  wire [2047:0] dataGroup_lo_1805 = {dataGroup_lo_hi_1805, dataGroup_lo_lo_1805};
  wire [2047:0] dataGroup_hi_1805 = {dataGroup_hi_hi_1805, dataGroup_hi_lo_1805};
  wire [7:0]    dataGroup_13_28 = dataGroup_lo_1805[839:832];
  wire [2047:0] dataGroup_lo_1806 = {dataGroup_lo_hi_1806, dataGroup_lo_lo_1806};
  wire [2047:0] dataGroup_hi_1806 = {dataGroup_hi_hi_1806, dataGroup_hi_lo_1806};
  wire [7:0]    dataGroup_14_28 = dataGroup_lo_1806[903:896];
  wire [2047:0] dataGroup_lo_1807 = {dataGroup_lo_hi_1807, dataGroup_lo_lo_1807};
  wire [2047:0] dataGroup_hi_1807 = {dataGroup_hi_hi_1807, dataGroup_hi_lo_1807};
  wire [7:0]    dataGroup_15_28 = dataGroup_lo_1807[967:960];
  wire [2047:0] dataGroup_lo_1808 = {dataGroup_lo_hi_1808, dataGroup_lo_lo_1808};
  wire [2047:0] dataGroup_hi_1808 = {dataGroup_hi_hi_1808, dataGroup_hi_lo_1808};
  wire [7:0]    dataGroup_16_28 = dataGroup_lo_1808[1031:1024];
  wire [2047:0] dataGroup_lo_1809 = {dataGroup_lo_hi_1809, dataGroup_lo_lo_1809};
  wire [2047:0] dataGroup_hi_1809 = {dataGroup_hi_hi_1809, dataGroup_hi_lo_1809};
  wire [7:0]    dataGroup_17_28 = dataGroup_lo_1809[1095:1088];
  wire [2047:0] dataGroup_lo_1810 = {dataGroup_lo_hi_1810, dataGroup_lo_lo_1810};
  wire [2047:0] dataGroup_hi_1810 = {dataGroup_hi_hi_1810, dataGroup_hi_lo_1810};
  wire [7:0]    dataGroup_18_28 = dataGroup_lo_1810[1159:1152];
  wire [2047:0] dataGroup_lo_1811 = {dataGroup_lo_hi_1811, dataGroup_lo_lo_1811};
  wire [2047:0] dataGroup_hi_1811 = {dataGroup_hi_hi_1811, dataGroup_hi_lo_1811};
  wire [7:0]    dataGroup_19_28 = dataGroup_lo_1811[1223:1216];
  wire [2047:0] dataGroup_lo_1812 = {dataGroup_lo_hi_1812, dataGroup_lo_lo_1812};
  wire [2047:0] dataGroup_hi_1812 = {dataGroup_hi_hi_1812, dataGroup_hi_lo_1812};
  wire [7:0]    dataGroup_20_28 = dataGroup_lo_1812[1287:1280];
  wire [2047:0] dataGroup_lo_1813 = {dataGroup_lo_hi_1813, dataGroup_lo_lo_1813};
  wire [2047:0] dataGroup_hi_1813 = {dataGroup_hi_hi_1813, dataGroup_hi_lo_1813};
  wire [7:0]    dataGroup_21_28 = dataGroup_lo_1813[1351:1344];
  wire [2047:0] dataGroup_lo_1814 = {dataGroup_lo_hi_1814, dataGroup_lo_lo_1814};
  wire [2047:0] dataGroup_hi_1814 = {dataGroup_hi_hi_1814, dataGroup_hi_lo_1814};
  wire [7:0]    dataGroup_22_28 = dataGroup_lo_1814[1415:1408];
  wire [2047:0] dataGroup_lo_1815 = {dataGroup_lo_hi_1815, dataGroup_lo_lo_1815};
  wire [2047:0] dataGroup_hi_1815 = {dataGroup_hi_hi_1815, dataGroup_hi_lo_1815};
  wire [7:0]    dataGroup_23_28 = dataGroup_lo_1815[1479:1472];
  wire [2047:0] dataGroup_lo_1816 = {dataGroup_lo_hi_1816, dataGroup_lo_lo_1816};
  wire [2047:0] dataGroup_hi_1816 = {dataGroup_hi_hi_1816, dataGroup_hi_lo_1816};
  wire [7:0]    dataGroup_24_28 = dataGroup_lo_1816[1543:1536];
  wire [2047:0] dataGroup_lo_1817 = {dataGroup_lo_hi_1817, dataGroup_lo_lo_1817};
  wire [2047:0] dataGroup_hi_1817 = {dataGroup_hi_hi_1817, dataGroup_hi_lo_1817};
  wire [7:0]    dataGroup_25_28 = dataGroup_lo_1817[1607:1600];
  wire [2047:0] dataGroup_lo_1818 = {dataGroup_lo_hi_1818, dataGroup_lo_lo_1818};
  wire [2047:0] dataGroup_hi_1818 = {dataGroup_hi_hi_1818, dataGroup_hi_lo_1818};
  wire [7:0]    dataGroup_26_28 = dataGroup_lo_1818[1671:1664];
  wire [2047:0] dataGroup_lo_1819 = {dataGroup_lo_hi_1819, dataGroup_lo_lo_1819};
  wire [2047:0] dataGroup_hi_1819 = {dataGroup_hi_hi_1819, dataGroup_hi_lo_1819};
  wire [7:0]    dataGroup_27_28 = dataGroup_lo_1819[1735:1728];
  wire [2047:0] dataGroup_lo_1820 = {dataGroup_lo_hi_1820, dataGroup_lo_lo_1820};
  wire [2047:0] dataGroup_hi_1820 = {dataGroup_hi_hi_1820, dataGroup_hi_lo_1820};
  wire [7:0]    dataGroup_28_28 = dataGroup_lo_1820[1799:1792];
  wire [2047:0] dataGroup_lo_1821 = {dataGroup_lo_hi_1821, dataGroup_lo_lo_1821};
  wire [2047:0] dataGroup_hi_1821 = {dataGroup_hi_hi_1821, dataGroup_hi_lo_1821};
  wire [7:0]    dataGroup_29_28 = dataGroup_lo_1821[1863:1856];
  wire [2047:0] dataGroup_lo_1822 = {dataGroup_lo_hi_1822, dataGroup_lo_lo_1822};
  wire [2047:0] dataGroup_hi_1822 = {dataGroup_hi_hi_1822, dataGroup_hi_lo_1822};
  wire [7:0]    dataGroup_30_28 = dataGroup_lo_1822[1927:1920];
  wire [2047:0] dataGroup_lo_1823 = {dataGroup_lo_hi_1823, dataGroup_lo_lo_1823};
  wire [2047:0] dataGroup_hi_1823 = {dataGroup_hi_hi_1823, dataGroup_hi_lo_1823};
  wire [7:0]    dataGroup_31_28 = dataGroup_lo_1823[1991:1984];
  wire [2047:0] dataGroup_lo_1824 = {dataGroup_lo_hi_1824, dataGroup_lo_lo_1824};
  wire [2047:0] dataGroup_hi_1824 = {dataGroup_hi_hi_1824, dataGroup_hi_lo_1824};
  wire [7:0]    dataGroup_32_28 = dataGroup_hi_1824[7:0];
  wire [2047:0] dataGroup_lo_1825 = {dataGroup_lo_hi_1825, dataGroup_lo_lo_1825};
  wire [2047:0] dataGroup_hi_1825 = {dataGroup_hi_hi_1825, dataGroup_hi_lo_1825};
  wire [7:0]    dataGroup_33_28 = dataGroup_hi_1825[71:64];
  wire [2047:0] dataGroup_lo_1826 = {dataGroup_lo_hi_1826, dataGroup_lo_lo_1826};
  wire [2047:0] dataGroup_hi_1826 = {dataGroup_hi_hi_1826, dataGroup_hi_lo_1826};
  wire [7:0]    dataGroup_34_28 = dataGroup_hi_1826[135:128];
  wire [2047:0] dataGroup_lo_1827 = {dataGroup_lo_hi_1827, dataGroup_lo_lo_1827};
  wire [2047:0] dataGroup_hi_1827 = {dataGroup_hi_hi_1827, dataGroup_hi_lo_1827};
  wire [7:0]    dataGroup_35_28 = dataGroup_hi_1827[199:192];
  wire [2047:0] dataGroup_lo_1828 = {dataGroup_lo_hi_1828, dataGroup_lo_lo_1828};
  wire [2047:0] dataGroup_hi_1828 = {dataGroup_hi_hi_1828, dataGroup_hi_lo_1828};
  wire [7:0]    dataGroup_36_28 = dataGroup_hi_1828[263:256];
  wire [2047:0] dataGroup_lo_1829 = {dataGroup_lo_hi_1829, dataGroup_lo_lo_1829};
  wire [2047:0] dataGroup_hi_1829 = {dataGroup_hi_hi_1829, dataGroup_hi_lo_1829};
  wire [7:0]    dataGroup_37_28 = dataGroup_hi_1829[327:320];
  wire [2047:0] dataGroup_lo_1830 = {dataGroup_lo_hi_1830, dataGroup_lo_lo_1830};
  wire [2047:0] dataGroup_hi_1830 = {dataGroup_hi_hi_1830, dataGroup_hi_lo_1830};
  wire [7:0]    dataGroup_38_28 = dataGroup_hi_1830[391:384];
  wire [2047:0] dataGroup_lo_1831 = {dataGroup_lo_hi_1831, dataGroup_lo_lo_1831};
  wire [2047:0] dataGroup_hi_1831 = {dataGroup_hi_hi_1831, dataGroup_hi_lo_1831};
  wire [7:0]    dataGroup_39_28 = dataGroup_hi_1831[455:448];
  wire [2047:0] dataGroup_lo_1832 = {dataGroup_lo_hi_1832, dataGroup_lo_lo_1832};
  wire [2047:0] dataGroup_hi_1832 = {dataGroup_hi_hi_1832, dataGroup_hi_lo_1832};
  wire [7:0]    dataGroup_40_28 = dataGroup_hi_1832[519:512];
  wire [2047:0] dataGroup_lo_1833 = {dataGroup_lo_hi_1833, dataGroup_lo_lo_1833};
  wire [2047:0] dataGroup_hi_1833 = {dataGroup_hi_hi_1833, dataGroup_hi_lo_1833};
  wire [7:0]    dataGroup_41_28 = dataGroup_hi_1833[583:576];
  wire [2047:0] dataGroup_lo_1834 = {dataGroup_lo_hi_1834, dataGroup_lo_lo_1834};
  wire [2047:0] dataGroup_hi_1834 = {dataGroup_hi_hi_1834, dataGroup_hi_lo_1834};
  wire [7:0]    dataGroup_42_28 = dataGroup_hi_1834[647:640];
  wire [2047:0] dataGroup_lo_1835 = {dataGroup_lo_hi_1835, dataGroup_lo_lo_1835};
  wire [2047:0] dataGroup_hi_1835 = {dataGroup_hi_hi_1835, dataGroup_hi_lo_1835};
  wire [7:0]    dataGroup_43_28 = dataGroup_hi_1835[711:704];
  wire [2047:0] dataGroup_lo_1836 = {dataGroup_lo_hi_1836, dataGroup_lo_lo_1836};
  wire [2047:0] dataGroup_hi_1836 = {dataGroup_hi_hi_1836, dataGroup_hi_lo_1836};
  wire [7:0]    dataGroup_44_28 = dataGroup_hi_1836[775:768];
  wire [2047:0] dataGroup_lo_1837 = {dataGroup_lo_hi_1837, dataGroup_lo_lo_1837};
  wire [2047:0] dataGroup_hi_1837 = {dataGroup_hi_hi_1837, dataGroup_hi_lo_1837};
  wire [7:0]    dataGroup_45_28 = dataGroup_hi_1837[839:832];
  wire [2047:0] dataGroup_lo_1838 = {dataGroup_lo_hi_1838, dataGroup_lo_lo_1838};
  wire [2047:0] dataGroup_hi_1838 = {dataGroup_hi_hi_1838, dataGroup_hi_lo_1838};
  wire [7:0]    dataGroup_46_28 = dataGroup_hi_1838[903:896];
  wire [2047:0] dataGroup_lo_1839 = {dataGroup_lo_hi_1839, dataGroup_lo_lo_1839};
  wire [2047:0] dataGroup_hi_1839 = {dataGroup_hi_hi_1839, dataGroup_hi_lo_1839};
  wire [7:0]    dataGroup_47_28 = dataGroup_hi_1839[967:960];
  wire [2047:0] dataGroup_lo_1840 = {dataGroup_lo_hi_1840, dataGroup_lo_lo_1840};
  wire [2047:0] dataGroup_hi_1840 = {dataGroup_hi_hi_1840, dataGroup_hi_lo_1840};
  wire [7:0]    dataGroup_48_28 = dataGroup_hi_1840[1031:1024];
  wire [2047:0] dataGroup_lo_1841 = {dataGroup_lo_hi_1841, dataGroup_lo_lo_1841};
  wire [2047:0] dataGroup_hi_1841 = {dataGroup_hi_hi_1841, dataGroup_hi_lo_1841};
  wire [7:0]    dataGroup_49_28 = dataGroup_hi_1841[1095:1088];
  wire [2047:0] dataGroup_lo_1842 = {dataGroup_lo_hi_1842, dataGroup_lo_lo_1842};
  wire [2047:0] dataGroup_hi_1842 = {dataGroup_hi_hi_1842, dataGroup_hi_lo_1842};
  wire [7:0]    dataGroup_50_28 = dataGroup_hi_1842[1159:1152];
  wire [2047:0] dataGroup_lo_1843 = {dataGroup_lo_hi_1843, dataGroup_lo_lo_1843};
  wire [2047:0] dataGroup_hi_1843 = {dataGroup_hi_hi_1843, dataGroup_hi_lo_1843};
  wire [7:0]    dataGroup_51_28 = dataGroup_hi_1843[1223:1216];
  wire [2047:0] dataGroup_lo_1844 = {dataGroup_lo_hi_1844, dataGroup_lo_lo_1844};
  wire [2047:0] dataGroup_hi_1844 = {dataGroup_hi_hi_1844, dataGroup_hi_lo_1844};
  wire [7:0]    dataGroup_52_28 = dataGroup_hi_1844[1287:1280];
  wire [2047:0] dataGroup_lo_1845 = {dataGroup_lo_hi_1845, dataGroup_lo_lo_1845};
  wire [2047:0] dataGroup_hi_1845 = {dataGroup_hi_hi_1845, dataGroup_hi_lo_1845};
  wire [7:0]    dataGroup_53_28 = dataGroup_hi_1845[1351:1344];
  wire [2047:0] dataGroup_lo_1846 = {dataGroup_lo_hi_1846, dataGroup_lo_lo_1846};
  wire [2047:0] dataGroup_hi_1846 = {dataGroup_hi_hi_1846, dataGroup_hi_lo_1846};
  wire [7:0]    dataGroup_54_28 = dataGroup_hi_1846[1415:1408];
  wire [2047:0] dataGroup_lo_1847 = {dataGroup_lo_hi_1847, dataGroup_lo_lo_1847};
  wire [2047:0] dataGroup_hi_1847 = {dataGroup_hi_hi_1847, dataGroup_hi_lo_1847};
  wire [7:0]    dataGroup_55_28 = dataGroup_hi_1847[1479:1472];
  wire [2047:0] dataGroup_lo_1848 = {dataGroup_lo_hi_1848, dataGroup_lo_lo_1848};
  wire [2047:0] dataGroup_hi_1848 = {dataGroup_hi_hi_1848, dataGroup_hi_lo_1848};
  wire [7:0]    dataGroup_56_28 = dataGroup_hi_1848[1543:1536];
  wire [2047:0] dataGroup_lo_1849 = {dataGroup_lo_hi_1849, dataGroup_lo_lo_1849};
  wire [2047:0] dataGroup_hi_1849 = {dataGroup_hi_hi_1849, dataGroup_hi_lo_1849};
  wire [7:0]    dataGroup_57_28 = dataGroup_hi_1849[1607:1600];
  wire [2047:0] dataGroup_lo_1850 = {dataGroup_lo_hi_1850, dataGroup_lo_lo_1850};
  wire [2047:0] dataGroup_hi_1850 = {dataGroup_hi_hi_1850, dataGroup_hi_lo_1850};
  wire [7:0]    dataGroup_58_28 = dataGroup_hi_1850[1671:1664];
  wire [2047:0] dataGroup_lo_1851 = {dataGroup_lo_hi_1851, dataGroup_lo_lo_1851};
  wire [2047:0] dataGroup_hi_1851 = {dataGroup_hi_hi_1851, dataGroup_hi_lo_1851};
  wire [7:0]    dataGroup_59_28 = dataGroup_hi_1851[1735:1728];
  wire [2047:0] dataGroup_lo_1852 = {dataGroup_lo_hi_1852, dataGroup_lo_lo_1852};
  wire [2047:0] dataGroup_hi_1852 = {dataGroup_hi_hi_1852, dataGroup_hi_lo_1852};
  wire [7:0]    dataGroup_60_28 = dataGroup_hi_1852[1799:1792];
  wire [2047:0] dataGroup_lo_1853 = {dataGroup_lo_hi_1853, dataGroup_lo_lo_1853};
  wire [2047:0] dataGroup_hi_1853 = {dataGroup_hi_hi_1853, dataGroup_hi_lo_1853};
  wire [7:0]    dataGroup_61_28 = dataGroup_hi_1853[1863:1856];
  wire [2047:0] dataGroup_lo_1854 = {dataGroup_lo_hi_1854, dataGroup_lo_lo_1854};
  wire [2047:0] dataGroup_hi_1854 = {dataGroup_hi_hi_1854, dataGroup_hi_lo_1854};
  wire [7:0]    dataGroup_62_28 = dataGroup_hi_1854[1927:1920];
  wire [2047:0] dataGroup_lo_1855 = {dataGroup_lo_hi_1855, dataGroup_lo_lo_1855};
  wire [2047:0] dataGroup_hi_1855 = {dataGroup_hi_hi_1855, dataGroup_hi_lo_1855};
  wire [7:0]    dataGroup_63_28 = dataGroup_hi_1855[1991:1984];
  wire [15:0]   res_lo_lo_lo_lo_lo_28 = {dataGroup_1_28, dataGroup_0_28};
  wire [15:0]   res_lo_lo_lo_lo_hi_28 = {dataGroup_3_28, dataGroup_2_28};
  wire [31:0]   res_lo_lo_lo_lo_28 = {res_lo_lo_lo_lo_hi_28, res_lo_lo_lo_lo_lo_28};
  wire [15:0]   res_lo_lo_lo_hi_lo_28 = {dataGroup_5_28, dataGroup_4_28};
  wire [15:0]   res_lo_lo_lo_hi_hi_28 = {dataGroup_7_28, dataGroup_6_28};
  wire [31:0]   res_lo_lo_lo_hi_28 = {res_lo_lo_lo_hi_hi_28, res_lo_lo_lo_hi_lo_28};
  wire [63:0]   res_lo_lo_lo_28 = {res_lo_lo_lo_hi_28, res_lo_lo_lo_lo_28};
  wire [15:0]   res_lo_lo_hi_lo_lo_28 = {dataGroup_9_28, dataGroup_8_28};
  wire [15:0]   res_lo_lo_hi_lo_hi_28 = {dataGroup_11_28, dataGroup_10_28};
  wire [31:0]   res_lo_lo_hi_lo_28 = {res_lo_lo_hi_lo_hi_28, res_lo_lo_hi_lo_lo_28};
  wire [15:0]   res_lo_lo_hi_hi_lo_28 = {dataGroup_13_28, dataGroup_12_28};
  wire [15:0]   res_lo_lo_hi_hi_hi_28 = {dataGroup_15_28, dataGroup_14_28};
  wire [31:0]   res_lo_lo_hi_hi_28 = {res_lo_lo_hi_hi_hi_28, res_lo_lo_hi_hi_lo_28};
  wire [63:0]   res_lo_lo_hi_28 = {res_lo_lo_hi_hi_28, res_lo_lo_hi_lo_28};
  wire [127:0]  res_lo_lo_28 = {res_lo_lo_hi_28, res_lo_lo_lo_28};
  wire [15:0]   res_lo_hi_lo_lo_lo_28 = {dataGroup_17_28, dataGroup_16_28};
  wire [15:0]   res_lo_hi_lo_lo_hi_28 = {dataGroup_19_28, dataGroup_18_28};
  wire [31:0]   res_lo_hi_lo_lo_28 = {res_lo_hi_lo_lo_hi_28, res_lo_hi_lo_lo_lo_28};
  wire [15:0]   res_lo_hi_lo_hi_lo_28 = {dataGroup_21_28, dataGroup_20_28};
  wire [15:0]   res_lo_hi_lo_hi_hi_28 = {dataGroup_23_28, dataGroup_22_28};
  wire [31:0]   res_lo_hi_lo_hi_28 = {res_lo_hi_lo_hi_hi_28, res_lo_hi_lo_hi_lo_28};
  wire [63:0]   res_lo_hi_lo_28 = {res_lo_hi_lo_hi_28, res_lo_hi_lo_lo_28};
  wire [15:0]   res_lo_hi_hi_lo_lo_28 = {dataGroup_25_28, dataGroup_24_28};
  wire [15:0]   res_lo_hi_hi_lo_hi_28 = {dataGroup_27_28, dataGroup_26_28};
  wire [31:0]   res_lo_hi_hi_lo_28 = {res_lo_hi_hi_lo_hi_28, res_lo_hi_hi_lo_lo_28};
  wire [15:0]   res_lo_hi_hi_hi_lo_28 = {dataGroup_29_28, dataGroup_28_28};
  wire [15:0]   res_lo_hi_hi_hi_hi_28 = {dataGroup_31_28, dataGroup_30_28};
  wire [31:0]   res_lo_hi_hi_hi_28 = {res_lo_hi_hi_hi_hi_28, res_lo_hi_hi_hi_lo_28};
  wire [63:0]   res_lo_hi_hi_28 = {res_lo_hi_hi_hi_28, res_lo_hi_hi_lo_28};
  wire [127:0]  res_lo_hi_28 = {res_lo_hi_hi_28, res_lo_hi_lo_28};
  wire [255:0]  res_lo_28 = {res_lo_hi_28, res_lo_lo_28};
  wire [15:0]   res_hi_lo_lo_lo_lo_28 = {dataGroup_33_28, dataGroup_32_28};
  wire [15:0]   res_hi_lo_lo_lo_hi_28 = {dataGroup_35_28, dataGroup_34_28};
  wire [31:0]   res_hi_lo_lo_lo_28 = {res_hi_lo_lo_lo_hi_28, res_hi_lo_lo_lo_lo_28};
  wire [15:0]   res_hi_lo_lo_hi_lo_28 = {dataGroup_37_28, dataGroup_36_28};
  wire [15:0]   res_hi_lo_lo_hi_hi_28 = {dataGroup_39_28, dataGroup_38_28};
  wire [31:0]   res_hi_lo_lo_hi_28 = {res_hi_lo_lo_hi_hi_28, res_hi_lo_lo_hi_lo_28};
  wire [63:0]   res_hi_lo_lo_28 = {res_hi_lo_lo_hi_28, res_hi_lo_lo_lo_28};
  wire [15:0]   res_hi_lo_hi_lo_lo_28 = {dataGroup_41_28, dataGroup_40_28};
  wire [15:0]   res_hi_lo_hi_lo_hi_28 = {dataGroup_43_28, dataGroup_42_28};
  wire [31:0]   res_hi_lo_hi_lo_28 = {res_hi_lo_hi_lo_hi_28, res_hi_lo_hi_lo_lo_28};
  wire [15:0]   res_hi_lo_hi_hi_lo_28 = {dataGroup_45_28, dataGroup_44_28};
  wire [15:0]   res_hi_lo_hi_hi_hi_28 = {dataGroup_47_28, dataGroup_46_28};
  wire [31:0]   res_hi_lo_hi_hi_28 = {res_hi_lo_hi_hi_hi_28, res_hi_lo_hi_hi_lo_28};
  wire [63:0]   res_hi_lo_hi_28 = {res_hi_lo_hi_hi_28, res_hi_lo_hi_lo_28};
  wire [127:0]  res_hi_lo_28 = {res_hi_lo_hi_28, res_hi_lo_lo_28};
  wire [15:0]   res_hi_hi_lo_lo_lo_28 = {dataGroup_49_28, dataGroup_48_28};
  wire [15:0]   res_hi_hi_lo_lo_hi_28 = {dataGroup_51_28, dataGroup_50_28};
  wire [31:0]   res_hi_hi_lo_lo_28 = {res_hi_hi_lo_lo_hi_28, res_hi_hi_lo_lo_lo_28};
  wire [15:0]   res_hi_hi_lo_hi_lo_28 = {dataGroup_53_28, dataGroup_52_28};
  wire [15:0]   res_hi_hi_lo_hi_hi_28 = {dataGroup_55_28, dataGroup_54_28};
  wire [31:0]   res_hi_hi_lo_hi_28 = {res_hi_hi_lo_hi_hi_28, res_hi_hi_lo_hi_lo_28};
  wire [63:0]   res_hi_hi_lo_28 = {res_hi_hi_lo_hi_28, res_hi_hi_lo_lo_28};
  wire [15:0]   res_hi_hi_hi_lo_lo_28 = {dataGroup_57_28, dataGroup_56_28};
  wire [15:0]   res_hi_hi_hi_lo_hi_28 = {dataGroup_59_28, dataGroup_58_28};
  wire [31:0]   res_hi_hi_hi_lo_28 = {res_hi_hi_hi_lo_hi_28, res_hi_hi_hi_lo_lo_28};
  wire [15:0]   res_hi_hi_hi_hi_lo_28 = {dataGroup_61_28, dataGroup_60_28};
  wire [15:0]   res_hi_hi_hi_hi_hi_28 = {dataGroup_63_28, dataGroup_62_28};
  wire [31:0]   res_hi_hi_hi_hi_28 = {res_hi_hi_hi_hi_hi_28, res_hi_hi_hi_hi_lo_28};
  wire [63:0]   res_hi_hi_hi_28 = {res_hi_hi_hi_hi_28, res_hi_hi_hi_lo_28};
  wire [127:0]  res_hi_hi_28 = {res_hi_hi_hi_28, res_hi_hi_lo_28};
  wire [255:0]  res_hi_28 = {res_hi_hi_28, res_hi_lo_28};
  wire [511:0]  res_56 = {res_hi_28, res_lo_28};
  wire [2047:0] dataGroup_lo_1856 = {dataGroup_lo_hi_1856, dataGroup_lo_lo_1856};
  wire [2047:0] dataGroup_hi_1856 = {dataGroup_hi_hi_1856, dataGroup_hi_lo_1856};
  wire [7:0]    dataGroup_0_29 = dataGroup_lo_1856[15:8];
  wire [2047:0] dataGroup_lo_1857 = {dataGroup_lo_hi_1857, dataGroup_lo_lo_1857};
  wire [2047:0] dataGroup_hi_1857 = {dataGroup_hi_hi_1857, dataGroup_hi_lo_1857};
  wire [7:0]    dataGroup_1_29 = dataGroup_lo_1857[79:72];
  wire [2047:0] dataGroup_lo_1858 = {dataGroup_lo_hi_1858, dataGroup_lo_lo_1858};
  wire [2047:0] dataGroup_hi_1858 = {dataGroup_hi_hi_1858, dataGroup_hi_lo_1858};
  wire [7:0]    dataGroup_2_29 = dataGroup_lo_1858[143:136];
  wire [2047:0] dataGroup_lo_1859 = {dataGroup_lo_hi_1859, dataGroup_lo_lo_1859};
  wire [2047:0] dataGroup_hi_1859 = {dataGroup_hi_hi_1859, dataGroup_hi_lo_1859};
  wire [7:0]    dataGroup_3_29 = dataGroup_lo_1859[207:200];
  wire [2047:0] dataGroup_lo_1860 = {dataGroup_lo_hi_1860, dataGroup_lo_lo_1860};
  wire [2047:0] dataGroup_hi_1860 = {dataGroup_hi_hi_1860, dataGroup_hi_lo_1860};
  wire [7:0]    dataGroup_4_29 = dataGroup_lo_1860[271:264];
  wire [2047:0] dataGroup_lo_1861 = {dataGroup_lo_hi_1861, dataGroup_lo_lo_1861};
  wire [2047:0] dataGroup_hi_1861 = {dataGroup_hi_hi_1861, dataGroup_hi_lo_1861};
  wire [7:0]    dataGroup_5_29 = dataGroup_lo_1861[335:328];
  wire [2047:0] dataGroup_lo_1862 = {dataGroup_lo_hi_1862, dataGroup_lo_lo_1862};
  wire [2047:0] dataGroup_hi_1862 = {dataGroup_hi_hi_1862, dataGroup_hi_lo_1862};
  wire [7:0]    dataGroup_6_29 = dataGroup_lo_1862[399:392];
  wire [2047:0] dataGroup_lo_1863 = {dataGroup_lo_hi_1863, dataGroup_lo_lo_1863};
  wire [2047:0] dataGroup_hi_1863 = {dataGroup_hi_hi_1863, dataGroup_hi_lo_1863};
  wire [7:0]    dataGroup_7_29 = dataGroup_lo_1863[463:456];
  wire [2047:0] dataGroup_lo_1864 = {dataGroup_lo_hi_1864, dataGroup_lo_lo_1864};
  wire [2047:0] dataGroup_hi_1864 = {dataGroup_hi_hi_1864, dataGroup_hi_lo_1864};
  wire [7:0]    dataGroup_8_29 = dataGroup_lo_1864[527:520];
  wire [2047:0] dataGroup_lo_1865 = {dataGroup_lo_hi_1865, dataGroup_lo_lo_1865};
  wire [2047:0] dataGroup_hi_1865 = {dataGroup_hi_hi_1865, dataGroup_hi_lo_1865};
  wire [7:0]    dataGroup_9_29 = dataGroup_lo_1865[591:584];
  wire [2047:0] dataGroup_lo_1866 = {dataGroup_lo_hi_1866, dataGroup_lo_lo_1866};
  wire [2047:0] dataGroup_hi_1866 = {dataGroup_hi_hi_1866, dataGroup_hi_lo_1866};
  wire [7:0]    dataGroup_10_29 = dataGroup_lo_1866[655:648];
  wire [2047:0] dataGroup_lo_1867 = {dataGroup_lo_hi_1867, dataGroup_lo_lo_1867};
  wire [2047:0] dataGroup_hi_1867 = {dataGroup_hi_hi_1867, dataGroup_hi_lo_1867};
  wire [7:0]    dataGroup_11_29 = dataGroup_lo_1867[719:712];
  wire [2047:0] dataGroup_lo_1868 = {dataGroup_lo_hi_1868, dataGroup_lo_lo_1868};
  wire [2047:0] dataGroup_hi_1868 = {dataGroup_hi_hi_1868, dataGroup_hi_lo_1868};
  wire [7:0]    dataGroup_12_29 = dataGroup_lo_1868[783:776];
  wire [2047:0] dataGroup_lo_1869 = {dataGroup_lo_hi_1869, dataGroup_lo_lo_1869};
  wire [2047:0] dataGroup_hi_1869 = {dataGroup_hi_hi_1869, dataGroup_hi_lo_1869};
  wire [7:0]    dataGroup_13_29 = dataGroup_lo_1869[847:840];
  wire [2047:0] dataGroup_lo_1870 = {dataGroup_lo_hi_1870, dataGroup_lo_lo_1870};
  wire [2047:0] dataGroup_hi_1870 = {dataGroup_hi_hi_1870, dataGroup_hi_lo_1870};
  wire [7:0]    dataGroup_14_29 = dataGroup_lo_1870[911:904];
  wire [2047:0] dataGroup_lo_1871 = {dataGroup_lo_hi_1871, dataGroup_lo_lo_1871};
  wire [2047:0] dataGroup_hi_1871 = {dataGroup_hi_hi_1871, dataGroup_hi_lo_1871};
  wire [7:0]    dataGroup_15_29 = dataGroup_lo_1871[975:968];
  wire [2047:0] dataGroup_lo_1872 = {dataGroup_lo_hi_1872, dataGroup_lo_lo_1872};
  wire [2047:0] dataGroup_hi_1872 = {dataGroup_hi_hi_1872, dataGroup_hi_lo_1872};
  wire [7:0]    dataGroup_16_29 = dataGroup_lo_1872[1039:1032];
  wire [2047:0] dataGroup_lo_1873 = {dataGroup_lo_hi_1873, dataGroup_lo_lo_1873};
  wire [2047:0] dataGroup_hi_1873 = {dataGroup_hi_hi_1873, dataGroup_hi_lo_1873};
  wire [7:0]    dataGroup_17_29 = dataGroup_lo_1873[1103:1096];
  wire [2047:0] dataGroup_lo_1874 = {dataGroup_lo_hi_1874, dataGroup_lo_lo_1874};
  wire [2047:0] dataGroup_hi_1874 = {dataGroup_hi_hi_1874, dataGroup_hi_lo_1874};
  wire [7:0]    dataGroup_18_29 = dataGroup_lo_1874[1167:1160];
  wire [2047:0] dataGroup_lo_1875 = {dataGroup_lo_hi_1875, dataGroup_lo_lo_1875};
  wire [2047:0] dataGroup_hi_1875 = {dataGroup_hi_hi_1875, dataGroup_hi_lo_1875};
  wire [7:0]    dataGroup_19_29 = dataGroup_lo_1875[1231:1224];
  wire [2047:0] dataGroup_lo_1876 = {dataGroup_lo_hi_1876, dataGroup_lo_lo_1876};
  wire [2047:0] dataGroup_hi_1876 = {dataGroup_hi_hi_1876, dataGroup_hi_lo_1876};
  wire [7:0]    dataGroup_20_29 = dataGroup_lo_1876[1295:1288];
  wire [2047:0] dataGroup_lo_1877 = {dataGroup_lo_hi_1877, dataGroup_lo_lo_1877};
  wire [2047:0] dataGroup_hi_1877 = {dataGroup_hi_hi_1877, dataGroup_hi_lo_1877};
  wire [7:0]    dataGroup_21_29 = dataGroup_lo_1877[1359:1352];
  wire [2047:0] dataGroup_lo_1878 = {dataGroup_lo_hi_1878, dataGroup_lo_lo_1878};
  wire [2047:0] dataGroup_hi_1878 = {dataGroup_hi_hi_1878, dataGroup_hi_lo_1878};
  wire [7:0]    dataGroup_22_29 = dataGroup_lo_1878[1423:1416];
  wire [2047:0] dataGroup_lo_1879 = {dataGroup_lo_hi_1879, dataGroup_lo_lo_1879};
  wire [2047:0] dataGroup_hi_1879 = {dataGroup_hi_hi_1879, dataGroup_hi_lo_1879};
  wire [7:0]    dataGroup_23_29 = dataGroup_lo_1879[1487:1480];
  wire [2047:0] dataGroup_lo_1880 = {dataGroup_lo_hi_1880, dataGroup_lo_lo_1880};
  wire [2047:0] dataGroup_hi_1880 = {dataGroup_hi_hi_1880, dataGroup_hi_lo_1880};
  wire [7:0]    dataGroup_24_29 = dataGroup_lo_1880[1551:1544];
  wire [2047:0] dataGroup_lo_1881 = {dataGroup_lo_hi_1881, dataGroup_lo_lo_1881};
  wire [2047:0] dataGroup_hi_1881 = {dataGroup_hi_hi_1881, dataGroup_hi_lo_1881};
  wire [7:0]    dataGroup_25_29 = dataGroup_lo_1881[1615:1608];
  wire [2047:0] dataGroup_lo_1882 = {dataGroup_lo_hi_1882, dataGroup_lo_lo_1882};
  wire [2047:0] dataGroup_hi_1882 = {dataGroup_hi_hi_1882, dataGroup_hi_lo_1882};
  wire [7:0]    dataGroup_26_29 = dataGroup_lo_1882[1679:1672];
  wire [2047:0] dataGroup_lo_1883 = {dataGroup_lo_hi_1883, dataGroup_lo_lo_1883};
  wire [2047:0] dataGroup_hi_1883 = {dataGroup_hi_hi_1883, dataGroup_hi_lo_1883};
  wire [7:0]    dataGroup_27_29 = dataGroup_lo_1883[1743:1736];
  wire [2047:0] dataGroup_lo_1884 = {dataGroup_lo_hi_1884, dataGroup_lo_lo_1884};
  wire [2047:0] dataGroup_hi_1884 = {dataGroup_hi_hi_1884, dataGroup_hi_lo_1884};
  wire [7:0]    dataGroup_28_29 = dataGroup_lo_1884[1807:1800];
  wire [2047:0] dataGroup_lo_1885 = {dataGroup_lo_hi_1885, dataGroup_lo_lo_1885};
  wire [2047:0] dataGroup_hi_1885 = {dataGroup_hi_hi_1885, dataGroup_hi_lo_1885};
  wire [7:0]    dataGroup_29_29 = dataGroup_lo_1885[1871:1864];
  wire [2047:0] dataGroup_lo_1886 = {dataGroup_lo_hi_1886, dataGroup_lo_lo_1886};
  wire [2047:0] dataGroup_hi_1886 = {dataGroup_hi_hi_1886, dataGroup_hi_lo_1886};
  wire [7:0]    dataGroup_30_29 = dataGroup_lo_1886[1935:1928];
  wire [2047:0] dataGroup_lo_1887 = {dataGroup_lo_hi_1887, dataGroup_lo_lo_1887};
  wire [2047:0] dataGroup_hi_1887 = {dataGroup_hi_hi_1887, dataGroup_hi_lo_1887};
  wire [7:0]    dataGroup_31_29 = dataGroup_lo_1887[1999:1992];
  wire [2047:0] dataGroup_lo_1888 = {dataGroup_lo_hi_1888, dataGroup_lo_lo_1888};
  wire [2047:0] dataGroup_hi_1888 = {dataGroup_hi_hi_1888, dataGroup_hi_lo_1888};
  wire [7:0]    dataGroup_32_29 = dataGroup_hi_1888[15:8];
  wire [2047:0] dataGroup_lo_1889 = {dataGroup_lo_hi_1889, dataGroup_lo_lo_1889};
  wire [2047:0] dataGroup_hi_1889 = {dataGroup_hi_hi_1889, dataGroup_hi_lo_1889};
  wire [7:0]    dataGroup_33_29 = dataGroup_hi_1889[79:72];
  wire [2047:0] dataGroup_lo_1890 = {dataGroup_lo_hi_1890, dataGroup_lo_lo_1890};
  wire [2047:0] dataGroup_hi_1890 = {dataGroup_hi_hi_1890, dataGroup_hi_lo_1890};
  wire [7:0]    dataGroup_34_29 = dataGroup_hi_1890[143:136];
  wire [2047:0] dataGroup_lo_1891 = {dataGroup_lo_hi_1891, dataGroup_lo_lo_1891};
  wire [2047:0] dataGroup_hi_1891 = {dataGroup_hi_hi_1891, dataGroup_hi_lo_1891};
  wire [7:0]    dataGroup_35_29 = dataGroup_hi_1891[207:200];
  wire [2047:0] dataGroup_lo_1892 = {dataGroup_lo_hi_1892, dataGroup_lo_lo_1892};
  wire [2047:0] dataGroup_hi_1892 = {dataGroup_hi_hi_1892, dataGroup_hi_lo_1892};
  wire [7:0]    dataGroup_36_29 = dataGroup_hi_1892[271:264];
  wire [2047:0] dataGroup_lo_1893 = {dataGroup_lo_hi_1893, dataGroup_lo_lo_1893};
  wire [2047:0] dataGroup_hi_1893 = {dataGroup_hi_hi_1893, dataGroup_hi_lo_1893};
  wire [7:0]    dataGroup_37_29 = dataGroup_hi_1893[335:328];
  wire [2047:0] dataGroup_lo_1894 = {dataGroup_lo_hi_1894, dataGroup_lo_lo_1894};
  wire [2047:0] dataGroup_hi_1894 = {dataGroup_hi_hi_1894, dataGroup_hi_lo_1894};
  wire [7:0]    dataGroup_38_29 = dataGroup_hi_1894[399:392];
  wire [2047:0] dataGroup_lo_1895 = {dataGroup_lo_hi_1895, dataGroup_lo_lo_1895};
  wire [2047:0] dataGroup_hi_1895 = {dataGroup_hi_hi_1895, dataGroup_hi_lo_1895};
  wire [7:0]    dataGroup_39_29 = dataGroup_hi_1895[463:456];
  wire [2047:0] dataGroup_lo_1896 = {dataGroup_lo_hi_1896, dataGroup_lo_lo_1896};
  wire [2047:0] dataGroup_hi_1896 = {dataGroup_hi_hi_1896, dataGroup_hi_lo_1896};
  wire [7:0]    dataGroup_40_29 = dataGroup_hi_1896[527:520];
  wire [2047:0] dataGroup_lo_1897 = {dataGroup_lo_hi_1897, dataGroup_lo_lo_1897};
  wire [2047:0] dataGroup_hi_1897 = {dataGroup_hi_hi_1897, dataGroup_hi_lo_1897};
  wire [7:0]    dataGroup_41_29 = dataGroup_hi_1897[591:584];
  wire [2047:0] dataGroup_lo_1898 = {dataGroup_lo_hi_1898, dataGroup_lo_lo_1898};
  wire [2047:0] dataGroup_hi_1898 = {dataGroup_hi_hi_1898, dataGroup_hi_lo_1898};
  wire [7:0]    dataGroup_42_29 = dataGroup_hi_1898[655:648];
  wire [2047:0] dataGroup_lo_1899 = {dataGroup_lo_hi_1899, dataGroup_lo_lo_1899};
  wire [2047:0] dataGroup_hi_1899 = {dataGroup_hi_hi_1899, dataGroup_hi_lo_1899};
  wire [7:0]    dataGroup_43_29 = dataGroup_hi_1899[719:712];
  wire [2047:0] dataGroup_lo_1900 = {dataGroup_lo_hi_1900, dataGroup_lo_lo_1900};
  wire [2047:0] dataGroup_hi_1900 = {dataGroup_hi_hi_1900, dataGroup_hi_lo_1900};
  wire [7:0]    dataGroup_44_29 = dataGroup_hi_1900[783:776];
  wire [2047:0] dataGroup_lo_1901 = {dataGroup_lo_hi_1901, dataGroup_lo_lo_1901};
  wire [2047:0] dataGroup_hi_1901 = {dataGroup_hi_hi_1901, dataGroup_hi_lo_1901};
  wire [7:0]    dataGroup_45_29 = dataGroup_hi_1901[847:840];
  wire [2047:0] dataGroup_lo_1902 = {dataGroup_lo_hi_1902, dataGroup_lo_lo_1902};
  wire [2047:0] dataGroup_hi_1902 = {dataGroup_hi_hi_1902, dataGroup_hi_lo_1902};
  wire [7:0]    dataGroup_46_29 = dataGroup_hi_1902[911:904];
  wire [2047:0] dataGroup_lo_1903 = {dataGroup_lo_hi_1903, dataGroup_lo_lo_1903};
  wire [2047:0] dataGroup_hi_1903 = {dataGroup_hi_hi_1903, dataGroup_hi_lo_1903};
  wire [7:0]    dataGroup_47_29 = dataGroup_hi_1903[975:968];
  wire [2047:0] dataGroup_lo_1904 = {dataGroup_lo_hi_1904, dataGroup_lo_lo_1904};
  wire [2047:0] dataGroup_hi_1904 = {dataGroup_hi_hi_1904, dataGroup_hi_lo_1904};
  wire [7:0]    dataGroup_48_29 = dataGroup_hi_1904[1039:1032];
  wire [2047:0] dataGroup_lo_1905 = {dataGroup_lo_hi_1905, dataGroup_lo_lo_1905};
  wire [2047:0] dataGroup_hi_1905 = {dataGroup_hi_hi_1905, dataGroup_hi_lo_1905};
  wire [7:0]    dataGroup_49_29 = dataGroup_hi_1905[1103:1096];
  wire [2047:0] dataGroup_lo_1906 = {dataGroup_lo_hi_1906, dataGroup_lo_lo_1906};
  wire [2047:0] dataGroup_hi_1906 = {dataGroup_hi_hi_1906, dataGroup_hi_lo_1906};
  wire [7:0]    dataGroup_50_29 = dataGroup_hi_1906[1167:1160];
  wire [2047:0] dataGroup_lo_1907 = {dataGroup_lo_hi_1907, dataGroup_lo_lo_1907};
  wire [2047:0] dataGroup_hi_1907 = {dataGroup_hi_hi_1907, dataGroup_hi_lo_1907};
  wire [7:0]    dataGroup_51_29 = dataGroup_hi_1907[1231:1224];
  wire [2047:0] dataGroup_lo_1908 = {dataGroup_lo_hi_1908, dataGroup_lo_lo_1908};
  wire [2047:0] dataGroup_hi_1908 = {dataGroup_hi_hi_1908, dataGroup_hi_lo_1908};
  wire [7:0]    dataGroup_52_29 = dataGroup_hi_1908[1295:1288];
  wire [2047:0] dataGroup_lo_1909 = {dataGroup_lo_hi_1909, dataGroup_lo_lo_1909};
  wire [2047:0] dataGroup_hi_1909 = {dataGroup_hi_hi_1909, dataGroup_hi_lo_1909};
  wire [7:0]    dataGroup_53_29 = dataGroup_hi_1909[1359:1352];
  wire [2047:0] dataGroup_lo_1910 = {dataGroup_lo_hi_1910, dataGroup_lo_lo_1910};
  wire [2047:0] dataGroup_hi_1910 = {dataGroup_hi_hi_1910, dataGroup_hi_lo_1910};
  wire [7:0]    dataGroup_54_29 = dataGroup_hi_1910[1423:1416];
  wire [2047:0] dataGroup_lo_1911 = {dataGroup_lo_hi_1911, dataGroup_lo_lo_1911};
  wire [2047:0] dataGroup_hi_1911 = {dataGroup_hi_hi_1911, dataGroup_hi_lo_1911};
  wire [7:0]    dataGroup_55_29 = dataGroup_hi_1911[1487:1480];
  wire [2047:0] dataGroup_lo_1912 = {dataGroup_lo_hi_1912, dataGroup_lo_lo_1912};
  wire [2047:0] dataGroup_hi_1912 = {dataGroup_hi_hi_1912, dataGroup_hi_lo_1912};
  wire [7:0]    dataGroup_56_29 = dataGroup_hi_1912[1551:1544];
  wire [2047:0] dataGroup_lo_1913 = {dataGroup_lo_hi_1913, dataGroup_lo_lo_1913};
  wire [2047:0] dataGroup_hi_1913 = {dataGroup_hi_hi_1913, dataGroup_hi_lo_1913};
  wire [7:0]    dataGroup_57_29 = dataGroup_hi_1913[1615:1608];
  wire [2047:0] dataGroup_lo_1914 = {dataGroup_lo_hi_1914, dataGroup_lo_lo_1914};
  wire [2047:0] dataGroup_hi_1914 = {dataGroup_hi_hi_1914, dataGroup_hi_lo_1914};
  wire [7:0]    dataGroup_58_29 = dataGroup_hi_1914[1679:1672];
  wire [2047:0] dataGroup_lo_1915 = {dataGroup_lo_hi_1915, dataGroup_lo_lo_1915};
  wire [2047:0] dataGroup_hi_1915 = {dataGroup_hi_hi_1915, dataGroup_hi_lo_1915};
  wire [7:0]    dataGroup_59_29 = dataGroup_hi_1915[1743:1736];
  wire [2047:0] dataGroup_lo_1916 = {dataGroup_lo_hi_1916, dataGroup_lo_lo_1916};
  wire [2047:0] dataGroup_hi_1916 = {dataGroup_hi_hi_1916, dataGroup_hi_lo_1916};
  wire [7:0]    dataGroup_60_29 = dataGroup_hi_1916[1807:1800];
  wire [2047:0] dataGroup_lo_1917 = {dataGroup_lo_hi_1917, dataGroup_lo_lo_1917};
  wire [2047:0] dataGroup_hi_1917 = {dataGroup_hi_hi_1917, dataGroup_hi_lo_1917};
  wire [7:0]    dataGroup_61_29 = dataGroup_hi_1917[1871:1864];
  wire [2047:0] dataGroup_lo_1918 = {dataGroup_lo_hi_1918, dataGroup_lo_lo_1918};
  wire [2047:0] dataGroup_hi_1918 = {dataGroup_hi_hi_1918, dataGroup_hi_lo_1918};
  wire [7:0]    dataGroup_62_29 = dataGroup_hi_1918[1935:1928];
  wire [2047:0] dataGroup_lo_1919 = {dataGroup_lo_hi_1919, dataGroup_lo_lo_1919};
  wire [2047:0] dataGroup_hi_1919 = {dataGroup_hi_hi_1919, dataGroup_hi_lo_1919};
  wire [7:0]    dataGroup_63_29 = dataGroup_hi_1919[1999:1992];
  wire [15:0]   res_lo_lo_lo_lo_lo_29 = {dataGroup_1_29, dataGroup_0_29};
  wire [15:0]   res_lo_lo_lo_lo_hi_29 = {dataGroup_3_29, dataGroup_2_29};
  wire [31:0]   res_lo_lo_lo_lo_29 = {res_lo_lo_lo_lo_hi_29, res_lo_lo_lo_lo_lo_29};
  wire [15:0]   res_lo_lo_lo_hi_lo_29 = {dataGroup_5_29, dataGroup_4_29};
  wire [15:0]   res_lo_lo_lo_hi_hi_29 = {dataGroup_7_29, dataGroup_6_29};
  wire [31:0]   res_lo_lo_lo_hi_29 = {res_lo_lo_lo_hi_hi_29, res_lo_lo_lo_hi_lo_29};
  wire [63:0]   res_lo_lo_lo_29 = {res_lo_lo_lo_hi_29, res_lo_lo_lo_lo_29};
  wire [15:0]   res_lo_lo_hi_lo_lo_29 = {dataGroup_9_29, dataGroup_8_29};
  wire [15:0]   res_lo_lo_hi_lo_hi_29 = {dataGroup_11_29, dataGroup_10_29};
  wire [31:0]   res_lo_lo_hi_lo_29 = {res_lo_lo_hi_lo_hi_29, res_lo_lo_hi_lo_lo_29};
  wire [15:0]   res_lo_lo_hi_hi_lo_29 = {dataGroup_13_29, dataGroup_12_29};
  wire [15:0]   res_lo_lo_hi_hi_hi_29 = {dataGroup_15_29, dataGroup_14_29};
  wire [31:0]   res_lo_lo_hi_hi_29 = {res_lo_lo_hi_hi_hi_29, res_lo_lo_hi_hi_lo_29};
  wire [63:0]   res_lo_lo_hi_29 = {res_lo_lo_hi_hi_29, res_lo_lo_hi_lo_29};
  wire [127:0]  res_lo_lo_29 = {res_lo_lo_hi_29, res_lo_lo_lo_29};
  wire [15:0]   res_lo_hi_lo_lo_lo_29 = {dataGroup_17_29, dataGroup_16_29};
  wire [15:0]   res_lo_hi_lo_lo_hi_29 = {dataGroup_19_29, dataGroup_18_29};
  wire [31:0]   res_lo_hi_lo_lo_29 = {res_lo_hi_lo_lo_hi_29, res_lo_hi_lo_lo_lo_29};
  wire [15:0]   res_lo_hi_lo_hi_lo_29 = {dataGroup_21_29, dataGroup_20_29};
  wire [15:0]   res_lo_hi_lo_hi_hi_29 = {dataGroup_23_29, dataGroup_22_29};
  wire [31:0]   res_lo_hi_lo_hi_29 = {res_lo_hi_lo_hi_hi_29, res_lo_hi_lo_hi_lo_29};
  wire [63:0]   res_lo_hi_lo_29 = {res_lo_hi_lo_hi_29, res_lo_hi_lo_lo_29};
  wire [15:0]   res_lo_hi_hi_lo_lo_29 = {dataGroup_25_29, dataGroup_24_29};
  wire [15:0]   res_lo_hi_hi_lo_hi_29 = {dataGroup_27_29, dataGroup_26_29};
  wire [31:0]   res_lo_hi_hi_lo_29 = {res_lo_hi_hi_lo_hi_29, res_lo_hi_hi_lo_lo_29};
  wire [15:0]   res_lo_hi_hi_hi_lo_29 = {dataGroup_29_29, dataGroup_28_29};
  wire [15:0]   res_lo_hi_hi_hi_hi_29 = {dataGroup_31_29, dataGroup_30_29};
  wire [31:0]   res_lo_hi_hi_hi_29 = {res_lo_hi_hi_hi_hi_29, res_lo_hi_hi_hi_lo_29};
  wire [63:0]   res_lo_hi_hi_29 = {res_lo_hi_hi_hi_29, res_lo_hi_hi_lo_29};
  wire [127:0]  res_lo_hi_29 = {res_lo_hi_hi_29, res_lo_hi_lo_29};
  wire [255:0]  res_lo_29 = {res_lo_hi_29, res_lo_lo_29};
  wire [15:0]   res_hi_lo_lo_lo_lo_29 = {dataGroup_33_29, dataGroup_32_29};
  wire [15:0]   res_hi_lo_lo_lo_hi_29 = {dataGroup_35_29, dataGroup_34_29};
  wire [31:0]   res_hi_lo_lo_lo_29 = {res_hi_lo_lo_lo_hi_29, res_hi_lo_lo_lo_lo_29};
  wire [15:0]   res_hi_lo_lo_hi_lo_29 = {dataGroup_37_29, dataGroup_36_29};
  wire [15:0]   res_hi_lo_lo_hi_hi_29 = {dataGroup_39_29, dataGroup_38_29};
  wire [31:0]   res_hi_lo_lo_hi_29 = {res_hi_lo_lo_hi_hi_29, res_hi_lo_lo_hi_lo_29};
  wire [63:0]   res_hi_lo_lo_29 = {res_hi_lo_lo_hi_29, res_hi_lo_lo_lo_29};
  wire [15:0]   res_hi_lo_hi_lo_lo_29 = {dataGroup_41_29, dataGroup_40_29};
  wire [15:0]   res_hi_lo_hi_lo_hi_29 = {dataGroup_43_29, dataGroup_42_29};
  wire [31:0]   res_hi_lo_hi_lo_29 = {res_hi_lo_hi_lo_hi_29, res_hi_lo_hi_lo_lo_29};
  wire [15:0]   res_hi_lo_hi_hi_lo_29 = {dataGroup_45_29, dataGroup_44_29};
  wire [15:0]   res_hi_lo_hi_hi_hi_29 = {dataGroup_47_29, dataGroup_46_29};
  wire [31:0]   res_hi_lo_hi_hi_29 = {res_hi_lo_hi_hi_hi_29, res_hi_lo_hi_hi_lo_29};
  wire [63:0]   res_hi_lo_hi_29 = {res_hi_lo_hi_hi_29, res_hi_lo_hi_lo_29};
  wire [127:0]  res_hi_lo_29 = {res_hi_lo_hi_29, res_hi_lo_lo_29};
  wire [15:0]   res_hi_hi_lo_lo_lo_29 = {dataGroup_49_29, dataGroup_48_29};
  wire [15:0]   res_hi_hi_lo_lo_hi_29 = {dataGroup_51_29, dataGroup_50_29};
  wire [31:0]   res_hi_hi_lo_lo_29 = {res_hi_hi_lo_lo_hi_29, res_hi_hi_lo_lo_lo_29};
  wire [15:0]   res_hi_hi_lo_hi_lo_29 = {dataGroup_53_29, dataGroup_52_29};
  wire [15:0]   res_hi_hi_lo_hi_hi_29 = {dataGroup_55_29, dataGroup_54_29};
  wire [31:0]   res_hi_hi_lo_hi_29 = {res_hi_hi_lo_hi_hi_29, res_hi_hi_lo_hi_lo_29};
  wire [63:0]   res_hi_hi_lo_29 = {res_hi_hi_lo_hi_29, res_hi_hi_lo_lo_29};
  wire [15:0]   res_hi_hi_hi_lo_lo_29 = {dataGroup_57_29, dataGroup_56_29};
  wire [15:0]   res_hi_hi_hi_lo_hi_29 = {dataGroup_59_29, dataGroup_58_29};
  wire [31:0]   res_hi_hi_hi_lo_29 = {res_hi_hi_hi_lo_hi_29, res_hi_hi_hi_lo_lo_29};
  wire [15:0]   res_hi_hi_hi_hi_lo_29 = {dataGroup_61_29, dataGroup_60_29};
  wire [15:0]   res_hi_hi_hi_hi_hi_29 = {dataGroup_63_29, dataGroup_62_29};
  wire [31:0]   res_hi_hi_hi_hi_29 = {res_hi_hi_hi_hi_hi_29, res_hi_hi_hi_hi_lo_29};
  wire [63:0]   res_hi_hi_hi_29 = {res_hi_hi_hi_hi_29, res_hi_hi_hi_lo_29};
  wire [127:0]  res_hi_hi_29 = {res_hi_hi_hi_29, res_hi_hi_lo_29};
  wire [255:0]  res_hi_29 = {res_hi_hi_29, res_hi_lo_29};
  wire [511:0]  res_57 = {res_hi_29, res_lo_29};
  wire [2047:0] dataGroup_lo_1920 = {dataGroup_lo_hi_1920, dataGroup_lo_lo_1920};
  wire [2047:0] dataGroup_hi_1920 = {dataGroup_hi_hi_1920, dataGroup_hi_lo_1920};
  wire [7:0]    dataGroup_0_30 = dataGroup_lo_1920[23:16];
  wire [2047:0] dataGroup_lo_1921 = {dataGroup_lo_hi_1921, dataGroup_lo_lo_1921};
  wire [2047:0] dataGroup_hi_1921 = {dataGroup_hi_hi_1921, dataGroup_hi_lo_1921};
  wire [7:0]    dataGroup_1_30 = dataGroup_lo_1921[87:80];
  wire [2047:0] dataGroup_lo_1922 = {dataGroup_lo_hi_1922, dataGroup_lo_lo_1922};
  wire [2047:0] dataGroup_hi_1922 = {dataGroup_hi_hi_1922, dataGroup_hi_lo_1922};
  wire [7:0]    dataGroup_2_30 = dataGroup_lo_1922[151:144];
  wire [2047:0] dataGroup_lo_1923 = {dataGroup_lo_hi_1923, dataGroup_lo_lo_1923};
  wire [2047:0] dataGroup_hi_1923 = {dataGroup_hi_hi_1923, dataGroup_hi_lo_1923};
  wire [7:0]    dataGroup_3_30 = dataGroup_lo_1923[215:208];
  wire [2047:0] dataGroup_lo_1924 = {dataGroup_lo_hi_1924, dataGroup_lo_lo_1924};
  wire [2047:0] dataGroup_hi_1924 = {dataGroup_hi_hi_1924, dataGroup_hi_lo_1924};
  wire [7:0]    dataGroup_4_30 = dataGroup_lo_1924[279:272];
  wire [2047:0] dataGroup_lo_1925 = {dataGroup_lo_hi_1925, dataGroup_lo_lo_1925};
  wire [2047:0] dataGroup_hi_1925 = {dataGroup_hi_hi_1925, dataGroup_hi_lo_1925};
  wire [7:0]    dataGroup_5_30 = dataGroup_lo_1925[343:336];
  wire [2047:0] dataGroup_lo_1926 = {dataGroup_lo_hi_1926, dataGroup_lo_lo_1926};
  wire [2047:0] dataGroup_hi_1926 = {dataGroup_hi_hi_1926, dataGroup_hi_lo_1926};
  wire [7:0]    dataGroup_6_30 = dataGroup_lo_1926[407:400];
  wire [2047:0] dataGroup_lo_1927 = {dataGroup_lo_hi_1927, dataGroup_lo_lo_1927};
  wire [2047:0] dataGroup_hi_1927 = {dataGroup_hi_hi_1927, dataGroup_hi_lo_1927};
  wire [7:0]    dataGroup_7_30 = dataGroup_lo_1927[471:464];
  wire [2047:0] dataGroup_lo_1928 = {dataGroup_lo_hi_1928, dataGroup_lo_lo_1928};
  wire [2047:0] dataGroup_hi_1928 = {dataGroup_hi_hi_1928, dataGroup_hi_lo_1928};
  wire [7:0]    dataGroup_8_30 = dataGroup_lo_1928[535:528];
  wire [2047:0] dataGroup_lo_1929 = {dataGroup_lo_hi_1929, dataGroup_lo_lo_1929};
  wire [2047:0] dataGroup_hi_1929 = {dataGroup_hi_hi_1929, dataGroup_hi_lo_1929};
  wire [7:0]    dataGroup_9_30 = dataGroup_lo_1929[599:592];
  wire [2047:0] dataGroup_lo_1930 = {dataGroup_lo_hi_1930, dataGroup_lo_lo_1930};
  wire [2047:0] dataGroup_hi_1930 = {dataGroup_hi_hi_1930, dataGroup_hi_lo_1930};
  wire [7:0]    dataGroup_10_30 = dataGroup_lo_1930[663:656];
  wire [2047:0] dataGroup_lo_1931 = {dataGroup_lo_hi_1931, dataGroup_lo_lo_1931};
  wire [2047:0] dataGroup_hi_1931 = {dataGroup_hi_hi_1931, dataGroup_hi_lo_1931};
  wire [7:0]    dataGroup_11_30 = dataGroup_lo_1931[727:720];
  wire [2047:0] dataGroup_lo_1932 = {dataGroup_lo_hi_1932, dataGroup_lo_lo_1932};
  wire [2047:0] dataGroup_hi_1932 = {dataGroup_hi_hi_1932, dataGroup_hi_lo_1932};
  wire [7:0]    dataGroup_12_30 = dataGroup_lo_1932[791:784];
  wire [2047:0] dataGroup_lo_1933 = {dataGroup_lo_hi_1933, dataGroup_lo_lo_1933};
  wire [2047:0] dataGroup_hi_1933 = {dataGroup_hi_hi_1933, dataGroup_hi_lo_1933};
  wire [7:0]    dataGroup_13_30 = dataGroup_lo_1933[855:848];
  wire [2047:0] dataGroup_lo_1934 = {dataGroup_lo_hi_1934, dataGroup_lo_lo_1934};
  wire [2047:0] dataGroup_hi_1934 = {dataGroup_hi_hi_1934, dataGroup_hi_lo_1934};
  wire [7:0]    dataGroup_14_30 = dataGroup_lo_1934[919:912];
  wire [2047:0] dataGroup_lo_1935 = {dataGroup_lo_hi_1935, dataGroup_lo_lo_1935};
  wire [2047:0] dataGroup_hi_1935 = {dataGroup_hi_hi_1935, dataGroup_hi_lo_1935};
  wire [7:0]    dataGroup_15_30 = dataGroup_lo_1935[983:976];
  wire [2047:0] dataGroup_lo_1936 = {dataGroup_lo_hi_1936, dataGroup_lo_lo_1936};
  wire [2047:0] dataGroup_hi_1936 = {dataGroup_hi_hi_1936, dataGroup_hi_lo_1936};
  wire [7:0]    dataGroup_16_30 = dataGroup_lo_1936[1047:1040];
  wire [2047:0] dataGroup_lo_1937 = {dataGroup_lo_hi_1937, dataGroup_lo_lo_1937};
  wire [2047:0] dataGroup_hi_1937 = {dataGroup_hi_hi_1937, dataGroup_hi_lo_1937};
  wire [7:0]    dataGroup_17_30 = dataGroup_lo_1937[1111:1104];
  wire [2047:0] dataGroup_lo_1938 = {dataGroup_lo_hi_1938, dataGroup_lo_lo_1938};
  wire [2047:0] dataGroup_hi_1938 = {dataGroup_hi_hi_1938, dataGroup_hi_lo_1938};
  wire [7:0]    dataGroup_18_30 = dataGroup_lo_1938[1175:1168];
  wire [2047:0] dataGroup_lo_1939 = {dataGroup_lo_hi_1939, dataGroup_lo_lo_1939};
  wire [2047:0] dataGroup_hi_1939 = {dataGroup_hi_hi_1939, dataGroup_hi_lo_1939};
  wire [7:0]    dataGroup_19_30 = dataGroup_lo_1939[1239:1232];
  wire [2047:0] dataGroup_lo_1940 = {dataGroup_lo_hi_1940, dataGroup_lo_lo_1940};
  wire [2047:0] dataGroup_hi_1940 = {dataGroup_hi_hi_1940, dataGroup_hi_lo_1940};
  wire [7:0]    dataGroup_20_30 = dataGroup_lo_1940[1303:1296];
  wire [2047:0] dataGroup_lo_1941 = {dataGroup_lo_hi_1941, dataGroup_lo_lo_1941};
  wire [2047:0] dataGroup_hi_1941 = {dataGroup_hi_hi_1941, dataGroup_hi_lo_1941};
  wire [7:0]    dataGroup_21_30 = dataGroup_lo_1941[1367:1360];
  wire [2047:0] dataGroup_lo_1942 = {dataGroup_lo_hi_1942, dataGroup_lo_lo_1942};
  wire [2047:0] dataGroup_hi_1942 = {dataGroup_hi_hi_1942, dataGroup_hi_lo_1942};
  wire [7:0]    dataGroup_22_30 = dataGroup_lo_1942[1431:1424];
  wire [2047:0] dataGroup_lo_1943 = {dataGroup_lo_hi_1943, dataGroup_lo_lo_1943};
  wire [2047:0] dataGroup_hi_1943 = {dataGroup_hi_hi_1943, dataGroup_hi_lo_1943};
  wire [7:0]    dataGroup_23_30 = dataGroup_lo_1943[1495:1488];
  wire [2047:0] dataGroup_lo_1944 = {dataGroup_lo_hi_1944, dataGroup_lo_lo_1944};
  wire [2047:0] dataGroup_hi_1944 = {dataGroup_hi_hi_1944, dataGroup_hi_lo_1944};
  wire [7:0]    dataGroup_24_30 = dataGroup_lo_1944[1559:1552];
  wire [2047:0] dataGroup_lo_1945 = {dataGroup_lo_hi_1945, dataGroup_lo_lo_1945};
  wire [2047:0] dataGroup_hi_1945 = {dataGroup_hi_hi_1945, dataGroup_hi_lo_1945};
  wire [7:0]    dataGroup_25_30 = dataGroup_lo_1945[1623:1616];
  wire [2047:0] dataGroup_lo_1946 = {dataGroup_lo_hi_1946, dataGroup_lo_lo_1946};
  wire [2047:0] dataGroup_hi_1946 = {dataGroup_hi_hi_1946, dataGroup_hi_lo_1946};
  wire [7:0]    dataGroup_26_30 = dataGroup_lo_1946[1687:1680];
  wire [2047:0] dataGroup_lo_1947 = {dataGroup_lo_hi_1947, dataGroup_lo_lo_1947};
  wire [2047:0] dataGroup_hi_1947 = {dataGroup_hi_hi_1947, dataGroup_hi_lo_1947};
  wire [7:0]    dataGroup_27_30 = dataGroup_lo_1947[1751:1744];
  wire [2047:0] dataGroup_lo_1948 = {dataGroup_lo_hi_1948, dataGroup_lo_lo_1948};
  wire [2047:0] dataGroup_hi_1948 = {dataGroup_hi_hi_1948, dataGroup_hi_lo_1948};
  wire [7:0]    dataGroup_28_30 = dataGroup_lo_1948[1815:1808];
  wire [2047:0] dataGroup_lo_1949 = {dataGroup_lo_hi_1949, dataGroup_lo_lo_1949};
  wire [2047:0] dataGroup_hi_1949 = {dataGroup_hi_hi_1949, dataGroup_hi_lo_1949};
  wire [7:0]    dataGroup_29_30 = dataGroup_lo_1949[1879:1872];
  wire [2047:0] dataGroup_lo_1950 = {dataGroup_lo_hi_1950, dataGroup_lo_lo_1950};
  wire [2047:0] dataGroup_hi_1950 = {dataGroup_hi_hi_1950, dataGroup_hi_lo_1950};
  wire [7:0]    dataGroup_30_30 = dataGroup_lo_1950[1943:1936];
  wire [2047:0] dataGroup_lo_1951 = {dataGroup_lo_hi_1951, dataGroup_lo_lo_1951};
  wire [2047:0] dataGroup_hi_1951 = {dataGroup_hi_hi_1951, dataGroup_hi_lo_1951};
  wire [7:0]    dataGroup_31_30 = dataGroup_lo_1951[2007:2000];
  wire [2047:0] dataGroup_lo_1952 = {dataGroup_lo_hi_1952, dataGroup_lo_lo_1952};
  wire [2047:0] dataGroup_hi_1952 = {dataGroup_hi_hi_1952, dataGroup_hi_lo_1952};
  wire [7:0]    dataGroup_32_30 = dataGroup_hi_1952[23:16];
  wire [2047:0] dataGroup_lo_1953 = {dataGroup_lo_hi_1953, dataGroup_lo_lo_1953};
  wire [2047:0] dataGroup_hi_1953 = {dataGroup_hi_hi_1953, dataGroup_hi_lo_1953};
  wire [7:0]    dataGroup_33_30 = dataGroup_hi_1953[87:80];
  wire [2047:0] dataGroup_lo_1954 = {dataGroup_lo_hi_1954, dataGroup_lo_lo_1954};
  wire [2047:0] dataGroup_hi_1954 = {dataGroup_hi_hi_1954, dataGroup_hi_lo_1954};
  wire [7:0]    dataGroup_34_30 = dataGroup_hi_1954[151:144];
  wire [2047:0] dataGroup_lo_1955 = {dataGroup_lo_hi_1955, dataGroup_lo_lo_1955};
  wire [2047:0] dataGroup_hi_1955 = {dataGroup_hi_hi_1955, dataGroup_hi_lo_1955};
  wire [7:0]    dataGroup_35_30 = dataGroup_hi_1955[215:208];
  wire [2047:0] dataGroup_lo_1956 = {dataGroup_lo_hi_1956, dataGroup_lo_lo_1956};
  wire [2047:0] dataGroup_hi_1956 = {dataGroup_hi_hi_1956, dataGroup_hi_lo_1956};
  wire [7:0]    dataGroup_36_30 = dataGroup_hi_1956[279:272];
  wire [2047:0] dataGroup_lo_1957 = {dataGroup_lo_hi_1957, dataGroup_lo_lo_1957};
  wire [2047:0] dataGroup_hi_1957 = {dataGroup_hi_hi_1957, dataGroup_hi_lo_1957};
  wire [7:0]    dataGroup_37_30 = dataGroup_hi_1957[343:336];
  wire [2047:0] dataGroup_lo_1958 = {dataGroup_lo_hi_1958, dataGroup_lo_lo_1958};
  wire [2047:0] dataGroup_hi_1958 = {dataGroup_hi_hi_1958, dataGroup_hi_lo_1958};
  wire [7:0]    dataGroup_38_30 = dataGroup_hi_1958[407:400];
  wire [2047:0] dataGroup_lo_1959 = {dataGroup_lo_hi_1959, dataGroup_lo_lo_1959};
  wire [2047:0] dataGroup_hi_1959 = {dataGroup_hi_hi_1959, dataGroup_hi_lo_1959};
  wire [7:0]    dataGroup_39_30 = dataGroup_hi_1959[471:464];
  wire [2047:0] dataGroup_lo_1960 = {dataGroup_lo_hi_1960, dataGroup_lo_lo_1960};
  wire [2047:0] dataGroup_hi_1960 = {dataGroup_hi_hi_1960, dataGroup_hi_lo_1960};
  wire [7:0]    dataGroup_40_30 = dataGroup_hi_1960[535:528];
  wire [2047:0] dataGroup_lo_1961 = {dataGroup_lo_hi_1961, dataGroup_lo_lo_1961};
  wire [2047:0] dataGroup_hi_1961 = {dataGroup_hi_hi_1961, dataGroup_hi_lo_1961};
  wire [7:0]    dataGroup_41_30 = dataGroup_hi_1961[599:592];
  wire [2047:0] dataGroup_lo_1962 = {dataGroup_lo_hi_1962, dataGroup_lo_lo_1962};
  wire [2047:0] dataGroup_hi_1962 = {dataGroup_hi_hi_1962, dataGroup_hi_lo_1962};
  wire [7:0]    dataGroup_42_30 = dataGroup_hi_1962[663:656];
  wire [2047:0] dataGroup_lo_1963 = {dataGroup_lo_hi_1963, dataGroup_lo_lo_1963};
  wire [2047:0] dataGroup_hi_1963 = {dataGroup_hi_hi_1963, dataGroup_hi_lo_1963};
  wire [7:0]    dataGroup_43_30 = dataGroup_hi_1963[727:720];
  wire [2047:0] dataGroup_lo_1964 = {dataGroup_lo_hi_1964, dataGroup_lo_lo_1964};
  wire [2047:0] dataGroup_hi_1964 = {dataGroup_hi_hi_1964, dataGroup_hi_lo_1964};
  wire [7:0]    dataGroup_44_30 = dataGroup_hi_1964[791:784];
  wire [2047:0] dataGroup_lo_1965 = {dataGroup_lo_hi_1965, dataGroup_lo_lo_1965};
  wire [2047:0] dataGroup_hi_1965 = {dataGroup_hi_hi_1965, dataGroup_hi_lo_1965};
  wire [7:0]    dataGroup_45_30 = dataGroup_hi_1965[855:848];
  wire [2047:0] dataGroup_lo_1966 = {dataGroup_lo_hi_1966, dataGroup_lo_lo_1966};
  wire [2047:0] dataGroup_hi_1966 = {dataGroup_hi_hi_1966, dataGroup_hi_lo_1966};
  wire [7:0]    dataGroup_46_30 = dataGroup_hi_1966[919:912];
  wire [2047:0] dataGroup_lo_1967 = {dataGroup_lo_hi_1967, dataGroup_lo_lo_1967};
  wire [2047:0] dataGroup_hi_1967 = {dataGroup_hi_hi_1967, dataGroup_hi_lo_1967};
  wire [7:0]    dataGroup_47_30 = dataGroup_hi_1967[983:976];
  wire [2047:0] dataGroup_lo_1968 = {dataGroup_lo_hi_1968, dataGroup_lo_lo_1968};
  wire [2047:0] dataGroup_hi_1968 = {dataGroup_hi_hi_1968, dataGroup_hi_lo_1968};
  wire [7:0]    dataGroup_48_30 = dataGroup_hi_1968[1047:1040];
  wire [2047:0] dataGroup_lo_1969 = {dataGroup_lo_hi_1969, dataGroup_lo_lo_1969};
  wire [2047:0] dataGroup_hi_1969 = {dataGroup_hi_hi_1969, dataGroup_hi_lo_1969};
  wire [7:0]    dataGroup_49_30 = dataGroup_hi_1969[1111:1104];
  wire [2047:0] dataGroup_lo_1970 = {dataGroup_lo_hi_1970, dataGroup_lo_lo_1970};
  wire [2047:0] dataGroup_hi_1970 = {dataGroup_hi_hi_1970, dataGroup_hi_lo_1970};
  wire [7:0]    dataGroup_50_30 = dataGroup_hi_1970[1175:1168];
  wire [2047:0] dataGroup_lo_1971 = {dataGroup_lo_hi_1971, dataGroup_lo_lo_1971};
  wire [2047:0] dataGroup_hi_1971 = {dataGroup_hi_hi_1971, dataGroup_hi_lo_1971};
  wire [7:0]    dataGroup_51_30 = dataGroup_hi_1971[1239:1232];
  wire [2047:0] dataGroup_lo_1972 = {dataGroup_lo_hi_1972, dataGroup_lo_lo_1972};
  wire [2047:0] dataGroup_hi_1972 = {dataGroup_hi_hi_1972, dataGroup_hi_lo_1972};
  wire [7:0]    dataGroup_52_30 = dataGroup_hi_1972[1303:1296];
  wire [2047:0] dataGroup_lo_1973 = {dataGroup_lo_hi_1973, dataGroup_lo_lo_1973};
  wire [2047:0] dataGroup_hi_1973 = {dataGroup_hi_hi_1973, dataGroup_hi_lo_1973};
  wire [7:0]    dataGroup_53_30 = dataGroup_hi_1973[1367:1360];
  wire [2047:0] dataGroup_lo_1974 = {dataGroup_lo_hi_1974, dataGroup_lo_lo_1974};
  wire [2047:0] dataGroup_hi_1974 = {dataGroup_hi_hi_1974, dataGroup_hi_lo_1974};
  wire [7:0]    dataGroup_54_30 = dataGroup_hi_1974[1431:1424];
  wire [2047:0] dataGroup_lo_1975 = {dataGroup_lo_hi_1975, dataGroup_lo_lo_1975};
  wire [2047:0] dataGroup_hi_1975 = {dataGroup_hi_hi_1975, dataGroup_hi_lo_1975};
  wire [7:0]    dataGroup_55_30 = dataGroup_hi_1975[1495:1488];
  wire [2047:0] dataGroup_lo_1976 = {dataGroup_lo_hi_1976, dataGroup_lo_lo_1976};
  wire [2047:0] dataGroup_hi_1976 = {dataGroup_hi_hi_1976, dataGroup_hi_lo_1976};
  wire [7:0]    dataGroup_56_30 = dataGroup_hi_1976[1559:1552];
  wire [2047:0] dataGroup_lo_1977 = {dataGroup_lo_hi_1977, dataGroup_lo_lo_1977};
  wire [2047:0] dataGroup_hi_1977 = {dataGroup_hi_hi_1977, dataGroup_hi_lo_1977};
  wire [7:0]    dataGroup_57_30 = dataGroup_hi_1977[1623:1616];
  wire [2047:0] dataGroup_lo_1978 = {dataGroup_lo_hi_1978, dataGroup_lo_lo_1978};
  wire [2047:0] dataGroup_hi_1978 = {dataGroup_hi_hi_1978, dataGroup_hi_lo_1978};
  wire [7:0]    dataGroup_58_30 = dataGroup_hi_1978[1687:1680];
  wire [2047:0] dataGroup_lo_1979 = {dataGroup_lo_hi_1979, dataGroup_lo_lo_1979};
  wire [2047:0] dataGroup_hi_1979 = {dataGroup_hi_hi_1979, dataGroup_hi_lo_1979};
  wire [7:0]    dataGroup_59_30 = dataGroup_hi_1979[1751:1744];
  wire [2047:0] dataGroup_lo_1980 = {dataGroup_lo_hi_1980, dataGroup_lo_lo_1980};
  wire [2047:0] dataGroup_hi_1980 = {dataGroup_hi_hi_1980, dataGroup_hi_lo_1980};
  wire [7:0]    dataGroup_60_30 = dataGroup_hi_1980[1815:1808];
  wire [2047:0] dataGroup_lo_1981 = {dataGroup_lo_hi_1981, dataGroup_lo_lo_1981};
  wire [2047:0] dataGroup_hi_1981 = {dataGroup_hi_hi_1981, dataGroup_hi_lo_1981};
  wire [7:0]    dataGroup_61_30 = dataGroup_hi_1981[1879:1872];
  wire [2047:0] dataGroup_lo_1982 = {dataGroup_lo_hi_1982, dataGroup_lo_lo_1982};
  wire [2047:0] dataGroup_hi_1982 = {dataGroup_hi_hi_1982, dataGroup_hi_lo_1982};
  wire [7:0]    dataGroup_62_30 = dataGroup_hi_1982[1943:1936];
  wire [2047:0] dataGroup_lo_1983 = {dataGroup_lo_hi_1983, dataGroup_lo_lo_1983};
  wire [2047:0] dataGroup_hi_1983 = {dataGroup_hi_hi_1983, dataGroup_hi_lo_1983};
  wire [7:0]    dataGroup_63_30 = dataGroup_hi_1983[2007:2000];
  wire [15:0]   res_lo_lo_lo_lo_lo_30 = {dataGroup_1_30, dataGroup_0_30};
  wire [15:0]   res_lo_lo_lo_lo_hi_30 = {dataGroup_3_30, dataGroup_2_30};
  wire [31:0]   res_lo_lo_lo_lo_30 = {res_lo_lo_lo_lo_hi_30, res_lo_lo_lo_lo_lo_30};
  wire [15:0]   res_lo_lo_lo_hi_lo_30 = {dataGroup_5_30, dataGroup_4_30};
  wire [15:0]   res_lo_lo_lo_hi_hi_30 = {dataGroup_7_30, dataGroup_6_30};
  wire [31:0]   res_lo_lo_lo_hi_30 = {res_lo_lo_lo_hi_hi_30, res_lo_lo_lo_hi_lo_30};
  wire [63:0]   res_lo_lo_lo_30 = {res_lo_lo_lo_hi_30, res_lo_lo_lo_lo_30};
  wire [15:0]   res_lo_lo_hi_lo_lo_30 = {dataGroup_9_30, dataGroup_8_30};
  wire [15:0]   res_lo_lo_hi_lo_hi_30 = {dataGroup_11_30, dataGroup_10_30};
  wire [31:0]   res_lo_lo_hi_lo_30 = {res_lo_lo_hi_lo_hi_30, res_lo_lo_hi_lo_lo_30};
  wire [15:0]   res_lo_lo_hi_hi_lo_30 = {dataGroup_13_30, dataGroup_12_30};
  wire [15:0]   res_lo_lo_hi_hi_hi_30 = {dataGroup_15_30, dataGroup_14_30};
  wire [31:0]   res_lo_lo_hi_hi_30 = {res_lo_lo_hi_hi_hi_30, res_lo_lo_hi_hi_lo_30};
  wire [63:0]   res_lo_lo_hi_30 = {res_lo_lo_hi_hi_30, res_lo_lo_hi_lo_30};
  wire [127:0]  res_lo_lo_30 = {res_lo_lo_hi_30, res_lo_lo_lo_30};
  wire [15:0]   res_lo_hi_lo_lo_lo_30 = {dataGroup_17_30, dataGroup_16_30};
  wire [15:0]   res_lo_hi_lo_lo_hi_30 = {dataGroup_19_30, dataGroup_18_30};
  wire [31:0]   res_lo_hi_lo_lo_30 = {res_lo_hi_lo_lo_hi_30, res_lo_hi_lo_lo_lo_30};
  wire [15:0]   res_lo_hi_lo_hi_lo_30 = {dataGroup_21_30, dataGroup_20_30};
  wire [15:0]   res_lo_hi_lo_hi_hi_30 = {dataGroup_23_30, dataGroup_22_30};
  wire [31:0]   res_lo_hi_lo_hi_30 = {res_lo_hi_lo_hi_hi_30, res_lo_hi_lo_hi_lo_30};
  wire [63:0]   res_lo_hi_lo_30 = {res_lo_hi_lo_hi_30, res_lo_hi_lo_lo_30};
  wire [15:0]   res_lo_hi_hi_lo_lo_30 = {dataGroup_25_30, dataGroup_24_30};
  wire [15:0]   res_lo_hi_hi_lo_hi_30 = {dataGroup_27_30, dataGroup_26_30};
  wire [31:0]   res_lo_hi_hi_lo_30 = {res_lo_hi_hi_lo_hi_30, res_lo_hi_hi_lo_lo_30};
  wire [15:0]   res_lo_hi_hi_hi_lo_30 = {dataGroup_29_30, dataGroup_28_30};
  wire [15:0]   res_lo_hi_hi_hi_hi_30 = {dataGroup_31_30, dataGroup_30_30};
  wire [31:0]   res_lo_hi_hi_hi_30 = {res_lo_hi_hi_hi_hi_30, res_lo_hi_hi_hi_lo_30};
  wire [63:0]   res_lo_hi_hi_30 = {res_lo_hi_hi_hi_30, res_lo_hi_hi_lo_30};
  wire [127:0]  res_lo_hi_30 = {res_lo_hi_hi_30, res_lo_hi_lo_30};
  wire [255:0]  res_lo_30 = {res_lo_hi_30, res_lo_lo_30};
  wire [15:0]   res_hi_lo_lo_lo_lo_30 = {dataGroup_33_30, dataGroup_32_30};
  wire [15:0]   res_hi_lo_lo_lo_hi_30 = {dataGroup_35_30, dataGroup_34_30};
  wire [31:0]   res_hi_lo_lo_lo_30 = {res_hi_lo_lo_lo_hi_30, res_hi_lo_lo_lo_lo_30};
  wire [15:0]   res_hi_lo_lo_hi_lo_30 = {dataGroup_37_30, dataGroup_36_30};
  wire [15:0]   res_hi_lo_lo_hi_hi_30 = {dataGroup_39_30, dataGroup_38_30};
  wire [31:0]   res_hi_lo_lo_hi_30 = {res_hi_lo_lo_hi_hi_30, res_hi_lo_lo_hi_lo_30};
  wire [63:0]   res_hi_lo_lo_30 = {res_hi_lo_lo_hi_30, res_hi_lo_lo_lo_30};
  wire [15:0]   res_hi_lo_hi_lo_lo_30 = {dataGroup_41_30, dataGroup_40_30};
  wire [15:0]   res_hi_lo_hi_lo_hi_30 = {dataGroup_43_30, dataGroup_42_30};
  wire [31:0]   res_hi_lo_hi_lo_30 = {res_hi_lo_hi_lo_hi_30, res_hi_lo_hi_lo_lo_30};
  wire [15:0]   res_hi_lo_hi_hi_lo_30 = {dataGroup_45_30, dataGroup_44_30};
  wire [15:0]   res_hi_lo_hi_hi_hi_30 = {dataGroup_47_30, dataGroup_46_30};
  wire [31:0]   res_hi_lo_hi_hi_30 = {res_hi_lo_hi_hi_hi_30, res_hi_lo_hi_hi_lo_30};
  wire [63:0]   res_hi_lo_hi_30 = {res_hi_lo_hi_hi_30, res_hi_lo_hi_lo_30};
  wire [127:0]  res_hi_lo_30 = {res_hi_lo_hi_30, res_hi_lo_lo_30};
  wire [15:0]   res_hi_hi_lo_lo_lo_30 = {dataGroup_49_30, dataGroup_48_30};
  wire [15:0]   res_hi_hi_lo_lo_hi_30 = {dataGroup_51_30, dataGroup_50_30};
  wire [31:0]   res_hi_hi_lo_lo_30 = {res_hi_hi_lo_lo_hi_30, res_hi_hi_lo_lo_lo_30};
  wire [15:0]   res_hi_hi_lo_hi_lo_30 = {dataGroup_53_30, dataGroup_52_30};
  wire [15:0]   res_hi_hi_lo_hi_hi_30 = {dataGroup_55_30, dataGroup_54_30};
  wire [31:0]   res_hi_hi_lo_hi_30 = {res_hi_hi_lo_hi_hi_30, res_hi_hi_lo_hi_lo_30};
  wire [63:0]   res_hi_hi_lo_30 = {res_hi_hi_lo_hi_30, res_hi_hi_lo_lo_30};
  wire [15:0]   res_hi_hi_hi_lo_lo_30 = {dataGroup_57_30, dataGroup_56_30};
  wire [15:0]   res_hi_hi_hi_lo_hi_30 = {dataGroup_59_30, dataGroup_58_30};
  wire [31:0]   res_hi_hi_hi_lo_30 = {res_hi_hi_hi_lo_hi_30, res_hi_hi_hi_lo_lo_30};
  wire [15:0]   res_hi_hi_hi_hi_lo_30 = {dataGroup_61_30, dataGroup_60_30};
  wire [15:0]   res_hi_hi_hi_hi_hi_30 = {dataGroup_63_30, dataGroup_62_30};
  wire [31:0]   res_hi_hi_hi_hi_30 = {res_hi_hi_hi_hi_hi_30, res_hi_hi_hi_hi_lo_30};
  wire [63:0]   res_hi_hi_hi_30 = {res_hi_hi_hi_hi_30, res_hi_hi_hi_lo_30};
  wire [127:0]  res_hi_hi_30 = {res_hi_hi_hi_30, res_hi_hi_lo_30};
  wire [255:0]  res_hi_30 = {res_hi_hi_30, res_hi_lo_30};
  wire [511:0]  res_58 = {res_hi_30, res_lo_30};
  wire [2047:0] dataGroup_lo_1984 = {dataGroup_lo_hi_1984, dataGroup_lo_lo_1984};
  wire [2047:0] dataGroup_hi_1984 = {dataGroup_hi_hi_1984, dataGroup_hi_lo_1984};
  wire [7:0]    dataGroup_0_31 = dataGroup_lo_1984[31:24];
  wire [2047:0] dataGroup_lo_1985 = {dataGroup_lo_hi_1985, dataGroup_lo_lo_1985};
  wire [2047:0] dataGroup_hi_1985 = {dataGroup_hi_hi_1985, dataGroup_hi_lo_1985};
  wire [7:0]    dataGroup_1_31 = dataGroup_lo_1985[95:88];
  wire [2047:0] dataGroup_lo_1986 = {dataGroup_lo_hi_1986, dataGroup_lo_lo_1986};
  wire [2047:0] dataGroup_hi_1986 = {dataGroup_hi_hi_1986, dataGroup_hi_lo_1986};
  wire [7:0]    dataGroup_2_31 = dataGroup_lo_1986[159:152];
  wire [2047:0] dataGroup_lo_1987 = {dataGroup_lo_hi_1987, dataGroup_lo_lo_1987};
  wire [2047:0] dataGroup_hi_1987 = {dataGroup_hi_hi_1987, dataGroup_hi_lo_1987};
  wire [7:0]    dataGroup_3_31 = dataGroup_lo_1987[223:216];
  wire [2047:0] dataGroup_lo_1988 = {dataGroup_lo_hi_1988, dataGroup_lo_lo_1988};
  wire [2047:0] dataGroup_hi_1988 = {dataGroup_hi_hi_1988, dataGroup_hi_lo_1988};
  wire [7:0]    dataGroup_4_31 = dataGroup_lo_1988[287:280];
  wire [2047:0] dataGroup_lo_1989 = {dataGroup_lo_hi_1989, dataGroup_lo_lo_1989};
  wire [2047:0] dataGroup_hi_1989 = {dataGroup_hi_hi_1989, dataGroup_hi_lo_1989};
  wire [7:0]    dataGroup_5_31 = dataGroup_lo_1989[351:344];
  wire [2047:0] dataGroup_lo_1990 = {dataGroup_lo_hi_1990, dataGroup_lo_lo_1990};
  wire [2047:0] dataGroup_hi_1990 = {dataGroup_hi_hi_1990, dataGroup_hi_lo_1990};
  wire [7:0]    dataGroup_6_31 = dataGroup_lo_1990[415:408];
  wire [2047:0] dataGroup_lo_1991 = {dataGroup_lo_hi_1991, dataGroup_lo_lo_1991};
  wire [2047:0] dataGroup_hi_1991 = {dataGroup_hi_hi_1991, dataGroup_hi_lo_1991};
  wire [7:0]    dataGroup_7_31 = dataGroup_lo_1991[479:472];
  wire [2047:0] dataGroup_lo_1992 = {dataGroup_lo_hi_1992, dataGroup_lo_lo_1992};
  wire [2047:0] dataGroup_hi_1992 = {dataGroup_hi_hi_1992, dataGroup_hi_lo_1992};
  wire [7:0]    dataGroup_8_31 = dataGroup_lo_1992[543:536];
  wire [2047:0] dataGroup_lo_1993 = {dataGroup_lo_hi_1993, dataGroup_lo_lo_1993};
  wire [2047:0] dataGroup_hi_1993 = {dataGroup_hi_hi_1993, dataGroup_hi_lo_1993};
  wire [7:0]    dataGroup_9_31 = dataGroup_lo_1993[607:600];
  wire [2047:0] dataGroup_lo_1994 = {dataGroup_lo_hi_1994, dataGroup_lo_lo_1994};
  wire [2047:0] dataGroup_hi_1994 = {dataGroup_hi_hi_1994, dataGroup_hi_lo_1994};
  wire [7:0]    dataGroup_10_31 = dataGroup_lo_1994[671:664];
  wire [2047:0] dataGroup_lo_1995 = {dataGroup_lo_hi_1995, dataGroup_lo_lo_1995};
  wire [2047:0] dataGroup_hi_1995 = {dataGroup_hi_hi_1995, dataGroup_hi_lo_1995};
  wire [7:0]    dataGroup_11_31 = dataGroup_lo_1995[735:728];
  wire [2047:0] dataGroup_lo_1996 = {dataGroup_lo_hi_1996, dataGroup_lo_lo_1996};
  wire [2047:0] dataGroup_hi_1996 = {dataGroup_hi_hi_1996, dataGroup_hi_lo_1996};
  wire [7:0]    dataGroup_12_31 = dataGroup_lo_1996[799:792];
  wire [2047:0] dataGroup_lo_1997 = {dataGroup_lo_hi_1997, dataGroup_lo_lo_1997};
  wire [2047:0] dataGroup_hi_1997 = {dataGroup_hi_hi_1997, dataGroup_hi_lo_1997};
  wire [7:0]    dataGroup_13_31 = dataGroup_lo_1997[863:856];
  wire [2047:0] dataGroup_lo_1998 = {dataGroup_lo_hi_1998, dataGroup_lo_lo_1998};
  wire [2047:0] dataGroup_hi_1998 = {dataGroup_hi_hi_1998, dataGroup_hi_lo_1998};
  wire [7:0]    dataGroup_14_31 = dataGroup_lo_1998[927:920];
  wire [2047:0] dataGroup_lo_1999 = {dataGroup_lo_hi_1999, dataGroup_lo_lo_1999};
  wire [2047:0] dataGroup_hi_1999 = {dataGroup_hi_hi_1999, dataGroup_hi_lo_1999};
  wire [7:0]    dataGroup_15_31 = dataGroup_lo_1999[991:984];
  wire [2047:0] dataGroup_lo_2000 = {dataGroup_lo_hi_2000, dataGroup_lo_lo_2000};
  wire [2047:0] dataGroup_hi_2000 = {dataGroup_hi_hi_2000, dataGroup_hi_lo_2000};
  wire [7:0]    dataGroup_16_31 = dataGroup_lo_2000[1055:1048];
  wire [2047:0] dataGroup_lo_2001 = {dataGroup_lo_hi_2001, dataGroup_lo_lo_2001};
  wire [2047:0] dataGroup_hi_2001 = {dataGroup_hi_hi_2001, dataGroup_hi_lo_2001};
  wire [7:0]    dataGroup_17_31 = dataGroup_lo_2001[1119:1112];
  wire [2047:0] dataGroup_lo_2002 = {dataGroup_lo_hi_2002, dataGroup_lo_lo_2002};
  wire [2047:0] dataGroup_hi_2002 = {dataGroup_hi_hi_2002, dataGroup_hi_lo_2002};
  wire [7:0]    dataGroup_18_31 = dataGroup_lo_2002[1183:1176];
  wire [2047:0] dataGroup_lo_2003 = {dataGroup_lo_hi_2003, dataGroup_lo_lo_2003};
  wire [2047:0] dataGroup_hi_2003 = {dataGroup_hi_hi_2003, dataGroup_hi_lo_2003};
  wire [7:0]    dataGroup_19_31 = dataGroup_lo_2003[1247:1240];
  wire [2047:0] dataGroup_lo_2004 = {dataGroup_lo_hi_2004, dataGroup_lo_lo_2004};
  wire [2047:0] dataGroup_hi_2004 = {dataGroup_hi_hi_2004, dataGroup_hi_lo_2004};
  wire [7:0]    dataGroup_20_31 = dataGroup_lo_2004[1311:1304];
  wire [2047:0] dataGroup_lo_2005 = {dataGroup_lo_hi_2005, dataGroup_lo_lo_2005};
  wire [2047:0] dataGroup_hi_2005 = {dataGroup_hi_hi_2005, dataGroup_hi_lo_2005};
  wire [7:0]    dataGroup_21_31 = dataGroup_lo_2005[1375:1368];
  wire [2047:0] dataGroup_lo_2006 = {dataGroup_lo_hi_2006, dataGroup_lo_lo_2006};
  wire [2047:0] dataGroup_hi_2006 = {dataGroup_hi_hi_2006, dataGroup_hi_lo_2006};
  wire [7:0]    dataGroup_22_31 = dataGroup_lo_2006[1439:1432];
  wire [2047:0] dataGroup_lo_2007 = {dataGroup_lo_hi_2007, dataGroup_lo_lo_2007};
  wire [2047:0] dataGroup_hi_2007 = {dataGroup_hi_hi_2007, dataGroup_hi_lo_2007};
  wire [7:0]    dataGroup_23_31 = dataGroup_lo_2007[1503:1496];
  wire [2047:0] dataGroup_lo_2008 = {dataGroup_lo_hi_2008, dataGroup_lo_lo_2008};
  wire [2047:0] dataGroup_hi_2008 = {dataGroup_hi_hi_2008, dataGroup_hi_lo_2008};
  wire [7:0]    dataGroup_24_31 = dataGroup_lo_2008[1567:1560];
  wire [2047:0] dataGroup_lo_2009 = {dataGroup_lo_hi_2009, dataGroup_lo_lo_2009};
  wire [2047:0] dataGroup_hi_2009 = {dataGroup_hi_hi_2009, dataGroup_hi_lo_2009};
  wire [7:0]    dataGroup_25_31 = dataGroup_lo_2009[1631:1624];
  wire [2047:0] dataGroup_lo_2010 = {dataGroup_lo_hi_2010, dataGroup_lo_lo_2010};
  wire [2047:0] dataGroup_hi_2010 = {dataGroup_hi_hi_2010, dataGroup_hi_lo_2010};
  wire [7:0]    dataGroup_26_31 = dataGroup_lo_2010[1695:1688];
  wire [2047:0] dataGroup_lo_2011 = {dataGroup_lo_hi_2011, dataGroup_lo_lo_2011};
  wire [2047:0] dataGroup_hi_2011 = {dataGroup_hi_hi_2011, dataGroup_hi_lo_2011};
  wire [7:0]    dataGroup_27_31 = dataGroup_lo_2011[1759:1752];
  wire [2047:0] dataGroup_lo_2012 = {dataGroup_lo_hi_2012, dataGroup_lo_lo_2012};
  wire [2047:0] dataGroup_hi_2012 = {dataGroup_hi_hi_2012, dataGroup_hi_lo_2012};
  wire [7:0]    dataGroup_28_31 = dataGroup_lo_2012[1823:1816];
  wire [2047:0] dataGroup_lo_2013 = {dataGroup_lo_hi_2013, dataGroup_lo_lo_2013};
  wire [2047:0] dataGroup_hi_2013 = {dataGroup_hi_hi_2013, dataGroup_hi_lo_2013};
  wire [7:0]    dataGroup_29_31 = dataGroup_lo_2013[1887:1880];
  wire [2047:0] dataGroup_lo_2014 = {dataGroup_lo_hi_2014, dataGroup_lo_lo_2014};
  wire [2047:0] dataGroup_hi_2014 = {dataGroup_hi_hi_2014, dataGroup_hi_lo_2014};
  wire [7:0]    dataGroup_30_31 = dataGroup_lo_2014[1951:1944];
  wire [2047:0] dataGroup_lo_2015 = {dataGroup_lo_hi_2015, dataGroup_lo_lo_2015};
  wire [2047:0] dataGroup_hi_2015 = {dataGroup_hi_hi_2015, dataGroup_hi_lo_2015};
  wire [7:0]    dataGroup_31_31 = dataGroup_lo_2015[2015:2008];
  wire [2047:0] dataGroup_lo_2016 = {dataGroup_lo_hi_2016, dataGroup_lo_lo_2016};
  wire [2047:0] dataGroup_hi_2016 = {dataGroup_hi_hi_2016, dataGroup_hi_lo_2016};
  wire [7:0]    dataGroup_32_31 = dataGroup_hi_2016[31:24];
  wire [2047:0] dataGroup_lo_2017 = {dataGroup_lo_hi_2017, dataGroup_lo_lo_2017};
  wire [2047:0] dataGroup_hi_2017 = {dataGroup_hi_hi_2017, dataGroup_hi_lo_2017};
  wire [7:0]    dataGroup_33_31 = dataGroup_hi_2017[95:88];
  wire [2047:0] dataGroup_lo_2018 = {dataGroup_lo_hi_2018, dataGroup_lo_lo_2018};
  wire [2047:0] dataGroup_hi_2018 = {dataGroup_hi_hi_2018, dataGroup_hi_lo_2018};
  wire [7:0]    dataGroup_34_31 = dataGroup_hi_2018[159:152];
  wire [2047:0] dataGroup_lo_2019 = {dataGroup_lo_hi_2019, dataGroup_lo_lo_2019};
  wire [2047:0] dataGroup_hi_2019 = {dataGroup_hi_hi_2019, dataGroup_hi_lo_2019};
  wire [7:0]    dataGroup_35_31 = dataGroup_hi_2019[223:216];
  wire [2047:0] dataGroup_lo_2020 = {dataGroup_lo_hi_2020, dataGroup_lo_lo_2020};
  wire [2047:0] dataGroup_hi_2020 = {dataGroup_hi_hi_2020, dataGroup_hi_lo_2020};
  wire [7:0]    dataGroup_36_31 = dataGroup_hi_2020[287:280];
  wire [2047:0] dataGroup_lo_2021 = {dataGroup_lo_hi_2021, dataGroup_lo_lo_2021};
  wire [2047:0] dataGroup_hi_2021 = {dataGroup_hi_hi_2021, dataGroup_hi_lo_2021};
  wire [7:0]    dataGroup_37_31 = dataGroup_hi_2021[351:344];
  wire [2047:0] dataGroup_lo_2022 = {dataGroup_lo_hi_2022, dataGroup_lo_lo_2022};
  wire [2047:0] dataGroup_hi_2022 = {dataGroup_hi_hi_2022, dataGroup_hi_lo_2022};
  wire [7:0]    dataGroup_38_31 = dataGroup_hi_2022[415:408];
  wire [2047:0] dataGroup_lo_2023 = {dataGroup_lo_hi_2023, dataGroup_lo_lo_2023};
  wire [2047:0] dataGroup_hi_2023 = {dataGroup_hi_hi_2023, dataGroup_hi_lo_2023};
  wire [7:0]    dataGroup_39_31 = dataGroup_hi_2023[479:472];
  wire [2047:0] dataGroup_lo_2024 = {dataGroup_lo_hi_2024, dataGroup_lo_lo_2024};
  wire [2047:0] dataGroup_hi_2024 = {dataGroup_hi_hi_2024, dataGroup_hi_lo_2024};
  wire [7:0]    dataGroup_40_31 = dataGroup_hi_2024[543:536];
  wire [2047:0] dataGroup_lo_2025 = {dataGroup_lo_hi_2025, dataGroup_lo_lo_2025};
  wire [2047:0] dataGroup_hi_2025 = {dataGroup_hi_hi_2025, dataGroup_hi_lo_2025};
  wire [7:0]    dataGroup_41_31 = dataGroup_hi_2025[607:600];
  wire [2047:0] dataGroup_lo_2026 = {dataGroup_lo_hi_2026, dataGroup_lo_lo_2026};
  wire [2047:0] dataGroup_hi_2026 = {dataGroup_hi_hi_2026, dataGroup_hi_lo_2026};
  wire [7:0]    dataGroup_42_31 = dataGroup_hi_2026[671:664];
  wire [2047:0] dataGroup_lo_2027 = {dataGroup_lo_hi_2027, dataGroup_lo_lo_2027};
  wire [2047:0] dataGroup_hi_2027 = {dataGroup_hi_hi_2027, dataGroup_hi_lo_2027};
  wire [7:0]    dataGroup_43_31 = dataGroup_hi_2027[735:728];
  wire [2047:0] dataGroup_lo_2028 = {dataGroup_lo_hi_2028, dataGroup_lo_lo_2028};
  wire [2047:0] dataGroup_hi_2028 = {dataGroup_hi_hi_2028, dataGroup_hi_lo_2028};
  wire [7:0]    dataGroup_44_31 = dataGroup_hi_2028[799:792];
  wire [2047:0] dataGroup_lo_2029 = {dataGroup_lo_hi_2029, dataGroup_lo_lo_2029};
  wire [2047:0] dataGroup_hi_2029 = {dataGroup_hi_hi_2029, dataGroup_hi_lo_2029};
  wire [7:0]    dataGroup_45_31 = dataGroup_hi_2029[863:856];
  wire [2047:0] dataGroup_lo_2030 = {dataGroup_lo_hi_2030, dataGroup_lo_lo_2030};
  wire [2047:0] dataGroup_hi_2030 = {dataGroup_hi_hi_2030, dataGroup_hi_lo_2030};
  wire [7:0]    dataGroup_46_31 = dataGroup_hi_2030[927:920];
  wire [2047:0] dataGroup_lo_2031 = {dataGroup_lo_hi_2031, dataGroup_lo_lo_2031};
  wire [2047:0] dataGroup_hi_2031 = {dataGroup_hi_hi_2031, dataGroup_hi_lo_2031};
  wire [7:0]    dataGroup_47_31 = dataGroup_hi_2031[991:984];
  wire [2047:0] dataGroup_lo_2032 = {dataGroup_lo_hi_2032, dataGroup_lo_lo_2032};
  wire [2047:0] dataGroup_hi_2032 = {dataGroup_hi_hi_2032, dataGroup_hi_lo_2032};
  wire [7:0]    dataGroup_48_31 = dataGroup_hi_2032[1055:1048];
  wire [2047:0] dataGroup_lo_2033 = {dataGroup_lo_hi_2033, dataGroup_lo_lo_2033};
  wire [2047:0] dataGroup_hi_2033 = {dataGroup_hi_hi_2033, dataGroup_hi_lo_2033};
  wire [7:0]    dataGroup_49_31 = dataGroup_hi_2033[1119:1112];
  wire [2047:0] dataGroup_lo_2034 = {dataGroup_lo_hi_2034, dataGroup_lo_lo_2034};
  wire [2047:0] dataGroup_hi_2034 = {dataGroup_hi_hi_2034, dataGroup_hi_lo_2034};
  wire [7:0]    dataGroup_50_31 = dataGroup_hi_2034[1183:1176];
  wire [2047:0] dataGroup_lo_2035 = {dataGroup_lo_hi_2035, dataGroup_lo_lo_2035};
  wire [2047:0] dataGroup_hi_2035 = {dataGroup_hi_hi_2035, dataGroup_hi_lo_2035};
  wire [7:0]    dataGroup_51_31 = dataGroup_hi_2035[1247:1240];
  wire [2047:0] dataGroup_lo_2036 = {dataGroup_lo_hi_2036, dataGroup_lo_lo_2036};
  wire [2047:0] dataGroup_hi_2036 = {dataGroup_hi_hi_2036, dataGroup_hi_lo_2036};
  wire [7:0]    dataGroup_52_31 = dataGroup_hi_2036[1311:1304];
  wire [2047:0] dataGroup_lo_2037 = {dataGroup_lo_hi_2037, dataGroup_lo_lo_2037};
  wire [2047:0] dataGroup_hi_2037 = {dataGroup_hi_hi_2037, dataGroup_hi_lo_2037};
  wire [7:0]    dataGroup_53_31 = dataGroup_hi_2037[1375:1368];
  wire [2047:0] dataGroup_lo_2038 = {dataGroup_lo_hi_2038, dataGroup_lo_lo_2038};
  wire [2047:0] dataGroup_hi_2038 = {dataGroup_hi_hi_2038, dataGroup_hi_lo_2038};
  wire [7:0]    dataGroup_54_31 = dataGroup_hi_2038[1439:1432];
  wire [2047:0] dataGroup_lo_2039 = {dataGroup_lo_hi_2039, dataGroup_lo_lo_2039};
  wire [2047:0] dataGroup_hi_2039 = {dataGroup_hi_hi_2039, dataGroup_hi_lo_2039};
  wire [7:0]    dataGroup_55_31 = dataGroup_hi_2039[1503:1496];
  wire [2047:0] dataGroup_lo_2040 = {dataGroup_lo_hi_2040, dataGroup_lo_lo_2040};
  wire [2047:0] dataGroup_hi_2040 = {dataGroup_hi_hi_2040, dataGroup_hi_lo_2040};
  wire [7:0]    dataGroup_56_31 = dataGroup_hi_2040[1567:1560];
  wire [2047:0] dataGroup_lo_2041 = {dataGroup_lo_hi_2041, dataGroup_lo_lo_2041};
  wire [2047:0] dataGroup_hi_2041 = {dataGroup_hi_hi_2041, dataGroup_hi_lo_2041};
  wire [7:0]    dataGroup_57_31 = dataGroup_hi_2041[1631:1624];
  wire [2047:0] dataGroup_lo_2042 = {dataGroup_lo_hi_2042, dataGroup_lo_lo_2042};
  wire [2047:0] dataGroup_hi_2042 = {dataGroup_hi_hi_2042, dataGroup_hi_lo_2042};
  wire [7:0]    dataGroup_58_31 = dataGroup_hi_2042[1695:1688];
  wire [2047:0] dataGroup_lo_2043 = {dataGroup_lo_hi_2043, dataGroup_lo_lo_2043};
  wire [2047:0] dataGroup_hi_2043 = {dataGroup_hi_hi_2043, dataGroup_hi_lo_2043};
  wire [7:0]    dataGroup_59_31 = dataGroup_hi_2043[1759:1752];
  wire [2047:0] dataGroup_lo_2044 = {dataGroup_lo_hi_2044, dataGroup_lo_lo_2044};
  wire [2047:0] dataGroup_hi_2044 = {dataGroup_hi_hi_2044, dataGroup_hi_lo_2044};
  wire [7:0]    dataGroup_60_31 = dataGroup_hi_2044[1823:1816];
  wire [2047:0] dataGroup_lo_2045 = {dataGroup_lo_hi_2045, dataGroup_lo_lo_2045};
  wire [2047:0] dataGroup_hi_2045 = {dataGroup_hi_hi_2045, dataGroup_hi_lo_2045};
  wire [7:0]    dataGroup_61_31 = dataGroup_hi_2045[1887:1880];
  wire [2047:0] dataGroup_lo_2046 = {dataGroup_lo_hi_2046, dataGroup_lo_lo_2046};
  wire [2047:0] dataGroup_hi_2046 = {dataGroup_hi_hi_2046, dataGroup_hi_lo_2046};
  wire [7:0]    dataGroup_62_31 = dataGroup_hi_2046[1951:1944];
  wire [2047:0] dataGroup_lo_2047 = {dataGroup_lo_hi_2047, dataGroup_lo_lo_2047};
  wire [2047:0] dataGroup_hi_2047 = {dataGroup_hi_hi_2047, dataGroup_hi_lo_2047};
  wire [7:0]    dataGroup_63_31 = dataGroup_hi_2047[2015:2008];
  wire [15:0]   res_lo_lo_lo_lo_lo_31 = {dataGroup_1_31, dataGroup_0_31};
  wire [15:0]   res_lo_lo_lo_lo_hi_31 = {dataGroup_3_31, dataGroup_2_31};
  wire [31:0]   res_lo_lo_lo_lo_31 = {res_lo_lo_lo_lo_hi_31, res_lo_lo_lo_lo_lo_31};
  wire [15:0]   res_lo_lo_lo_hi_lo_31 = {dataGroup_5_31, dataGroup_4_31};
  wire [15:0]   res_lo_lo_lo_hi_hi_31 = {dataGroup_7_31, dataGroup_6_31};
  wire [31:0]   res_lo_lo_lo_hi_31 = {res_lo_lo_lo_hi_hi_31, res_lo_lo_lo_hi_lo_31};
  wire [63:0]   res_lo_lo_lo_31 = {res_lo_lo_lo_hi_31, res_lo_lo_lo_lo_31};
  wire [15:0]   res_lo_lo_hi_lo_lo_31 = {dataGroup_9_31, dataGroup_8_31};
  wire [15:0]   res_lo_lo_hi_lo_hi_31 = {dataGroup_11_31, dataGroup_10_31};
  wire [31:0]   res_lo_lo_hi_lo_31 = {res_lo_lo_hi_lo_hi_31, res_lo_lo_hi_lo_lo_31};
  wire [15:0]   res_lo_lo_hi_hi_lo_31 = {dataGroup_13_31, dataGroup_12_31};
  wire [15:0]   res_lo_lo_hi_hi_hi_31 = {dataGroup_15_31, dataGroup_14_31};
  wire [31:0]   res_lo_lo_hi_hi_31 = {res_lo_lo_hi_hi_hi_31, res_lo_lo_hi_hi_lo_31};
  wire [63:0]   res_lo_lo_hi_31 = {res_lo_lo_hi_hi_31, res_lo_lo_hi_lo_31};
  wire [127:0]  res_lo_lo_31 = {res_lo_lo_hi_31, res_lo_lo_lo_31};
  wire [15:0]   res_lo_hi_lo_lo_lo_31 = {dataGroup_17_31, dataGroup_16_31};
  wire [15:0]   res_lo_hi_lo_lo_hi_31 = {dataGroup_19_31, dataGroup_18_31};
  wire [31:0]   res_lo_hi_lo_lo_31 = {res_lo_hi_lo_lo_hi_31, res_lo_hi_lo_lo_lo_31};
  wire [15:0]   res_lo_hi_lo_hi_lo_31 = {dataGroup_21_31, dataGroup_20_31};
  wire [15:0]   res_lo_hi_lo_hi_hi_31 = {dataGroup_23_31, dataGroup_22_31};
  wire [31:0]   res_lo_hi_lo_hi_31 = {res_lo_hi_lo_hi_hi_31, res_lo_hi_lo_hi_lo_31};
  wire [63:0]   res_lo_hi_lo_31 = {res_lo_hi_lo_hi_31, res_lo_hi_lo_lo_31};
  wire [15:0]   res_lo_hi_hi_lo_lo_31 = {dataGroup_25_31, dataGroup_24_31};
  wire [15:0]   res_lo_hi_hi_lo_hi_31 = {dataGroup_27_31, dataGroup_26_31};
  wire [31:0]   res_lo_hi_hi_lo_31 = {res_lo_hi_hi_lo_hi_31, res_lo_hi_hi_lo_lo_31};
  wire [15:0]   res_lo_hi_hi_hi_lo_31 = {dataGroup_29_31, dataGroup_28_31};
  wire [15:0]   res_lo_hi_hi_hi_hi_31 = {dataGroup_31_31, dataGroup_30_31};
  wire [31:0]   res_lo_hi_hi_hi_31 = {res_lo_hi_hi_hi_hi_31, res_lo_hi_hi_hi_lo_31};
  wire [63:0]   res_lo_hi_hi_31 = {res_lo_hi_hi_hi_31, res_lo_hi_hi_lo_31};
  wire [127:0]  res_lo_hi_31 = {res_lo_hi_hi_31, res_lo_hi_lo_31};
  wire [255:0]  res_lo_31 = {res_lo_hi_31, res_lo_lo_31};
  wire [15:0]   res_hi_lo_lo_lo_lo_31 = {dataGroup_33_31, dataGroup_32_31};
  wire [15:0]   res_hi_lo_lo_lo_hi_31 = {dataGroup_35_31, dataGroup_34_31};
  wire [31:0]   res_hi_lo_lo_lo_31 = {res_hi_lo_lo_lo_hi_31, res_hi_lo_lo_lo_lo_31};
  wire [15:0]   res_hi_lo_lo_hi_lo_31 = {dataGroup_37_31, dataGroup_36_31};
  wire [15:0]   res_hi_lo_lo_hi_hi_31 = {dataGroup_39_31, dataGroup_38_31};
  wire [31:0]   res_hi_lo_lo_hi_31 = {res_hi_lo_lo_hi_hi_31, res_hi_lo_lo_hi_lo_31};
  wire [63:0]   res_hi_lo_lo_31 = {res_hi_lo_lo_hi_31, res_hi_lo_lo_lo_31};
  wire [15:0]   res_hi_lo_hi_lo_lo_31 = {dataGroup_41_31, dataGroup_40_31};
  wire [15:0]   res_hi_lo_hi_lo_hi_31 = {dataGroup_43_31, dataGroup_42_31};
  wire [31:0]   res_hi_lo_hi_lo_31 = {res_hi_lo_hi_lo_hi_31, res_hi_lo_hi_lo_lo_31};
  wire [15:0]   res_hi_lo_hi_hi_lo_31 = {dataGroup_45_31, dataGroup_44_31};
  wire [15:0]   res_hi_lo_hi_hi_hi_31 = {dataGroup_47_31, dataGroup_46_31};
  wire [31:0]   res_hi_lo_hi_hi_31 = {res_hi_lo_hi_hi_hi_31, res_hi_lo_hi_hi_lo_31};
  wire [63:0]   res_hi_lo_hi_31 = {res_hi_lo_hi_hi_31, res_hi_lo_hi_lo_31};
  wire [127:0]  res_hi_lo_31 = {res_hi_lo_hi_31, res_hi_lo_lo_31};
  wire [15:0]   res_hi_hi_lo_lo_lo_31 = {dataGroup_49_31, dataGroup_48_31};
  wire [15:0]   res_hi_hi_lo_lo_hi_31 = {dataGroup_51_31, dataGroup_50_31};
  wire [31:0]   res_hi_hi_lo_lo_31 = {res_hi_hi_lo_lo_hi_31, res_hi_hi_lo_lo_lo_31};
  wire [15:0]   res_hi_hi_lo_hi_lo_31 = {dataGroup_53_31, dataGroup_52_31};
  wire [15:0]   res_hi_hi_lo_hi_hi_31 = {dataGroup_55_31, dataGroup_54_31};
  wire [31:0]   res_hi_hi_lo_hi_31 = {res_hi_hi_lo_hi_hi_31, res_hi_hi_lo_hi_lo_31};
  wire [63:0]   res_hi_hi_lo_31 = {res_hi_hi_lo_hi_31, res_hi_hi_lo_lo_31};
  wire [15:0]   res_hi_hi_hi_lo_lo_31 = {dataGroup_57_31, dataGroup_56_31};
  wire [15:0]   res_hi_hi_hi_lo_hi_31 = {dataGroup_59_31, dataGroup_58_31};
  wire [31:0]   res_hi_hi_hi_lo_31 = {res_hi_hi_hi_lo_hi_31, res_hi_hi_hi_lo_lo_31};
  wire [15:0]   res_hi_hi_hi_hi_lo_31 = {dataGroup_61_31, dataGroup_60_31};
  wire [15:0]   res_hi_hi_hi_hi_hi_31 = {dataGroup_63_31, dataGroup_62_31};
  wire [31:0]   res_hi_hi_hi_hi_31 = {res_hi_hi_hi_hi_hi_31, res_hi_hi_hi_hi_lo_31};
  wire [63:0]   res_hi_hi_hi_31 = {res_hi_hi_hi_hi_31, res_hi_hi_hi_lo_31};
  wire [127:0]  res_hi_hi_31 = {res_hi_hi_hi_31, res_hi_hi_lo_31};
  wire [255:0]  res_hi_31 = {res_hi_hi_31, res_hi_lo_31};
  wire [511:0]  res_59 = {res_hi_31, res_lo_31};
  wire [2047:0] dataGroup_lo_2048 = {dataGroup_lo_hi_2048, dataGroup_lo_lo_2048};
  wire [2047:0] dataGroup_hi_2048 = {dataGroup_hi_hi_2048, dataGroup_hi_lo_2048};
  wire [7:0]    dataGroup_0_32 = dataGroup_lo_2048[39:32];
  wire [2047:0] dataGroup_lo_2049 = {dataGroup_lo_hi_2049, dataGroup_lo_lo_2049};
  wire [2047:0] dataGroup_hi_2049 = {dataGroup_hi_hi_2049, dataGroup_hi_lo_2049};
  wire [7:0]    dataGroup_1_32 = dataGroup_lo_2049[103:96];
  wire [2047:0] dataGroup_lo_2050 = {dataGroup_lo_hi_2050, dataGroup_lo_lo_2050};
  wire [2047:0] dataGroup_hi_2050 = {dataGroup_hi_hi_2050, dataGroup_hi_lo_2050};
  wire [7:0]    dataGroup_2_32 = dataGroup_lo_2050[167:160];
  wire [2047:0] dataGroup_lo_2051 = {dataGroup_lo_hi_2051, dataGroup_lo_lo_2051};
  wire [2047:0] dataGroup_hi_2051 = {dataGroup_hi_hi_2051, dataGroup_hi_lo_2051};
  wire [7:0]    dataGroup_3_32 = dataGroup_lo_2051[231:224];
  wire [2047:0] dataGroup_lo_2052 = {dataGroup_lo_hi_2052, dataGroup_lo_lo_2052};
  wire [2047:0] dataGroup_hi_2052 = {dataGroup_hi_hi_2052, dataGroup_hi_lo_2052};
  wire [7:0]    dataGroup_4_32 = dataGroup_lo_2052[295:288];
  wire [2047:0] dataGroup_lo_2053 = {dataGroup_lo_hi_2053, dataGroup_lo_lo_2053};
  wire [2047:0] dataGroup_hi_2053 = {dataGroup_hi_hi_2053, dataGroup_hi_lo_2053};
  wire [7:0]    dataGroup_5_32 = dataGroup_lo_2053[359:352];
  wire [2047:0] dataGroup_lo_2054 = {dataGroup_lo_hi_2054, dataGroup_lo_lo_2054};
  wire [2047:0] dataGroup_hi_2054 = {dataGroup_hi_hi_2054, dataGroup_hi_lo_2054};
  wire [7:0]    dataGroup_6_32 = dataGroup_lo_2054[423:416];
  wire [2047:0] dataGroup_lo_2055 = {dataGroup_lo_hi_2055, dataGroup_lo_lo_2055};
  wire [2047:0] dataGroup_hi_2055 = {dataGroup_hi_hi_2055, dataGroup_hi_lo_2055};
  wire [7:0]    dataGroup_7_32 = dataGroup_lo_2055[487:480];
  wire [2047:0] dataGroup_lo_2056 = {dataGroup_lo_hi_2056, dataGroup_lo_lo_2056};
  wire [2047:0] dataGroup_hi_2056 = {dataGroup_hi_hi_2056, dataGroup_hi_lo_2056};
  wire [7:0]    dataGroup_8_32 = dataGroup_lo_2056[551:544];
  wire [2047:0] dataGroup_lo_2057 = {dataGroup_lo_hi_2057, dataGroup_lo_lo_2057};
  wire [2047:0] dataGroup_hi_2057 = {dataGroup_hi_hi_2057, dataGroup_hi_lo_2057};
  wire [7:0]    dataGroup_9_32 = dataGroup_lo_2057[615:608];
  wire [2047:0] dataGroup_lo_2058 = {dataGroup_lo_hi_2058, dataGroup_lo_lo_2058};
  wire [2047:0] dataGroup_hi_2058 = {dataGroup_hi_hi_2058, dataGroup_hi_lo_2058};
  wire [7:0]    dataGroup_10_32 = dataGroup_lo_2058[679:672];
  wire [2047:0] dataGroup_lo_2059 = {dataGroup_lo_hi_2059, dataGroup_lo_lo_2059};
  wire [2047:0] dataGroup_hi_2059 = {dataGroup_hi_hi_2059, dataGroup_hi_lo_2059};
  wire [7:0]    dataGroup_11_32 = dataGroup_lo_2059[743:736];
  wire [2047:0] dataGroup_lo_2060 = {dataGroup_lo_hi_2060, dataGroup_lo_lo_2060};
  wire [2047:0] dataGroup_hi_2060 = {dataGroup_hi_hi_2060, dataGroup_hi_lo_2060};
  wire [7:0]    dataGroup_12_32 = dataGroup_lo_2060[807:800];
  wire [2047:0] dataGroup_lo_2061 = {dataGroup_lo_hi_2061, dataGroup_lo_lo_2061};
  wire [2047:0] dataGroup_hi_2061 = {dataGroup_hi_hi_2061, dataGroup_hi_lo_2061};
  wire [7:0]    dataGroup_13_32 = dataGroup_lo_2061[871:864];
  wire [2047:0] dataGroup_lo_2062 = {dataGroup_lo_hi_2062, dataGroup_lo_lo_2062};
  wire [2047:0] dataGroup_hi_2062 = {dataGroup_hi_hi_2062, dataGroup_hi_lo_2062};
  wire [7:0]    dataGroup_14_32 = dataGroup_lo_2062[935:928];
  wire [2047:0] dataGroup_lo_2063 = {dataGroup_lo_hi_2063, dataGroup_lo_lo_2063};
  wire [2047:0] dataGroup_hi_2063 = {dataGroup_hi_hi_2063, dataGroup_hi_lo_2063};
  wire [7:0]    dataGroup_15_32 = dataGroup_lo_2063[999:992];
  wire [2047:0] dataGroup_lo_2064 = {dataGroup_lo_hi_2064, dataGroup_lo_lo_2064};
  wire [2047:0] dataGroup_hi_2064 = {dataGroup_hi_hi_2064, dataGroup_hi_lo_2064};
  wire [7:0]    dataGroup_16_32 = dataGroup_lo_2064[1063:1056];
  wire [2047:0] dataGroup_lo_2065 = {dataGroup_lo_hi_2065, dataGroup_lo_lo_2065};
  wire [2047:0] dataGroup_hi_2065 = {dataGroup_hi_hi_2065, dataGroup_hi_lo_2065};
  wire [7:0]    dataGroup_17_32 = dataGroup_lo_2065[1127:1120];
  wire [2047:0] dataGroup_lo_2066 = {dataGroup_lo_hi_2066, dataGroup_lo_lo_2066};
  wire [2047:0] dataGroup_hi_2066 = {dataGroup_hi_hi_2066, dataGroup_hi_lo_2066};
  wire [7:0]    dataGroup_18_32 = dataGroup_lo_2066[1191:1184];
  wire [2047:0] dataGroup_lo_2067 = {dataGroup_lo_hi_2067, dataGroup_lo_lo_2067};
  wire [2047:0] dataGroup_hi_2067 = {dataGroup_hi_hi_2067, dataGroup_hi_lo_2067};
  wire [7:0]    dataGroup_19_32 = dataGroup_lo_2067[1255:1248];
  wire [2047:0] dataGroup_lo_2068 = {dataGroup_lo_hi_2068, dataGroup_lo_lo_2068};
  wire [2047:0] dataGroup_hi_2068 = {dataGroup_hi_hi_2068, dataGroup_hi_lo_2068};
  wire [7:0]    dataGroup_20_32 = dataGroup_lo_2068[1319:1312];
  wire [2047:0] dataGroup_lo_2069 = {dataGroup_lo_hi_2069, dataGroup_lo_lo_2069};
  wire [2047:0] dataGroup_hi_2069 = {dataGroup_hi_hi_2069, dataGroup_hi_lo_2069};
  wire [7:0]    dataGroup_21_32 = dataGroup_lo_2069[1383:1376];
  wire [2047:0] dataGroup_lo_2070 = {dataGroup_lo_hi_2070, dataGroup_lo_lo_2070};
  wire [2047:0] dataGroup_hi_2070 = {dataGroup_hi_hi_2070, dataGroup_hi_lo_2070};
  wire [7:0]    dataGroup_22_32 = dataGroup_lo_2070[1447:1440];
  wire [2047:0] dataGroup_lo_2071 = {dataGroup_lo_hi_2071, dataGroup_lo_lo_2071};
  wire [2047:0] dataGroup_hi_2071 = {dataGroup_hi_hi_2071, dataGroup_hi_lo_2071};
  wire [7:0]    dataGroup_23_32 = dataGroup_lo_2071[1511:1504];
  wire [2047:0] dataGroup_lo_2072 = {dataGroup_lo_hi_2072, dataGroup_lo_lo_2072};
  wire [2047:0] dataGroup_hi_2072 = {dataGroup_hi_hi_2072, dataGroup_hi_lo_2072};
  wire [7:0]    dataGroup_24_32 = dataGroup_lo_2072[1575:1568];
  wire [2047:0] dataGroup_lo_2073 = {dataGroup_lo_hi_2073, dataGroup_lo_lo_2073};
  wire [2047:0] dataGroup_hi_2073 = {dataGroup_hi_hi_2073, dataGroup_hi_lo_2073};
  wire [7:0]    dataGroup_25_32 = dataGroup_lo_2073[1639:1632];
  wire [2047:0] dataGroup_lo_2074 = {dataGroup_lo_hi_2074, dataGroup_lo_lo_2074};
  wire [2047:0] dataGroup_hi_2074 = {dataGroup_hi_hi_2074, dataGroup_hi_lo_2074};
  wire [7:0]    dataGroup_26_32 = dataGroup_lo_2074[1703:1696];
  wire [2047:0] dataGroup_lo_2075 = {dataGroup_lo_hi_2075, dataGroup_lo_lo_2075};
  wire [2047:0] dataGroup_hi_2075 = {dataGroup_hi_hi_2075, dataGroup_hi_lo_2075};
  wire [7:0]    dataGroup_27_32 = dataGroup_lo_2075[1767:1760];
  wire [2047:0] dataGroup_lo_2076 = {dataGroup_lo_hi_2076, dataGroup_lo_lo_2076};
  wire [2047:0] dataGroup_hi_2076 = {dataGroup_hi_hi_2076, dataGroup_hi_lo_2076};
  wire [7:0]    dataGroup_28_32 = dataGroup_lo_2076[1831:1824];
  wire [2047:0] dataGroup_lo_2077 = {dataGroup_lo_hi_2077, dataGroup_lo_lo_2077};
  wire [2047:0] dataGroup_hi_2077 = {dataGroup_hi_hi_2077, dataGroup_hi_lo_2077};
  wire [7:0]    dataGroup_29_32 = dataGroup_lo_2077[1895:1888];
  wire [2047:0] dataGroup_lo_2078 = {dataGroup_lo_hi_2078, dataGroup_lo_lo_2078};
  wire [2047:0] dataGroup_hi_2078 = {dataGroup_hi_hi_2078, dataGroup_hi_lo_2078};
  wire [7:0]    dataGroup_30_32 = dataGroup_lo_2078[1959:1952];
  wire [2047:0] dataGroup_lo_2079 = {dataGroup_lo_hi_2079, dataGroup_lo_lo_2079};
  wire [2047:0] dataGroup_hi_2079 = {dataGroup_hi_hi_2079, dataGroup_hi_lo_2079};
  wire [7:0]    dataGroup_31_32 = dataGroup_lo_2079[2023:2016];
  wire [2047:0] dataGroup_lo_2080 = {dataGroup_lo_hi_2080, dataGroup_lo_lo_2080};
  wire [2047:0] dataGroup_hi_2080 = {dataGroup_hi_hi_2080, dataGroup_hi_lo_2080};
  wire [7:0]    dataGroup_32_32 = dataGroup_hi_2080[39:32];
  wire [2047:0] dataGroup_lo_2081 = {dataGroup_lo_hi_2081, dataGroup_lo_lo_2081};
  wire [2047:0] dataGroup_hi_2081 = {dataGroup_hi_hi_2081, dataGroup_hi_lo_2081};
  wire [7:0]    dataGroup_33_32 = dataGroup_hi_2081[103:96];
  wire [2047:0] dataGroup_lo_2082 = {dataGroup_lo_hi_2082, dataGroup_lo_lo_2082};
  wire [2047:0] dataGroup_hi_2082 = {dataGroup_hi_hi_2082, dataGroup_hi_lo_2082};
  wire [7:0]    dataGroup_34_32 = dataGroup_hi_2082[167:160];
  wire [2047:0] dataGroup_lo_2083 = {dataGroup_lo_hi_2083, dataGroup_lo_lo_2083};
  wire [2047:0] dataGroup_hi_2083 = {dataGroup_hi_hi_2083, dataGroup_hi_lo_2083};
  wire [7:0]    dataGroup_35_32 = dataGroup_hi_2083[231:224];
  wire [2047:0] dataGroup_lo_2084 = {dataGroup_lo_hi_2084, dataGroup_lo_lo_2084};
  wire [2047:0] dataGroup_hi_2084 = {dataGroup_hi_hi_2084, dataGroup_hi_lo_2084};
  wire [7:0]    dataGroup_36_32 = dataGroup_hi_2084[295:288];
  wire [2047:0] dataGroup_lo_2085 = {dataGroup_lo_hi_2085, dataGroup_lo_lo_2085};
  wire [2047:0] dataGroup_hi_2085 = {dataGroup_hi_hi_2085, dataGroup_hi_lo_2085};
  wire [7:0]    dataGroup_37_32 = dataGroup_hi_2085[359:352];
  wire [2047:0] dataGroup_lo_2086 = {dataGroup_lo_hi_2086, dataGroup_lo_lo_2086};
  wire [2047:0] dataGroup_hi_2086 = {dataGroup_hi_hi_2086, dataGroup_hi_lo_2086};
  wire [7:0]    dataGroup_38_32 = dataGroup_hi_2086[423:416];
  wire [2047:0] dataGroup_lo_2087 = {dataGroup_lo_hi_2087, dataGroup_lo_lo_2087};
  wire [2047:0] dataGroup_hi_2087 = {dataGroup_hi_hi_2087, dataGroup_hi_lo_2087};
  wire [7:0]    dataGroup_39_32 = dataGroup_hi_2087[487:480];
  wire [2047:0] dataGroup_lo_2088 = {dataGroup_lo_hi_2088, dataGroup_lo_lo_2088};
  wire [2047:0] dataGroup_hi_2088 = {dataGroup_hi_hi_2088, dataGroup_hi_lo_2088};
  wire [7:0]    dataGroup_40_32 = dataGroup_hi_2088[551:544];
  wire [2047:0] dataGroup_lo_2089 = {dataGroup_lo_hi_2089, dataGroup_lo_lo_2089};
  wire [2047:0] dataGroup_hi_2089 = {dataGroup_hi_hi_2089, dataGroup_hi_lo_2089};
  wire [7:0]    dataGroup_41_32 = dataGroup_hi_2089[615:608];
  wire [2047:0] dataGroup_lo_2090 = {dataGroup_lo_hi_2090, dataGroup_lo_lo_2090};
  wire [2047:0] dataGroup_hi_2090 = {dataGroup_hi_hi_2090, dataGroup_hi_lo_2090};
  wire [7:0]    dataGroup_42_32 = dataGroup_hi_2090[679:672];
  wire [2047:0] dataGroup_lo_2091 = {dataGroup_lo_hi_2091, dataGroup_lo_lo_2091};
  wire [2047:0] dataGroup_hi_2091 = {dataGroup_hi_hi_2091, dataGroup_hi_lo_2091};
  wire [7:0]    dataGroup_43_32 = dataGroup_hi_2091[743:736];
  wire [2047:0] dataGroup_lo_2092 = {dataGroup_lo_hi_2092, dataGroup_lo_lo_2092};
  wire [2047:0] dataGroup_hi_2092 = {dataGroup_hi_hi_2092, dataGroup_hi_lo_2092};
  wire [7:0]    dataGroup_44_32 = dataGroup_hi_2092[807:800];
  wire [2047:0] dataGroup_lo_2093 = {dataGroup_lo_hi_2093, dataGroup_lo_lo_2093};
  wire [2047:0] dataGroup_hi_2093 = {dataGroup_hi_hi_2093, dataGroup_hi_lo_2093};
  wire [7:0]    dataGroup_45_32 = dataGroup_hi_2093[871:864];
  wire [2047:0] dataGroup_lo_2094 = {dataGroup_lo_hi_2094, dataGroup_lo_lo_2094};
  wire [2047:0] dataGroup_hi_2094 = {dataGroup_hi_hi_2094, dataGroup_hi_lo_2094};
  wire [7:0]    dataGroup_46_32 = dataGroup_hi_2094[935:928];
  wire [2047:0] dataGroup_lo_2095 = {dataGroup_lo_hi_2095, dataGroup_lo_lo_2095};
  wire [2047:0] dataGroup_hi_2095 = {dataGroup_hi_hi_2095, dataGroup_hi_lo_2095};
  wire [7:0]    dataGroup_47_32 = dataGroup_hi_2095[999:992];
  wire [2047:0] dataGroup_lo_2096 = {dataGroup_lo_hi_2096, dataGroup_lo_lo_2096};
  wire [2047:0] dataGroup_hi_2096 = {dataGroup_hi_hi_2096, dataGroup_hi_lo_2096};
  wire [7:0]    dataGroup_48_32 = dataGroup_hi_2096[1063:1056];
  wire [2047:0] dataGroup_lo_2097 = {dataGroup_lo_hi_2097, dataGroup_lo_lo_2097};
  wire [2047:0] dataGroup_hi_2097 = {dataGroup_hi_hi_2097, dataGroup_hi_lo_2097};
  wire [7:0]    dataGroup_49_32 = dataGroup_hi_2097[1127:1120];
  wire [2047:0] dataGroup_lo_2098 = {dataGroup_lo_hi_2098, dataGroup_lo_lo_2098};
  wire [2047:0] dataGroup_hi_2098 = {dataGroup_hi_hi_2098, dataGroup_hi_lo_2098};
  wire [7:0]    dataGroup_50_32 = dataGroup_hi_2098[1191:1184];
  wire [2047:0] dataGroup_lo_2099 = {dataGroup_lo_hi_2099, dataGroup_lo_lo_2099};
  wire [2047:0] dataGroup_hi_2099 = {dataGroup_hi_hi_2099, dataGroup_hi_lo_2099};
  wire [7:0]    dataGroup_51_32 = dataGroup_hi_2099[1255:1248];
  wire [2047:0] dataGroup_lo_2100 = {dataGroup_lo_hi_2100, dataGroup_lo_lo_2100};
  wire [2047:0] dataGroup_hi_2100 = {dataGroup_hi_hi_2100, dataGroup_hi_lo_2100};
  wire [7:0]    dataGroup_52_32 = dataGroup_hi_2100[1319:1312];
  wire [2047:0] dataGroup_lo_2101 = {dataGroup_lo_hi_2101, dataGroup_lo_lo_2101};
  wire [2047:0] dataGroup_hi_2101 = {dataGroup_hi_hi_2101, dataGroup_hi_lo_2101};
  wire [7:0]    dataGroup_53_32 = dataGroup_hi_2101[1383:1376];
  wire [2047:0] dataGroup_lo_2102 = {dataGroup_lo_hi_2102, dataGroup_lo_lo_2102};
  wire [2047:0] dataGroup_hi_2102 = {dataGroup_hi_hi_2102, dataGroup_hi_lo_2102};
  wire [7:0]    dataGroup_54_32 = dataGroup_hi_2102[1447:1440];
  wire [2047:0] dataGroup_lo_2103 = {dataGroup_lo_hi_2103, dataGroup_lo_lo_2103};
  wire [2047:0] dataGroup_hi_2103 = {dataGroup_hi_hi_2103, dataGroup_hi_lo_2103};
  wire [7:0]    dataGroup_55_32 = dataGroup_hi_2103[1511:1504];
  wire [2047:0] dataGroup_lo_2104 = {dataGroup_lo_hi_2104, dataGroup_lo_lo_2104};
  wire [2047:0] dataGroup_hi_2104 = {dataGroup_hi_hi_2104, dataGroup_hi_lo_2104};
  wire [7:0]    dataGroup_56_32 = dataGroup_hi_2104[1575:1568];
  wire [2047:0] dataGroup_lo_2105 = {dataGroup_lo_hi_2105, dataGroup_lo_lo_2105};
  wire [2047:0] dataGroup_hi_2105 = {dataGroup_hi_hi_2105, dataGroup_hi_lo_2105};
  wire [7:0]    dataGroup_57_32 = dataGroup_hi_2105[1639:1632];
  wire [2047:0] dataGroup_lo_2106 = {dataGroup_lo_hi_2106, dataGroup_lo_lo_2106};
  wire [2047:0] dataGroup_hi_2106 = {dataGroup_hi_hi_2106, dataGroup_hi_lo_2106};
  wire [7:0]    dataGroup_58_32 = dataGroup_hi_2106[1703:1696];
  wire [2047:0] dataGroup_lo_2107 = {dataGroup_lo_hi_2107, dataGroup_lo_lo_2107};
  wire [2047:0] dataGroup_hi_2107 = {dataGroup_hi_hi_2107, dataGroup_hi_lo_2107};
  wire [7:0]    dataGroup_59_32 = dataGroup_hi_2107[1767:1760];
  wire [2047:0] dataGroup_lo_2108 = {dataGroup_lo_hi_2108, dataGroup_lo_lo_2108};
  wire [2047:0] dataGroup_hi_2108 = {dataGroup_hi_hi_2108, dataGroup_hi_lo_2108};
  wire [7:0]    dataGroup_60_32 = dataGroup_hi_2108[1831:1824];
  wire [2047:0] dataGroup_lo_2109 = {dataGroup_lo_hi_2109, dataGroup_lo_lo_2109};
  wire [2047:0] dataGroup_hi_2109 = {dataGroup_hi_hi_2109, dataGroup_hi_lo_2109};
  wire [7:0]    dataGroup_61_32 = dataGroup_hi_2109[1895:1888];
  wire [2047:0] dataGroup_lo_2110 = {dataGroup_lo_hi_2110, dataGroup_lo_lo_2110};
  wire [2047:0] dataGroup_hi_2110 = {dataGroup_hi_hi_2110, dataGroup_hi_lo_2110};
  wire [7:0]    dataGroup_62_32 = dataGroup_hi_2110[1959:1952];
  wire [2047:0] dataGroup_lo_2111 = {dataGroup_lo_hi_2111, dataGroup_lo_lo_2111};
  wire [2047:0] dataGroup_hi_2111 = {dataGroup_hi_hi_2111, dataGroup_hi_lo_2111};
  wire [7:0]    dataGroup_63_32 = dataGroup_hi_2111[2023:2016];
  wire [15:0]   res_lo_lo_lo_lo_lo_32 = {dataGroup_1_32, dataGroup_0_32};
  wire [15:0]   res_lo_lo_lo_lo_hi_32 = {dataGroup_3_32, dataGroup_2_32};
  wire [31:0]   res_lo_lo_lo_lo_32 = {res_lo_lo_lo_lo_hi_32, res_lo_lo_lo_lo_lo_32};
  wire [15:0]   res_lo_lo_lo_hi_lo_32 = {dataGroup_5_32, dataGroup_4_32};
  wire [15:0]   res_lo_lo_lo_hi_hi_32 = {dataGroup_7_32, dataGroup_6_32};
  wire [31:0]   res_lo_lo_lo_hi_32 = {res_lo_lo_lo_hi_hi_32, res_lo_lo_lo_hi_lo_32};
  wire [63:0]   res_lo_lo_lo_32 = {res_lo_lo_lo_hi_32, res_lo_lo_lo_lo_32};
  wire [15:0]   res_lo_lo_hi_lo_lo_32 = {dataGroup_9_32, dataGroup_8_32};
  wire [15:0]   res_lo_lo_hi_lo_hi_32 = {dataGroup_11_32, dataGroup_10_32};
  wire [31:0]   res_lo_lo_hi_lo_32 = {res_lo_lo_hi_lo_hi_32, res_lo_lo_hi_lo_lo_32};
  wire [15:0]   res_lo_lo_hi_hi_lo_32 = {dataGroup_13_32, dataGroup_12_32};
  wire [15:0]   res_lo_lo_hi_hi_hi_32 = {dataGroup_15_32, dataGroup_14_32};
  wire [31:0]   res_lo_lo_hi_hi_32 = {res_lo_lo_hi_hi_hi_32, res_lo_lo_hi_hi_lo_32};
  wire [63:0]   res_lo_lo_hi_32 = {res_lo_lo_hi_hi_32, res_lo_lo_hi_lo_32};
  wire [127:0]  res_lo_lo_32 = {res_lo_lo_hi_32, res_lo_lo_lo_32};
  wire [15:0]   res_lo_hi_lo_lo_lo_32 = {dataGroup_17_32, dataGroup_16_32};
  wire [15:0]   res_lo_hi_lo_lo_hi_32 = {dataGroup_19_32, dataGroup_18_32};
  wire [31:0]   res_lo_hi_lo_lo_32 = {res_lo_hi_lo_lo_hi_32, res_lo_hi_lo_lo_lo_32};
  wire [15:0]   res_lo_hi_lo_hi_lo_32 = {dataGroup_21_32, dataGroup_20_32};
  wire [15:0]   res_lo_hi_lo_hi_hi_32 = {dataGroup_23_32, dataGroup_22_32};
  wire [31:0]   res_lo_hi_lo_hi_32 = {res_lo_hi_lo_hi_hi_32, res_lo_hi_lo_hi_lo_32};
  wire [63:0]   res_lo_hi_lo_32 = {res_lo_hi_lo_hi_32, res_lo_hi_lo_lo_32};
  wire [15:0]   res_lo_hi_hi_lo_lo_32 = {dataGroup_25_32, dataGroup_24_32};
  wire [15:0]   res_lo_hi_hi_lo_hi_32 = {dataGroup_27_32, dataGroup_26_32};
  wire [31:0]   res_lo_hi_hi_lo_32 = {res_lo_hi_hi_lo_hi_32, res_lo_hi_hi_lo_lo_32};
  wire [15:0]   res_lo_hi_hi_hi_lo_32 = {dataGroup_29_32, dataGroup_28_32};
  wire [15:0]   res_lo_hi_hi_hi_hi_32 = {dataGroup_31_32, dataGroup_30_32};
  wire [31:0]   res_lo_hi_hi_hi_32 = {res_lo_hi_hi_hi_hi_32, res_lo_hi_hi_hi_lo_32};
  wire [63:0]   res_lo_hi_hi_32 = {res_lo_hi_hi_hi_32, res_lo_hi_hi_lo_32};
  wire [127:0]  res_lo_hi_32 = {res_lo_hi_hi_32, res_lo_hi_lo_32};
  wire [255:0]  res_lo_32 = {res_lo_hi_32, res_lo_lo_32};
  wire [15:0]   res_hi_lo_lo_lo_lo_32 = {dataGroup_33_32, dataGroup_32_32};
  wire [15:0]   res_hi_lo_lo_lo_hi_32 = {dataGroup_35_32, dataGroup_34_32};
  wire [31:0]   res_hi_lo_lo_lo_32 = {res_hi_lo_lo_lo_hi_32, res_hi_lo_lo_lo_lo_32};
  wire [15:0]   res_hi_lo_lo_hi_lo_32 = {dataGroup_37_32, dataGroup_36_32};
  wire [15:0]   res_hi_lo_lo_hi_hi_32 = {dataGroup_39_32, dataGroup_38_32};
  wire [31:0]   res_hi_lo_lo_hi_32 = {res_hi_lo_lo_hi_hi_32, res_hi_lo_lo_hi_lo_32};
  wire [63:0]   res_hi_lo_lo_32 = {res_hi_lo_lo_hi_32, res_hi_lo_lo_lo_32};
  wire [15:0]   res_hi_lo_hi_lo_lo_32 = {dataGroup_41_32, dataGroup_40_32};
  wire [15:0]   res_hi_lo_hi_lo_hi_32 = {dataGroup_43_32, dataGroup_42_32};
  wire [31:0]   res_hi_lo_hi_lo_32 = {res_hi_lo_hi_lo_hi_32, res_hi_lo_hi_lo_lo_32};
  wire [15:0]   res_hi_lo_hi_hi_lo_32 = {dataGroup_45_32, dataGroup_44_32};
  wire [15:0]   res_hi_lo_hi_hi_hi_32 = {dataGroup_47_32, dataGroup_46_32};
  wire [31:0]   res_hi_lo_hi_hi_32 = {res_hi_lo_hi_hi_hi_32, res_hi_lo_hi_hi_lo_32};
  wire [63:0]   res_hi_lo_hi_32 = {res_hi_lo_hi_hi_32, res_hi_lo_hi_lo_32};
  wire [127:0]  res_hi_lo_32 = {res_hi_lo_hi_32, res_hi_lo_lo_32};
  wire [15:0]   res_hi_hi_lo_lo_lo_32 = {dataGroup_49_32, dataGroup_48_32};
  wire [15:0]   res_hi_hi_lo_lo_hi_32 = {dataGroup_51_32, dataGroup_50_32};
  wire [31:0]   res_hi_hi_lo_lo_32 = {res_hi_hi_lo_lo_hi_32, res_hi_hi_lo_lo_lo_32};
  wire [15:0]   res_hi_hi_lo_hi_lo_32 = {dataGroup_53_32, dataGroup_52_32};
  wire [15:0]   res_hi_hi_lo_hi_hi_32 = {dataGroup_55_32, dataGroup_54_32};
  wire [31:0]   res_hi_hi_lo_hi_32 = {res_hi_hi_lo_hi_hi_32, res_hi_hi_lo_hi_lo_32};
  wire [63:0]   res_hi_hi_lo_32 = {res_hi_hi_lo_hi_32, res_hi_hi_lo_lo_32};
  wire [15:0]   res_hi_hi_hi_lo_lo_32 = {dataGroup_57_32, dataGroup_56_32};
  wire [15:0]   res_hi_hi_hi_lo_hi_32 = {dataGroup_59_32, dataGroup_58_32};
  wire [31:0]   res_hi_hi_hi_lo_32 = {res_hi_hi_hi_lo_hi_32, res_hi_hi_hi_lo_lo_32};
  wire [15:0]   res_hi_hi_hi_hi_lo_32 = {dataGroup_61_32, dataGroup_60_32};
  wire [15:0]   res_hi_hi_hi_hi_hi_32 = {dataGroup_63_32, dataGroup_62_32};
  wire [31:0]   res_hi_hi_hi_hi_32 = {res_hi_hi_hi_hi_hi_32, res_hi_hi_hi_hi_lo_32};
  wire [63:0]   res_hi_hi_hi_32 = {res_hi_hi_hi_hi_32, res_hi_hi_hi_lo_32};
  wire [127:0]  res_hi_hi_32 = {res_hi_hi_hi_32, res_hi_hi_lo_32};
  wire [255:0]  res_hi_32 = {res_hi_hi_32, res_hi_lo_32};
  wire [511:0]  res_60 = {res_hi_32, res_lo_32};
  wire [2047:0] dataGroup_lo_2112 = {dataGroup_lo_hi_2112, dataGroup_lo_lo_2112};
  wire [2047:0] dataGroup_hi_2112 = {dataGroup_hi_hi_2112, dataGroup_hi_lo_2112};
  wire [7:0]    dataGroup_0_33 = dataGroup_lo_2112[47:40];
  wire [2047:0] dataGroup_lo_2113 = {dataGroup_lo_hi_2113, dataGroup_lo_lo_2113};
  wire [2047:0] dataGroup_hi_2113 = {dataGroup_hi_hi_2113, dataGroup_hi_lo_2113};
  wire [7:0]    dataGroup_1_33 = dataGroup_lo_2113[111:104];
  wire [2047:0] dataGroup_lo_2114 = {dataGroup_lo_hi_2114, dataGroup_lo_lo_2114};
  wire [2047:0] dataGroup_hi_2114 = {dataGroup_hi_hi_2114, dataGroup_hi_lo_2114};
  wire [7:0]    dataGroup_2_33 = dataGroup_lo_2114[175:168];
  wire [2047:0] dataGroup_lo_2115 = {dataGroup_lo_hi_2115, dataGroup_lo_lo_2115};
  wire [2047:0] dataGroup_hi_2115 = {dataGroup_hi_hi_2115, dataGroup_hi_lo_2115};
  wire [7:0]    dataGroup_3_33 = dataGroup_lo_2115[239:232];
  wire [2047:0] dataGroup_lo_2116 = {dataGroup_lo_hi_2116, dataGroup_lo_lo_2116};
  wire [2047:0] dataGroup_hi_2116 = {dataGroup_hi_hi_2116, dataGroup_hi_lo_2116};
  wire [7:0]    dataGroup_4_33 = dataGroup_lo_2116[303:296];
  wire [2047:0] dataGroup_lo_2117 = {dataGroup_lo_hi_2117, dataGroup_lo_lo_2117};
  wire [2047:0] dataGroup_hi_2117 = {dataGroup_hi_hi_2117, dataGroup_hi_lo_2117};
  wire [7:0]    dataGroup_5_33 = dataGroup_lo_2117[367:360];
  wire [2047:0] dataGroup_lo_2118 = {dataGroup_lo_hi_2118, dataGroup_lo_lo_2118};
  wire [2047:0] dataGroup_hi_2118 = {dataGroup_hi_hi_2118, dataGroup_hi_lo_2118};
  wire [7:0]    dataGroup_6_33 = dataGroup_lo_2118[431:424];
  wire [2047:0] dataGroup_lo_2119 = {dataGroup_lo_hi_2119, dataGroup_lo_lo_2119};
  wire [2047:0] dataGroup_hi_2119 = {dataGroup_hi_hi_2119, dataGroup_hi_lo_2119};
  wire [7:0]    dataGroup_7_33 = dataGroup_lo_2119[495:488];
  wire [2047:0] dataGroup_lo_2120 = {dataGroup_lo_hi_2120, dataGroup_lo_lo_2120};
  wire [2047:0] dataGroup_hi_2120 = {dataGroup_hi_hi_2120, dataGroup_hi_lo_2120};
  wire [7:0]    dataGroup_8_33 = dataGroup_lo_2120[559:552];
  wire [2047:0] dataGroup_lo_2121 = {dataGroup_lo_hi_2121, dataGroup_lo_lo_2121};
  wire [2047:0] dataGroup_hi_2121 = {dataGroup_hi_hi_2121, dataGroup_hi_lo_2121};
  wire [7:0]    dataGroup_9_33 = dataGroup_lo_2121[623:616];
  wire [2047:0] dataGroup_lo_2122 = {dataGroup_lo_hi_2122, dataGroup_lo_lo_2122};
  wire [2047:0] dataGroup_hi_2122 = {dataGroup_hi_hi_2122, dataGroup_hi_lo_2122};
  wire [7:0]    dataGroup_10_33 = dataGroup_lo_2122[687:680];
  wire [2047:0] dataGroup_lo_2123 = {dataGroup_lo_hi_2123, dataGroup_lo_lo_2123};
  wire [2047:0] dataGroup_hi_2123 = {dataGroup_hi_hi_2123, dataGroup_hi_lo_2123};
  wire [7:0]    dataGroup_11_33 = dataGroup_lo_2123[751:744];
  wire [2047:0] dataGroup_lo_2124 = {dataGroup_lo_hi_2124, dataGroup_lo_lo_2124};
  wire [2047:0] dataGroup_hi_2124 = {dataGroup_hi_hi_2124, dataGroup_hi_lo_2124};
  wire [7:0]    dataGroup_12_33 = dataGroup_lo_2124[815:808];
  wire [2047:0] dataGroup_lo_2125 = {dataGroup_lo_hi_2125, dataGroup_lo_lo_2125};
  wire [2047:0] dataGroup_hi_2125 = {dataGroup_hi_hi_2125, dataGroup_hi_lo_2125};
  wire [7:0]    dataGroup_13_33 = dataGroup_lo_2125[879:872];
  wire [2047:0] dataGroup_lo_2126 = {dataGroup_lo_hi_2126, dataGroup_lo_lo_2126};
  wire [2047:0] dataGroup_hi_2126 = {dataGroup_hi_hi_2126, dataGroup_hi_lo_2126};
  wire [7:0]    dataGroup_14_33 = dataGroup_lo_2126[943:936];
  wire [2047:0] dataGroup_lo_2127 = {dataGroup_lo_hi_2127, dataGroup_lo_lo_2127};
  wire [2047:0] dataGroup_hi_2127 = {dataGroup_hi_hi_2127, dataGroup_hi_lo_2127};
  wire [7:0]    dataGroup_15_33 = dataGroup_lo_2127[1007:1000];
  wire [2047:0] dataGroup_lo_2128 = {dataGroup_lo_hi_2128, dataGroup_lo_lo_2128};
  wire [2047:0] dataGroup_hi_2128 = {dataGroup_hi_hi_2128, dataGroup_hi_lo_2128};
  wire [7:0]    dataGroup_16_33 = dataGroup_lo_2128[1071:1064];
  wire [2047:0] dataGroup_lo_2129 = {dataGroup_lo_hi_2129, dataGroup_lo_lo_2129};
  wire [2047:0] dataGroup_hi_2129 = {dataGroup_hi_hi_2129, dataGroup_hi_lo_2129};
  wire [7:0]    dataGroup_17_33 = dataGroup_lo_2129[1135:1128];
  wire [2047:0] dataGroup_lo_2130 = {dataGroup_lo_hi_2130, dataGroup_lo_lo_2130};
  wire [2047:0] dataGroup_hi_2130 = {dataGroup_hi_hi_2130, dataGroup_hi_lo_2130};
  wire [7:0]    dataGroup_18_33 = dataGroup_lo_2130[1199:1192];
  wire [2047:0] dataGroup_lo_2131 = {dataGroup_lo_hi_2131, dataGroup_lo_lo_2131};
  wire [2047:0] dataGroup_hi_2131 = {dataGroup_hi_hi_2131, dataGroup_hi_lo_2131};
  wire [7:0]    dataGroup_19_33 = dataGroup_lo_2131[1263:1256];
  wire [2047:0] dataGroup_lo_2132 = {dataGroup_lo_hi_2132, dataGroup_lo_lo_2132};
  wire [2047:0] dataGroup_hi_2132 = {dataGroup_hi_hi_2132, dataGroup_hi_lo_2132};
  wire [7:0]    dataGroup_20_33 = dataGroup_lo_2132[1327:1320];
  wire [2047:0] dataGroup_lo_2133 = {dataGroup_lo_hi_2133, dataGroup_lo_lo_2133};
  wire [2047:0] dataGroup_hi_2133 = {dataGroup_hi_hi_2133, dataGroup_hi_lo_2133};
  wire [7:0]    dataGroup_21_33 = dataGroup_lo_2133[1391:1384];
  wire [2047:0] dataGroup_lo_2134 = {dataGroup_lo_hi_2134, dataGroup_lo_lo_2134};
  wire [2047:0] dataGroup_hi_2134 = {dataGroup_hi_hi_2134, dataGroup_hi_lo_2134};
  wire [7:0]    dataGroup_22_33 = dataGroup_lo_2134[1455:1448];
  wire [2047:0] dataGroup_lo_2135 = {dataGroup_lo_hi_2135, dataGroup_lo_lo_2135};
  wire [2047:0] dataGroup_hi_2135 = {dataGroup_hi_hi_2135, dataGroup_hi_lo_2135};
  wire [7:0]    dataGroup_23_33 = dataGroup_lo_2135[1519:1512];
  wire [2047:0] dataGroup_lo_2136 = {dataGroup_lo_hi_2136, dataGroup_lo_lo_2136};
  wire [2047:0] dataGroup_hi_2136 = {dataGroup_hi_hi_2136, dataGroup_hi_lo_2136};
  wire [7:0]    dataGroup_24_33 = dataGroup_lo_2136[1583:1576];
  wire [2047:0] dataGroup_lo_2137 = {dataGroup_lo_hi_2137, dataGroup_lo_lo_2137};
  wire [2047:0] dataGroup_hi_2137 = {dataGroup_hi_hi_2137, dataGroup_hi_lo_2137};
  wire [7:0]    dataGroup_25_33 = dataGroup_lo_2137[1647:1640];
  wire [2047:0] dataGroup_lo_2138 = {dataGroup_lo_hi_2138, dataGroup_lo_lo_2138};
  wire [2047:0] dataGroup_hi_2138 = {dataGroup_hi_hi_2138, dataGroup_hi_lo_2138};
  wire [7:0]    dataGroup_26_33 = dataGroup_lo_2138[1711:1704];
  wire [2047:0] dataGroup_lo_2139 = {dataGroup_lo_hi_2139, dataGroup_lo_lo_2139};
  wire [2047:0] dataGroup_hi_2139 = {dataGroup_hi_hi_2139, dataGroup_hi_lo_2139};
  wire [7:0]    dataGroup_27_33 = dataGroup_lo_2139[1775:1768];
  wire [2047:0] dataGroup_lo_2140 = {dataGroup_lo_hi_2140, dataGroup_lo_lo_2140};
  wire [2047:0] dataGroup_hi_2140 = {dataGroup_hi_hi_2140, dataGroup_hi_lo_2140};
  wire [7:0]    dataGroup_28_33 = dataGroup_lo_2140[1839:1832];
  wire [2047:0] dataGroup_lo_2141 = {dataGroup_lo_hi_2141, dataGroup_lo_lo_2141};
  wire [2047:0] dataGroup_hi_2141 = {dataGroup_hi_hi_2141, dataGroup_hi_lo_2141};
  wire [7:0]    dataGroup_29_33 = dataGroup_lo_2141[1903:1896];
  wire [2047:0] dataGroup_lo_2142 = {dataGroup_lo_hi_2142, dataGroup_lo_lo_2142};
  wire [2047:0] dataGroup_hi_2142 = {dataGroup_hi_hi_2142, dataGroup_hi_lo_2142};
  wire [7:0]    dataGroup_30_33 = dataGroup_lo_2142[1967:1960];
  wire [2047:0] dataGroup_lo_2143 = {dataGroup_lo_hi_2143, dataGroup_lo_lo_2143};
  wire [2047:0] dataGroup_hi_2143 = {dataGroup_hi_hi_2143, dataGroup_hi_lo_2143};
  wire [7:0]    dataGroup_31_33 = dataGroup_lo_2143[2031:2024];
  wire [2047:0] dataGroup_lo_2144 = {dataGroup_lo_hi_2144, dataGroup_lo_lo_2144};
  wire [2047:0] dataGroup_hi_2144 = {dataGroup_hi_hi_2144, dataGroup_hi_lo_2144};
  wire [7:0]    dataGroup_32_33 = dataGroup_hi_2144[47:40];
  wire [2047:0] dataGroup_lo_2145 = {dataGroup_lo_hi_2145, dataGroup_lo_lo_2145};
  wire [2047:0] dataGroup_hi_2145 = {dataGroup_hi_hi_2145, dataGroup_hi_lo_2145};
  wire [7:0]    dataGroup_33_33 = dataGroup_hi_2145[111:104];
  wire [2047:0] dataGroup_lo_2146 = {dataGroup_lo_hi_2146, dataGroup_lo_lo_2146};
  wire [2047:0] dataGroup_hi_2146 = {dataGroup_hi_hi_2146, dataGroup_hi_lo_2146};
  wire [7:0]    dataGroup_34_33 = dataGroup_hi_2146[175:168];
  wire [2047:0] dataGroup_lo_2147 = {dataGroup_lo_hi_2147, dataGroup_lo_lo_2147};
  wire [2047:0] dataGroup_hi_2147 = {dataGroup_hi_hi_2147, dataGroup_hi_lo_2147};
  wire [7:0]    dataGroup_35_33 = dataGroup_hi_2147[239:232];
  wire [2047:0] dataGroup_lo_2148 = {dataGroup_lo_hi_2148, dataGroup_lo_lo_2148};
  wire [2047:0] dataGroup_hi_2148 = {dataGroup_hi_hi_2148, dataGroup_hi_lo_2148};
  wire [7:0]    dataGroup_36_33 = dataGroup_hi_2148[303:296];
  wire [2047:0] dataGroup_lo_2149 = {dataGroup_lo_hi_2149, dataGroup_lo_lo_2149};
  wire [2047:0] dataGroup_hi_2149 = {dataGroup_hi_hi_2149, dataGroup_hi_lo_2149};
  wire [7:0]    dataGroup_37_33 = dataGroup_hi_2149[367:360];
  wire [2047:0] dataGroup_lo_2150 = {dataGroup_lo_hi_2150, dataGroup_lo_lo_2150};
  wire [2047:0] dataGroup_hi_2150 = {dataGroup_hi_hi_2150, dataGroup_hi_lo_2150};
  wire [7:0]    dataGroup_38_33 = dataGroup_hi_2150[431:424];
  wire [2047:0] dataGroup_lo_2151 = {dataGroup_lo_hi_2151, dataGroup_lo_lo_2151};
  wire [2047:0] dataGroup_hi_2151 = {dataGroup_hi_hi_2151, dataGroup_hi_lo_2151};
  wire [7:0]    dataGroup_39_33 = dataGroup_hi_2151[495:488];
  wire [2047:0] dataGroup_lo_2152 = {dataGroup_lo_hi_2152, dataGroup_lo_lo_2152};
  wire [2047:0] dataGroup_hi_2152 = {dataGroup_hi_hi_2152, dataGroup_hi_lo_2152};
  wire [7:0]    dataGroup_40_33 = dataGroup_hi_2152[559:552];
  wire [2047:0] dataGroup_lo_2153 = {dataGroup_lo_hi_2153, dataGroup_lo_lo_2153};
  wire [2047:0] dataGroup_hi_2153 = {dataGroup_hi_hi_2153, dataGroup_hi_lo_2153};
  wire [7:0]    dataGroup_41_33 = dataGroup_hi_2153[623:616];
  wire [2047:0] dataGroup_lo_2154 = {dataGroup_lo_hi_2154, dataGroup_lo_lo_2154};
  wire [2047:0] dataGroup_hi_2154 = {dataGroup_hi_hi_2154, dataGroup_hi_lo_2154};
  wire [7:0]    dataGroup_42_33 = dataGroup_hi_2154[687:680];
  wire [2047:0] dataGroup_lo_2155 = {dataGroup_lo_hi_2155, dataGroup_lo_lo_2155};
  wire [2047:0] dataGroup_hi_2155 = {dataGroup_hi_hi_2155, dataGroup_hi_lo_2155};
  wire [7:0]    dataGroup_43_33 = dataGroup_hi_2155[751:744];
  wire [2047:0] dataGroup_lo_2156 = {dataGroup_lo_hi_2156, dataGroup_lo_lo_2156};
  wire [2047:0] dataGroup_hi_2156 = {dataGroup_hi_hi_2156, dataGroup_hi_lo_2156};
  wire [7:0]    dataGroup_44_33 = dataGroup_hi_2156[815:808];
  wire [2047:0] dataGroup_lo_2157 = {dataGroup_lo_hi_2157, dataGroup_lo_lo_2157};
  wire [2047:0] dataGroup_hi_2157 = {dataGroup_hi_hi_2157, dataGroup_hi_lo_2157};
  wire [7:0]    dataGroup_45_33 = dataGroup_hi_2157[879:872];
  wire [2047:0] dataGroup_lo_2158 = {dataGroup_lo_hi_2158, dataGroup_lo_lo_2158};
  wire [2047:0] dataGroup_hi_2158 = {dataGroup_hi_hi_2158, dataGroup_hi_lo_2158};
  wire [7:0]    dataGroup_46_33 = dataGroup_hi_2158[943:936];
  wire [2047:0] dataGroup_lo_2159 = {dataGroup_lo_hi_2159, dataGroup_lo_lo_2159};
  wire [2047:0] dataGroup_hi_2159 = {dataGroup_hi_hi_2159, dataGroup_hi_lo_2159};
  wire [7:0]    dataGroup_47_33 = dataGroup_hi_2159[1007:1000];
  wire [2047:0] dataGroup_lo_2160 = {dataGroup_lo_hi_2160, dataGroup_lo_lo_2160};
  wire [2047:0] dataGroup_hi_2160 = {dataGroup_hi_hi_2160, dataGroup_hi_lo_2160};
  wire [7:0]    dataGroup_48_33 = dataGroup_hi_2160[1071:1064];
  wire [2047:0] dataGroup_lo_2161 = {dataGroup_lo_hi_2161, dataGroup_lo_lo_2161};
  wire [2047:0] dataGroup_hi_2161 = {dataGroup_hi_hi_2161, dataGroup_hi_lo_2161};
  wire [7:0]    dataGroup_49_33 = dataGroup_hi_2161[1135:1128];
  wire [2047:0] dataGroup_lo_2162 = {dataGroup_lo_hi_2162, dataGroup_lo_lo_2162};
  wire [2047:0] dataGroup_hi_2162 = {dataGroup_hi_hi_2162, dataGroup_hi_lo_2162};
  wire [7:0]    dataGroup_50_33 = dataGroup_hi_2162[1199:1192];
  wire [2047:0] dataGroup_lo_2163 = {dataGroup_lo_hi_2163, dataGroup_lo_lo_2163};
  wire [2047:0] dataGroup_hi_2163 = {dataGroup_hi_hi_2163, dataGroup_hi_lo_2163};
  wire [7:0]    dataGroup_51_33 = dataGroup_hi_2163[1263:1256];
  wire [2047:0] dataGroup_lo_2164 = {dataGroup_lo_hi_2164, dataGroup_lo_lo_2164};
  wire [2047:0] dataGroup_hi_2164 = {dataGroup_hi_hi_2164, dataGroup_hi_lo_2164};
  wire [7:0]    dataGroup_52_33 = dataGroup_hi_2164[1327:1320];
  wire [2047:0] dataGroup_lo_2165 = {dataGroup_lo_hi_2165, dataGroup_lo_lo_2165};
  wire [2047:0] dataGroup_hi_2165 = {dataGroup_hi_hi_2165, dataGroup_hi_lo_2165};
  wire [7:0]    dataGroup_53_33 = dataGroup_hi_2165[1391:1384];
  wire [2047:0] dataGroup_lo_2166 = {dataGroup_lo_hi_2166, dataGroup_lo_lo_2166};
  wire [2047:0] dataGroup_hi_2166 = {dataGroup_hi_hi_2166, dataGroup_hi_lo_2166};
  wire [7:0]    dataGroup_54_33 = dataGroup_hi_2166[1455:1448];
  wire [2047:0] dataGroup_lo_2167 = {dataGroup_lo_hi_2167, dataGroup_lo_lo_2167};
  wire [2047:0] dataGroup_hi_2167 = {dataGroup_hi_hi_2167, dataGroup_hi_lo_2167};
  wire [7:0]    dataGroup_55_33 = dataGroup_hi_2167[1519:1512];
  wire [2047:0] dataGroup_lo_2168 = {dataGroup_lo_hi_2168, dataGroup_lo_lo_2168};
  wire [2047:0] dataGroup_hi_2168 = {dataGroup_hi_hi_2168, dataGroup_hi_lo_2168};
  wire [7:0]    dataGroup_56_33 = dataGroup_hi_2168[1583:1576];
  wire [2047:0] dataGroup_lo_2169 = {dataGroup_lo_hi_2169, dataGroup_lo_lo_2169};
  wire [2047:0] dataGroup_hi_2169 = {dataGroup_hi_hi_2169, dataGroup_hi_lo_2169};
  wire [7:0]    dataGroup_57_33 = dataGroup_hi_2169[1647:1640];
  wire [2047:0] dataGroup_lo_2170 = {dataGroup_lo_hi_2170, dataGroup_lo_lo_2170};
  wire [2047:0] dataGroup_hi_2170 = {dataGroup_hi_hi_2170, dataGroup_hi_lo_2170};
  wire [7:0]    dataGroup_58_33 = dataGroup_hi_2170[1711:1704];
  wire [2047:0] dataGroup_lo_2171 = {dataGroup_lo_hi_2171, dataGroup_lo_lo_2171};
  wire [2047:0] dataGroup_hi_2171 = {dataGroup_hi_hi_2171, dataGroup_hi_lo_2171};
  wire [7:0]    dataGroup_59_33 = dataGroup_hi_2171[1775:1768];
  wire [2047:0] dataGroup_lo_2172 = {dataGroup_lo_hi_2172, dataGroup_lo_lo_2172};
  wire [2047:0] dataGroup_hi_2172 = {dataGroup_hi_hi_2172, dataGroup_hi_lo_2172};
  wire [7:0]    dataGroup_60_33 = dataGroup_hi_2172[1839:1832];
  wire [2047:0] dataGroup_lo_2173 = {dataGroup_lo_hi_2173, dataGroup_lo_lo_2173};
  wire [2047:0] dataGroup_hi_2173 = {dataGroup_hi_hi_2173, dataGroup_hi_lo_2173};
  wire [7:0]    dataGroup_61_33 = dataGroup_hi_2173[1903:1896];
  wire [2047:0] dataGroup_lo_2174 = {dataGroup_lo_hi_2174, dataGroup_lo_lo_2174};
  wire [2047:0] dataGroup_hi_2174 = {dataGroup_hi_hi_2174, dataGroup_hi_lo_2174};
  wire [7:0]    dataGroup_62_33 = dataGroup_hi_2174[1967:1960];
  wire [2047:0] dataGroup_lo_2175 = {dataGroup_lo_hi_2175, dataGroup_lo_lo_2175};
  wire [2047:0] dataGroup_hi_2175 = {dataGroup_hi_hi_2175, dataGroup_hi_lo_2175};
  wire [7:0]    dataGroup_63_33 = dataGroup_hi_2175[2031:2024];
  wire [15:0]   res_lo_lo_lo_lo_lo_33 = {dataGroup_1_33, dataGroup_0_33};
  wire [15:0]   res_lo_lo_lo_lo_hi_33 = {dataGroup_3_33, dataGroup_2_33};
  wire [31:0]   res_lo_lo_lo_lo_33 = {res_lo_lo_lo_lo_hi_33, res_lo_lo_lo_lo_lo_33};
  wire [15:0]   res_lo_lo_lo_hi_lo_33 = {dataGroup_5_33, dataGroup_4_33};
  wire [15:0]   res_lo_lo_lo_hi_hi_33 = {dataGroup_7_33, dataGroup_6_33};
  wire [31:0]   res_lo_lo_lo_hi_33 = {res_lo_lo_lo_hi_hi_33, res_lo_lo_lo_hi_lo_33};
  wire [63:0]   res_lo_lo_lo_33 = {res_lo_lo_lo_hi_33, res_lo_lo_lo_lo_33};
  wire [15:0]   res_lo_lo_hi_lo_lo_33 = {dataGroup_9_33, dataGroup_8_33};
  wire [15:0]   res_lo_lo_hi_lo_hi_33 = {dataGroup_11_33, dataGroup_10_33};
  wire [31:0]   res_lo_lo_hi_lo_33 = {res_lo_lo_hi_lo_hi_33, res_lo_lo_hi_lo_lo_33};
  wire [15:0]   res_lo_lo_hi_hi_lo_33 = {dataGroup_13_33, dataGroup_12_33};
  wire [15:0]   res_lo_lo_hi_hi_hi_33 = {dataGroup_15_33, dataGroup_14_33};
  wire [31:0]   res_lo_lo_hi_hi_33 = {res_lo_lo_hi_hi_hi_33, res_lo_lo_hi_hi_lo_33};
  wire [63:0]   res_lo_lo_hi_33 = {res_lo_lo_hi_hi_33, res_lo_lo_hi_lo_33};
  wire [127:0]  res_lo_lo_33 = {res_lo_lo_hi_33, res_lo_lo_lo_33};
  wire [15:0]   res_lo_hi_lo_lo_lo_33 = {dataGroup_17_33, dataGroup_16_33};
  wire [15:0]   res_lo_hi_lo_lo_hi_33 = {dataGroup_19_33, dataGroup_18_33};
  wire [31:0]   res_lo_hi_lo_lo_33 = {res_lo_hi_lo_lo_hi_33, res_lo_hi_lo_lo_lo_33};
  wire [15:0]   res_lo_hi_lo_hi_lo_33 = {dataGroup_21_33, dataGroup_20_33};
  wire [15:0]   res_lo_hi_lo_hi_hi_33 = {dataGroup_23_33, dataGroup_22_33};
  wire [31:0]   res_lo_hi_lo_hi_33 = {res_lo_hi_lo_hi_hi_33, res_lo_hi_lo_hi_lo_33};
  wire [63:0]   res_lo_hi_lo_33 = {res_lo_hi_lo_hi_33, res_lo_hi_lo_lo_33};
  wire [15:0]   res_lo_hi_hi_lo_lo_33 = {dataGroup_25_33, dataGroup_24_33};
  wire [15:0]   res_lo_hi_hi_lo_hi_33 = {dataGroup_27_33, dataGroup_26_33};
  wire [31:0]   res_lo_hi_hi_lo_33 = {res_lo_hi_hi_lo_hi_33, res_lo_hi_hi_lo_lo_33};
  wire [15:0]   res_lo_hi_hi_hi_lo_33 = {dataGroup_29_33, dataGroup_28_33};
  wire [15:0]   res_lo_hi_hi_hi_hi_33 = {dataGroup_31_33, dataGroup_30_33};
  wire [31:0]   res_lo_hi_hi_hi_33 = {res_lo_hi_hi_hi_hi_33, res_lo_hi_hi_hi_lo_33};
  wire [63:0]   res_lo_hi_hi_33 = {res_lo_hi_hi_hi_33, res_lo_hi_hi_lo_33};
  wire [127:0]  res_lo_hi_33 = {res_lo_hi_hi_33, res_lo_hi_lo_33};
  wire [255:0]  res_lo_33 = {res_lo_hi_33, res_lo_lo_33};
  wire [15:0]   res_hi_lo_lo_lo_lo_33 = {dataGroup_33_33, dataGroup_32_33};
  wire [15:0]   res_hi_lo_lo_lo_hi_33 = {dataGroup_35_33, dataGroup_34_33};
  wire [31:0]   res_hi_lo_lo_lo_33 = {res_hi_lo_lo_lo_hi_33, res_hi_lo_lo_lo_lo_33};
  wire [15:0]   res_hi_lo_lo_hi_lo_33 = {dataGroup_37_33, dataGroup_36_33};
  wire [15:0]   res_hi_lo_lo_hi_hi_33 = {dataGroup_39_33, dataGroup_38_33};
  wire [31:0]   res_hi_lo_lo_hi_33 = {res_hi_lo_lo_hi_hi_33, res_hi_lo_lo_hi_lo_33};
  wire [63:0]   res_hi_lo_lo_33 = {res_hi_lo_lo_hi_33, res_hi_lo_lo_lo_33};
  wire [15:0]   res_hi_lo_hi_lo_lo_33 = {dataGroup_41_33, dataGroup_40_33};
  wire [15:0]   res_hi_lo_hi_lo_hi_33 = {dataGroup_43_33, dataGroup_42_33};
  wire [31:0]   res_hi_lo_hi_lo_33 = {res_hi_lo_hi_lo_hi_33, res_hi_lo_hi_lo_lo_33};
  wire [15:0]   res_hi_lo_hi_hi_lo_33 = {dataGroup_45_33, dataGroup_44_33};
  wire [15:0]   res_hi_lo_hi_hi_hi_33 = {dataGroup_47_33, dataGroup_46_33};
  wire [31:0]   res_hi_lo_hi_hi_33 = {res_hi_lo_hi_hi_hi_33, res_hi_lo_hi_hi_lo_33};
  wire [63:0]   res_hi_lo_hi_33 = {res_hi_lo_hi_hi_33, res_hi_lo_hi_lo_33};
  wire [127:0]  res_hi_lo_33 = {res_hi_lo_hi_33, res_hi_lo_lo_33};
  wire [15:0]   res_hi_hi_lo_lo_lo_33 = {dataGroup_49_33, dataGroup_48_33};
  wire [15:0]   res_hi_hi_lo_lo_hi_33 = {dataGroup_51_33, dataGroup_50_33};
  wire [31:0]   res_hi_hi_lo_lo_33 = {res_hi_hi_lo_lo_hi_33, res_hi_hi_lo_lo_lo_33};
  wire [15:0]   res_hi_hi_lo_hi_lo_33 = {dataGroup_53_33, dataGroup_52_33};
  wire [15:0]   res_hi_hi_lo_hi_hi_33 = {dataGroup_55_33, dataGroup_54_33};
  wire [31:0]   res_hi_hi_lo_hi_33 = {res_hi_hi_lo_hi_hi_33, res_hi_hi_lo_hi_lo_33};
  wire [63:0]   res_hi_hi_lo_33 = {res_hi_hi_lo_hi_33, res_hi_hi_lo_lo_33};
  wire [15:0]   res_hi_hi_hi_lo_lo_33 = {dataGroup_57_33, dataGroup_56_33};
  wire [15:0]   res_hi_hi_hi_lo_hi_33 = {dataGroup_59_33, dataGroup_58_33};
  wire [31:0]   res_hi_hi_hi_lo_33 = {res_hi_hi_hi_lo_hi_33, res_hi_hi_hi_lo_lo_33};
  wire [15:0]   res_hi_hi_hi_hi_lo_33 = {dataGroup_61_33, dataGroup_60_33};
  wire [15:0]   res_hi_hi_hi_hi_hi_33 = {dataGroup_63_33, dataGroup_62_33};
  wire [31:0]   res_hi_hi_hi_hi_33 = {res_hi_hi_hi_hi_hi_33, res_hi_hi_hi_hi_lo_33};
  wire [63:0]   res_hi_hi_hi_33 = {res_hi_hi_hi_hi_33, res_hi_hi_hi_lo_33};
  wire [127:0]  res_hi_hi_33 = {res_hi_hi_hi_33, res_hi_hi_lo_33};
  wire [255:0]  res_hi_33 = {res_hi_hi_33, res_hi_lo_33};
  wire [511:0]  res_61 = {res_hi_33, res_lo_33};
  wire [2047:0] dataGroup_lo_2176 = {dataGroup_lo_hi_2176, dataGroup_lo_lo_2176};
  wire [2047:0] dataGroup_hi_2176 = {dataGroup_hi_hi_2176, dataGroup_hi_lo_2176};
  wire [7:0]    dataGroup_0_34 = dataGroup_lo_2176[55:48];
  wire [2047:0] dataGroup_lo_2177 = {dataGroup_lo_hi_2177, dataGroup_lo_lo_2177};
  wire [2047:0] dataGroup_hi_2177 = {dataGroup_hi_hi_2177, dataGroup_hi_lo_2177};
  wire [7:0]    dataGroup_1_34 = dataGroup_lo_2177[119:112];
  wire [2047:0] dataGroup_lo_2178 = {dataGroup_lo_hi_2178, dataGroup_lo_lo_2178};
  wire [2047:0] dataGroup_hi_2178 = {dataGroup_hi_hi_2178, dataGroup_hi_lo_2178};
  wire [7:0]    dataGroup_2_34 = dataGroup_lo_2178[183:176];
  wire [2047:0] dataGroup_lo_2179 = {dataGroup_lo_hi_2179, dataGroup_lo_lo_2179};
  wire [2047:0] dataGroup_hi_2179 = {dataGroup_hi_hi_2179, dataGroup_hi_lo_2179};
  wire [7:0]    dataGroup_3_34 = dataGroup_lo_2179[247:240];
  wire [2047:0] dataGroup_lo_2180 = {dataGroup_lo_hi_2180, dataGroup_lo_lo_2180};
  wire [2047:0] dataGroup_hi_2180 = {dataGroup_hi_hi_2180, dataGroup_hi_lo_2180};
  wire [7:0]    dataGroup_4_34 = dataGroup_lo_2180[311:304];
  wire [2047:0] dataGroup_lo_2181 = {dataGroup_lo_hi_2181, dataGroup_lo_lo_2181};
  wire [2047:0] dataGroup_hi_2181 = {dataGroup_hi_hi_2181, dataGroup_hi_lo_2181};
  wire [7:0]    dataGroup_5_34 = dataGroup_lo_2181[375:368];
  wire [2047:0] dataGroup_lo_2182 = {dataGroup_lo_hi_2182, dataGroup_lo_lo_2182};
  wire [2047:0] dataGroup_hi_2182 = {dataGroup_hi_hi_2182, dataGroup_hi_lo_2182};
  wire [7:0]    dataGroup_6_34 = dataGroup_lo_2182[439:432];
  wire [2047:0] dataGroup_lo_2183 = {dataGroup_lo_hi_2183, dataGroup_lo_lo_2183};
  wire [2047:0] dataGroup_hi_2183 = {dataGroup_hi_hi_2183, dataGroup_hi_lo_2183};
  wire [7:0]    dataGroup_7_34 = dataGroup_lo_2183[503:496];
  wire [2047:0] dataGroup_lo_2184 = {dataGroup_lo_hi_2184, dataGroup_lo_lo_2184};
  wire [2047:0] dataGroup_hi_2184 = {dataGroup_hi_hi_2184, dataGroup_hi_lo_2184};
  wire [7:0]    dataGroup_8_34 = dataGroup_lo_2184[567:560];
  wire [2047:0] dataGroup_lo_2185 = {dataGroup_lo_hi_2185, dataGroup_lo_lo_2185};
  wire [2047:0] dataGroup_hi_2185 = {dataGroup_hi_hi_2185, dataGroup_hi_lo_2185};
  wire [7:0]    dataGroup_9_34 = dataGroup_lo_2185[631:624];
  wire [2047:0] dataGroup_lo_2186 = {dataGroup_lo_hi_2186, dataGroup_lo_lo_2186};
  wire [2047:0] dataGroup_hi_2186 = {dataGroup_hi_hi_2186, dataGroup_hi_lo_2186};
  wire [7:0]    dataGroup_10_34 = dataGroup_lo_2186[695:688];
  wire [2047:0] dataGroup_lo_2187 = {dataGroup_lo_hi_2187, dataGroup_lo_lo_2187};
  wire [2047:0] dataGroup_hi_2187 = {dataGroup_hi_hi_2187, dataGroup_hi_lo_2187};
  wire [7:0]    dataGroup_11_34 = dataGroup_lo_2187[759:752];
  wire [2047:0] dataGroup_lo_2188 = {dataGroup_lo_hi_2188, dataGroup_lo_lo_2188};
  wire [2047:0] dataGroup_hi_2188 = {dataGroup_hi_hi_2188, dataGroup_hi_lo_2188};
  wire [7:0]    dataGroup_12_34 = dataGroup_lo_2188[823:816];
  wire [2047:0] dataGroup_lo_2189 = {dataGroup_lo_hi_2189, dataGroup_lo_lo_2189};
  wire [2047:0] dataGroup_hi_2189 = {dataGroup_hi_hi_2189, dataGroup_hi_lo_2189};
  wire [7:0]    dataGroup_13_34 = dataGroup_lo_2189[887:880];
  wire [2047:0] dataGroup_lo_2190 = {dataGroup_lo_hi_2190, dataGroup_lo_lo_2190};
  wire [2047:0] dataGroup_hi_2190 = {dataGroup_hi_hi_2190, dataGroup_hi_lo_2190};
  wire [7:0]    dataGroup_14_34 = dataGroup_lo_2190[951:944];
  wire [2047:0] dataGroup_lo_2191 = {dataGroup_lo_hi_2191, dataGroup_lo_lo_2191};
  wire [2047:0] dataGroup_hi_2191 = {dataGroup_hi_hi_2191, dataGroup_hi_lo_2191};
  wire [7:0]    dataGroup_15_34 = dataGroup_lo_2191[1015:1008];
  wire [2047:0] dataGroup_lo_2192 = {dataGroup_lo_hi_2192, dataGroup_lo_lo_2192};
  wire [2047:0] dataGroup_hi_2192 = {dataGroup_hi_hi_2192, dataGroup_hi_lo_2192};
  wire [7:0]    dataGroup_16_34 = dataGroup_lo_2192[1079:1072];
  wire [2047:0] dataGroup_lo_2193 = {dataGroup_lo_hi_2193, dataGroup_lo_lo_2193};
  wire [2047:0] dataGroup_hi_2193 = {dataGroup_hi_hi_2193, dataGroup_hi_lo_2193};
  wire [7:0]    dataGroup_17_34 = dataGroup_lo_2193[1143:1136];
  wire [2047:0] dataGroup_lo_2194 = {dataGroup_lo_hi_2194, dataGroup_lo_lo_2194};
  wire [2047:0] dataGroup_hi_2194 = {dataGroup_hi_hi_2194, dataGroup_hi_lo_2194};
  wire [7:0]    dataGroup_18_34 = dataGroup_lo_2194[1207:1200];
  wire [2047:0] dataGroup_lo_2195 = {dataGroup_lo_hi_2195, dataGroup_lo_lo_2195};
  wire [2047:0] dataGroup_hi_2195 = {dataGroup_hi_hi_2195, dataGroup_hi_lo_2195};
  wire [7:0]    dataGroup_19_34 = dataGroup_lo_2195[1271:1264];
  wire [2047:0] dataGroup_lo_2196 = {dataGroup_lo_hi_2196, dataGroup_lo_lo_2196};
  wire [2047:0] dataGroup_hi_2196 = {dataGroup_hi_hi_2196, dataGroup_hi_lo_2196};
  wire [7:0]    dataGroup_20_34 = dataGroup_lo_2196[1335:1328];
  wire [2047:0] dataGroup_lo_2197 = {dataGroup_lo_hi_2197, dataGroup_lo_lo_2197};
  wire [2047:0] dataGroup_hi_2197 = {dataGroup_hi_hi_2197, dataGroup_hi_lo_2197};
  wire [7:0]    dataGroup_21_34 = dataGroup_lo_2197[1399:1392];
  wire [2047:0] dataGroup_lo_2198 = {dataGroup_lo_hi_2198, dataGroup_lo_lo_2198};
  wire [2047:0] dataGroup_hi_2198 = {dataGroup_hi_hi_2198, dataGroup_hi_lo_2198};
  wire [7:0]    dataGroup_22_34 = dataGroup_lo_2198[1463:1456];
  wire [2047:0] dataGroup_lo_2199 = {dataGroup_lo_hi_2199, dataGroup_lo_lo_2199};
  wire [2047:0] dataGroup_hi_2199 = {dataGroup_hi_hi_2199, dataGroup_hi_lo_2199};
  wire [7:0]    dataGroup_23_34 = dataGroup_lo_2199[1527:1520];
  wire [2047:0] dataGroup_lo_2200 = {dataGroup_lo_hi_2200, dataGroup_lo_lo_2200};
  wire [2047:0] dataGroup_hi_2200 = {dataGroup_hi_hi_2200, dataGroup_hi_lo_2200};
  wire [7:0]    dataGroup_24_34 = dataGroup_lo_2200[1591:1584];
  wire [2047:0] dataGroup_lo_2201 = {dataGroup_lo_hi_2201, dataGroup_lo_lo_2201};
  wire [2047:0] dataGroup_hi_2201 = {dataGroup_hi_hi_2201, dataGroup_hi_lo_2201};
  wire [7:0]    dataGroup_25_34 = dataGroup_lo_2201[1655:1648];
  wire [2047:0] dataGroup_lo_2202 = {dataGroup_lo_hi_2202, dataGroup_lo_lo_2202};
  wire [2047:0] dataGroup_hi_2202 = {dataGroup_hi_hi_2202, dataGroup_hi_lo_2202};
  wire [7:0]    dataGroup_26_34 = dataGroup_lo_2202[1719:1712];
  wire [2047:0] dataGroup_lo_2203 = {dataGroup_lo_hi_2203, dataGroup_lo_lo_2203};
  wire [2047:0] dataGroup_hi_2203 = {dataGroup_hi_hi_2203, dataGroup_hi_lo_2203};
  wire [7:0]    dataGroup_27_34 = dataGroup_lo_2203[1783:1776];
  wire [2047:0] dataGroup_lo_2204 = {dataGroup_lo_hi_2204, dataGroup_lo_lo_2204};
  wire [2047:0] dataGroup_hi_2204 = {dataGroup_hi_hi_2204, dataGroup_hi_lo_2204};
  wire [7:0]    dataGroup_28_34 = dataGroup_lo_2204[1847:1840];
  wire [2047:0] dataGroup_lo_2205 = {dataGroup_lo_hi_2205, dataGroup_lo_lo_2205};
  wire [2047:0] dataGroup_hi_2205 = {dataGroup_hi_hi_2205, dataGroup_hi_lo_2205};
  wire [7:0]    dataGroup_29_34 = dataGroup_lo_2205[1911:1904];
  wire [2047:0] dataGroup_lo_2206 = {dataGroup_lo_hi_2206, dataGroup_lo_lo_2206};
  wire [2047:0] dataGroup_hi_2206 = {dataGroup_hi_hi_2206, dataGroup_hi_lo_2206};
  wire [7:0]    dataGroup_30_34 = dataGroup_lo_2206[1975:1968];
  wire [2047:0] dataGroup_lo_2207 = {dataGroup_lo_hi_2207, dataGroup_lo_lo_2207};
  wire [2047:0] dataGroup_hi_2207 = {dataGroup_hi_hi_2207, dataGroup_hi_lo_2207};
  wire [7:0]    dataGroup_31_34 = dataGroup_lo_2207[2039:2032];
  wire [2047:0] dataGroup_lo_2208 = {dataGroup_lo_hi_2208, dataGroup_lo_lo_2208};
  wire [2047:0] dataGroup_hi_2208 = {dataGroup_hi_hi_2208, dataGroup_hi_lo_2208};
  wire [7:0]    dataGroup_32_34 = dataGroup_hi_2208[55:48];
  wire [2047:0] dataGroup_lo_2209 = {dataGroup_lo_hi_2209, dataGroup_lo_lo_2209};
  wire [2047:0] dataGroup_hi_2209 = {dataGroup_hi_hi_2209, dataGroup_hi_lo_2209};
  wire [7:0]    dataGroup_33_34 = dataGroup_hi_2209[119:112];
  wire [2047:0] dataGroup_lo_2210 = {dataGroup_lo_hi_2210, dataGroup_lo_lo_2210};
  wire [2047:0] dataGroup_hi_2210 = {dataGroup_hi_hi_2210, dataGroup_hi_lo_2210};
  wire [7:0]    dataGroup_34_34 = dataGroup_hi_2210[183:176];
  wire [2047:0] dataGroup_lo_2211 = {dataGroup_lo_hi_2211, dataGroup_lo_lo_2211};
  wire [2047:0] dataGroup_hi_2211 = {dataGroup_hi_hi_2211, dataGroup_hi_lo_2211};
  wire [7:0]    dataGroup_35_34 = dataGroup_hi_2211[247:240];
  wire [2047:0] dataGroup_lo_2212 = {dataGroup_lo_hi_2212, dataGroup_lo_lo_2212};
  wire [2047:0] dataGroup_hi_2212 = {dataGroup_hi_hi_2212, dataGroup_hi_lo_2212};
  wire [7:0]    dataGroup_36_34 = dataGroup_hi_2212[311:304];
  wire [2047:0] dataGroup_lo_2213 = {dataGroup_lo_hi_2213, dataGroup_lo_lo_2213};
  wire [2047:0] dataGroup_hi_2213 = {dataGroup_hi_hi_2213, dataGroup_hi_lo_2213};
  wire [7:0]    dataGroup_37_34 = dataGroup_hi_2213[375:368];
  wire [2047:0] dataGroup_lo_2214 = {dataGroup_lo_hi_2214, dataGroup_lo_lo_2214};
  wire [2047:0] dataGroup_hi_2214 = {dataGroup_hi_hi_2214, dataGroup_hi_lo_2214};
  wire [7:0]    dataGroup_38_34 = dataGroup_hi_2214[439:432];
  wire [2047:0] dataGroup_lo_2215 = {dataGroup_lo_hi_2215, dataGroup_lo_lo_2215};
  wire [2047:0] dataGroup_hi_2215 = {dataGroup_hi_hi_2215, dataGroup_hi_lo_2215};
  wire [7:0]    dataGroup_39_34 = dataGroup_hi_2215[503:496];
  wire [2047:0] dataGroup_lo_2216 = {dataGroup_lo_hi_2216, dataGroup_lo_lo_2216};
  wire [2047:0] dataGroup_hi_2216 = {dataGroup_hi_hi_2216, dataGroup_hi_lo_2216};
  wire [7:0]    dataGroup_40_34 = dataGroup_hi_2216[567:560];
  wire [2047:0] dataGroup_lo_2217 = {dataGroup_lo_hi_2217, dataGroup_lo_lo_2217};
  wire [2047:0] dataGroup_hi_2217 = {dataGroup_hi_hi_2217, dataGroup_hi_lo_2217};
  wire [7:0]    dataGroup_41_34 = dataGroup_hi_2217[631:624];
  wire [2047:0] dataGroup_lo_2218 = {dataGroup_lo_hi_2218, dataGroup_lo_lo_2218};
  wire [2047:0] dataGroup_hi_2218 = {dataGroup_hi_hi_2218, dataGroup_hi_lo_2218};
  wire [7:0]    dataGroup_42_34 = dataGroup_hi_2218[695:688];
  wire [2047:0] dataGroup_lo_2219 = {dataGroup_lo_hi_2219, dataGroup_lo_lo_2219};
  wire [2047:0] dataGroup_hi_2219 = {dataGroup_hi_hi_2219, dataGroup_hi_lo_2219};
  wire [7:0]    dataGroup_43_34 = dataGroup_hi_2219[759:752];
  wire [2047:0] dataGroup_lo_2220 = {dataGroup_lo_hi_2220, dataGroup_lo_lo_2220};
  wire [2047:0] dataGroup_hi_2220 = {dataGroup_hi_hi_2220, dataGroup_hi_lo_2220};
  wire [7:0]    dataGroup_44_34 = dataGroup_hi_2220[823:816];
  wire [2047:0] dataGroup_lo_2221 = {dataGroup_lo_hi_2221, dataGroup_lo_lo_2221};
  wire [2047:0] dataGroup_hi_2221 = {dataGroup_hi_hi_2221, dataGroup_hi_lo_2221};
  wire [7:0]    dataGroup_45_34 = dataGroup_hi_2221[887:880];
  wire [2047:0] dataGroup_lo_2222 = {dataGroup_lo_hi_2222, dataGroup_lo_lo_2222};
  wire [2047:0] dataGroup_hi_2222 = {dataGroup_hi_hi_2222, dataGroup_hi_lo_2222};
  wire [7:0]    dataGroup_46_34 = dataGroup_hi_2222[951:944];
  wire [2047:0] dataGroup_lo_2223 = {dataGroup_lo_hi_2223, dataGroup_lo_lo_2223};
  wire [2047:0] dataGroup_hi_2223 = {dataGroup_hi_hi_2223, dataGroup_hi_lo_2223};
  wire [7:0]    dataGroup_47_34 = dataGroup_hi_2223[1015:1008];
  wire [2047:0] dataGroup_lo_2224 = {dataGroup_lo_hi_2224, dataGroup_lo_lo_2224};
  wire [2047:0] dataGroup_hi_2224 = {dataGroup_hi_hi_2224, dataGroup_hi_lo_2224};
  wire [7:0]    dataGroup_48_34 = dataGroup_hi_2224[1079:1072];
  wire [2047:0] dataGroup_lo_2225 = {dataGroup_lo_hi_2225, dataGroup_lo_lo_2225};
  wire [2047:0] dataGroup_hi_2225 = {dataGroup_hi_hi_2225, dataGroup_hi_lo_2225};
  wire [7:0]    dataGroup_49_34 = dataGroup_hi_2225[1143:1136];
  wire [2047:0] dataGroup_lo_2226 = {dataGroup_lo_hi_2226, dataGroup_lo_lo_2226};
  wire [2047:0] dataGroup_hi_2226 = {dataGroup_hi_hi_2226, dataGroup_hi_lo_2226};
  wire [7:0]    dataGroup_50_34 = dataGroup_hi_2226[1207:1200];
  wire [2047:0] dataGroup_lo_2227 = {dataGroup_lo_hi_2227, dataGroup_lo_lo_2227};
  wire [2047:0] dataGroup_hi_2227 = {dataGroup_hi_hi_2227, dataGroup_hi_lo_2227};
  wire [7:0]    dataGroup_51_34 = dataGroup_hi_2227[1271:1264];
  wire [2047:0] dataGroup_lo_2228 = {dataGroup_lo_hi_2228, dataGroup_lo_lo_2228};
  wire [2047:0] dataGroup_hi_2228 = {dataGroup_hi_hi_2228, dataGroup_hi_lo_2228};
  wire [7:0]    dataGroup_52_34 = dataGroup_hi_2228[1335:1328];
  wire [2047:0] dataGroup_lo_2229 = {dataGroup_lo_hi_2229, dataGroup_lo_lo_2229};
  wire [2047:0] dataGroup_hi_2229 = {dataGroup_hi_hi_2229, dataGroup_hi_lo_2229};
  wire [7:0]    dataGroup_53_34 = dataGroup_hi_2229[1399:1392];
  wire [2047:0] dataGroup_lo_2230 = {dataGroup_lo_hi_2230, dataGroup_lo_lo_2230};
  wire [2047:0] dataGroup_hi_2230 = {dataGroup_hi_hi_2230, dataGroup_hi_lo_2230};
  wire [7:0]    dataGroup_54_34 = dataGroup_hi_2230[1463:1456];
  wire [2047:0] dataGroup_lo_2231 = {dataGroup_lo_hi_2231, dataGroup_lo_lo_2231};
  wire [2047:0] dataGroup_hi_2231 = {dataGroup_hi_hi_2231, dataGroup_hi_lo_2231};
  wire [7:0]    dataGroup_55_34 = dataGroup_hi_2231[1527:1520];
  wire [2047:0] dataGroup_lo_2232 = {dataGroup_lo_hi_2232, dataGroup_lo_lo_2232};
  wire [2047:0] dataGroup_hi_2232 = {dataGroup_hi_hi_2232, dataGroup_hi_lo_2232};
  wire [7:0]    dataGroup_56_34 = dataGroup_hi_2232[1591:1584];
  wire [2047:0] dataGroup_lo_2233 = {dataGroup_lo_hi_2233, dataGroup_lo_lo_2233};
  wire [2047:0] dataGroup_hi_2233 = {dataGroup_hi_hi_2233, dataGroup_hi_lo_2233};
  wire [7:0]    dataGroup_57_34 = dataGroup_hi_2233[1655:1648];
  wire [2047:0] dataGroup_lo_2234 = {dataGroup_lo_hi_2234, dataGroup_lo_lo_2234};
  wire [2047:0] dataGroup_hi_2234 = {dataGroup_hi_hi_2234, dataGroup_hi_lo_2234};
  wire [7:0]    dataGroup_58_34 = dataGroup_hi_2234[1719:1712];
  wire [2047:0] dataGroup_lo_2235 = {dataGroup_lo_hi_2235, dataGroup_lo_lo_2235};
  wire [2047:0] dataGroup_hi_2235 = {dataGroup_hi_hi_2235, dataGroup_hi_lo_2235};
  wire [7:0]    dataGroup_59_34 = dataGroup_hi_2235[1783:1776];
  wire [2047:0] dataGroup_lo_2236 = {dataGroup_lo_hi_2236, dataGroup_lo_lo_2236};
  wire [2047:0] dataGroup_hi_2236 = {dataGroup_hi_hi_2236, dataGroup_hi_lo_2236};
  wire [7:0]    dataGroup_60_34 = dataGroup_hi_2236[1847:1840];
  wire [2047:0] dataGroup_lo_2237 = {dataGroup_lo_hi_2237, dataGroup_lo_lo_2237};
  wire [2047:0] dataGroup_hi_2237 = {dataGroup_hi_hi_2237, dataGroup_hi_lo_2237};
  wire [7:0]    dataGroup_61_34 = dataGroup_hi_2237[1911:1904];
  wire [2047:0] dataGroup_lo_2238 = {dataGroup_lo_hi_2238, dataGroup_lo_lo_2238};
  wire [2047:0] dataGroup_hi_2238 = {dataGroup_hi_hi_2238, dataGroup_hi_lo_2238};
  wire [7:0]    dataGroup_62_34 = dataGroup_hi_2238[1975:1968];
  wire [2047:0] dataGroup_lo_2239 = {dataGroup_lo_hi_2239, dataGroup_lo_lo_2239};
  wire [2047:0] dataGroup_hi_2239 = {dataGroup_hi_hi_2239, dataGroup_hi_lo_2239};
  wire [7:0]    dataGroup_63_34 = dataGroup_hi_2239[2039:2032];
  wire [15:0]   res_lo_lo_lo_lo_lo_34 = {dataGroup_1_34, dataGroup_0_34};
  wire [15:0]   res_lo_lo_lo_lo_hi_34 = {dataGroup_3_34, dataGroup_2_34};
  wire [31:0]   res_lo_lo_lo_lo_34 = {res_lo_lo_lo_lo_hi_34, res_lo_lo_lo_lo_lo_34};
  wire [15:0]   res_lo_lo_lo_hi_lo_34 = {dataGroup_5_34, dataGroup_4_34};
  wire [15:0]   res_lo_lo_lo_hi_hi_34 = {dataGroup_7_34, dataGroup_6_34};
  wire [31:0]   res_lo_lo_lo_hi_34 = {res_lo_lo_lo_hi_hi_34, res_lo_lo_lo_hi_lo_34};
  wire [63:0]   res_lo_lo_lo_34 = {res_lo_lo_lo_hi_34, res_lo_lo_lo_lo_34};
  wire [15:0]   res_lo_lo_hi_lo_lo_34 = {dataGroup_9_34, dataGroup_8_34};
  wire [15:0]   res_lo_lo_hi_lo_hi_34 = {dataGroup_11_34, dataGroup_10_34};
  wire [31:0]   res_lo_lo_hi_lo_34 = {res_lo_lo_hi_lo_hi_34, res_lo_lo_hi_lo_lo_34};
  wire [15:0]   res_lo_lo_hi_hi_lo_34 = {dataGroup_13_34, dataGroup_12_34};
  wire [15:0]   res_lo_lo_hi_hi_hi_34 = {dataGroup_15_34, dataGroup_14_34};
  wire [31:0]   res_lo_lo_hi_hi_34 = {res_lo_lo_hi_hi_hi_34, res_lo_lo_hi_hi_lo_34};
  wire [63:0]   res_lo_lo_hi_34 = {res_lo_lo_hi_hi_34, res_lo_lo_hi_lo_34};
  wire [127:0]  res_lo_lo_34 = {res_lo_lo_hi_34, res_lo_lo_lo_34};
  wire [15:0]   res_lo_hi_lo_lo_lo_34 = {dataGroup_17_34, dataGroup_16_34};
  wire [15:0]   res_lo_hi_lo_lo_hi_34 = {dataGroup_19_34, dataGroup_18_34};
  wire [31:0]   res_lo_hi_lo_lo_34 = {res_lo_hi_lo_lo_hi_34, res_lo_hi_lo_lo_lo_34};
  wire [15:0]   res_lo_hi_lo_hi_lo_34 = {dataGroup_21_34, dataGroup_20_34};
  wire [15:0]   res_lo_hi_lo_hi_hi_34 = {dataGroup_23_34, dataGroup_22_34};
  wire [31:0]   res_lo_hi_lo_hi_34 = {res_lo_hi_lo_hi_hi_34, res_lo_hi_lo_hi_lo_34};
  wire [63:0]   res_lo_hi_lo_34 = {res_lo_hi_lo_hi_34, res_lo_hi_lo_lo_34};
  wire [15:0]   res_lo_hi_hi_lo_lo_34 = {dataGroup_25_34, dataGroup_24_34};
  wire [15:0]   res_lo_hi_hi_lo_hi_34 = {dataGroup_27_34, dataGroup_26_34};
  wire [31:0]   res_lo_hi_hi_lo_34 = {res_lo_hi_hi_lo_hi_34, res_lo_hi_hi_lo_lo_34};
  wire [15:0]   res_lo_hi_hi_hi_lo_34 = {dataGroup_29_34, dataGroup_28_34};
  wire [15:0]   res_lo_hi_hi_hi_hi_34 = {dataGroup_31_34, dataGroup_30_34};
  wire [31:0]   res_lo_hi_hi_hi_34 = {res_lo_hi_hi_hi_hi_34, res_lo_hi_hi_hi_lo_34};
  wire [63:0]   res_lo_hi_hi_34 = {res_lo_hi_hi_hi_34, res_lo_hi_hi_lo_34};
  wire [127:0]  res_lo_hi_34 = {res_lo_hi_hi_34, res_lo_hi_lo_34};
  wire [255:0]  res_lo_34 = {res_lo_hi_34, res_lo_lo_34};
  wire [15:0]   res_hi_lo_lo_lo_lo_34 = {dataGroup_33_34, dataGroup_32_34};
  wire [15:0]   res_hi_lo_lo_lo_hi_34 = {dataGroup_35_34, dataGroup_34_34};
  wire [31:0]   res_hi_lo_lo_lo_34 = {res_hi_lo_lo_lo_hi_34, res_hi_lo_lo_lo_lo_34};
  wire [15:0]   res_hi_lo_lo_hi_lo_34 = {dataGroup_37_34, dataGroup_36_34};
  wire [15:0]   res_hi_lo_lo_hi_hi_34 = {dataGroup_39_34, dataGroup_38_34};
  wire [31:0]   res_hi_lo_lo_hi_34 = {res_hi_lo_lo_hi_hi_34, res_hi_lo_lo_hi_lo_34};
  wire [63:0]   res_hi_lo_lo_34 = {res_hi_lo_lo_hi_34, res_hi_lo_lo_lo_34};
  wire [15:0]   res_hi_lo_hi_lo_lo_34 = {dataGroup_41_34, dataGroup_40_34};
  wire [15:0]   res_hi_lo_hi_lo_hi_34 = {dataGroup_43_34, dataGroup_42_34};
  wire [31:0]   res_hi_lo_hi_lo_34 = {res_hi_lo_hi_lo_hi_34, res_hi_lo_hi_lo_lo_34};
  wire [15:0]   res_hi_lo_hi_hi_lo_34 = {dataGroup_45_34, dataGroup_44_34};
  wire [15:0]   res_hi_lo_hi_hi_hi_34 = {dataGroup_47_34, dataGroup_46_34};
  wire [31:0]   res_hi_lo_hi_hi_34 = {res_hi_lo_hi_hi_hi_34, res_hi_lo_hi_hi_lo_34};
  wire [63:0]   res_hi_lo_hi_34 = {res_hi_lo_hi_hi_34, res_hi_lo_hi_lo_34};
  wire [127:0]  res_hi_lo_34 = {res_hi_lo_hi_34, res_hi_lo_lo_34};
  wire [15:0]   res_hi_hi_lo_lo_lo_34 = {dataGroup_49_34, dataGroup_48_34};
  wire [15:0]   res_hi_hi_lo_lo_hi_34 = {dataGroup_51_34, dataGroup_50_34};
  wire [31:0]   res_hi_hi_lo_lo_34 = {res_hi_hi_lo_lo_hi_34, res_hi_hi_lo_lo_lo_34};
  wire [15:0]   res_hi_hi_lo_hi_lo_34 = {dataGroup_53_34, dataGroup_52_34};
  wire [15:0]   res_hi_hi_lo_hi_hi_34 = {dataGroup_55_34, dataGroup_54_34};
  wire [31:0]   res_hi_hi_lo_hi_34 = {res_hi_hi_lo_hi_hi_34, res_hi_hi_lo_hi_lo_34};
  wire [63:0]   res_hi_hi_lo_34 = {res_hi_hi_lo_hi_34, res_hi_hi_lo_lo_34};
  wire [15:0]   res_hi_hi_hi_lo_lo_34 = {dataGroup_57_34, dataGroup_56_34};
  wire [15:0]   res_hi_hi_hi_lo_hi_34 = {dataGroup_59_34, dataGroup_58_34};
  wire [31:0]   res_hi_hi_hi_lo_34 = {res_hi_hi_hi_lo_hi_34, res_hi_hi_hi_lo_lo_34};
  wire [15:0]   res_hi_hi_hi_hi_lo_34 = {dataGroup_61_34, dataGroup_60_34};
  wire [15:0]   res_hi_hi_hi_hi_hi_34 = {dataGroup_63_34, dataGroup_62_34};
  wire [31:0]   res_hi_hi_hi_hi_34 = {res_hi_hi_hi_hi_hi_34, res_hi_hi_hi_hi_lo_34};
  wire [63:0]   res_hi_hi_hi_34 = {res_hi_hi_hi_hi_34, res_hi_hi_hi_lo_34};
  wire [127:0]  res_hi_hi_34 = {res_hi_hi_hi_34, res_hi_hi_lo_34};
  wire [255:0]  res_hi_34 = {res_hi_hi_34, res_hi_lo_34};
  wire [511:0]  res_62 = {res_hi_34, res_lo_34};
  wire [2047:0] dataGroup_lo_2240 = {dataGroup_lo_hi_2240, dataGroup_lo_lo_2240};
  wire [2047:0] dataGroup_hi_2240 = {dataGroup_hi_hi_2240, dataGroup_hi_lo_2240};
  wire [7:0]    dataGroup_0_35 = dataGroup_lo_2240[63:56];
  wire [2047:0] dataGroup_lo_2241 = {dataGroup_lo_hi_2241, dataGroup_lo_lo_2241};
  wire [2047:0] dataGroup_hi_2241 = {dataGroup_hi_hi_2241, dataGroup_hi_lo_2241};
  wire [7:0]    dataGroup_1_35 = dataGroup_lo_2241[127:120];
  wire [2047:0] dataGroup_lo_2242 = {dataGroup_lo_hi_2242, dataGroup_lo_lo_2242};
  wire [2047:0] dataGroup_hi_2242 = {dataGroup_hi_hi_2242, dataGroup_hi_lo_2242};
  wire [7:0]    dataGroup_2_35 = dataGroup_lo_2242[191:184];
  wire [2047:0] dataGroup_lo_2243 = {dataGroup_lo_hi_2243, dataGroup_lo_lo_2243};
  wire [2047:0] dataGroup_hi_2243 = {dataGroup_hi_hi_2243, dataGroup_hi_lo_2243};
  wire [7:0]    dataGroup_3_35 = dataGroup_lo_2243[255:248];
  wire [2047:0] dataGroup_lo_2244 = {dataGroup_lo_hi_2244, dataGroup_lo_lo_2244};
  wire [2047:0] dataGroup_hi_2244 = {dataGroup_hi_hi_2244, dataGroup_hi_lo_2244};
  wire [7:0]    dataGroup_4_35 = dataGroup_lo_2244[319:312];
  wire [2047:0] dataGroup_lo_2245 = {dataGroup_lo_hi_2245, dataGroup_lo_lo_2245};
  wire [2047:0] dataGroup_hi_2245 = {dataGroup_hi_hi_2245, dataGroup_hi_lo_2245};
  wire [7:0]    dataGroup_5_35 = dataGroup_lo_2245[383:376];
  wire [2047:0] dataGroup_lo_2246 = {dataGroup_lo_hi_2246, dataGroup_lo_lo_2246};
  wire [2047:0] dataGroup_hi_2246 = {dataGroup_hi_hi_2246, dataGroup_hi_lo_2246};
  wire [7:0]    dataGroup_6_35 = dataGroup_lo_2246[447:440];
  wire [2047:0] dataGroup_lo_2247 = {dataGroup_lo_hi_2247, dataGroup_lo_lo_2247};
  wire [2047:0] dataGroup_hi_2247 = {dataGroup_hi_hi_2247, dataGroup_hi_lo_2247};
  wire [7:0]    dataGroup_7_35 = dataGroup_lo_2247[511:504];
  wire [2047:0] dataGroup_lo_2248 = {dataGroup_lo_hi_2248, dataGroup_lo_lo_2248};
  wire [2047:0] dataGroup_hi_2248 = {dataGroup_hi_hi_2248, dataGroup_hi_lo_2248};
  wire [7:0]    dataGroup_8_35 = dataGroup_lo_2248[575:568];
  wire [2047:0] dataGroup_lo_2249 = {dataGroup_lo_hi_2249, dataGroup_lo_lo_2249};
  wire [2047:0] dataGroup_hi_2249 = {dataGroup_hi_hi_2249, dataGroup_hi_lo_2249};
  wire [7:0]    dataGroup_9_35 = dataGroup_lo_2249[639:632];
  wire [2047:0] dataGroup_lo_2250 = {dataGroup_lo_hi_2250, dataGroup_lo_lo_2250};
  wire [2047:0] dataGroup_hi_2250 = {dataGroup_hi_hi_2250, dataGroup_hi_lo_2250};
  wire [7:0]    dataGroup_10_35 = dataGroup_lo_2250[703:696];
  wire [2047:0] dataGroup_lo_2251 = {dataGroup_lo_hi_2251, dataGroup_lo_lo_2251};
  wire [2047:0] dataGroup_hi_2251 = {dataGroup_hi_hi_2251, dataGroup_hi_lo_2251};
  wire [7:0]    dataGroup_11_35 = dataGroup_lo_2251[767:760];
  wire [2047:0] dataGroup_lo_2252 = {dataGroup_lo_hi_2252, dataGroup_lo_lo_2252};
  wire [2047:0] dataGroup_hi_2252 = {dataGroup_hi_hi_2252, dataGroup_hi_lo_2252};
  wire [7:0]    dataGroup_12_35 = dataGroup_lo_2252[831:824];
  wire [2047:0] dataGroup_lo_2253 = {dataGroup_lo_hi_2253, dataGroup_lo_lo_2253};
  wire [2047:0] dataGroup_hi_2253 = {dataGroup_hi_hi_2253, dataGroup_hi_lo_2253};
  wire [7:0]    dataGroup_13_35 = dataGroup_lo_2253[895:888];
  wire [2047:0] dataGroup_lo_2254 = {dataGroup_lo_hi_2254, dataGroup_lo_lo_2254};
  wire [2047:0] dataGroup_hi_2254 = {dataGroup_hi_hi_2254, dataGroup_hi_lo_2254};
  wire [7:0]    dataGroup_14_35 = dataGroup_lo_2254[959:952];
  wire [2047:0] dataGroup_lo_2255 = {dataGroup_lo_hi_2255, dataGroup_lo_lo_2255};
  wire [2047:0] dataGroup_hi_2255 = {dataGroup_hi_hi_2255, dataGroup_hi_lo_2255};
  wire [7:0]    dataGroup_15_35 = dataGroup_lo_2255[1023:1016];
  wire [2047:0] dataGroup_lo_2256 = {dataGroup_lo_hi_2256, dataGroup_lo_lo_2256};
  wire [2047:0] dataGroup_hi_2256 = {dataGroup_hi_hi_2256, dataGroup_hi_lo_2256};
  wire [7:0]    dataGroup_16_35 = dataGroup_lo_2256[1087:1080];
  wire [2047:0] dataGroup_lo_2257 = {dataGroup_lo_hi_2257, dataGroup_lo_lo_2257};
  wire [2047:0] dataGroup_hi_2257 = {dataGroup_hi_hi_2257, dataGroup_hi_lo_2257};
  wire [7:0]    dataGroup_17_35 = dataGroup_lo_2257[1151:1144];
  wire [2047:0] dataGroup_lo_2258 = {dataGroup_lo_hi_2258, dataGroup_lo_lo_2258};
  wire [2047:0] dataGroup_hi_2258 = {dataGroup_hi_hi_2258, dataGroup_hi_lo_2258};
  wire [7:0]    dataGroup_18_35 = dataGroup_lo_2258[1215:1208];
  wire [2047:0] dataGroup_lo_2259 = {dataGroup_lo_hi_2259, dataGroup_lo_lo_2259};
  wire [2047:0] dataGroup_hi_2259 = {dataGroup_hi_hi_2259, dataGroup_hi_lo_2259};
  wire [7:0]    dataGroup_19_35 = dataGroup_lo_2259[1279:1272];
  wire [2047:0] dataGroup_lo_2260 = {dataGroup_lo_hi_2260, dataGroup_lo_lo_2260};
  wire [2047:0] dataGroup_hi_2260 = {dataGroup_hi_hi_2260, dataGroup_hi_lo_2260};
  wire [7:0]    dataGroup_20_35 = dataGroup_lo_2260[1343:1336];
  wire [2047:0] dataGroup_lo_2261 = {dataGroup_lo_hi_2261, dataGroup_lo_lo_2261};
  wire [2047:0] dataGroup_hi_2261 = {dataGroup_hi_hi_2261, dataGroup_hi_lo_2261};
  wire [7:0]    dataGroup_21_35 = dataGroup_lo_2261[1407:1400];
  wire [2047:0] dataGroup_lo_2262 = {dataGroup_lo_hi_2262, dataGroup_lo_lo_2262};
  wire [2047:0] dataGroup_hi_2262 = {dataGroup_hi_hi_2262, dataGroup_hi_lo_2262};
  wire [7:0]    dataGroup_22_35 = dataGroup_lo_2262[1471:1464];
  wire [2047:0] dataGroup_lo_2263 = {dataGroup_lo_hi_2263, dataGroup_lo_lo_2263};
  wire [2047:0] dataGroup_hi_2263 = {dataGroup_hi_hi_2263, dataGroup_hi_lo_2263};
  wire [7:0]    dataGroup_23_35 = dataGroup_lo_2263[1535:1528];
  wire [2047:0] dataGroup_lo_2264 = {dataGroup_lo_hi_2264, dataGroup_lo_lo_2264};
  wire [2047:0] dataGroup_hi_2264 = {dataGroup_hi_hi_2264, dataGroup_hi_lo_2264};
  wire [7:0]    dataGroup_24_35 = dataGroup_lo_2264[1599:1592];
  wire [2047:0] dataGroup_lo_2265 = {dataGroup_lo_hi_2265, dataGroup_lo_lo_2265};
  wire [2047:0] dataGroup_hi_2265 = {dataGroup_hi_hi_2265, dataGroup_hi_lo_2265};
  wire [7:0]    dataGroup_25_35 = dataGroup_lo_2265[1663:1656];
  wire [2047:0] dataGroup_lo_2266 = {dataGroup_lo_hi_2266, dataGroup_lo_lo_2266};
  wire [2047:0] dataGroup_hi_2266 = {dataGroup_hi_hi_2266, dataGroup_hi_lo_2266};
  wire [7:0]    dataGroup_26_35 = dataGroup_lo_2266[1727:1720];
  wire [2047:0] dataGroup_lo_2267 = {dataGroup_lo_hi_2267, dataGroup_lo_lo_2267};
  wire [2047:0] dataGroup_hi_2267 = {dataGroup_hi_hi_2267, dataGroup_hi_lo_2267};
  wire [7:0]    dataGroup_27_35 = dataGroup_lo_2267[1791:1784];
  wire [2047:0] dataGroup_lo_2268 = {dataGroup_lo_hi_2268, dataGroup_lo_lo_2268};
  wire [2047:0] dataGroup_hi_2268 = {dataGroup_hi_hi_2268, dataGroup_hi_lo_2268};
  wire [7:0]    dataGroup_28_35 = dataGroup_lo_2268[1855:1848];
  wire [2047:0] dataGroup_lo_2269 = {dataGroup_lo_hi_2269, dataGroup_lo_lo_2269};
  wire [2047:0] dataGroup_hi_2269 = {dataGroup_hi_hi_2269, dataGroup_hi_lo_2269};
  wire [7:0]    dataGroup_29_35 = dataGroup_lo_2269[1919:1912];
  wire [2047:0] dataGroup_lo_2270 = {dataGroup_lo_hi_2270, dataGroup_lo_lo_2270};
  wire [2047:0] dataGroup_hi_2270 = {dataGroup_hi_hi_2270, dataGroup_hi_lo_2270};
  wire [7:0]    dataGroup_30_35 = dataGroup_lo_2270[1983:1976];
  wire [2047:0] dataGroup_lo_2271 = {dataGroup_lo_hi_2271, dataGroup_lo_lo_2271};
  wire [2047:0] dataGroup_hi_2271 = {dataGroup_hi_hi_2271, dataGroup_hi_lo_2271};
  wire [7:0]    dataGroup_31_35 = dataGroup_lo_2271[2047:2040];
  wire [2047:0] dataGroup_lo_2272 = {dataGroup_lo_hi_2272, dataGroup_lo_lo_2272};
  wire [2047:0] dataGroup_hi_2272 = {dataGroup_hi_hi_2272, dataGroup_hi_lo_2272};
  wire [7:0]    dataGroup_32_35 = dataGroup_hi_2272[63:56];
  wire [2047:0] dataGroup_lo_2273 = {dataGroup_lo_hi_2273, dataGroup_lo_lo_2273};
  wire [2047:0] dataGroup_hi_2273 = {dataGroup_hi_hi_2273, dataGroup_hi_lo_2273};
  wire [7:0]    dataGroup_33_35 = dataGroup_hi_2273[127:120];
  wire [2047:0] dataGroup_lo_2274 = {dataGroup_lo_hi_2274, dataGroup_lo_lo_2274};
  wire [2047:0] dataGroup_hi_2274 = {dataGroup_hi_hi_2274, dataGroup_hi_lo_2274};
  wire [7:0]    dataGroup_34_35 = dataGroup_hi_2274[191:184];
  wire [2047:0] dataGroup_lo_2275 = {dataGroup_lo_hi_2275, dataGroup_lo_lo_2275};
  wire [2047:0] dataGroup_hi_2275 = {dataGroup_hi_hi_2275, dataGroup_hi_lo_2275};
  wire [7:0]    dataGroup_35_35 = dataGroup_hi_2275[255:248];
  wire [2047:0] dataGroup_lo_2276 = {dataGroup_lo_hi_2276, dataGroup_lo_lo_2276};
  wire [2047:0] dataGroup_hi_2276 = {dataGroup_hi_hi_2276, dataGroup_hi_lo_2276};
  wire [7:0]    dataGroup_36_35 = dataGroup_hi_2276[319:312];
  wire [2047:0] dataGroup_lo_2277 = {dataGroup_lo_hi_2277, dataGroup_lo_lo_2277};
  wire [2047:0] dataGroup_hi_2277 = {dataGroup_hi_hi_2277, dataGroup_hi_lo_2277};
  wire [7:0]    dataGroup_37_35 = dataGroup_hi_2277[383:376];
  wire [2047:0] dataGroup_lo_2278 = {dataGroup_lo_hi_2278, dataGroup_lo_lo_2278};
  wire [2047:0] dataGroup_hi_2278 = {dataGroup_hi_hi_2278, dataGroup_hi_lo_2278};
  wire [7:0]    dataGroup_38_35 = dataGroup_hi_2278[447:440];
  wire [2047:0] dataGroup_lo_2279 = {dataGroup_lo_hi_2279, dataGroup_lo_lo_2279};
  wire [2047:0] dataGroup_hi_2279 = {dataGroup_hi_hi_2279, dataGroup_hi_lo_2279};
  wire [7:0]    dataGroup_39_35 = dataGroup_hi_2279[511:504];
  wire [2047:0] dataGroup_lo_2280 = {dataGroup_lo_hi_2280, dataGroup_lo_lo_2280};
  wire [2047:0] dataGroup_hi_2280 = {dataGroup_hi_hi_2280, dataGroup_hi_lo_2280};
  wire [7:0]    dataGroup_40_35 = dataGroup_hi_2280[575:568];
  wire [2047:0] dataGroup_lo_2281 = {dataGroup_lo_hi_2281, dataGroup_lo_lo_2281};
  wire [2047:0] dataGroup_hi_2281 = {dataGroup_hi_hi_2281, dataGroup_hi_lo_2281};
  wire [7:0]    dataGroup_41_35 = dataGroup_hi_2281[639:632];
  wire [2047:0] dataGroup_lo_2282 = {dataGroup_lo_hi_2282, dataGroup_lo_lo_2282};
  wire [2047:0] dataGroup_hi_2282 = {dataGroup_hi_hi_2282, dataGroup_hi_lo_2282};
  wire [7:0]    dataGroup_42_35 = dataGroup_hi_2282[703:696];
  wire [2047:0] dataGroup_lo_2283 = {dataGroup_lo_hi_2283, dataGroup_lo_lo_2283};
  wire [2047:0] dataGroup_hi_2283 = {dataGroup_hi_hi_2283, dataGroup_hi_lo_2283};
  wire [7:0]    dataGroup_43_35 = dataGroup_hi_2283[767:760];
  wire [2047:0] dataGroup_lo_2284 = {dataGroup_lo_hi_2284, dataGroup_lo_lo_2284};
  wire [2047:0] dataGroup_hi_2284 = {dataGroup_hi_hi_2284, dataGroup_hi_lo_2284};
  wire [7:0]    dataGroup_44_35 = dataGroup_hi_2284[831:824];
  wire [2047:0] dataGroup_lo_2285 = {dataGroup_lo_hi_2285, dataGroup_lo_lo_2285};
  wire [2047:0] dataGroup_hi_2285 = {dataGroup_hi_hi_2285, dataGroup_hi_lo_2285};
  wire [7:0]    dataGroup_45_35 = dataGroup_hi_2285[895:888];
  wire [2047:0] dataGroup_lo_2286 = {dataGroup_lo_hi_2286, dataGroup_lo_lo_2286};
  wire [2047:0] dataGroup_hi_2286 = {dataGroup_hi_hi_2286, dataGroup_hi_lo_2286};
  wire [7:0]    dataGroup_46_35 = dataGroup_hi_2286[959:952];
  wire [2047:0] dataGroup_lo_2287 = {dataGroup_lo_hi_2287, dataGroup_lo_lo_2287};
  wire [2047:0] dataGroup_hi_2287 = {dataGroup_hi_hi_2287, dataGroup_hi_lo_2287};
  wire [7:0]    dataGroup_47_35 = dataGroup_hi_2287[1023:1016];
  wire [2047:0] dataGroup_lo_2288 = {dataGroup_lo_hi_2288, dataGroup_lo_lo_2288};
  wire [2047:0] dataGroup_hi_2288 = {dataGroup_hi_hi_2288, dataGroup_hi_lo_2288};
  wire [7:0]    dataGroup_48_35 = dataGroup_hi_2288[1087:1080];
  wire [2047:0] dataGroup_lo_2289 = {dataGroup_lo_hi_2289, dataGroup_lo_lo_2289};
  wire [2047:0] dataGroup_hi_2289 = {dataGroup_hi_hi_2289, dataGroup_hi_lo_2289};
  wire [7:0]    dataGroup_49_35 = dataGroup_hi_2289[1151:1144];
  wire [2047:0] dataGroup_lo_2290 = {dataGroup_lo_hi_2290, dataGroup_lo_lo_2290};
  wire [2047:0] dataGroup_hi_2290 = {dataGroup_hi_hi_2290, dataGroup_hi_lo_2290};
  wire [7:0]    dataGroup_50_35 = dataGroup_hi_2290[1215:1208];
  wire [2047:0] dataGroup_lo_2291 = {dataGroup_lo_hi_2291, dataGroup_lo_lo_2291};
  wire [2047:0] dataGroup_hi_2291 = {dataGroup_hi_hi_2291, dataGroup_hi_lo_2291};
  wire [7:0]    dataGroup_51_35 = dataGroup_hi_2291[1279:1272];
  wire [2047:0] dataGroup_lo_2292 = {dataGroup_lo_hi_2292, dataGroup_lo_lo_2292};
  wire [2047:0] dataGroup_hi_2292 = {dataGroup_hi_hi_2292, dataGroup_hi_lo_2292};
  wire [7:0]    dataGroup_52_35 = dataGroup_hi_2292[1343:1336];
  wire [2047:0] dataGroup_lo_2293 = {dataGroup_lo_hi_2293, dataGroup_lo_lo_2293};
  wire [2047:0] dataGroup_hi_2293 = {dataGroup_hi_hi_2293, dataGroup_hi_lo_2293};
  wire [7:0]    dataGroup_53_35 = dataGroup_hi_2293[1407:1400];
  wire [2047:0] dataGroup_lo_2294 = {dataGroup_lo_hi_2294, dataGroup_lo_lo_2294};
  wire [2047:0] dataGroup_hi_2294 = {dataGroup_hi_hi_2294, dataGroup_hi_lo_2294};
  wire [7:0]    dataGroup_54_35 = dataGroup_hi_2294[1471:1464];
  wire [2047:0] dataGroup_lo_2295 = {dataGroup_lo_hi_2295, dataGroup_lo_lo_2295};
  wire [2047:0] dataGroup_hi_2295 = {dataGroup_hi_hi_2295, dataGroup_hi_lo_2295};
  wire [7:0]    dataGroup_55_35 = dataGroup_hi_2295[1535:1528];
  wire [2047:0] dataGroup_lo_2296 = {dataGroup_lo_hi_2296, dataGroup_lo_lo_2296};
  wire [2047:0] dataGroup_hi_2296 = {dataGroup_hi_hi_2296, dataGroup_hi_lo_2296};
  wire [7:0]    dataGroup_56_35 = dataGroup_hi_2296[1599:1592];
  wire [2047:0] dataGroup_lo_2297 = {dataGroup_lo_hi_2297, dataGroup_lo_lo_2297};
  wire [2047:0] dataGroup_hi_2297 = {dataGroup_hi_hi_2297, dataGroup_hi_lo_2297};
  wire [7:0]    dataGroup_57_35 = dataGroup_hi_2297[1663:1656];
  wire [2047:0] dataGroup_lo_2298 = {dataGroup_lo_hi_2298, dataGroup_lo_lo_2298};
  wire [2047:0] dataGroup_hi_2298 = {dataGroup_hi_hi_2298, dataGroup_hi_lo_2298};
  wire [7:0]    dataGroup_58_35 = dataGroup_hi_2298[1727:1720];
  wire [2047:0] dataGroup_lo_2299 = {dataGroup_lo_hi_2299, dataGroup_lo_lo_2299};
  wire [2047:0] dataGroup_hi_2299 = {dataGroup_hi_hi_2299, dataGroup_hi_lo_2299};
  wire [7:0]    dataGroup_59_35 = dataGroup_hi_2299[1791:1784];
  wire [2047:0] dataGroup_lo_2300 = {dataGroup_lo_hi_2300, dataGroup_lo_lo_2300};
  wire [2047:0] dataGroup_hi_2300 = {dataGroup_hi_hi_2300, dataGroup_hi_lo_2300};
  wire [7:0]    dataGroup_60_35 = dataGroup_hi_2300[1855:1848];
  wire [2047:0] dataGroup_lo_2301 = {dataGroup_lo_hi_2301, dataGroup_lo_lo_2301};
  wire [2047:0] dataGroup_hi_2301 = {dataGroup_hi_hi_2301, dataGroup_hi_lo_2301};
  wire [7:0]    dataGroup_61_35 = dataGroup_hi_2301[1919:1912];
  wire [2047:0] dataGroup_lo_2302 = {dataGroup_lo_hi_2302, dataGroup_lo_lo_2302};
  wire [2047:0] dataGroup_hi_2302 = {dataGroup_hi_hi_2302, dataGroup_hi_lo_2302};
  wire [7:0]    dataGroup_62_35 = dataGroup_hi_2302[1983:1976];
  wire [2047:0] dataGroup_lo_2303 = {dataGroup_lo_hi_2303, dataGroup_lo_lo_2303};
  wire [2047:0] dataGroup_hi_2303 = {dataGroup_hi_hi_2303, dataGroup_hi_lo_2303};
  wire [7:0]    dataGroup_63_35 = dataGroup_hi_2303[2047:2040];
  wire [15:0]   res_lo_lo_lo_lo_lo_35 = {dataGroup_1_35, dataGroup_0_35};
  wire [15:0]   res_lo_lo_lo_lo_hi_35 = {dataGroup_3_35, dataGroup_2_35};
  wire [31:0]   res_lo_lo_lo_lo_35 = {res_lo_lo_lo_lo_hi_35, res_lo_lo_lo_lo_lo_35};
  wire [15:0]   res_lo_lo_lo_hi_lo_35 = {dataGroup_5_35, dataGroup_4_35};
  wire [15:0]   res_lo_lo_lo_hi_hi_35 = {dataGroup_7_35, dataGroup_6_35};
  wire [31:0]   res_lo_lo_lo_hi_35 = {res_lo_lo_lo_hi_hi_35, res_lo_lo_lo_hi_lo_35};
  wire [63:0]   res_lo_lo_lo_35 = {res_lo_lo_lo_hi_35, res_lo_lo_lo_lo_35};
  wire [15:0]   res_lo_lo_hi_lo_lo_35 = {dataGroup_9_35, dataGroup_8_35};
  wire [15:0]   res_lo_lo_hi_lo_hi_35 = {dataGroup_11_35, dataGroup_10_35};
  wire [31:0]   res_lo_lo_hi_lo_35 = {res_lo_lo_hi_lo_hi_35, res_lo_lo_hi_lo_lo_35};
  wire [15:0]   res_lo_lo_hi_hi_lo_35 = {dataGroup_13_35, dataGroup_12_35};
  wire [15:0]   res_lo_lo_hi_hi_hi_35 = {dataGroup_15_35, dataGroup_14_35};
  wire [31:0]   res_lo_lo_hi_hi_35 = {res_lo_lo_hi_hi_hi_35, res_lo_lo_hi_hi_lo_35};
  wire [63:0]   res_lo_lo_hi_35 = {res_lo_lo_hi_hi_35, res_lo_lo_hi_lo_35};
  wire [127:0]  res_lo_lo_35 = {res_lo_lo_hi_35, res_lo_lo_lo_35};
  wire [15:0]   res_lo_hi_lo_lo_lo_35 = {dataGroup_17_35, dataGroup_16_35};
  wire [15:0]   res_lo_hi_lo_lo_hi_35 = {dataGroup_19_35, dataGroup_18_35};
  wire [31:0]   res_lo_hi_lo_lo_35 = {res_lo_hi_lo_lo_hi_35, res_lo_hi_lo_lo_lo_35};
  wire [15:0]   res_lo_hi_lo_hi_lo_35 = {dataGroup_21_35, dataGroup_20_35};
  wire [15:0]   res_lo_hi_lo_hi_hi_35 = {dataGroup_23_35, dataGroup_22_35};
  wire [31:0]   res_lo_hi_lo_hi_35 = {res_lo_hi_lo_hi_hi_35, res_lo_hi_lo_hi_lo_35};
  wire [63:0]   res_lo_hi_lo_35 = {res_lo_hi_lo_hi_35, res_lo_hi_lo_lo_35};
  wire [15:0]   res_lo_hi_hi_lo_lo_35 = {dataGroup_25_35, dataGroup_24_35};
  wire [15:0]   res_lo_hi_hi_lo_hi_35 = {dataGroup_27_35, dataGroup_26_35};
  wire [31:0]   res_lo_hi_hi_lo_35 = {res_lo_hi_hi_lo_hi_35, res_lo_hi_hi_lo_lo_35};
  wire [15:0]   res_lo_hi_hi_hi_lo_35 = {dataGroup_29_35, dataGroup_28_35};
  wire [15:0]   res_lo_hi_hi_hi_hi_35 = {dataGroup_31_35, dataGroup_30_35};
  wire [31:0]   res_lo_hi_hi_hi_35 = {res_lo_hi_hi_hi_hi_35, res_lo_hi_hi_hi_lo_35};
  wire [63:0]   res_lo_hi_hi_35 = {res_lo_hi_hi_hi_35, res_lo_hi_hi_lo_35};
  wire [127:0]  res_lo_hi_35 = {res_lo_hi_hi_35, res_lo_hi_lo_35};
  wire [255:0]  res_lo_35 = {res_lo_hi_35, res_lo_lo_35};
  wire [15:0]   res_hi_lo_lo_lo_lo_35 = {dataGroup_33_35, dataGroup_32_35};
  wire [15:0]   res_hi_lo_lo_lo_hi_35 = {dataGroup_35_35, dataGroup_34_35};
  wire [31:0]   res_hi_lo_lo_lo_35 = {res_hi_lo_lo_lo_hi_35, res_hi_lo_lo_lo_lo_35};
  wire [15:0]   res_hi_lo_lo_hi_lo_35 = {dataGroup_37_35, dataGroup_36_35};
  wire [15:0]   res_hi_lo_lo_hi_hi_35 = {dataGroup_39_35, dataGroup_38_35};
  wire [31:0]   res_hi_lo_lo_hi_35 = {res_hi_lo_lo_hi_hi_35, res_hi_lo_lo_hi_lo_35};
  wire [63:0]   res_hi_lo_lo_35 = {res_hi_lo_lo_hi_35, res_hi_lo_lo_lo_35};
  wire [15:0]   res_hi_lo_hi_lo_lo_35 = {dataGroup_41_35, dataGroup_40_35};
  wire [15:0]   res_hi_lo_hi_lo_hi_35 = {dataGroup_43_35, dataGroup_42_35};
  wire [31:0]   res_hi_lo_hi_lo_35 = {res_hi_lo_hi_lo_hi_35, res_hi_lo_hi_lo_lo_35};
  wire [15:0]   res_hi_lo_hi_hi_lo_35 = {dataGroup_45_35, dataGroup_44_35};
  wire [15:0]   res_hi_lo_hi_hi_hi_35 = {dataGroup_47_35, dataGroup_46_35};
  wire [31:0]   res_hi_lo_hi_hi_35 = {res_hi_lo_hi_hi_hi_35, res_hi_lo_hi_hi_lo_35};
  wire [63:0]   res_hi_lo_hi_35 = {res_hi_lo_hi_hi_35, res_hi_lo_hi_lo_35};
  wire [127:0]  res_hi_lo_35 = {res_hi_lo_hi_35, res_hi_lo_lo_35};
  wire [15:0]   res_hi_hi_lo_lo_lo_35 = {dataGroup_49_35, dataGroup_48_35};
  wire [15:0]   res_hi_hi_lo_lo_hi_35 = {dataGroup_51_35, dataGroup_50_35};
  wire [31:0]   res_hi_hi_lo_lo_35 = {res_hi_hi_lo_lo_hi_35, res_hi_hi_lo_lo_lo_35};
  wire [15:0]   res_hi_hi_lo_hi_lo_35 = {dataGroup_53_35, dataGroup_52_35};
  wire [15:0]   res_hi_hi_lo_hi_hi_35 = {dataGroup_55_35, dataGroup_54_35};
  wire [31:0]   res_hi_hi_lo_hi_35 = {res_hi_hi_lo_hi_hi_35, res_hi_hi_lo_hi_lo_35};
  wire [63:0]   res_hi_hi_lo_35 = {res_hi_hi_lo_hi_35, res_hi_hi_lo_lo_35};
  wire [15:0]   res_hi_hi_hi_lo_lo_35 = {dataGroup_57_35, dataGroup_56_35};
  wire [15:0]   res_hi_hi_hi_lo_hi_35 = {dataGroup_59_35, dataGroup_58_35};
  wire [31:0]   res_hi_hi_hi_lo_35 = {res_hi_hi_hi_lo_hi_35, res_hi_hi_hi_lo_lo_35};
  wire [15:0]   res_hi_hi_hi_hi_lo_35 = {dataGroup_61_35, dataGroup_60_35};
  wire [15:0]   res_hi_hi_hi_hi_hi_35 = {dataGroup_63_35, dataGroup_62_35};
  wire [31:0]   res_hi_hi_hi_hi_35 = {res_hi_hi_hi_hi_hi_35, res_hi_hi_hi_hi_lo_35};
  wire [63:0]   res_hi_hi_hi_35 = {res_hi_hi_hi_hi_35, res_hi_hi_hi_lo_35};
  wire [127:0]  res_hi_hi_35 = {res_hi_hi_hi_35, res_hi_hi_lo_35};
  wire [255:0]  res_hi_35 = {res_hi_hi_35, res_hi_lo_35};
  wire [511:0]  res_63 = {res_hi_35, res_lo_35};
  wire [1023:0] lo_lo_7 = {res_57, res_56};
  wire [1023:0] lo_hi_7 = {res_59, res_58};
  wire [2047:0] lo_7 = {lo_hi_7, lo_lo_7};
  wire [1023:0] hi_lo_7 = {res_61, res_60};
  wire [1023:0] hi_hi_7 = {res_63, res_62};
  wire [2047:0] hi_7 = {hi_hi_7, hi_lo_7};
  wire [4095:0] regroupLoadData_0_7 = {hi_7, lo_7};
  wire [2047:0] dataGroup_lo_2304 = {dataGroup_lo_hi_2304, dataGroup_lo_lo_2304};
  wire [2047:0] dataGroup_hi_2304 = {dataGroup_hi_hi_2304, dataGroup_hi_lo_2304};
  wire [15:0]   dataGroup_0_36 = dataGroup_lo_2304[15:0];
  wire [2047:0] dataGroup_lo_2305 = {dataGroup_lo_hi_2305, dataGroup_lo_lo_2305};
  wire [2047:0] dataGroup_hi_2305 = {dataGroup_hi_hi_2305, dataGroup_hi_lo_2305};
  wire [15:0]   dataGroup_1_36 = dataGroup_lo_2305[31:16];
  wire [2047:0] dataGroup_lo_2306 = {dataGroup_lo_hi_2306, dataGroup_lo_lo_2306};
  wire [2047:0] dataGroup_hi_2306 = {dataGroup_hi_hi_2306, dataGroup_hi_lo_2306};
  wire [15:0]   dataGroup_2_36 = dataGroup_lo_2306[47:32];
  wire [2047:0] dataGroup_lo_2307 = {dataGroup_lo_hi_2307, dataGroup_lo_lo_2307};
  wire [2047:0] dataGroup_hi_2307 = {dataGroup_hi_hi_2307, dataGroup_hi_lo_2307};
  wire [15:0]   dataGroup_3_36 = dataGroup_lo_2307[63:48];
  wire [2047:0] dataGroup_lo_2308 = {dataGroup_lo_hi_2308, dataGroup_lo_lo_2308};
  wire [2047:0] dataGroup_hi_2308 = {dataGroup_hi_hi_2308, dataGroup_hi_lo_2308};
  wire [15:0]   dataGroup_4_36 = dataGroup_lo_2308[79:64];
  wire [2047:0] dataGroup_lo_2309 = {dataGroup_lo_hi_2309, dataGroup_lo_lo_2309};
  wire [2047:0] dataGroup_hi_2309 = {dataGroup_hi_hi_2309, dataGroup_hi_lo_2309};
  wire [15:0]   dataGroup_5_36 = dataGroup_lo_2309[95:80];
  wire [2047:0] dataGroup_lo_2310 = {dataGroup_lo_hi_2310, dataGroup_lo_lo_2310};
  wire [2047:0] dataGroup_hi_2310 = {dataGroup_hi_hi_2310, dataGroup_hi_lo_2310};
  wire [15:0]   dataGroup_6_36 = dataGroup_lo_2310[111:96];
  wire [2047:0] dataGroup_lo_2311 = {dataGroup_lo_hi_2311, dataGroup_lo_lo_2311};
  wire [2047:0] dataGroup_hi_2311 = {dataGroup_hi_hi_2311, dataGroup_hi_lo_2311};
  wire [15:0]   dataGroup_7_36 = dataGroup_lo_2311[127:112];
  wire [2047:0] dataGroup_lo_2312 = {dataGroup_lo_hi_2312, dataGroup_lo_lo_2312};
  wire [2047:0] dataGroup_hi_2312 = {dataGroup_hi_hi_2312, dataGroup_hi_lo_2312};
  wire [15:0]   dataGroup_8_36 = dataGroup_lo_2312[143:128];
  wire [2047:0] dataGroup_lo_2313 = {dataGroup_lo_hi_2313, dataGroup_lo_lo_2313};
  wire [2047:0] dataGroup_hi_2313 = {dataGroup_hi_hi_2313, dataGroup_hi_lo_2313};
  wire [15:0]   dataGroup_9_36 = dataGroup_lo_2313[159:144];
  wire [2047:0] dataGroup_lo_2314 = {dataGroup_lo_hi_2314, dataGroup_lo_lo_2314};
  wire [2047:0] dataGroup_hi_2314 = {dataGroup_hi_hi_2314, dataGroup_hi_lo_2314};
  wire [15:0]   dataGroup_10_36 = dataGroup_lo_2314[175:160];
  wire [2047:0] dataGroup_lo_2315 = {dataGroup_lo_hi_2315, dataGroup_lo_lo_2315};
  wire [2047:0] dataGroup_hi_2315 = {dataGroup_hi_hi_2315, dataGroup_hi_lo_2315};
  wire [15:0]   dataGroup_11_36 = dataGroup_lo_2315[191:176];
  wire [2047:0] dataGroup_lo_2316 = {dataGroup_lo_hi_2316, dataGroup_lo_lo_2316};
  wire [2047:0] dataGroup_hi_2316 = {dataGroup_hi_hi_2316, dataGroup_hi_lo_2316};
  wire [15:0]   dataGroup_12_36 = dataGroup_lo_2316[207:192];
  wire [2047:0] dataGroup_lo_2317 = {dataGroup_lo_hi_2317, dataGroup_lo_lo_2317};
  wire [2047:0] dataGroup_hi_2317 = {dataGroup_hi_hi_2317, dataGroup_hi_lo_2317};
  wire [15:0]   dataGroup_13_36 = dataGroup_lo_2317[223:208];
  wire [2047:0] dataGroup_lo_2318 = {dataGroup_lo_hi_2318, dataGroup_lo_lo_2318};
  wire [2047:0] dataGroup_hi_2318 = {dataGroup_hi_hi_2318, dataGroup_hi_lo_2318};
  wire [15:0]   dataGroup_14_36 = dataGroup_lo_2318[239:224];
  wire [2047:0] dataGroup_lo_2319 = {dataGroup_lo_hi_2319, dataGroup_lo_lo_2319};
  wire [2047:0] dataGroup_hi_2319 = {dataGroup_hi_hi_2319, dataGroup_hi_lo_2319};
  wire [15:0]   dataGroup_15_36 = dataGroup_lo_2319[255:240];
  wire [2047:0] dataGroup_lo_2320 = {dataGroup_lo_hi_2320, dataGroup_lo_lo_2320};
  wire [2047:0] dataGroup_hi_2320 = {dataGroup_hi_hi_2320, dataGroup_hi_lo_2320};
  wire [15:0]   dataGroup_16_36 = dataGroup_lo_2320[271:256];
  wire [2047:0] dataGroup_lo_2321 = {dataGroup_lo_hi_2321, dataGroup_lo_lo_2321};
  wire [2047:0] dataGroup_hi_2321 = {dataGroup_hi_hi_2321, dataGroup_hi_lo_2321};
  wire [15:0]   dataGroup_17_36 = dataGroup_lo_2321[287:272];
  wire [2047:0] dataGroup_lo_2322 = {dataGroup_lo_hi_2322, dataGroup_lo_lo_2322};
  wire [2047:0] dataGroup_hi_2322 = {dataGroup_hi_hi_2322, dataGroup_hi_lo_2322};
  wire [15:0]   dataGroup_18_36 = dataGroup_lo_2322[303:288];
  wire [2047:0] dataGroup_lo_2323 = {dataGroup_lo_hi_2323, dataGroup_lo_lo_2323};
  wire [2047:0] dataGroup_hi_2323 = {dataGroup_hi_hi_2323, dataGroup_hi_lo_2323};
  wire [15:0]   dataGroup_19_36 = dataGroup_lo_2323[319:304];
  wire [2047:0] dataGroup_lo_2324 = {dataGroup_lo_hi_2324, dataGroup_lo_lo_2324};
  wire [2047:0] dataGroup_hi_2324 = {dataGroup_hi_hi_2324, dataGroup_hi_lo_2324};
  wire [15:0]   dataGroup_20_36 = dataGroup_lo_2324[335:320];
  wire [2047:0] dataGroup_lo_2325 = {dataGroup_lo_hi_2325, dataGroup_lo_lo_2325};
  wire [2047:0] dataGroup_hi_2325 = {dataGroup_hi_hi_2325, dataGroup_hi_lo_2325};
  wire [15:0]   dataGroup_21_36 = dataGroup_lo_2325[351:336];
  wire [2047:0] dataGroup_lo_2326 = {dataGroup_lo_hi_2326, dataGroup_lo_lo_2326};
  wire [2047:0] dataGroup_hi_2326 = {dataGroup_hi_hi_2326, dataGroup_hi_lo_2326};
  wire [15:0]   dataGroup_22_36 = dataGroup_lo_2326[367:352];
  wire [2047:0] dataGroup_lo_2327 = {dataGroup_lo_hi_2327, dataGroup_lo_lo_2327};
  wire [2047:0] dataGroup_hi_2327 = {dataGroup_hi_hi_2327, dataGroup_hi_lo_2327};
  wire [15:0]   dataGroup_23_36 = dataGroup_lo_2327[383:368];
  wire [2047:0] dataGroup_lo_2328 = {dataGroup_lo_hi_2328, dataGroup_lo_lo_2328};
  wire [2047:0] dataGroup_hi_2328 = {dataGroup_hi_hi_2328, dataGroup_hi_lo_2328};
  wire [15:0]   dataGroup_24_36 = dataGroup_lo_2328[399:384];
  wire [2047:0] dataGroup_lo_2329 = {dataGroup_lo_hi_2329, dataGroup_lo_lo_2329};
  wire [2047:0] dataGroup_hi_2329 = {dataGroup_hi_hi_2329, dataGroup_hi_lo_2329};
  wire [15:0]   dataGroup_25_36 = dataGroup_lo_2329[415:400];
  wire [2047:0] dataGroup_lo_2330 = {dataGroup_lo_hi_2330, dataGroup_lo_lo_2330};
  wire [2047:0] dataGroup_hi_2330 = {dataGroup_hi_hi_2330, dataGroup_hi_lo_2330};
  wire [15:0]   dataGroup_26_36 = dataGroup_lo_2330[431:416];
  wire [2047:0] dataGroup_lo_2331 = {dataGroup_lo_hi_2331, dataGroup_lo_lo_2331};
  wire [2047:0] dataGroup_hi_2331 = {dataGroup_hi_hi_2331, dataGroup_hi_lo_2331};
  wire [15:0]   dataGroup_27_36 = dataGroup_lo_2331[447:432];
  wire [2047:0] dataGroup_lo_2332 = {dataGroup_lo_hi_2332, dataGroup_lo_lo_2332};
  wire [2047:0] dataGroup_hi_2332 = {dataGroup_hi_hi_2332, dataGroup_hi_lo_2332};
  wire [15:0]   dataGroup_28_36 = dataGroup_lo_2332[463:448];
  wire [2047:0] dataGroup_lo_2333 = {dataGroup_lo_hi_2333, dataGroup_lo_lo_2333};
  wire [2047:0] dataGroup_hi_2333 = {dataGroup_hi_hi_2333, dataGroup_hi_lo_2333};
  wire [15:0]   dataGroup_29_36 = dataGroup_lo_2333[479:464];
  wire [2047:0] dataGroup_lo_2334 = {dataGroup_lo_hi_2334, dataGroup_lo_lo_2334};
  wire [2047:0] dataGroup_hi_2334 = {dataGroup_hi_hi_2334, dataGroup_hi_lo_2334};
  wire [15:0]   dataGroup_30_36 = dataGroup_lo_2334[495:480];
  wire [2047:0] dataGroup_lo_2335 = {dataGroup_lo_hi_2335, dataGroup_lo_lo_2335};
  wire [2047:0] dataGroup_hi_2335 = {dataGroup_hi_hi_2335, dataGroup_hi_lo_2335};
  wire [15:0]   dataGroup_31_36 = dataGroup_lo_2335[511:496];
  wire [31:0]   res_lo_lo_lo_lo_36 = {dataGroup_1_36, dataGroup_0_36};
  wire [31:0]   res_lo_lo_lo_hi_36 = {dataGroup_3_36, dataGroup_2_36};
  wire [63:0]   res_lo_lo_lo_36 = {res_lo_lo_lo_hi_36, res_lo_lo_lo_lo_36};
  wire [31:0]   res_lo_lo_hi_lo_36 = {dataGroup_5_36, dataGroup_4_36};
  wire [31:0]   res_lo_lo_hi_hi_36 = {dataGroup_7_36, dataGroup_6_36};
  wire [63:0]   res_lo_lo_hi_36 = {res_lo_lo_hi_hi_36, res_lo_lo_hi_lo_36};
  wire [127:0]  res_lo_lo_36 = {res_lo_lo_hi_36, res_lo_lo_lo_36};
  wire [31:0]   res_lo_hi_lo_lo_36 = {dataGroup_9_36, dataGroup_8_36};
  wire [31:0]   res_lo_hi_lo_hi_36 = {dataGroup_11_36, dataGroup_10_36};
  wire [63:0]   res_lo_hi_lo_36 = {res_lo_hi_lo_hi_36, res_lo_hi_lo_lo_36};
  wire [31:0]   res_lo_hi_hi_lo_36 = {dataGroup_13_36, dataGroup_12_36};
  wire [31:0]   res_lo_hi_hi_hi_36 = {dataGroup_15_36, dataGroup_14_36};
  wire [63:0]   res_lo_hi_hi_36 = {res_lo_hi_hi_hi_36, res_lo_hi_hi_lo_36};
  wire [127:0]  res_lo_hi_36 = {res_lo_hi_hi_36, res_lo_hi_lo_36};
  wire [255:0]  res_lo_36 = {res_lo_hi_36, res_lo_lo_36};
  wire [31:0]   res_hi_lo_lo_lo_36 = {dataGroup_17_36, dataGroup_16_36};
  wire [31:0]   res_hi_lo_lo_hi_36 = {dataGroup_19_36, dataGroup_18_36};
  wire [63:0]   res_hi_lo_lo_36 = {res_hi_lo_lo_hi_36, res_hi_lo_lo_lo_36};
  wire [31:0]   res_hi_lo_hi_lo_36 = {dataGroup_21_36, dataGroup_20_36};
  wire [31:0]   res_hi_lo_hi_hi_36 = {dataGroup_23_36, dataGroup_22_36};
  wire [63:0]   res_hi_lo_hi_36 = {res_hi_lo_hi_hi_36, res_hi_lo_hi_lo_36};
  wire [127:0]  res_hi_lo_36 = {res_hi_lo_hi_36, res_hi_lo_lo_36};
  wire [31:0]   res_hi_hi_lo_lo_36 = {dataGroup_25_36, dataGroup_24_36};
  wire [31:0]   res_hi_hi_lo_hi_36 = {dataGroup_27_36, dataGroup_26_36};
  wire [63:0]   res_hi_hi_lo_36 = {res_hi_hi_lo_hi_36, res_hi_hi_lo_lo_36};
  wire [31:0]   res_hi_hi_hi_lo_36 = {dataGroup_29_36, dataGroup_28_36};
  wire [31:0]   res_hi_hi_hi_hi_36 = {dataGroup_31_36, dataGroup_30_36};
  wire [63:0]   res_hi_hi_hi_36 = {res_hi_hi_hi_hi_36, res_hi_hi_hi_lo_36};
  wire [127:0]  res_hi_hi_36 = {res_hi_hi_hi_36, res_hi_hi_lo_36};
  wire [255:0]  res_hi_36 = {res_hi_hi_36, res_hi_lo_36};
  wire [511:0]  res_64 = {res_hi_36, res_lo_36};
  wire [1023:0] lo_lo_8 = {512'h0, res_64};
  wire [2047:0] lo_8 = {1024'h0, lo_lo_8};
  wire [4095:0] regroupLoadData_1_0 = {2048'h0, lo_8};
  wire [2047:0] dataGroup_lo_2336 = {dataGroup_lo_hi_2336, dataGroup_lo_lo_2336};
  wire [2047:0] dataGroup_hi_2336 = {dataGroup_hi_hi_2336, dataGroup_hi_lo_2336};
  wire [15:0]   dataGroup_0_37 = dataGroup_lo_2336[15:0];
  wire [2047:0] dataGroup_lo_2337 = {dataGroup_lo_hi_2337, dataGroup_lo_lo_2337};
  wire [2047:0] dataGroup_hi_2337 = {dataGroup_hi_hi_2337, dataGroup_hi_lo_2337};
  wire [15:0]   dataGroup_1_37 = dataGroup_lo_2337[47:32];
  wire [2047:0] dataGroup_lo_2338 = {dataGroup_lo_hi_2338, dataGroup_lo_lo_2338};
  wire [2047:0] dataGroup_hi_2338 = {dataGroup_hi_hi_2338, dataGroup_hi_lo_2338};
  wire [15:0]   dataGroup_2_37 = dataGroup_lo_2338[79:64];
  wire [2047:0] dataGroup_lo_2339 = {dataGroup_lo_hi_2339, dataGroup_lo_lo_2339};
  wire [2047:0] dataGroup_hi_2339 = {dataGroup_hi_hi_2339, dataGroup_hi_lo_2339};
  wire [15:0]   dataGroup_3_37 = dataGroup_lo_2339[111:96];
  wire [2047:0] dataGroup_lo_2340 = {dataGroup_lo_hi_2340, dataGroup_lo_lo_2340};
  wire [2047:0] dataGroup_hi_2340 = {dataGroup_hi_hi_2340, dataGroup_hi_lo_2340};
  wire [15:0]   dataGroup_4_37 = dataGroup_lo_2340[143:128];
  wire [2047:0] dataGroup_lo_2341 = {dataGroup_lo_hi_2341, dataGroup_lo_lo_2341};
  wire [2047:0] dataGroup_hi_2341 = {dataGroup_hi_hi_2341, dataGroup_hi_lo_2341};
  wire [15:0]   dataGroup_5_37 = dataGroup_lo_2341[175:160];
  wire [2047:0] dataGroup_lo_2342 = {dataGroup_lo_hi_2342, dataGroup_lo_lo_2342};
  wire [2047:0] dataGroup_hi_2342 = {dataGroup_hi_hi_2342, dataGroup_hi_lo_2342};
  wire [15:0]   dataGroup_6_37 = dataGroup_lo_2342[207:192];
  wire [2047:0] dataGroup_lo_2343 = {dataGroup_lo_hi_2343, dataGroup_lo_lo_2343};
  wire [2047:0] dataGroup_hi_2343 = {dataGroup_hi_hi_2343, dataGroup_hi_lo_2343};
  wire [15:0]   dataGroup_7_37 = dataGroup_lo_2343[239:224];
  wire [2047:0] dataGroup_lo_2344 = {dataGroup_lo_hi_2344, dataGroup_lo_lo_2344};
  wire [2047:0] dataGroup_hi_2344 = {dataGroup_hi_hi_2344, dataGroup_hi_lo_2344};
  wire [15:0]   dataGroup_8_37 = dataGroup_lo_2344[271:256];
  wire [2047:0] dataGroup_lo_2345 = {dataGroup_lo_hi_2345, dataGroup_lo_lo_2345};
  wire [2047:0] dataGroup_hi_2345 = {dataGroup_hi_hi_2345, dataGroup_hi_lo_2345};
  wire [15:0]   dataGroup_9_37 = dataGroup_lo_2345[303:288];
  wire [2047:0] dataGroup_lo_2346 = {dataGroup_lo_hi_2346, dataGroup_lo_lo_2346};
  wire [2047:0] dataGroup_hi_2346 = {dataGroup_hi_hi_2346, dataGroup_hi_lo_2346};
  wire [15:0]   dataGroup_10_37 = dataGroup_lo_2346[335:320];
  wire [2047:0] dataGroup_lo_2347 = {dataGroup_lo_hi_2347, dataGroup_lo_lo_2347};
  wire [2047:0] dataGroup_hi_2347 = {dataGroup_hi_hi_2347, dataGroup_hi_lo_2347};
  wire [15:0]   dataGroup_11_37 = dataGroup_lo_2347[367:352];
  wire [2047:0] dataGroup_lo_2348 = {dataGroup_lo_hi_2348, dataGroup_lo_lo_2348};
  wire [2047:0] dataGroup_hi_2348 = {dataGroup_hi_hi_2348, dataGroup_hi_lo_2348};
  wire [15:0]   dataGroup_12_37 = dataGroup_lo_2348[399:384];
  wire [2047:0] dataGroup_lo_2349 = {dataGroup_lo_hi_2349, dataGroup_lo_lo_2349};
  wire [2047:0] dataGroup_hi_2349 = {dataGroup_hi_hi_2349, dataGroup_hi_lo_2349};
  wire [15:0]   dataGroup_13_37 = dataGroup_lo_2349[431:416];
  wire [2047:0] dataGroup_lo_2350 = {dataGroup_lo_hi_2350, dataGroup_lo_lo_2350};
  wire [2047:0] dataGroup_hi_2350 = {dataGroup_hi_hi_2350, dataGroup_hi_lo_2350};
  wire [15:0]   dataGroup_14_37 = dataGroup_lo_2350[463:448];
  wire [2047:0] dataGroup_lo_2351 = {dataGroup_lo_hi_2351, dataGroup_lo_lo_2351};
  wire [2047:0] dataGroup_hi_2351 = {dataGroup_hi_hi_2351, dataGroup_hi_lo_2351};
  wire [15:0]   dataGroup_15_37 = dataGroup_lo_2351[495:480];
  wire [2047:0] dataGroup_lo_2352 = {dataGroup_lo_hi_2352, dataGroup_lo_lo_2352};
  wire [2047:0] dataGroup_hi_2352 = {dataGroup_hi_hi_2352, dataGroup_hi_lo_2352};
  wire [15:0]   dataGroup_16_37 = dataGroup_lo_2352[527:512];
  wire [2047:0] dataGroup_lo_2353 = {dataGroup_lo_hi_2353, dataGroup_lo_lo_2353};
  wire [2047:0] dataGroup_hi_2353 = {dataGroup_hi_hi_2353, dataGroup_hi_lo_2353};
  wire [15:0]   dataGroup_17_37 = dataGroup_lo_2353[559:544];
  wire [2047:0] dataGroup_lo_2354 = {dataGroup_lo_hi_2354, dataGroup_lo_lo_2354};
  wire [2047:0] dataGroup_hi_2354 = {dataGroup_hi_hi_2354, dataGroup_hi_lo_2354};
  wire [15:0]   dataGroup_18_37 = dataGroup_lo_2354[591:576];
  wire [2047:0] dataGroup_lo_2355 = {dataGroup_lo_hi_2355, dataGroup_lo_lo_2355};
  wire [2047:0] dataGroup_hi_2355 = {dataGroup_hi_hi_2355, dataGroup_hi_lo_2355};
  wire [15:0]   dataGroup_19_37 = dataGroup_lo_2355[623:608];
  wire [2047:0] dataGroup_lo_2356 = {dataGroup_lo_hi_2356, dataGroup_lo_lo_2356};
  wire [2047:0] dataGroup_hi_2356 = {dataGroup_hi_hi_2356, dataGroup_hi_lo_2356};
  wire [15:0]   dataGroup_20_37 = dataGroup_lo_2356[655:640];
  wire [2047:0] dataGroup_lo_2357 = {dataGroup_lo_hi_2357, dataGroup_lo_lo_2357};
  wire [2047:0] dataGroup_hi_2357 = {dataGroup_hi_hi_2357, dataGroup_hi_lo_2357};
  wire [15:0]   dataGroup_21_37 = dataGroup_lo_2357[687:672];
  wire [2047:0] dataGroup_lo_2358 = {dataGroup_lo_hi_2358, dataGroup_lo_lo_2358};
  wire [2047:0] dataGroup_hi_2358 = {dataGroup_hi_hi_2358, dataGroup_hi_lo_2358};
  wire [15:0]   dataGroup_22_37 = dataGroup_lo_2358[719:704];
  wire [2047:0] dataGroup_lo_2359 = {dataGroup_lo_hi_2359, dataGroup_lo_lo_2359};
  wire [2047:0] dataGroup_hi_2359 = {dataGroup_hi_hi_2359, dataGroup_hi_lo_2359};
  wire [15:0]   dataGroup_23_37 = dataGroup_lo_2359[751:736];
  wire [2047:0] dataGroup_lo_2360 = {dataGroup_lo_hi_2360, dataGroup_lo_lo_2360};
  wire [2047:0] dataGroup_hi_2360 = {dataGroup_hi_hi_2360, dataGroup_hi_lo_2360};
  wire [15:0]   dataGroup_24_37 = dataGroup_lo_2360[783:768];
  wire [2047:0] dataGroup_lo_2361 = {dataGroup_lo_hi_2361, dataGroup_lo_lo_2361};
  wire [2047:0] dataGroup_hi_2361 = {dataGroup_hi_hi_2361, dataGroup_hi_lo_2361};
  wire [15:0]   dataGroup_25_37 = dataGroup_lo_2361[815:800];
  wire [2047:0] dataGroup_lo_2362 = {dataGroup_lo_hi_2362, dataGroup_lo_lo_2362};
  wire [2047:0] dataGroup_hi_2362 = {dataGroup_hi_hi_2362, dataGroup_hi_lo_2362};
  wire [15:0]   dataGroup_26_37 = dataGroup_lo_2362[847:832];
  wire [2047:0] dataGroup_lo_2363 = {dataGroup_lo_hi_2363, dataGroup_lo_lo_2363};
  wire [2047:0] dataGroup_hi_2363 = {dataGroup_hi_hi_2363, dataGroup_hi_lo_2363};
  wire [15:0]   dataGroup_27_37 = dataGroup_lo_2363[879:864];
  wire [2047:0] dataGroup_lo_2364 = {dataGroup_lo_hi_2364, dataGroup_lo_lo_2364};
  wire [2047:0] dataGroup_hi_2364 = {dataGroup_hi_hi_2364, dataGroup_hi_lo_2364};
  wire [15:0]   dataGroup_28_37 = dataGroup_lo_2364[911:896];
  wire [2047:0] dataGroup_lo_2365 = {dataGroup_lo_hi_2365, dataGroup_lo_lo_2365};
  wire [2047:0] dataGroup_hi_2365 = {dataGroup_hi_hi_2365, dataGroup_hi_lo_2365};
  wire [15:0]   dataGroup_29_37 = dataGroup_lo_2365[943:928];
  wire [2047:0] dataGroup_lo_2366 = {dataGroup_lo_hi_2366, dataGroup_lo_lo_2366};
  wire [2047:0] dataGroup_hi_2366 = {dataGroup_hi_hi_2366, dataGroup_hi_lo_2366};
  wire [15:0]   dataGroup_30_37 = dataGroup_lo_2366[975:960];
  wire [2047:0] dataGroup_lo_2367 = {dataGroup_lo_hi_2367, dataGroup_lo_lo_2367};
  wire [2047:0] dataGroup_hi_2367 = {dataGroup_hi_hi_2367, dataGroup_hi_lo_2367};
  wire [15:0]   dataGroup_31_37 = dataGroup_lo_2367[1007:992];
  wire [31:0]   res_lo_lo_lo_lo_37 = {dataGroup_1_37, dataGroup_0_37};
  wire [31:0]   res_lo_lo_lo_hi_37 = {dataGroup_3_37, dataGroup_2_37};
  wire [63:0]   res_lo_lo_lo_37 = {res_lo_lo_lo_hi_37, res_lo_lo_lo_lo_37};
  wire [31:0]   res_lo_lo_hi_lo_37 = {dataGroup_5_37, dataGroup_4_37};
  wire [31:0]   res_lo_lo_hi_hi_37 = {dataGroup_7_37, dataGroup_6_37};
  wire [63:0]   res_lo_lo_hi_37 = {res_lo_lo_hi_hi_37, res_lo_lo_hi_lo_37};
  wire [127:0]  res_lo_lo_37 = {res_lo_lo_hi_37, res_lo_lo_lo_37};
  wire [31:0]   res_lo_hi_lo_lo_37 = {dataGroup_9_37, dataGroup_8_37};
  wire [31:0]   res_lo_hi_lo_hi_37 = {dataGroup_11_37, dataGroup_10_37};
  wire [63:0]   res_lo_hi_lo_37 = {res_lo_hi_lo_hi_37, res_lo_hi_lo_lo_37};
  wire [31:0]   res_lo_hi_hi_lo_37 = {dataGroup_13_37, dataGroup_12_37};
  wire [31:0]   res_lo_hi_hi_hi_37 = {dataGroup_15_37, dataGroup_14_37};
  wire [63:0]   res_lo_hi_hi_37 = {res_lo_hi_hi_hi_37, res_lo_hi_hi_lo_37};
  wire [127:0]  res_lo_hi_37 = {res_lo_hi_hi_37, res_lo_hi_lo_37};
  wire [255:0]  res_lo_37 = {res_lo_hi_37, res_lo_lo_37};
  wire [31:0]   res_hi_lo_lo_lo_37 = {dataGroup_17_37, dataGroup_16_37};
  wire [31:0]   res_hi_lo_lo_hi_37 = {dataGroup_19_37, dataGroup_18_37};
  wire [63:0]   res_hi_lo_lo_37 = {res_hi_lo_lo_hi_37, res_hi_lo_lo_lo_37};
  wire [31:0]   res_hi_lo_hi_lo_37 = {dataGroup_21_37, dataGroup_20_37};
  wire [31:0]   res_hi_lo_hi_hi_37 = {dataGroup_23_37, dataGroup_22_37};
  wire [63:0]   res_hi_lo_hi_37 = {res_hi_lo_hi_hi_37, res_hi_lo_hi_lo_37};
  wire [127:0]  res_hi_lo_37 = {res_hi_lo_hi_37, res_hi_lo_lo_37};
  wire [31:0]   res_hi_hi_lo_lo_37 = {dataGroup_25_37, dataGroup_24_37};
  wire [31:0]   res_hi_hi_lo_hi_37 = {dataGroup_27_37, dataGroup_26_37};
  wire [63:0]   res_hi_hi_lo_37 = {res_hi_hi_lo_hi_37, res_hi_hi_lo_lo_37};
  wire [31:0]   res_hi_hi_hi_lo_37 = {dataGroup_29_37, dataGroup_28_37};
  wire [31:0]   res_hi_hi_hi_hi_37 = {dataGroup_31_37, dataGroup_30_37};
  wire [63:0]   res_hi_hi_hi_37 = {res_hi_hi_hi_hi_37, res_hi_hi_hi_lo_37};
  wire [127:0]  res_hi_hi_37 = {res_hi_hi_hi_37, res_hi_hi_lo_37};
  wire [255:0]  res_hi_37 = {res_hi_hi_37, res_hi_lo_37};
  wire [511:0]  res_72 = {res_hi_37, res_lo_37};
  wire [2047:0] dataGroup_lo_2368 = {dataGroup_lo_hi_2368, dataGroup_lo_lo_2368};
  wire [2047:0] dataGroup_hi_2368 = {dataGroup_hi_hi_2368, dataGroup_hi_lo_2368};
  wire [15:0]   dataGroup_0_38 = dataGroup_lo_2368[31:16];
  wire [2047:0] dataGroup_lo_2369 = {dataGroup_lo_hi_2369, dataGroup_lo_lo_2369};
  wire [2047:0] dataGroup_hi_2369 = {dataGroup_hi_hi_2369, dataGroup_hi_lo_2369};
  wire [15:0]   dataGroup_1_38 = dataGroup_lo_2369[63:48];
  wire [2047:0] dataGroup_lo_2370 = {dataGroup_lo_hi_2370, dataGroup_lo_lo_2370};
  wire [2047:0] dataGroup_hi_2370 = {dataGroup_hi_hi_2370, dataGroup_hi_lo_2370};
  wire [15:0]   dataGroup_2_38 = dataGroup_lo_2370[95:80];
  wire [2047:0] dataGroup_lo_2371 = {dataGroup_lo_hi_2371, dataGroup_lo_lo_2371};
  wire [2047:0] dataGroup_hi_2371 = {dataGroup_hi_hi_2371, dataGroup_hi_lo_2371};
  wire [15:0]   dataGroup_3_38 = dataGroup_lo_2371[127:112];
  wire [2047:0] dataGroup_lo_2372 = {dataGroup_lo_hi_2372, dataGroup_lo_lo_2372};
  wire [2047:0] dataGroup_hi_2372 = {dataGroup_hi_hi_2372, dataGroup_hi_lo_2372};
  wire [15:0]   dataGroup_4_38 = dataGroup_lo_2372[159:144];
  wire [2047:0] dataGroup_lo_2373 = {dataGroup_lo_hi_2373, dataGroup_lo_lo_2373};
  wire [2047:0] dataGroup_hi_2373 = {dataGroup_hi_hi_2373, dataGroup_hi_lo_2373};
  wire [15:0]   dataGroup_5_38 = dataGroup_lo_2373[191:176];
  wire [2047:0] dataGroup_lo_2374 = {dataGroup_lo_hi_2374, dataGroup_lo_lo_2374};
  wire [2047:0] dataGroup_hi_2374 = {dataGroup_hi_hi_2374, dataGroup_hi_lo_2374};
  wire [15:0]   dataGroup_6_38 = dataGroup_lo_2374[223:208];
  wire [2047:0] dataGroup_lo_2375 = {dataGroup_lo_hi_2375, dataGroup_lo_lo_2375};
  wire [2047:0] dataGroup_hi_2375 = {dataGroup_hi_hi_2375, dataGroup_hi_lo_2375};
  wire [15:0]   dataGroup_7_38 = dataGroup_lo_2375[255:240];
  wire [2047:0] dataGroup_lo_2376 = {dataGroup_lo_hi_2376, dataGroup_lo_lo_2376};
  wire [2047:0] dataGroup_hi_2376 = {dataGroup_hi_hi_2376, dataGroup_hi_lo_2376};
  wire [15:0]   dataGroup_8_38 = dataGroup_lo_2376[287:272];
  wire [2047:0] dataGroup_lo_2377 = {dataGroup_lo_hi_2377, dataGroup_lo_lo_2377};
  wire [2047:0] dataGroup_hi_2377 = {dataGroup_hi_hi_2377, dataGroup_hi_lo_2377};
  wire [15:0]   dataGroup_9_38 = dataGroup_lo_2377[319:304];
  wire [2047:0] dataGroup_lo_2378 = {dataGroup_lo_hi_2378, dataGroup_lo_lo_2378};
  wire [2047:0] dataGroup_hi_2378 = {dataGroup_hi_hi_2378, dataGroup_hi_lo_2378};
  wire [15:0]   dataGroup_10_38 = dataGroup_lo_2378[351:336];
  wire [2047:0] dataGroup_lo_2379 = {dataGroup_lo_hi_2379, dataGroup_lo_lo_2379};
  wire [2047:0] dataGroup_hi_2379 = {dataGroup_hi_hi_2379, dataGroup_hi_lo_2379};
  wire [15:0]   dataGroup_11_38 = dataGroup_lo_2379[383:368];
  wire [2047:0] dataGroup_lo_2380 = {dataGroup_lo_hi_2380, dataGroup_lo_lo_2380};
  wire [2047:0] dataGroup_hi_2380 = {dataGroup_hi_hi_2380, dataGroup_hi_lo_2380};
  wire [15:0]   dataGroup_12_38 = dataGroup_lo_2380[415:400];
  wire [2047:0] dataGroup_lo_2381 = {dataGroup_lo_hi_2381, dataGroup_lo_lo_2381};
  wire [2047:0] dataGroup_hi_2381 = {dataGroup_hi_hi_2381, dataGroup_hi_lo_2381};
  wire [15:0]   dataGroup_13_38 = dataGroup_lo_2381[447:432];
  wire [2047:0] dataGroup_lo_2382 = {dataGroup_lo_hi_2382, dataGroup_lo_lo_2382};
  wire [2047:0] dataGroup_hi_2382 = {dataGroup_hi_hi_2382, dataGroup_hi_lo_2382};
  wire [15:0]   dataGroup_14_38 = dataGroup_lo_2382[479:464];
  wire [2047:0] dataGroup_lo_2383 = {dataGroup_lo_hi_2383, dataGroup_lo_lo_2383};
  wire [2047:0] dataGroup_hi_2383 = {dataGroup_hi_hi_2383, dataGroup_hi_lo_2383};
  wire [15:0]   dataGroup_15_38 = dataGroup_lo_2383[511:496];
  wire [2047:0] dataGroup_lo_2384 = {dataGroup_lo_hi_2384, dataGroup_lo_lo_2384};
  wire [2047:0] dataGroup_hi_2384 = {dataGroup_hi_hi_2384, dataGroup_hi_lo_2384};
  wire [15:0]   dataGroup_16_38 = dataGroup_lo_2384[543:528];
  wire [2047:0] dataGroup_lo_2385 = {dataGroup_lo_hi_2385, dataGroup_lo_lo_2385};
  wire [2047:0] dataGroup_hi_2385 = {dataGroup_hi_hi_2385, dataGroup_hi_lo_2385};
  wire [15:0]   dataGroup_17_38 = dataGroup_lo_2385[575:560];
  wire [2047:0] dataGroup_lo_2386 = {dataGroup_lo_hi_2386, dataGroup_lo_lo_2386};
  wire [2047:0] dataGroup_hi_2386 = {dataGroup_hi_hi_2386, dataGroup_hi_lo_2386};
  wire [15:0]   dataGroup_18_38 = dataGroup_lo_2386[607:592];
  wire [2047:0] dataGroup_lo_2387 = {dataGroup_lo_hi_2387, dataGroup_lo_lo_2387};
  wire [2047:0] dataGroup_hi_2387 = {dataGroup_hi_hi_2387, dataGroup_hi_lo_2387};
  wire [15:0]   dataGroup_19_38 = dataGroup_lo_2387[639:624];
  wire [2047:0] dataGroup_lo_2388 = {dataGroup_lo_hi_2388, dataGroup_lo_lo_2388};
  wire [2047:0] dataGroup_hi_2388 = {dataGroup_hi_hi_2388, dataGroup_hi_lo_2388};
  wire [15:0]   dataGroup_20_38 = dataGroup_lo_2388[671:656];
  wire [2047:0] dataGroup_lo_2389 = {dataGroup_lo_hi_2389, dataGroup_lo_lo_2389};
  wire [2047:0] dataGroup_hi_2389 = {dataGroup_hi_hi_2389, dataGroup_hi_lo_2389};
  wire [15:0]   dataGroup_21_38 = dataGroup_lo_2389[703:688];
  wire [2047:0] dataGroup_lo_2390 = {dataGroup_lo_hi_2390, dataGroup_lo_lo_2390};
  wire [2047:0] dataGroup_hi_2390 = {dataGroup_hi_hi_2390, dataGroup_hi_lo_2390};
  wire [15:0]   dataGroup_22_38 = dataGroup_lo_2390[735:720];
  wire [2047:0] dataGroup_lo_2391 = {dataGroup_lo_hi_2391, dataGroup_lo_lo_2391};
  wire [2047:0] dataGroup_hi_2391 = {dataGroup_hi_hi_2391, dataGroup_hi_lo_2391};
  wire [15:0]   dataGroup_23_38 = dataGroup_lo_2391[767:752];
  wire [2047:0] dataGroup_lo_2392 = {dataGroup_lo_hi_2392, dataGroup_lo_lo_2392};
  wire [2047:0] dataGroup_hi_2392 = {dataGroup_hi_hi_2392, dataGroup_hi_lo_2392};
  wire [15:0]   dataGroup_24_38 = dataGroup_lo_2392[799:784];
  wire [2047:0] dataGroup_lo_2393 = {dataGroup_lo_hi_2393, dataGroup_lo_lo_2393};
  wire [2047:0] dataGroup_hi_2393 = {dataGroup_hi_hi_2393, dataGroup_hi_lo_2393};
  wire [15:0]   dataGroup_25_38 = dataGroup_lo_2393[831:816];
  wire [2047:0] dataGroup_lo_2394 = {dataGroup_lo_hi_2394, dataGroup_lo_lo_2394};
  wire [2047:0] dataGroup_hi_2394 = {dataGroup_hi_hi_2394, dataGroup_hi_lo_2394};
  wire [15:0]   dataGroup_26_38 = dataGroup_lo_2394[863:848];
  wire [2047:0] dataGroup_lo_2395 = {dataGroup_lo_hi_2395, dataGroup_lo_lo_2395};
  wire [2047:0] dataGroup_hi_2395 = {dataGroup_hi_hi_2395, dataGroup_hi_lo_2395};
  wire [15:0]   dataGroup_27_38 = dataGroup_lo_2395[895:880];
  wire [2047:0] dataGroup_lo_2396 = {dataGroup_lo_hi_2396, dataGroup_lo_lo_2396};
  wire [2047:0] dataGroup_hi_2396 = {dataGroup_hi_hi_2396, dataGroup_hi_lo_2396};
  wire [15:0]   dataGroup_28_38 = dataGroup_lo_2396[927:912];
  wire [2047:0] dataGroup_lo_2397 = {dataGroup_lo_hi_2397, dataGroup_lo_lo_2397};
  wire [2047:0] dataGroup_hi_2397 = {dataGroup_hi_hi_2397, dataGroup_hi_lo_2397};
  wire [15:0]   dataGroup_29_38 = dataGroup_lo_2397[959:944];
  wire [2047:0] dataGroup_lo_2398 = {dataGroup_lo_hi_2398, dataGroup_lo_lo_2398};
  wire [2047:0] dataGroup_hi_2398 = {dataGroup_hi_hi_2398, dataGroup_hi_lo_2398};
  wire [15:0]   dataGroup_30_38 = dataGroup_lo_2398[991:976];
  wire [2047:0] dataGroup_lo_2399 = {dataGroup_lo_hi_2399, dataGroup_lo_lo_2399};
  wire [2047:0] dataGroup_hi_2399 = {dataGroup_hi_hi_2399, dataGroup_hi_lo_2399};
  wire [15:0]   dataGroup_31_38 = dataGroup_lo_2399[1023:1008];
  wire [31:0]   res_lo_lo_lo_lo_38 = {dataGroup_1_38, dataGroup_0_38};
  wire [31:0]   res_lo_lo_lo_hi_38 = {dataGroup_3_38, dataGroup_2_38};
  wire [63:0]   res_lo_lo_lo_38 = {res_lo_lo_lo_hi_38, res_lo_lo_lo_lo_38};
  wire [31:0]   res_lo_lo_hi_lo_38 = {dataGroup_5_38, dataGroup_4_38};
  wire [31:0]   res_lo_lo_hi_hi_38 = {dataGroup_7_38, dataGroup_6_38};
  wire [63:0]   res_lo_lo_hi_38 = {res_lo_lo_hi_hi_38, res_lo_lo_hi_lo_38};
  wire [127:0]  res_lo_lo_38 = {res_lo_lo_hi_38, res_lo_lo_lo_38};
  wire [31:0]   res_lo_hi_lo_lo_38 = {dataGroup_9_38, dataGroup_8_38};
  wire [31:0]   res_lo_hi_lo_hi_38 = {dataGroup_11_38, dataGroup_10_38};
  wire [63:0]   res_lo_hi_lo_38 = {res_lo_hi_lo_hi_38, res_lo_hi_lo_lo_38};
  wire [31:0]   res_lo_hi_hi_lo_38 = {dataGroup_13_38, dataGroup_12_38};
  wire [31:0]   res_lo_hi_hi_hi_38 = {dataGroup_15_38, dataGroup_14_38};
  wire [63:0]   res_lo_hi_hi_38 = {res_lo_hi_hi_hi_38, res_lo_hi_hi_lo_38};
  wire [127:0]  res_lo_hi_38 = {res_lo_hi_hi_38, res_lo_hi_lo_38};
  wire [255:0]  res_lo_38 = {res_lo_hi_38, res_lo_lo_38};
  wire [31:0]   res_hi_lo_lo_lo_38 = {dataGroup_17_38, dataGroup_16_38};
  wire [31:0]   res_hi_lo_lo_hi_38 = {dataGroup_19_38, dataGroup_18_38};
  wire [63:0]   res_hi_lo_lo_38 = {res_hi_lo_lo_hi_38, res_hi_lo_lo_lo_38};
  wire [31:0]   res_hi_lo_hi_lo_38 = {dataGroup_21_38, dataGroup_20_38};
  wire [31:0]   res_hi_lo_hi_hi_38 = {dataGroup_23_38, dataGroup_22_38};
  wire [63:0]   res_hi_lo_hi_38 = {res_hi_lo_hi_hi_38, res_hi_lo_hi_lo_38};
  wire [127:0]  res_hi_lo_38 = {res_hi_lo_hi_38, res_hi_lo_lo_38};
  wire [31:0]   res_hi_hi_lo_lo_38 = {dataGroup_25_38, dataGroup_24_38};
  wire [31:0]   res_hi_hi_lo_hi_38 = {dataGroup_27_38, dataGroup_26_38};
  wire [63:0]   res_hi_hi_lo_38 = {res_hi_hi_lo_hi_38, res_hi_hi_lo_lo_38};
  wire [31:0]   res_hi_hi_hi_lo_38 = {dataGroup_29_38, dataGroup_28_38};
  wire [31:0]   res_hi_hi_hi_hi_38 = {dataGroup_31_38, dataGroup_30_38};
  wire [63:0]   res_hi_hi_hi_38 = {res_hi_hi_hi_hi_38, res_hi_hi_hi_lo_38};
  wire [127:0]  res_hi_hi_38 = {res_hi_hi_hi_38, res_hi_hi_lo_38};
  wire [255:0]  res_hi_38 = {res_hi_hi_38, res_hi_lo_38};
  wire [511:0]  res_73 = {res_hi_38, res_lo_38};
  wire [1023:0] lo_lo_9 = {res_73, res_72};
  wire [2047:0] lo_9 = {1024'h0, lo_lo_9};
  wire [4095:0] regroupLoadData_1_1 = {2048'h0, lo_9};
  wire [2047:0] dataGroup_lo_2400 = {dataGroup_lo_hi_2400, dataGroup_lo_lo_2400};
  wire [2047:0] dataGroup_hi_2400 = {dataGroup_hi_hi_2400, dataGroup_hi_lo_2400};
  wire [15:0]   dataGroup_0_39 = dataGroup_lo_2400[15:0];
  wire [2047:0] dataGroup_lo_2401 = {dataGroup_lo_hi_2401, dataGroup_lo_lo_2401};
  wire [2047:0] dataGroup_hi_2401 = {dataGroup_hi_hi_2401, dataGroup_hi_lo_2401};
  wire [15:0]   dataGroup_1_39 = dataGroup_lo_2401[63:48];
  wire [2047:0] dataGroup_lo_2402 = {dataGroup_lo_hi_2402, dataGroup_lo_lo_2402};
  wire [2047:0] dataGroup_hi_2402 = {dataGroup_hi_hi_2402, dataGroup_hi_lo_2402};
  wire [15:0]   dataGroup_2_39 = dataGroup_lo_2402[111:96];
  wire [2047:0] dataGroup_lo_2403 = {dataGroup_lo_hi_2403, dataGroup_lo_lo_2403};
  wire [2047:0] dataGroup_hi_2403 = {dataGroup_hi_hi_2403, dataGroup_hi_lo_2403};
  wire [15:0]   dataGroup_3_39 = dataGroup_lo_2403[159:144];
  wire [2047:0] dataGroup_lo_2404 = {dataGroup_lo_hi_2404, dataGroup_lo_lo_2404};
  wire [2047:0] dataGroup_hi_2404 = {dataGroup_hi_hi_2404, dataGroup_hi_lo_2404};
  wire [15:0]   dataGroup_4_39 = dataGroup_lo_2404[207:192];
  wire [2047:0] dataGroup_lo_2405 = {dataGroup_lo_hi_2405, dataGroup_lo_lo_2405};
  wire [2047:0] dataGroup_hi_2405 = {dataGroup_hi_hi_2405, dataGroup_hi_lo_2405};
  wire [15:0]   dataGroup_5_39 = dataGroup_lo_2405[255:240];
  wire [2047:0] dataGroup_lo_2406 = {dataGroup_lo_hi_2406, dataGroup_lo_lo_2406};
  wire [2047:0] dataGroup_hi_2406 = {dataGroup_hi_hi_2406, dataGroup_hi_lo_2406};
  wire [15:0]   dataGroup_6_39 = dataGroup_lo_2406[303:288];
  wire [2047:0] dataGroup_lo_2407 = {dataGroup_lo_hi_2407, dataGroup_lo_lo_2407};
  wire [2047:0] dataGroup_hi_2407 = {dataGroup_hi_hi_2407, dataGroup_hi_lo_2407};
  wire [15:0]   dataGroup_7_39 = dataGroup_lo_2407[351:336];
  wire [2047:0] dataGroup_lo_2408 = {dataGroup_lo_hi_2408, dataGroup_lo_lo_2408};
  wire [2047:0] dataGroup_hi_2408 = {dataGroup_hi_hi_2408, dataGroup_hi_lo_2408};
  wire [15:0]   dataGroup_8_39 = dataGroup_lo_2408[399:384];
  wire [2047:0] dataGroup_lo_2409 = {dataGroup_lo_hi_2409, dataGroup_lo_lo_2409};
  wire [2047:0] dataGroup_hi_2409 = {dataGroup_hi_hi_2409, dataGroup_hi_lo_2409};
  wire [15:0]   dataGroup_9_39 = dataGroup_lo_2409[447:432];
  wire [2047:0] dataGroup_lo_2410 = {dataGroup_lo_hi_2410, dataGroup_lo_lo_2410};
  wire [2047:0] dataGroup_hi_2410 = {dataGroup_hi_hi_2410, dataGroup_hi_lo_2410};
  wire [15:0]   dataGroup_10_39 = dataGroup_lo_2410[495:480];
  wire [2047:0] dataGroup_lo_2411 = {dataGroup_lo_hi_2411, dataGroup_lo_lo_2411};
  wire [2047:0] dataGroup_hi_2411 = {dataGroup_hi_hi_2411, dataGroup_hi_lo_2411};
  wire [15:0]   dataGroup_11_39 = dataGroup_lo_2411[543:528];
  wire [2047:0] dataGroup_lo_2412 = {dataGroup_lo_hi_2412, dataGroup_lo_lo_2412};
  wire [2047:0] dataGroup_hi_2412 = {dataGroup_hi_hi_2412, dataGroup_hi_lo_2412};
  wire [15:0]   dataGroup_12_39 = dataGroup_lo_2412[591:576];
  wire [2047:0] dataGroup_lo_2413 = {dataGroup_lo_hi_2413, dataGroup_lo_lo_2413};
  wire [2047:0] dataGroup_hi_2413 = {dataGroup_hi_hi_2413, dataGroup_hi_lo_2413};
  wire [15:0]   dataGroup_13_39 = dataGroup_lo_2413[639:624];
  wire [2047:0] dataGroup_lo_2414 = {dataGroup_lo_hi_2414, dataGroup_lo_lo_2414};
  wire [2047:0] dataGroup_hi_2414 = {dataGroup_hi_hi_2414, dataGroup_hi_lo_2414};
  wire [15:0]   dataGroup_14_39 = dataGroup_lo_2414[687:672];
  wire [2047:0] dataGroup_lo_2415 = {dataGroup_lo_hi_2415, dataGroup_lo_lo_2415};
  wire [2047:0] dataGroup_hi_2415 = {dataGroup_hi_hi_2415, dataGroup_hi_lo_2415};
  wire [15:0]   dataGroup_15_39 = dataGroup_lo_2415[735:720];
  wire [2047:0] dataGroup_lo_2416 = {dataGroup_lo_hi_2416, dataGroup_lo_lo_2416};
  wire [2047:0] dataGroup_hi_2416 = {dataGroup_hi_hi_2416, dataGroup_hi_lo_2416};
  wire [15:0]   dataGroup_16_39 = dataGroup_lo_2416[783:768];
  wire [2047:0] dataGroup_lo_2417 = {dataGroup_lo_hi_2417, dataGroup_lo_lo_2417};
  wire [2047:0] dataGroup_hi_2417 = {dataGroup_hi_hi_2417, dataGroup_hi_lo_2417};
  wire [15:0]   dataGroup_17_39 = dataGroup_lo_2417[831:816];
  wire [2047:0] dataGroup_lo_2418 = {dataGroup_lo_hi_2418, dataGroup_lo_lo_2418};
  wire [2047:0] dataGroup_hi_2418 = {dataGroup_hi_hi_2418, dataGroup_hi_lo_2418};
  wire [15:0]   dataGroup_18_39 = dataGroup_lo_2418[879:864];
  wire [2047:0] dataGroup_lo_2419 = {dataGroup_lo_hi_2419, dataGroup_lo_lo_2419};
  wire [2047:0] dataGroup_hi_2419 = {dataGroup_hi_hi_2419, dataGroup_hi_lo_2419};
  wire [15:0]   dataGroup_19_39 = dataGroup_lo_2419[927:912];
  wire [2047:0] dataGroup_lo_2420 = {dataGroup_lo_hi_2420, dataGroup_lo_lo_2420};
  wire [2047:0] dataGroup_hi_2420 = {dataGroup_hi_hi_2420, dataGroup_hi_lo_2420};
  wire [15:0]   dataGroup_20_39 = dataGroup_lo_2420[975:960];
  wire [2047:0] dataGroup_lo_2421 = {dataGroup_lo_hi_2421, dataGroup_lo_lo_2421};
  wire [2047:0] dataGroup_hi_2421 = {dataGroup_hi_hi_2421, dataGroup_hi_lo_2421};
  wire [15:0]   dataGroup_21_39 = dataGroup_lo_2421[1023:1008];
  wire [2047:0] dataGroup_lo_2422 = {dataGroup_lo_hi_2422, dataGroup_lo_lo_2422};
  wire [2047:0] dataGroup_hi_2422 = {dataGroup_hi_hi_2422, dataGroup_hi_lo_2422};
  wire [15:0]   dataGroup_22_39 = dataGroup_lo_2422[1071:1056];
  wire [2047:0] dataGroup_lo_2423 = {dataGroup_lo_hi_2423, dataGroup_lo_lo_2423};
  wire [2047:0] dataGroup_hi_2423 = {dataGroup_hi_hi_2423, dataGroup_hi_lo_2423};
  wire [15:0]   dataGroup_23_39 = dataGroup_lo_2423[1119:1104];
  wire [2047:0] dataGroup_lo_2424 = {dataGroup_lo_hi_2424, dataGroup_lo_lo_2424};
  wire [2047:0] dataGroup_hi_2424 = {dataGroup_hi_hi_2424, dataGroup_hi_lo_2424};
  wire [15:0]   dataGroup_24_39 = dataGroup_lo_2424[1167:1152];
  wire [2047:0] dataGroup_lo_2425 = {dataGroup_lo_hi_2425, dataGroup_lo_lo_2425};
  wire [2047:0] dataGroup_hi_2425 = {dataGroup_hi_hi_2425, dataGroup_hi_lo_2425};
  wire [15:0]   dataGroup_25_39 = dataGroup_lo_2425[1215:1200];
  wire [2047:0] dataGroup_lo_2426 = {dataGroup_lo_hi_2426, dataGroup_lo_lo_2426};
  wire [2047:0] dataGroup_hi_2426 = {dataGroup_hi_hi_2426, dataGroup_hi_lo_2426};
  wire [15:0]   dataGroup_26_39 = dataGroup_lo_2426[1263:1248];
  wire [2047:0] dataGroup_lo_2427 = {dataGroup_lo_hi_2427, dataGroup_lo_lo_2427};
  wire [2047:0] dataGroup_hi_2427 = {dataGroup_hi_hi_2427, dataGroup_hi_lo_2427};
  wire [15:0]   dataGroup_27_39 = dataGroup_lo_2427[1311:1296];
  wire [2047:0] dataGroup_lo_2428 = {dataGroup_lo_hi_2428, dataGroup_lo_lo_2428};
  wire [2047:0] dataGroup_hi_2428 = {dataGroup_hi_hi_2428, dataGroup_hi_lo_2428};
  wire [15:0]   dataGroup_28_39 = dataGroup_lo_2428[1359:1344];
  wire [2047:0] dataGroup_lo_2429 = {dataGroup_lo_hi_2429, dataGroup_lo_lo_2429};
  wire [2047:0] dataGroup_hi_2429 = {dataGroup_hi_hi_2429, dataGroup_hi_lo_2429};
  wire [15:0]   dataGroup_29_39 = dataGroup_lo_2429[1407:1392];
  wire [2047:0] dataGroup_lo_2430 = {dataGroup_lo_hi_2430, dataGroup_lo_lo_2430};
  wire [2047:0] dataGroup_hi_2430 = {dataGroup_hi_hi_2430, dataGroup_hi_lo_2430};
  wire [15:0]   dataGroup_30_39 = dataGroup_lo_2430[1455:1440];
  wire [2047:0] dataGroup_lo_2431 = {dataGroup_lo_hi_2431, dataGroup_lo_lo_2431};
  wire [2047:0] dataGroup_hi_2431 = {dataGroup_hi_hi_2431, dataGroup_hi_lo_2431};
  wire [15:0]   dataGroup_31_39 = dataGroup_lo_2431[1503:1488];
  wire [31:0]   res_lo_lo_lo_lo_39 = {dataGroup_1_39, dataGroup_0_39};
  wire [31:0]   res_lo_lo_lo_hi_39 = {dataGroup_3_39, dataGroup_2_39};
  wire [63:0]   res_lo_lo_lo_39 = {res_lo_lo_lo_hi_39, res_lo_lo_lo_lo_39};
  wire [31:0]   res_lo_lo_hi_lo_39 = {dataGroup_5_39, dataGroup_4_39};
  wire [31:0]   res_lo_lo_hi_hi_39 = {dataGroup_7_39, dataGroup_6_39};
  wire [63:0]   res_lo_lo_hi_39 = {res_lo_lo_hi_hi_39, res_lo_lo_hi_lo_39};
  wire [127:0]  res_lo_lo_39 = {res_lo_lo_hi_39, res_lo_lo_lo_39};
  wire [31:0]   res_lo_hi_lo_lo_39 = {dataGroup_9_39, dataGroup_8_39};
  wire [31:0]   res_lo_hi_lo_hi_39 = {dataGroup_11_39, dataGroup_10_39};
  wire [63:0]   res_lo_hi_lo_39 = {res_lo_hi_lo_hi_39, res_lo_hi_lo_lo_39};
  wire [31:0]   res_lo_hi_hi_lo_39 = {dataGroup_13_39, dataGroup_12_39};
  wire [31:0]   res_lo_hi_hi_hi_39 = {dataGroup_15_39, dataGroup_14_39};
  wire [63:0]   res_lo_hi_hi_39 = {res_lo_hi_hi_hi_39, res_lo_hi_hi_lo_39};
  wire [127:0]  res_lo_hi_39 = {res_lo_hi_hi_39, res_lo_hi_lo_39};
  wire [255:0]  res_lo_39 = {res_lo_hi_39, res_lo_lo_39};
  wire [31:0]   res_hi_lo_lo_lo_39 = {dataGroup_17_39, dataGroup_16_39};
  wire [31:0]   res_hi_lo_lo_hi_39 = {dataGroup_19_39, dataGroup_18_39};
  wire [63:0]   res_hi_lo_lo_39 = {res_hi_lo_lo_hi_39, res_hi_lo_lo_lo_39};
  wire [31:0]   res_hi_lo_hi_lo_39 = {dataGroup_21_39, dataGroup_20_39};
  wire [31:0]   res_hi_lo_hi_hi_39 = {dataGroup_23_39, dataGroup_22_39};
  wire [63:0]   res_hi_lo_hi_39 = {res_hi_lo_hi_hi_39, res_hi_lo_hi_lo_39};
  wire [127:0]  res_hi_lo_39 = {res_hi_lo_hi_39, res_hi_lo_lo_39};
  wire [31:0]   res_hi_hi_lo_lo_39 = {dataGroup_25_39, dataGroup_24_39};
  wire [31:0]   res_hi_hi_lo_hi_39 = {dataGroup_27_39, dataGroup_26_39};
  wire [63:0]   res_hi_hi_lo_39 = {res_hi_hi_lo_hi_39, res_hi_hi_lo_lo_39};
  wire [31:0]   res_hi_hi_hi_lo_39 = {dataGroup_29_39, dataGroup_28_39};
  wire [31:0]   res_hi_hi_hi_hi_39 = {dataGroup_31_39, dataGroup_30_39};
  wire [63:0]   res_hi_hi_hi_39 = {res_hi_hi_hi_hi_39, res_hi_hi_hi_lo_39};
  wire [127:0]  res_hi_hi_39 = {res_hi_hi_hi_39, res_hi_hi_lo_39};
  wire [255:0]  res_hi_39 = {res_hi_hi_39, res_hi_lo_39};
  wire [511:0]  res_80 = {res_hi_39, res_lo_39};
  wire [2047:0] dataGroup_lo_2432 = {dataGroup_lo_hi_2432, dataGroup_lo_lo_2432};
  wire [2047:0] dataGroup_hi_2432 = {dataGroup_hi_hi_2432, dataGroup_hi_lo_2432};
  wire [15:0]   dataGroup_0_40 = dataGroup_lo_2432[31:16];
  wire [2047:0] dataGroup_lo_2433 = {dataGroup_lo_hi_2433, dataGroup_lo_lo_2433};
  wire [2047:0] dataGroup_hi_2433 = {dataGroup_hi_hi_2433, dataGroup_hi_lo_2433};
  wire [15:0]   dataGroup_1_40 = dataGroup_lo_2433[79:64];
  wire [2047:0] dataGroup_lo_2434 = {dataGroup_lo_hi_2434, dataGroup_lo_lo_2434};
  wire [2047:0] dataGroup_hi_2434 = {dataGroup_hi_hi_2434, dataGroup_hi_lo_2434};
  wire [15:0]   dataGroup_2_40 = dataGroup_lo_2434[127:112];
  wire [2047:0] dataGroup_lo_2435 = {dataGroup_lo_hi_2435, dataGroup_lo_lo_2435};
  wire [2047:0] dataGroup_hi_2435 = {dataGroup_hi_hi_2435, dataGroup_hi_lo_2435};
  wire [15:0]   dataGroup_3_40 = dataGroup_lo_2435[175:160];
  wire [2047:0] dataGroup_lo_2436 = {dataGroup_lo_hi_2436, dataGroup_lo_lo_2436};
  wire [2047:0] dataGroup_hi_2436 = {dataGroup_hi_hi_2436, dataGroup_hi_lo_2436};
  wire [15:0]   dataGroup_4_40 = dataGroup_lo_2436[223:208];
  wire [2047:0] dataGroup_lo_2437 = {dataGroup_lo_hi_2437, dataGroup_lo_lo_2437};
  wire [2047:0] dataGroup_hi_2437 = {dataGroup_hi_hi_2437, dataGroup_hi_lo_2437};
  wire [15:0]   dataGroup_5_40 = dataGroup_lo_2437[271:256];
  wire [2047:0] dataGroup_lo_2438 = {dataGroup_lo_hi_2438, dataGroup_lo_lo_2438};
  wire [2047:0] dataGroup_hi_2438 = {dataGroup_hi_hi_2438, dataGroup_hi_lo_2438};
  wire [15:0]   dataGroup_6_40 = dataGroup_lo_2438[319:304];
  wire [2047:0] dataGroup_lo_2439 = {dataGroup_lo_hi_2439, dataGroup_lo_lo_2439};
  wire [2047:0] dataGroup_hi_2439 = {dataGroup_hi_hi_2439, dataGroup_hi_lo_2439};
  wire [15:0]   dataGroup_7_40 = dataGroup_lo_2439[367:352];
  wire [2047:0] dataGroup_lo_2440 = {dataGroup_lo_hi_2440, dataGroup_lo_lo_2440};
  wire [2047:0] dataGroup_hi_2440 = {dataGroup_hi_hi_2440, dataGroup_hi_lo_2440};
  wire [15:0]   dataGroup_8_40 = dataGroup_lo_2440[415:400];
  wire [2047:0] dataGroup_lo_2441 = {dataGroup_lo_hi_2441, dataGroup_lo_lo_2441};
  wire [2047:0] dataGroup_hi_2441 = {dataGroup_hi_hi_2441, dataGroup_hi_lo_2441};
  wire [15:0]   dataGroup_9_40 = dataGroup_lo_2441[463:448];
  wire [2047:0] dataGroup_lo_2442 = {dataGroup_lo_hi_2442, dataGroup_lo_lo_2442};
  wire [2047:0] dataGroup_hi_2442 = {dataGroup_hi_hi_2442, dataGroup_hi_lo_2442};
  wire [15:0]   dataGroup_10_40 = dataGroup_lo_2442[511:496];
  wire [2047:0] dataGroup_lo_2443 = {dataGroup_lo_hi_2443, dataGroup_lo_lo_2443};
  wire [2047:0] dataGroup_hi_2443 = {dataGroup_hi_hi_2443, dataGroup_hi_lo_2443};
  wire [15:0]   dataGroup_11_40 = dataGroup_lo_2443[559:544];
  wire [2047:0] dataGroup_lo_2444 = {dataGroup_lo_hi_2444, dataGroup_lo_lo_2444};
  wire [2047:0] dataGroup_hi_2444 = {dataGroup_hi_hi_2444, dataGroup_hi_lo_2444};
  wire [15:0]   dataGroup_12_40 = dataGroup_lo_2444[607:592];
  wire [2047:0] dataGroup_lo_2445 = {dataGroup_lo_hi_2445, dataGroup_lo_lo_2445};
  wire [2047:0] dataGroup_hi_2445 = {dataGroup_hi_hi_2445, dataGroup_hi_lo_2445};
  wire [15:0]   dataGroup_13_40 = dataGroup_lo_2445[655:640];
  wire [2047:0] dataGroup_lo_2446 = {dataGroup_lo_hi_2446, dataGroup_lo_lo_2446};
  wire [2047:0] dataGroup_hi_2446 = {dataGroup_hi_hi_2446, dataGroup_hi_lo_2446};
  wire [15:0]   dataGroup_14_40 = dataGroup_lo_2446[703:688];
  wire [2047:0] dataGroup_lo_2447 = {dataGroup_lo_hi_2447, dataGroup_lo_lo_2447};
  wire [2047:0] dataGroup_hi_2447 = {dataGroup_hi_hi_2447, dataGroup_hi_lo_2447};
  wire [15:0]   dataGroup_15_40 = dataGroup_lo_2447[751:736];
  wire [2047:0] dataGroup_lo_2448 = {dataGroup_lo_hi_2448, dataGroup_lo_lo_2448};
  wire [2047:0] dataGroup_hi_2448 = {dataGroup_hi_hi_2448, dataGroup_hi_lo_2448};
  wire [15:0]   dataGroup_16_40 = dataGroup_lo_2448[799:784];
  wire [2047:0] dataGroup_lo_2449 = {dataGroup_lo_hi_2449, dataGroup_lo_lo_2449};
  wire [2047:0] dataGroup_hi_2449 = {dataGroup_hi_hi_2449, dataGroup_hi_lo_2449};
  wire [15:0]   dataGroup_17_40 = dataGroup_lo_2449[847:832];
  wire [2047:0] dataGroup_lo_2450 = {dataGroup_lo_hi_2450, dataGroup_lo_lo_2450};
  wire [2047:0] dataGroup_hi_2450 = {dataGroup_hi_hi_2450, dataGroup_hi_lo_2450};
  wire [15:0]   dataGroup_18_40 = dataGroup_lo_2450[895:880];
  wire [2047:0] dataGroup_lo_2451 = {dataGroup_lo_hi_2451, dataGroup_lo_lo_2451};
  wire [2047:0] dataGroup_hi_2451 = {dataGroup_hi_hi_2451, dataGroup_hi_lo_2451};
  wire [15:0]   dataGroup_19_40 = dataGroup_lo_2451[943:928];
  wire [2047:0] dataGroup_lo_2452 = {dataGroup_lo_hi_2452, dataGroup_lo_lo_2452};
  wire [2047:0] dataGroup_hi_2452 = {dataGroup_hi_hi_2452, dataGroup_hi_lo_2452};
  wire [15:0]   dataGroup_20_40 = dataGroup_lo_2452[991:976];
  wire [2047:0] dataGroup_lo_2453 = {dataGroup_lo_hi_2453, dataGroup_lo_lo_2453};
  wire [2047:0] dataGroup_hi_2453 = {dataGroup_hi_hi_2453, dataGroup_hi_lo_2453};
  wire [15:0]   dataGroup_21_40 = dataGroup_lo_2453[1039:1024];
  wire [2047:0] dataGroup_lo_2454 = {dataGroup_lo_hi_2454, dataGroup_lo_lo_2454};
  wire [2047:0] dataGroup_hi_2454 = {dataGroup_hi_hi_2454, dataGroup_hi_lo_2454};
  wire [15:0]   dataGroup_22_40 = dataGroup_lo_2454[1087:1072];
  wire [2047:0] dataGroup_lo_2455 = {dataGroup_lo_hi_2455, dataGroup_lo_lo_2455};
  wire [2047:0] dataGroup_hi_2455 = {dataGroup_hi_hi_2455, dataGroup_hi_lo_2455};
  wire [15:0]   dataGroup_23_40 = dataGroup_lo_2455[1135:1120];
  wire [2047:0] dataGroup_lo_2456 = {dataGroup_lo_hi_2456, dataGroup_lo_lo_2456};
  wire [2047:0] dataGroup_hi_2456 = {dataGroup_hi_hi_2456, dataGroup_hi_lo_2456};
  wire [15:0]   dataGroup_24_40 = dataGroup_lo_2456[1183:1168];
  wire [2047:0] dataGroup_lo_2457 = {dataGroup_lo_hi_2457, dataGroup_lo_lo_2457};
  wire [2047:0] dataGroup_hi_2457 = {dataGroup_hi_hi_2457, dataGroup_hi_lo_2457};
  wire [15:0]   dataGroup_25_40 = dataGroup_lo_2457[1231:1216];
  wire [2047:0] dataGroup_lo_2458 = {dataGroup_lo_hi_2458, dataGroup_lo_lo_2458};
  wire [2047:0] dataGroup_hi_2458 = {dataGroup_hi_hi_2458, dataGroup_hi_lo_2458};
  wire [15:0]   dataGroup_26_40 = dataGroup_lo_2458[1279:1264];
  wire [2047:0] dataGroup_lo_2459 = {dataGroup_lo_hi_2459, dataGroup_lo_lo_2459};
  wire [2047:0] dataGroup_hi_2459 = {dataGroup_hi_hi_2459, dataGroup_hi_lo_2459};
  wire [15:0]   dataGroup_27_40 = dataGroup_lo_2459[1327:1312];
  wire [2047:0] dataGroup_lo_2460 = {dataGroup_lo_hi_2460, dataGroup_lo_lo_2460};
  wire [2047:0] dataGroup_hi_2460 = {dataGroup_hi_hi_2460, dataGroup_hi_lo_2460};
  wire [15:0]   dataGroup_28_40 = dataGroup_lo_2460[1375:1360];
  wire [2047:0] dataGroup_lo_2461 = {dataGroup_lo_hi_2461, dataGroup_lo_lo_2461};
  wire [2047:0] dataGroup_hi_2461 = {dataGroup_hi_hi_2461, dataGroup_hi_lo_2461};
  wire [15:0]   dataGroup_29_40 = dataGroup_lo_2461[1423:1408];
  wire [2047:0] dataGroup_lo_2462 = {dataGroup_lo_hi_2462, dataGroup_lo_lo_2462};
  wire [2047:0] dataGroup_hi_2462 = {dataGroup_hi_hi_2462, dataGroup_hi_lo_2462};
  wire [15:0]   dataGroup_30_40 = dataGroup_lo_2462[1471:1456];
  wire [2047:0] dataGroup_lo_2463 = {dataGroup_lo_hi_2463, dataGroup_lo_lo_2463};
  wire [2047:0] dataGroup_hi_2463 = {dataGroup_hi_hi_2463, dataGroup_hi_lo_2463};
  wire [15:0]   dataGroup_31_40 = dataGroup_lo_2463[1519:1504];
  wire [31:0]   res_lo_lo_lo_lo_40 = {dataGroup_1_40, dataGroup_0_40};
  wire [31:0]   res_lo_lo_lo_hi_40 = {dataGroup_3_40, dataGroup_2_40};
  wire [63:0]   res_lo_lo_lo_40 = {res_lo_lo_lo_hi_40, res_lo_lo_lo_lo_40};
  wire [31:0]   res_lo_lo_hi_lo_40 = {dataGroup_5_40, dataGroup_4_40};
  wire [31:0]   res_lo_lo_hi_hi_40 = {dataGroup_7_40, dataGroup_6_40};
  wire [63:0]   res_lo_lo_hi_40 = {res_lo_lo_hi_hi_40, res_lo_lo_hi_lo_40};
  wire [127:0]  res_lo_lo_40 = {res_lo_lo_hi_40, res_lo_lo_lo_40};
  wire [31:0]   res_lo_hi_lo_lo_40 = {dataGroup_9_40, dataGroup_8_40};
  wire [31:0]   res_lo_hi_lo_hi_40 = {dataGroup_11_40, dataGroup_10_40};
  wire [63:0]   res_lo_hi_lo_40 = {res_lo_hi_lo_hi_40, res_lo_hi_lo_lo_40};
  wire [31:0]   res_lo_hi_hi_lo_40 = {dataGroup_13_40, dataGroup_12_40};
  wire [31:0]   res_lo_hi_hi_hi_40 = {dataGroup_15_40, dataGroup_14_40};
  wire [63:0]   res_lo_hi_hi_40 = {res_lo_hi_hi_hi_40, res_lo_hi_hi_lo_40};
  wire [127:0]  res_lo_hi_40 = {res_lo_hi_hi_40, res_lo_hi_lo_40};
  wire [255:0]  res_lo_40 = {res_lo_hi_40, res_lo_lo_40};
  wire [31:0]   res_hi_lo_lo_lo_40 = {dataGroup_17_40, dataGroup_16_40};
  wire [31:0]   res_hi_lo_lo_hi_40 = {dataGroup_19_40, dataGroup_18_40};
  wire [63:0]   res_hi_lo_lo_40 = {res_hi_lo_lo_hi_40, res_hi_lo_lo_lo_40};
  wire [31:0]   res_hi_lo_hi_lo_40 = {dataGroup_21_40, dataGroup_20_40};
  wire [31:0]   res_hi_lo_hi_hi_40 = {dataGroup_23_40, dataGroup_22_40};
  wire [63:0]   res_hi_lo_hi_40 = {res_hi_lo_hi_hi_40, res_hi_lo_hi_lo_40};
  wire [127:0]  res_hi_lo_40 = {res_hi_lo_hi_40, res_hi_lo_lo_40};
  wire [31:0]   res_hi_hi_lo_lo_40 = {dataGroup_25_40, dataGroup_24_40};
  wire [31:0]   res_hi_hi_lo_hi_40 = {dataGroup_27_40, dataGroup_26_40};
  wire [63:0]   res_hi_hi_lo_40 = {res_hi_hi_lo_hi_40, res_hi_hi_lo_lo_40};
  wire [31:0]   res_hi_hi_hi_lo_40 = {dataGroup_29_40, dataGroup_28_40};
  wire [31:0]   res_hi_hi_hi_hi_40 = {dataGroup_31_40, dataGroup_30_40};
  wire [63:0]   res_hi_hi_hi_40 = {res_hi_hi_hi_hi_40, res_hi_hi_hi_lo_40};
  wire [127:0]  res_hi_hi_40 = {res_hi_hi_hi_40, res_hi_hi_lo_40};
  wire [255:0]  res_hi_40 = {res_hi_hi_40, res_hi_lo_40};
  wire [511:0]  res_81 = {res_hi_40, res_lo_40};
  wire [2047:0] dataGroup_lo_2464 = {dataGroup_lo_hi_2464, dataGroup_lo_lo_2464};
  wire [2047:0] dataGroup_hi_2464 = {dataGroup_hi_hi_2464, dataGroup_hi_lo_2464};
  wire [15:0]   dataGroup_0_41 = dataGroup_lo_2464[47:32];
  wire [2047:0] dataGroup_lo_2465 = {dataGroup_lo_hi_2465, dataGroup_lo_lo_2465};
  wire [2047:0] dataGroup_hi_2465 = {dataGroup_hi_hi_2465, dataGroup_hi_lo_2465};
  wire [15:0]   dataGroup_1_41 = dataGroup_lo_2465[95:80];
  wire [2047:0] dataGroup_lo_2466 = {dataGroup_lo_hi_2466, dataGroup_lo_lo_2466};
  wire [2047:0] dataGroup_hi_2466 = {dataGroup_hi_hi_2466, dataGroup_hi_lo_2466};
  wire [15:0]   dataGroup_2_41 = dataGroup_lo_2466[143:128];
  wire [2047:0] dataGroup_lo_2467 = {dataGroup_lo_hi_2467, dataGroup_lo_lo_2467};
  wire [2047:0] dataGroup_hi_2467 = {dataGroup_hi_hi_2467, dataGroup_hi_lo_2467};
  wire [15:0]   dataGroup_3_41 = dataGroup_lo_2467[191:176];
  wire [2047:0] dataGroup_lo_2468 = {dataGroup_lo_hi_2468, dataGroup_lo_lo_2468};
  wire [2047:0] dataGroup_hi_2468 = {dataGroup_hi_hi_2468, dataGroup_hi_lo_2468};
  wire [15:0]   dataGroup_4_41 = dataGroup_lo_2468[239:224];
  wire [2047:0] dataGroup_lo_2469 = {dataGroup_lo_hi_2469, dataGroup_lo_lo_2469};
  wire [2047:0] dataGroup_hi_2469 = {dataGroup_hi_hi_2469, dataGroup_hi_lo_2469};
  wire [15:0]   dataGroup_5_41 = dataGroup_lo_2469[287:272];
  wire [2047:0] dataGroup_lo_2470 = {dataGroup_lo_hi_2470, dataGroup_lo_lo_2470};
  wire [2047:0] dataGroup_hi_2470 = {dataGroup_hi_hi_2470, dataGroup_hi_lo_2470};
  wire [15:0]   dataGroup_6_41 = dataGroup_lo_2470[335:320];
  wire [2047:0] dataGroup_lo_2471 = {dataGroup_lo_hi_2471, dataGroup_lo_lo_2471};
  wire [2047:0] dataGroup_hi_2471 = {dataGroup_hi_hi_2471, dataGroup_hi_lo_2471};
  wire [15:0]   dataGroup_7_41 = dataGroup_lo_2471[383:368];
  wire [2047:0] dataGroup_lo_2472 = {dataGroup_lo_hi_2472, dataGroup_lo_lo_2472};
  wire [2047:0] dataGroup_hi_2472 = {dataGroup_hi_hi_2472, dataGroup_hi_lo_2472};
  wire [15:0]   dataGroup_8_41 = dataGroup_lo_2472[431:416];
  wire [2047:0] dataGroup_lo_2473 = {dataGroup_lo_hi_2473, dataGroup_lo_lo_2473};
  wire [2047:0] dataGroup_hi_2473 = {dataGroup_hi_hi_2473, dataGroup_hi_lo_2473};
  wire [15:0]   dataGroup_9_41 = dataGroup_lo_2473[479:464];
  wire [2047:0] dataGroup_lo_2474 = {dataGroup_lo_hi_2474, dataGroup_lo_lo_2474};
  wire [2047:0] dataGroup_hi_2474 = {dataGroup_hi_hi_2474, dataGroup_hi_lo_2474};
  wire [15:0]   dataGroup_10_41 = dataGroup_lo_2474[527:512];
  wire [2047:0] dataGroup_lo_2475 = {dataGroup_lo_hi_2475, dataGroup_lo_lo_2475};
  wire [2047:0] dataGroup_hi_2475 = {dataGroup_hi_hi_2475, dataGroup_hi_lo_2475};
  wire [15:0]   dataGroup_11_41 = dataGroup_lo_2475[575:560];
  wire [2047:0] dataGroup_lo_2476 = {dataGroup_lo_hi_2476, dataGroup_lo_lo_2476};
  wire [2047:0] dataGroup_hi_2476 = {dataGroup_hi_hi_2476, dataGroup_hi_lo_2476};
  wire [15:0]   dataGroup_12_41 = dataGroup_lo_2476[623:608];
  wire [2047:0] dataGroup_lo_2477 = {dataGroup_lo_hi_2477, dataGroup_lo_lo_2477};
  wire [2047:0] dataGroup_hi_2477 = {dataGroup_hi_hi_2477, dataGroup_hi_lo_2477};
  wire [15:0]   dataGroup_13_41 = dataGroup_lo_2477[671:656];
  wire [2047:0] dataGroup_lo_2478 = {dataGroup_lo_hi_2478, dataGroup_lo_lo_2478};
  wire [2047:0] dataGroup_hi_2478 = {dataGroup_hi_hi_2478, dataGroup_hi_lo_2478};
  wire [15:0]   dataGroup_14_41 = dataGroup_lo_2478[719:704];
  wire [2047:0] dataGroup_lo_2479 = {dataGroup_lo_hi_2479, dataGroup_lo_lo_2479};
  wire [2047:0] dataGroup_hi_2479 = {dataGroup_hi_hi_2479, dataGroup_hi_lo_2479};
  wire [15:0]   dataGroup_15_41 = dataGroup_lo_2479[767:752];
  wire [2047:0] dataGroup_lo_2480 = {dataGroup_lo_hi_2480, dataGroup_lo_lo_2480};
  wire [2047:0] dataGroup_hi_2480 = {dataGroup_hi_hi_2480, dataGroup_hi_lo_2480};
  wire [15:0]   dataGroup_16_41 = dataGroup_lo_2480[815:800];
  wire [2047:0] dataGroup_lo_2481 = {dataGroup_lo_hi_2481, dataGroup_lo_lo_2481};
  wire [2047:0] dataGroup_hi_2481 = {dataGroup_hi_hi_2481, dataGroup_hi_lo_2481};
  wire [15:0]   dataGroup_17_41 = dataGroup_lo_2481[863:848];
  wire [2047:0] dataGroup_lo_2482 = {dataGroup_lo_hi_2482, dataGroup_lo_lo_2482};
  wire [2047:0] dataGroup_hi_2482 = {dataGroup_hi_hi_2482, dataGroup_hi_lo_2482};
  wire [15:0]   dataGroup_18_41 = dataGroup_lo_2482[911:896];
  wire [2047:0] dataGroup_lo_2483 = {dataGroup_lo_hi_2483, dataGroup_lo_lo_2483};
  wire [2047:0] dataGroup_hi_2483 = {dataGroup_hi_hi_2483, dataGroup_hi_lo_2483};
  wire [15:0]   dataGroup_19_41 = dataGroup_lo_2483[959:944];
  wire [2047:0] dataGroup_lo_2484 = {dataGroup_lo_hi_2484, dataGroup_lo_lo_2484};
  wire [2047:0] dataGroup_hi_2484 = {dataGroup_hi_hi_2484, dataGroup_hi_lo_2484};
  wire [15:0]   dataGroup_20_41 = dataGroup_lo_2484[1007:992];
  wire [2047:0] dataGroup_lo_2485 = {dataGroup_lo_hi_2485, dataGroup_lo_lo_2485};
  wire [2047:0] dataGroup_hi_2485 = {dataGroup_hi_hi_2485, dataGroup_hi_lo_2485};
  wire [15:0]   dataGroup_21_41 = dataGroup_lo_2485[1055:1040];
  wire [2047:0] dataGroup_lo_2486 = {dataGroup_lo_hi_2486, dataGroup_lo_lo_2486};
  wire [2047:0] dataGroup_hi_2486 = {dataGroup_hi_hi_2486, dataGroup_hi_lo_2486};
  wire [15:0]   dataGroup_22_41 = dataGroup_lo_2486[1103:1088];
  wire [2047:0] dataGroup_lo_2487 = {dataGroup_lo_hi_2487, dataGroup_lo_lo_2487};
  wire [2047:0] dataGroup_hi_2487 = {dataGroup_hi_hi_2487, dataGroup_hi_lo_2487};
  wire [15:0]   dataGroup_23_41 = dataGroup_lo_2487[1151:1136];
  wire [2047:0] dataGroup_lo_2488 = {dataGroup_lo_hi_2488, dataGroup_lo_lo_2488};
  wire [2047:0] dataGroup_hi_2488 = {dataGroup_hi_hi_2488, dataGroup_hi_lo_2488};
  wire [15:0]   dataGroup_24_41 = dataGroup_lo_2488[1199:1184];
  wire [2047:0] dataGroup_lo_2489 = {dataGroup_lo_hi_2489, dataGroup_lo_lo_2489};
  wire [2047:0] dataGroup_hi_2489 = {dataGroup_hi_hi_2489, dataGroup_hi_lo_2489};
  wire [15:0]   dataGroup_25_41 = dataGroup_lo_2489[1247:1232];
  wire [2047:0] dataGroup_lo_2490 = {dataGroup_lo_hi_2490, dataGroup_lo_lo_2490};
  wire [2047:0] dataGroup_hi_2490 = {dataGroup_hi_hi_2490, dataGroup_hi_lo_2490};
  wire [15:0]   dataGroup_26_41 = dataGroup_lo_2490[1295:1280];
  wire [2047:0] dataGroup_lo_2491 = {dataGroup_lo_hi_2491, dataGroup_lo_lo_2491};
  wire [2047:0] dataGroup_hi_2491 = {dataGroup_hi_hi_2491, dataGroup_hi_lo_2491};
  wire [15:0]   dataGroup_27_41 = dataGroup_lo_2491[1343:1328];
  wire [2047:0] dataGroup_lo_2492 = {dataGroup_lo_hi_2492, dataGroup_lo_lo_2492};
  wire [2047:0] dataGroup_hi_2492 = {dataGroup_hi_hi_2492, dataGroup_hi_lo_2492};
  wire [15:0]   dataGroup_28_41 = dataGroup_lo_2492[1391:1376];
  wire [2047:0] dataGroup_lo_2493 = {dataGroup_lo_hi_2493, dataGroup_lo_lo_2493};
  wire [2047:0] dataGroup_hi_2493 = {dataGroup_hi_hi_2493, dataGroup_hi_lo_2493};
  wire [15:0]   dataGroup_29_41 = dataGroup_lo_2493[1439:1424];
  wire [2047:0] dataGroup_lo_2494 = {dataGroup_lo_hi_2494, dataGroup_lo_lo_2494};
  wire [2047:0] dataGroup_hi_2494 = {dataGroup_hi_hi_2494, dataGroup_hi_lo_2494};
  wire [15:0]   dataGroup_30_41 = dataGroup_lo_2494[1487:1472];
  wire [2047:0] dataGroup_lo_2495 = {dataGroup_lo_hi_2495, dataGroup_lo_lo_2495};
  wire [2047:0] dataGroup_hi_2495 = {dataGroup_hi_hi_2495, dataGroup_hi_lo_2495};
  wire [15:0]   dataGroup_31_41 = dataGroup_lo_2495[1535:1520];
  wire [31:0]   res_lo_lo_lo_lo_41 = {dataGroup_1_41, dataGroup_0_41};
  wire [31:0]   res_lo_lo_lo_hi_41 = {dataGroup_3_41, dataGroup_2_41};
  wire [63:0]   res_lo_lo_lo_41 = {res_lo_lo_lo_hi_41, res_lo_lo_lo_lo_41};
  wire [31:0]   res_lo_lo_hi_lo_41 = {dataGroup_5_41, dataGroup_4_41};
  wire [31:0]   res_lo_lo_hi_hi_41 = {dataGroup_7_41, dataGroup_6_41};
  wire [63:0]   res_lo_lo_hi_41 = {res_lo_lo_hi_hi_41, res_lo_lo_hi_lo_41};
  wire [127:0]  res_lo_lo_41 = {res_lo_lo_hi_41, res_lo_lo_lo_41};
  wire [31:0]   res_lo_hi_lo_lo_41 = {dataGroup_9_41, dataGroup_8_41};
  wire [31:0]   res_lo_hi_lo_hi_41 = {dataGroup_11_41, dataGroup_10_41};
  wire [63:0]   res_lo_hi_lo_41 = {res_lo_hi_lo_hi_41, res_lo_hi_lo_lo_41};
  wire [31:0]   res_lo_hi_hi_lo_41 = {dataGroup_13_41, dataGroup_12_41};
  wire [31:0]   res_lo_hi_hi_hi_41 = {dataGroup_15_41, dataGroup_14_41};
  wire [63:0]   res_lo_hi_hi_41 = {res_lo_hi_hi_hi_41, res_lo_hi_hi_lo_41};
  wire [127:0]  res_lo_hi_41 = {res_lo_hi_hi_41, res_lo_hi_lo_41};
  wire [255:0]  res_lo_41 = {res_lo_hi_41, res_lo_lo_41};
  wire [31:0]   res_hi_lo_lo_lo_41 = {dataGroup_17_41, dataGroup_16_41};
  wire [31:0]   res_hi_lo_lo_hi_41 = {dataGroup_19_41, dataGroup_18_41};
  wire [63:0]   res_hi_lo_lo_41 = {res_hi_lo_lo_hi_41, res_hi_lo_lo_lo_41};
  wire [31:0]   res_hi_lo_hi_lo_41 = {dataGroup_21_41, dataGroup_20_41};
  wire [31:0]   res_hi_lo_hi_hi_41 = {dataGroup_23_41, dataGroup_22_41};
  wire [63:0]   res_hi_lo_hi_41 = {res_hi_lo_hi_hi_41, res_hi_lo_hi_lo_41};
  wire [127:0]  res_hi_lo_41 = {res_hi_lo_hi_41, res_hi_lo_lo_41};
  wire [31:0]   res_hi_hi_lo_lo_41 = {dataGroup_25_41, dataGroup_24_41};
  wire [31:0]   res_hi_hi_lo_hi_41 = {dataGroup_27_41, dataGroup_26_41};
  wire [63:0]   res_hi_hi_lo_41 = {res_hi_hi_lo_hi_41, res_hi_hi_lo_lo_41};
  wire [31:0]   res_hi_hi_hi_lo_41 = {dataGroup_29_41, dataGroup_28_41};
  wire [31:0]   res_hi_hi_hi_hi_41 = {dataGroup_31_41, dataGroup_30_41};
  wire [63:0]   res_hi_hi_hi_41 = {res_hi_hi_hi_hi_41, res_hi_hi_hi_lo_41};
  wire [127:0]  res_hi_hi_41 = {res_hi_hi_hi_41, res_hi_hi_lo_41};
  wire [255:0]  res_hi_41 = {res_hi_hi_41, res_hi_lo_41};
  wire [511:0]  res_82 = {res_hi_41, res_lo_41};
  wire [1023:0] lo_lo_10 = {res_81, res_80};
  wire [1023:0] lo_hi_10 = {512'h0, res_82};
  wire [2047:0] lo_10 = {lo_hi_10, lo_lo_10};
  wire [4095:0] regroupLoadData_1_2 = {2048'h0, lo_10};
  wire [2047:0] dataGroup_lo_2496 = {dataGroup_lo_hi_2496, dataGroup_lo_lo_2496};
  wire [2047:0] dataGroup_hi_2496 = {dataGroup_hi_hi_2496, dataGroup_hi_lo_2496};
  wire [15:0]   dataGroup_0_42 = dataGroup_lo_2496[15:0];
  wire [2047:0] dataGroup_lo_2497 = {dataGroup_lo_hi_2497, dataGroup_lo_lo_2497};
  wire [2047:0] dataGroup_hi_2497 = {dataGroup_hi_hi_2497, dataGroup_hi_lo_2497};
  wire [15:0]   dataGroup_1_42 = dataGroup_lo_2497[79:64];
  wire [2047:0] dataGroup_lo_2498 = {dataGroup_lo_hi_2498, dataGroup_lo_lo_2498};
  wire [2047:0] dataGroup_hi_2498 = {dataGroup_hi_hi_2498, dataGroup_hi_lo_2498};
  wire [15:0]   dataGroup_2_42 = dataGroup_lo_2498[143:128];
  wire [2047:0] dataGroup_lo_2499 = {dataGroup_lo_hi_2499, dataGroup_lo_lo_2499};
  wire [2047:0] dataGroup_hi_2499 = {dataGroup_hi_hi_2499, dataGroup_hi_lo_2499};
  wire [15:0]   dataGroup_3_42 = dataGroup_lo_2499[207:192];
  wire [2047:0] dataGroup_lo_2500 = {dataGroup_lo_hi_2500, dataGroup_lo_lo_2500};
  wire [2047:0] dataGroup_hi_2500 = {dataGroup_hi_hi_2500, dataGroup_hi_lo_2500};
  wire [15:0]   dataGroup_4_42 = dataGroup_lo_2500[271:256];
  wire [2047:0] dataGroup_lo_2501 = {dataGroup_lo_hi_2501, dataGroup_lo_lo_2501};
  wire [2047:0] dataGroup_hi_2501 = {dataGroup_hi_hi_2501, dataGroup_hi_lo_2501};
  wire [15:0]   dataGroup_5_42 = dataGroup_lo_2501[335:320];
  wire [2047:0] dataGroup_lo_2502 = {dataGroup_lo_hi_2502, dataGroup_lo_lo_2502};
  wire [2047:0] dataGroup_hi_2502 = {dataGroup_hi_hi_2502, dataGroup_hi_lo_2502};
  wire [15:0]   dataGroup_6_42 = dataGroup_lo_2502[399:384];
  wire [2047:0] dataGroup_lo_2503 = {dataGroup_lo_hi_2503, dataGroup_lo_lo_2503};
  wire [2047:0] dataGroup_hi_2503 = {dataGroup_hi_hi_2503, dataGroup_hi_lo_2503};
  wire [15:0]   dataGroup_7_42 = dataGroup_lo_2503[463:448];
  wire [2047:0] dataGroup_lo_2504 = {dataGroup_lo_hi_2504, dataGroup_lo_lo_2504};
  wire [2047:0] dataGroup_hi_2504 = {dataGroup_hi_hi_2504, dataGroup_hi_lo_2504};
  wire [15:0]   dataGroup_8_42 = dataGroup_lo_2504[527:512];
  wire [2047:0] dataGroup_lo_2505 = {dataGroup_lo_hi_2505, dataGroup_lo_lo_2505};
  wire [2047:0] dataGroup_hi_2505 = {dataGroup_hi_hi_2505, dataGroup_hi_lo_2505};
  wire [15:0]   dataGroup_9_42 = dataGroup_lo_2505[591:576];
  wire [2047:0] dataGroup_lo_2506 = {dataGroup_lo_hi_2506, dataGroup_lo_lo_2506};
  wire [2047:0] dataGroup_hi_2506 = {dataGroup_hi_hi_2506, dataGroup_hi_lo_2506};
  wire [15:0]   dataGroup_10_42 = dataGroup_lo_2506[655:640];
  wire [2047:0] dataGroup_lo_2507 = {dataGroup_lo_hi_2507, dataGroup_lo_lo_2507};
  wire [2047:0] dataGroup_hi_2507 = {dataGroup_hi_hi_2507, dataGroup_hi_lo_2507};
  wire [15:0]   dataGroup_11_42 = dataGroup_lo_2507[719:704];
  wire [2047:0] dataGroup_lo_2508 = {dataGroup_lo_hi_2508, dataGroup_lo_lo_2508};
  wire [2047:0] dataGroup_hi_2508 = {dataGroup_hi_hi_2508, dataGroup_hi_lo_2508};
  wire [15:0]   dataGroup_12_42 = dataGroup_lo_2508[783:768];
  wire [2047:0] dataGroup_lo_2509 = {dataGroup_lo_hi_2509, dataGroup_lo_lo_2509};
  wire [2047:0] dataGroup_hi_2509 = {dataGroup_hi_hi_2509, dataGroup_hi_lo_2509};
  wire [15:0]   dataGroup_13_42 = dataGroup_lo_2509[847:832];
  wire [2047:0] dataGroup_lo_2510 = {dataGroup_lo_hi_2510, dataGroup_lo_lo_2510};
  wire [2047:0] dataGroup_hi_2510 = {dataGroup_hi_hi_2510, dataGroup_hi_lo_2510};
  wire [15:0]   dataGroup_14_42 = dataGroup_lo_2510[911:896];
  wire [2047:0] dataGroup_lo_2511 = {dataGroup_lo_hi_2511, dataGroup_lo_lo_2511};
  wire [2047:0] dataGroup_hi_2511 = {dataGroup_hi_hi_2511, dataGroup_hi_lo_2511};
  wire [15:0]   dataGroup_15_42 = dataGroup_lo_2511[975:960];
  wire [2047:0] dataGroup_lo_2512 = {dataGroup_lo_hi_2512, dataGroup_lo_lo_2512};
  wire [2047:0] dataGroup_hi_2512 = {dataGroup_hi_hi_2512, dataGroup_hi_lo_2512};
  wire [15:0]   dataGroup_16_42 = dataGroup_lo_2512[1039:1024];
  wire [2047:0] dataGroup_lo_2513 = {dataGroup_lo_hi_2513, dataGroup_lo_lo_2513};
  wire [2047:0] dataGroup_hi_2513 = {dataGroup_hi_hi_2513, dataGroup_hi_lo_2513};
  wire [15:0]   dataGroup_17_42 = dataGroup_lo_2513[1103:1088];
  wire [2047:0] dataGroup_lo_2514 = {dataGroup_lo_hi_2514, dataGroup_lo_lo_2514};
  wire [2047:0] dataGroup_hi_2514 = {dataGroup_hi_hi_2514, dataGroup_hi_lo_2514};
  wire [15:0]   dataGroup_18_42 = dataGroup_lo_2514[1167:1152];
  wire [2047:0] dataGroup_lo_2515 = {dataGroup_lo_hi_2515, dataGroup_lo_lo_2515};
  wire [2047:0] dataGroup_hi_2515 = {dataGroup_hi_hi_2515, dataGroup_hi_lo_2515};
  wire [15:0]   dataGroup_19_42 = dataGroup_lo_2515[1231:1216];
  wire [2047:0] dataGroup_lo_2516 = {dataGroup_lo_hi_2516, dataGroup_lo_lo_2516};
  wire [2047:0] dataGroup_hi_2516 = {dataGroup_hi_hi_2516, dataGroup_hi_lo_2516};
  wire [15:0]   dataGroup_20_42 = dataGroup_lo_2516[1295:1280];
  wire [2047:0] dataGroup_lo_2517 = {dataGroup_lo_hi_2517, dataGroup_lo_lo_2517};
  wire [2047:0] dataGroup_hi_2517 = {dataGroup_hi_hi_2517, dataGroup_hi_lo_2517};
  wire [15:0]   dataGroup_21_42 = dataGroup_lo_2517[1359:1344];
  wire [2047:0] dataGroup_lo_2518 = {dataGroup_lo_hi_2518, dataGroup_lo_lo_2518};
  wire [2047:0] dataGroup_hi_2518 = {dataGroup_hi_hi_2518, dataGroup_hi_lo_2518};
  wire [15:0]   dataGroup_22_42 = dataGroup_lo_2518[1423:1408];
  wire [2047:0] dataGroup_lo_2519 = {dataGroup_lo_hi_2519, dataGroup_lo_lo_2519};
  wire [2047:0] dataGroup_hi_2519 = {dataGroup_hi_hi_2519, dataGroup_hi_lo_2519};
  wire [15:0]   dataGroup_23_42 = dataGroup_lo_2519[1487:1472];
  wire [2047:0] dataGroup_lo_2520 = {dataGroup_lo_hi_2520, dataGroup_lo_lo_2520};
  wire [2047:0] dataGroup_hi_2520 = {dataGroup_hi_hi_2520, dataGroup_hi_lo_2520};
  wire [15:0]   dataGroup_24_42 = dataGroup_lo_2520[1551:1536];
  wire [2047:0] dataGroup_lo_2521 = {dataGroup_lo_hi_2521, dataGroup_lo_lo_2521};
  wire [2047:0] dataGroup_hi_2521 = {dataGroup_hi_hi_2521, dataGroup_hi_lo_2521};
  wire [15:0]   dataGroup_25_42 = dataGroup_lo_2521[1615:1600];
  wire [2047:0] dataGroup_lo_2522 = {dataGroup_lo_hi_2522, dataGroup_lo_lo_2522};
  wire [2047:0] dataGroup_hi_2522 = {dataGroup_hi_hi_2522, dataGroup_hi_lo_2522};
  wire [15:0]   dataGroup_26_42 = dataGroup_lo_2522[1679:1664];
  wire [2047:0] dataGroup_lo_2523 = {dataGroup_lo_hi_2523, dataGroup_lo_lo_2523};
  wire [2047:0] dataGroup_hi_2523 = {dataGroup_hi_hi_2523, dataGroup_hi_lo_2523};
  wire [15:0]   dataGroup_27_42 = dataGroup_lo_2523[1743:1728];
  wire [2047:0] dataGroup_lo_2524 = {dataGroup_lo_hi_2524, dataGroup_lo_lo_2524};
  wire [2047:0] dataGroup_hi_2524 = {dataGroup_hi_hi_2524, dataGroup_hi_lo_2524};
  wire [15:0]   dataGroup_28_42 = dataGroup_lo_2524[1807:1792];
  wire [2047:0] dataGroup_lo_2525 = {dataGroup_lo_hi_2525, dataGroup_lo_lo_2525};
  wire [2047:0] dataGroup_hi_2525 = {dataGroup_hi_hi_2525, dataGroup_hi_lo_2525};
  wire [15:0]   dataGroup_29_42 = dataGroup_lo_2525[1871:1856];
  wire [2047:0] dataGroup_lo_2526 = {dataGroup_lo_hi_2526, dataGroup_lo_lo_2526};
  wire [2047:0] dataGroup_hi_2526 = {dataGroup_hi_hi_2526, dataGroup_hi_lo_2526};
  wire [15:0]   dataGroup_30_42 = dataGroup_lo_2526[1935:1920];
  wire [2047:0] dataGroup_lo_2527 = {dataGroup_lo_hi_2527, dataGroup_lo_lo_2527};
  wire [2047:0] dataGroup_hi_2527 = {dataGroup_hi_hi_2527, dataGroup_hi_lo_2527};
  wire [15:0]   dataGroup_31_42 = dataGroup_lo_2527[1999:1984];
  wire [31:0]   res_lo_lo_lo_lo_42 = {dataGroup_1_42, dataGroup_0_42};
  wire [31:0]   res_lo_lo_lo_hi_42 = {dataGroup_3_42, dataGroup_2_42};
  wire [63:0]   res_lo_lo_lo_42 = {res_lo_lo_lo_hi_42, res_lo_lo_lo_lo_42};
  wire [31:0]   res_lo_lo_hi_lo_42 = {dataGroup_5_42, dataGroup_4_42};
  wire [31:0]   res_lo_lo_hi_hi_42 = {dataGroup_7_42, dataGroup_6_42};
  wire [63:0]   res_lo_lo_hi_42 = {res_lo_lo_hi_hi_42, res_lo_lo_hi_lo_42};
  wire [127:0]  res_lo_lo_42 = {res_lo_lo_hi_42, res_lo_lo_lo_42};
  wire [31:0]   res_lo_hi_lo_lo_42 = {dataGroup_9_42, dataGroup_8_42};
  wire [31:0]   res_lo_hi_lo_hi_42 = {dataGroup_11_42, dataGroup_10_42};
  wire [63:0]   res_lo_hi_lo_42 = {res_lo_hi_lo_hi_42, res_lo_hi_lo_lo_42};
  wire [31:0]   res_lo_hi_hi_lo_42 = {dataGroup_13_42, dataGroup_12_42};
  wire [31:0]   res_lo_hi_hi_hi_42 = {dataGroup_15_42, dataGroup_14_42};
  wire [63:0]   res_lo_hi_hi_42 = {res_lo_hi_hi_hi_42, res_lo_hi_hi_lo_42};
  wire [127:0]  res_lo_hi_42 = {res_lo_hi_hi_42, res_lo_hi_lo_42};
  wire [255:0]  res_lo_42 = {res_lo_hi_42, res_lo_lo_42};
  wire [31:0]   res_hi_lo_lo_lo_42 = {dataGroup_17_42, dataGroup_16_42};
  wire [31:0]   res_hi_lo_lo_hi_42 = {dataGroup_19_42, dataGroup_18_42};
  wire [63:0]   res_hi_lo_lo_42 = {res_hi_lo_lo_hi_42, res_hi_lo_lo_lo_42};
  wire [31:0]   res_hi_lo_hi_lo_42 = {dataGroup_21_42, dataGroup_20_42};
  wire [31:0]   res_hi_lo_hi_hi_42 = {dataGroup_23_42, dataGroup_22_42};
  wire [63:0]   res_hi_lo_hi_42 = {res_hi_lo_hi_hi_42, res_hi_lo_hi_lo_42};
  wire [127:0]  res_hi_lo_42 = {res_hi_lo_hi_42, res_hi_lo_lo_42};
  wire [31:0]   res_hi_hi_lo_lo_42 = {dataGroup_25_42, dataGroup_24_42};
  wire [31:0]   res_hi_hi_lo_hi_42 = {dataGroup_27_42, dataGroup_26_42};
  wire [63:0]   res_hi_hi_lo_42 = {res_hi_hi_lo_hi_42, res_hi_hi_lo_lo_42};
  wire [31:0]   res_hi_hi_hi_lo_42 = {dataGroup_29_42, dataGroup_28_42};
  wire [31:0]   res_hi_hi_hi_hi_42 = {dataGroup_31_42, dataGroup_30_42};
  wire [63:0]   res_hi_hi_hi_42 = {res_hi_hi_hi_hi_42, res_hi_hi_hi_lo_42};
  wire [127:0]  res_hi_hi_42 = {res_hi_hi_hi_42, res_hi_hi_lo_42};
  wire [255:0]  res_hi_42 = {res_hi_hi_42, res_hi_lo_42};
  wire [511:0]  res_88 = {res_hi_42, res_lo_42};
  wire [2047:0] dataGroup_lo_2528 = {dataGroup_lo_hi_2528, dataGroup_lo_lo_2528};
  wire [2047:0] dataGroup_hi_2528 = {dataGroup_hi_hi_2528, dataGroup_hi_lo_2528};
  wire [15:0]   dataGroup_0_43 = dataGroup_lo_2528[31:16];
  wire [2047:0] dataGroup_lo_2529 = {dataGroup_lo_hi_2529, dataGroup_lo_lo_2529};
  wire [2047:0] dataGroup_hi_2529 = {dataGroup_hi_hi_2529, dataGroup_hi_lo_2529};
  wire [15:0]   dataGroup_1_43 = dataGroup_lo_2529[95:80];
  wire [2047:0] dataGroup_lo_2530 = {dataGroup_lo_hi_2530, dataGroup_lo_lo_2530};
  wire [2047:0] dataGroup_hi_2530 = {dataGroup_hi_hi_2530, dataGroup_hi_lo_2530};
  wire [15:0]   dataGroup_2_43 = dataGroup_lo_2530[159:144];
  wire [2047:0] dataGroup_lo_2531 = {dataGroup_lo_hi_2531, dataGroup_lo_lo_2531};
  wire [2047:0] dataGroup_hi_2531 = {dataGroup_hi_hi_2531, dataGroup_hi_lo_2531};
  wire [15:0]   dataGroup_3_43 = dataGroup_lo_2531[223:208];
  wire [2047:0] dataGroup_lo_2532 = {dataGroup_lo_hi_2532, dataGroup_lo_lo_2532};
  wire [2047:0] dataGroup_hi_2532 = {dataGroup_hi_hi_2532, dataGroup_hi_lo_2532};
  wire [15:0]   dataGroup_4_43 = dataGroup_lo_2532[287:272];
  wire [2047:0] dataGroup_lo_2533 = {dataGroup_lo_hi_2533, dataGroup_lo_lo_2533};
  wire [2047:0] dataGroup_hi_2533 = {dataGroup_hi_hi_2533, dataGroup_hi_lo_2533};
  wire [15:0]   dataGroup_5_43 = dataGroup_lo_2533[351:336];
  wire [2047:0] dataGroup_lo_2534 = {dataGroup_lo_hi_2534, dataGroup_lo_lo_2534};
  wire [2047:0] dataGroup_hi_2534 = {dataGroup_hi_hi_2534, dataGroup_hi_lo_2534};
  wire [15:0]   dataGroup_6_43 = dataGroup_lo_2534[415:400];
  wire [2047:0] dataGroup_lo_2535 = {dataGroup_lo_hi_2535, dataGroup_lo_lo_2535};
  wire [2047:0] dataGroup_hi_2535 = {dataGroup_hi_hi_2535, dataGroup_hi_lo_2535};
  wire [15:0]   dataGroup_7_43 = dataGroup_lo_2535[479:464];
  wire [2047:0] dataGroup_lo_2536 = {dataGroup_lo_hi_2536, dataGroup_lo_lo_2536};
  wire [2047:0] dataGroup_hi_2536 = {dataGroup_hi_hi_2536, dataGroup_hi_lo_2536};
  wire [15:0]   dataGroup_8_43 = dataGroup_lo_2536[543:528];
  wire [2047:0] dataGroup_lo_2537 = {dataGroup_lo_hi_2537, dataGroup_lo_lo_2537};
  wire [2047:0] dataGroup_hi_2537 = {dataGroup_hi_hi_2537, dataGroup_hi_lo_2537};
  wire [15:0]   dataGroup_9_43 = dataGroup_lo_2537[607:592];
  wire [2047:0] dataGroup_lo_2538 = {dataGroup_lo_hi_2538, dataGroup_lo_lo_2538};
  wire [2047:0] dataGroup_hi_2538 = {dataGroup_hi_hi_2538, dataGroup_hi_lo_2538};
  wire [15:0]   dataGroup_10_43 = dataGroup_lo_2538[671:656];
  wire [2047:0] dataGroup_lo_2539 = {dataGroup_lo_hi_2539, dataGroup_lo_lo_2539};
  wire [2047:0] dataGroup_hi_2539 = {dataGroup_hi_hi_2539, dataGroup_hi_lo_2539};
  wire [15:0]   dataGroup_11_43 = dataGroup_lo_2539[735:720];
  wire [2047:0] dataGroup_lo_2540 = {dataGroup_lo_hi_2540, dataGroup_lo_lo_2540};
  wire [2047:0] dataGroup_hi_2540 = {dataGroup_hi_hi_2540, dataGroup_hi_lo_2540};
  wire [15:0]   dataGroup_12_43 = dataGroup_lo_2540[799:784];
  wire [2047:0] dataGroup_lo_2541 = {dataGroup_lo_hi_2541, dataGroup_lo_lo_2541};
  wire [2047:0] dataGroup_hi_2541 = {dataGroup_hi_hi_2541, dataGroup_hi_lo_2541};
  wire [15:0]   dataGroup_13_43 = dataGroup_lo_2541[863:848];
  wire [2047:0] dataGroup_lo_2542 = {dataGroup_lo_hi_2542, dataGroup_lo_lo_2542};
  wire [2047:0] dataGroup_hi_2542 = {dataGroup_hi_hi_2542, dataGroup_hi_lo_2542};
  wire [15:0]   dataGroup_14_43 = dataGroup_lo_2542[927:912];
  wire [2047:0] dataGroup_lo_2543 = {dataGroup_lo_hi_2543, dataGroup_lo_lo_2543};
  wire [2047:0] dataGroup_hi_2543 = {dataGroup_hi_hi_2543, dataGroup_hi_lo_2543};
  wire [15:0]   dataGroup_15_43 = dataGroup_lo_2543[991:976];
  wire [2047:0] dataGroup_lo_2544 = {dataGroup_lo_hi_2544, dataGroup_lo_lo_2544};
  wire [2047:0] dataGroup_hi_2544 = {dataGroup_hi_hi_2544, dataGroup_hi_lo_2544};
  wire [15:0]   dataGroup_16_43 = dataGroup_lo_2544[1055:1040];
  wire [2047:0] dataGroup_lo_2545 = {dataGroup_lo_hi_2545, dataGroup_lo_lo_2545};
  wire [2047:0] dataGroup_hi_2545 = {dataGroup_hi_hi_2545, dataGroup_hi_lo_2545};
  wire [15:0]   dataGroup_17_43 = dataGroup_lo_2545[1119:1104];
  wire [2047:0] dataGroup_lo_2546 = {dataGroup_lo_hi_2546, dataGroup_lo_lo_2546};
  wire [2047:0] dataGroup_hi_2546 = {dataGroup_hi_hi_2546, dataGroup_hi_lo_2546};
  wire [15:0]   dataGroup_18_43 = dataGroup_lo_2546[1183:1168];
  wire [2047:0] dataGroup_lo_2547 = {dataGroup_lo_hi_2547, dataGroup_lo_lo_2547};
  wire [2047:0] dataGroup_hi_2547 = {dataGroup_hi_hi_2547, dataGroup_hi_lo_2547};
  wire [15:0]   dataGroup_19_43 = dataGroup_lo_2547[1247:1232];
  wire [2047:0] dataGroup_lo_2548 = {dataGroup_lo_hi_2548, dataGroup_lo_lo_2548};
  wire [2047:0] dataGroup_hi_2548 = {dataGroup_hi_hi_2548, dataGroup_hi_lo_2548};
  wire [15:0]   dataGroup_20_43 = dataGroup_lo_2548[1311:1296];
  wire [2047:0] dataGroup_lo_2549 = {dataGroup_lo_hi_2549, dataGroup_lo_lo_2549};
  wire [2047:0] dataGroup_hi_2549 = {dataGroup_hi_hi_2549, dataGroup_hi_lo_2549};
  wire [15:0]   dataGroup_21_43 = dataGroup_lo_2549[1375:1360];
  wire [2047:0] dataGroup_lo_2550 = {dataGroup_lo_hi_2550, dataGroup_lo_lo_2550};
  wire [2047:0] dataGroup_hi_2550 = {dataGroup_hi_hi_2550, dataGroup_hi_lo_2550};
  wire [15:0]   dataGroup_22_43 = dataGroup_lo_2550[1439:1424];
  wire [2047:0] dataGroup_lo_2551 = {dataGroup_lo_hi_2551, dataGroup_lo_lo_2551};
  wire [2047:0] dataGroup_hi_2551 = {dataGroup_hi_hi_2551, dataGroup_hi_lo_2551};
  wire [15:0]   dataGroup_23_43 = dataGroup_lo_2551[1503:1488];
  wire [2047:0] dataGroup_lo_2552 = {dataGroup_lo_hi_2552, dataGroup_lo_lo_2552};
  wire [2047:0] dataGroup_hi_2552 = {dataGroup_hi_hi_2552, dataGroup_hi_lo_2552};
  wire [15:0]   dataGroup_24_43 = dataGroup_lo_2552[1567:1552];
  wire [2047:0] dataGroup_lo_2553 = {dataGroup_lo_hi_2553, dataGroup_lo_lo_2553};
  wire [2047:0] dataGroup_hi_2553 = {dataGroup_hi_hi_2553, dataGroup_hi_lo_2553};
  wire [15:0]   dataGroup_25_43 = dataGroup_lo_2553[1631:1616];
  wire [2047:0] dataGroup_lo_2554 = {dataGroup_lo_hi_2554, dataGroup_lo_lo_2554};
  wire [2047:0] dataGroup_hi_2554 = {dataGroup_hi_hi_2554, dataGroup_hi_lo_2554};
  wire [15:0]   dataGroup_26_43 = dataGroup_lo_2554[1695:1680];
  wire [2047:0] dataGroup_lo_2555 = {dataGroup_lo_hi_2555, dataGroup_lo_lo_2555};
  wire [2047:0] dataGroup_hi_2555 = {dataGroup_hi_hi_2555, dataGroup_hi_lo_2555};
  wire [15:0]   dataGroup_27_43 = dataGroup_lo_2555[1759:1744];
  wire [2047:0] dataGroup_lo_2556 = {dataGroup_lo_hi_2556, dataGroup_lo_lo_2556};
  wire [2047:0] dataGroup_hi_2556 = {dataGroup_hi_hi_2556, dataGroup_hi_lo_2556};
  wire [15:0]   dataGroup_28_43 = dataGroup_lo_2556[1823:1808];
  wire [2047:0] dataGroup_lo_2557 = {dataGroup_lo_hi_2557, dataGroup_lo_lo_2557};
  wire [2047:0] dataGroup_hi_2557 = {dataGroup_hi_hi_2557, dataGroup_hi_lo_2557};
  wire [15:0]   dataGroup_29_43 = dataGroup_lo_2557[1887:1872];
  wire [2047:0] dataGroup_lo_2558 = {dataGroup_lo_hi_2558, dataGroup_lo_lo_2558};
  wire [2047:0] dataGroup_hi_2558 = {dataGroup_hi_hi_2558, dataGroup_hi_lo_2558};
  wire [15:0]   dataGroup_30_43 = dataGroup_lo_2558[1951:1936];
  wire [2047:0] dataGroup_lo_2559 = {dataGroup_lo_hi_2559, dataGroup_lo_lo_2559};
  wire [2047:0] dataGroup_hi_2559 = {dataGroup_hi_hi_2559, dataGroup_hi_lo_2559};
  wire [15:0]   dataGroup_31_43 = dataGroup_lo_2559[2015:2000];
  wire [31:0]   res_lo_lo_lo_lo_43 = {dataGroup_1_43, dataGroup_0_43};
  wire [31:0]   res_lo_lo_lo_hi_43 = {dataGroup_3_43, dataGroup_2_43};
  wire [63:0]   res_lo_lo_lo_43 = {res_lo_lo_lo_hi_43, res_lo_lo_lo_lo_43};
  wire [31:0]   res_lo_lo_hi_lo_43 = {dataGroup_5_43, dataGroup_4_43};
  wire [31:0]   res_lo_lo_hi_hi_43 = {dataGroup_7_43, dataGroup_6_43};
  wire [63:0]   res_lo_lo_hi_43 = {res_lo_lo_hi_hi_43, res_lo_lo_hi_lo_43};
  wire [127:0]  res_lo_lo_43 = {res_lo_lo_hi_43, res_lo_lo_lo_43};
  wire [31:0]   res_lo_hi_lo_lo_43 = {dataGroup_9_43, dataGroup_8_43};
  wire [31:0]   res_lo_hi_lo_hi_43 = {dataGroup_11_43, dataGroup_10_43};
  wire [63:0]   res_lo_hi_lo_43 = {res_lo_hi_lo_hi_43, res_lo_hi_lo_lo_43};
  wire [31:0]   res_lo_hi_hi_lo_43 = {dataGroup_13_43, dataGroup_12_43};
  wire [31:0]   res_lo_hi_hi_hi_43 = {dataGroup_15_43, dataGroup_14_43};
  wire [63:0]   res_lo_hi_hi_43 = {res_lo_hi_hi_hi_43, res_lo_hi_hi_lo_43};
  wire [127:0]  res_lo_hi_43 = {res_lo_hi_hi_43, res_lo_hi_lo_43};
  wire [255:0]  res_lo_43 = {res_lo_hi_43, res_lo_lo_43};
  wire [31:0]   res_hi_lo_lo_lo_43 = {dataGroup_17_43, dataGroup_16_43};
  wire [31:0]   res_hi_lo_lo_hi_43 = {dataGroup_19_43, dataGroup_18_43};
  wire [63:0]   res_hi_lo_lo_43 = {res_hi_lo_lo_hi_43, res_hi_lo_lo_lo_43};
  wire [31:0]   res_hi_lo_hi_lo_43 = {dataGroup_21_43, dataGroup_20_43};
  wire [31:0]   res_hi_lo_hi_hi_43 = {dataGroup_23_43, dataGroup_22_43};
  wire [63:0]   res_hi_lo_hi_43 = {res_hi_lo_hi_hi_43, res_hi_lo_hi_lo_43};
  wire [127:0]  res_hi_lo_43 = {res_hi_lo_hi_43, res_hi_lo_lo_43};
  wire [31:0]   res_hi_hi_lo_lo_43 = {dataGroup_25_43, dataGroup_24_43};
  wire [31:0]   res_hi_hi_lo_hi_43 = {dataGroup_27_43, dataGroup_26_43};
  wire [63:0]   res_hi_hi_lo_43 = {res_hi_hi_lo_hi_43, res_hi_hi_lo_lo_43};
  wire [31:0]   res_hi_hi_hi_lo_43 = {dataGroup_29_43, dataGroup_28_43};
  wire [31:0]   res_hi_hi_hi_hi_43 = {dataGroup_31_43, dataGroup_30_43};
  wire [63:0]   res_hi_hi_hi_43 = {res_hi_hi_hi_hi_43, res_hi_hi_hi_lo_43};
  wire [127:0]  res_hi_hi_43 = {res_hi_hi_hi_43, res_hi_hi_lo_43};
  wire [255:0]  res_hi_43 = {res_hi_hi_43, res_hi_lo_43};
  wire [511:0]  res_89 = {res_hi_43, res_lo_43};
  wire [2047:0] dataGroup_lo_2560 = {dataGroup_lo_hi_2560, dataGroup_lo_lo_2560};
  wire [2047:0] dataGroup_hi_2560 = {dataGroup_hi_hi_2560, dataGroup_hi_lo_2560};
  wire [15:0]   dataGroup_0_44 = dataGroup_lo_2560[47:32];
  wire [2047:0] dataGroup_lo_2561 = {dataGroup_lo_hi_2561, dataGroup_lo_lo_2561};
  wire [2047:0] dataGroup_hi_2561 = {dataGroup_hi_hi_2561, dataGroup_hi_lo_2561};
  wire [15:0]   dataGroup_1_44 = dataGroup_lo_2561[111:96];
  wire [2047:0] dataGroup_lo_2562 = {dataGroup_lo_hi_2562, dataGroup_lo_lo_2562};
  wire [2047:0] dataGroup_hi_2562 = {dataGroup_hi_hi_2562, dataGroup_hi_lo_2562};
  wire [15:0]   dataGroup_2_44 = dataGroup_lo_2562[175:160];
  wire [2047:0] dataGroup_lo_2563 = {dataGroup_lo_hi_2563, dataGroup_lo_lo_2563};
  wire [2047:0] dataGroup_hi_2563 = {dataGroup_hi_hi_2563, dataGroup_hi_lo_2563};
  wire [15:0]   dataGroup_3_44 = dataGroup_lo_2563[239:224];
  wire [2047:0] dataGroup_lo_2564 = {dataGroup_lo_hi_2564, dataGroup_lo_lo_2564};
  wire [2047:0] dataGroup_hi_2564 = {dataGroup_hi_hi_2564, dataGroup_hi_lo_2564};
  wire [15:0]   dataGroup_4_44 = dataGroup_lo_2564[303:288];
  wire [2047:0] dataGroup_lo_2565 = {dataGroup_lo_hi_2565, dataGroup_lo_lo_2565};
  wire [2047:0] dataGroup_hi_2565 = {dataGroup_hi_hi_2565, dataGroup_hi_lo_2565};
  wire [15:0]   dataGroup_5_44 = dataGroup_lo_2565[367:352];
  wire [2047:0] dataGroup_lo_2566 = {dataGroup_lo_hi_2566, dataGroup_lo_lo_2566};
  wire [2047:0] dataGroup_hi_2566 = {dataGroup_hi_hi_2566, dataGroup_hi_lo_2566};
  wire [15:0]   dataGroup_6_44 = dataGroup_lo_2566[431:416];
  wire [2047:0] dataGroup_lo_2567 = {dataGroup_lo_hi_2567, dataGroup_lo_lo_2567};
  wire [2047:0] dataGroup_hi_2567 = {dataGroup_hi_hi_2567, dataGroup_hi_lo_2567};
  wire [15:0]   dataGroup_7_44 = dataGroup_lo_2567[495:480];
  wire [2047:0] dataGroup_lo_2568 = {dataGroup_lo_hi_2568, dataGroup_lo_lo_2568};
  wire [2047:0] dataGroup_hi_2568 = {dataGroup_hi_hi_2568, dataGroup_hi_lo_2568};
  wire [15:0]   dataGroup_8_44 = dataGroup_lo_2568[559:544];
  wire [2047:0] dataGroup_lo_2569 = {dataGroup_lo_hi_2569, dataGroup_lo_lo_2569};
  wire [2047:0] dataGroup_hi_2569 = {dataGroup_hi_hi_2569, dataGroup_hi_lo_2569};
  wire [15:0]   dataGroup_9_44 = dataGroup_lo_2569[623:608];
  wire [2047:0] dataGroup_lo_2570 = {dataGroup_lo_hi_2570, dataGroup_lo_lo_2570};
  wire [2047:0] dataGroup_hi_2570 = {dataGroup_hi_hi_2570, dataGroup_hi_lo_2570};
  wire [15:0]   dataGroup_10_44 = dataGroup_lo_2570[687:672];
  wire [2047:0] dataGroup_lo_2571 = {dataGroup_lo_hi_2571, dataGroup_lo_lo_2571};
  wire [2047:0] dataGroup_hi_2571 = {dataGroup_hi_hi_2571, dataGroup_hi_lo_2571};
  wire [15:0]   dataGroup_11_44 = dataGroup_lo_2571[751:736];
  wire [2047:0] dataGroup_lo_2572 = {dataGroup_lo_hi_2572, dataGroup_lo_lo_2572};
  wire [2047:0] dataGroup_hi_2572 = {dataGroup_hi_hi_2572, dataGroup_hi_lo_2572};
  wire [15:0]   dataGroup_12_44 = dataGroup_lo_2572[815:800];
  wire [2047:0] dataGroup_lo_2573 = {dataGroup_lo_hi_2573, dataGroup_lo_lo_2573};
  wire [2047:0] dataGroup_hi_2573 = {dataGroup_hi_hi_2573, dataGroup_hi_lo_2573};
  wire [15:0]   dataGroup_13_44 = dataGroup_lo_2573[879:864];
  wire [2047:0] dataGroup_lo_2574 = {dataGroup_lo_hi_2574, dataGroup_lo_lo_2574};
  wire [2047:0] dataGroup_hi_2574 = {dataGroup_hi_hi_2574, dataGroup_hi_lo_2574};
  wire [15:0]   dataGroup_14_44 = dataGroup_lo_2574[943:928];
  wire [2047:0] dataGroup_lo_2575 = {dataGroup_lo_hi_2575, dataGroup_lo_lo_2575};
  wire [2047:0] dataGroup_hi_2575 = {dataGroup_hi_hi_2575, dataGroup_hi_lo_2575};
  wire [15:0]   dataGroup_15_44 = dataGroup_lo_2575[1007:992];
  wire [2047:0] dataGroup_lo_2576 = {dataGroup_lo_hi_2576, dataGroup_lo_lo_2576};
  wire [2047:0] dataGroup_hi_2576 = {dataGroup_hi_hi_2576, dataGroup_hi_lo_2576};
  wire [15:0]   dataGroup_16_44 = dataGroup_lo_2576[1071:1056];
  wire [2047:0] dataGroup_lo_2577 = {dataGroup_lo_hi_2577, dataGroup_lo_lo_2577};
  wire [2047:0] dataGroup_hi_2577 = {dataGroup_hi_hi_2577, dataGroup_hi_lo_2577};
  wire [15:0]   dataGroup_17_44 = dataGroup_lo_2577[1135:1120];
  wire [2047:0] dataGroup_lo_2578 = {dataGroup_lo_hi_2578, dataGroup_lo_lo_2578};
  wire [2047:0] dataGroup_hi_2578 = {dataGroup_hi_hi_2578, dataGroup_hi_lo_2578};
  wire [15:0]   dataGroup_18_44 = dataGroup_lo_2578[1199:1184];
  wire [2047:0] dataGroup_lo_2579 = {dataGroup_lo_hi_2579, dataGroup_lo_lo_2579};
  wire [2047:0] dataGroup_hi_2579 = {dataGroup_hi_hi_2579, dataGroup_hi_lo_2579};
  wire [15:0]   dataGroup_19_44 = dataGroup_lo_2579[1263:1248];
  wire [2047:0] dataGroup_lo_2580 = {dataGroup_lo_hi_2580, dataGroup_lo_lo_2580};
  wire [2047:0] dataGroup_hi_2580 = {dataGroup_hi_hi_2580, dataGroup_hi_lo_2580};
  wire [15:0]   dataGroup_20_44 = dataGroup_lo_2580[1327:1312];
  wire [2047:0] dataGroup_lo_2581 = {dataGroup_lo_hi_2581, dataGroup_lo_lo_2581};
  wire [2047:0] dataGroup_hi_2581 = {dataGroup_hi_hi_2581, dataGroup_hi_lo_2581};
  wire [15:0]   dataGroup_21_44 = dataGroup_lo_2581[1391:1376];
  wire [2047:0] dataGroup_lo_2582 = {dataGroup_lo_hi_2582, dataGroup_lo_lo_2582};
  wire [2047:0] dataGroup_hi_2582 = {dataGroup_hi_hi_2582, dataGroup_hi_lo_2582};
  wire [15:0]   dataGroup_22_44 = dataGroup_lo_2582[1455:1440];
  wire [2047:0] dataGroup_lo_2583 = {dataGroup_lo_hi_2583, dataGroup_lo_lo_2583};
  wire [2047:0] dataGroup_hi_2583 = {dataGroup_hi_hi_2583, dataGroup_hi_lo_2583};
  wire [15:0]   dataGroup_23_44 = dataGroup_lo_2583[1519:1504];
  wire [2047:0] dataGroup_lo_2584 = {dataGroup_lo_hi_2584, dataGroup_lo_lo_2584};
  wire [2047:0] dataGroup_hi_2584 = {dataGroup_hi_hi_2584, dataGroup_hi_lo_2584};
  wire [15:0]   dataGroup_24_44 = dataGroup_lo_2584[1583:1568];
  wire [2047:0] dataGroup_lo_2585 = {dataGroup_lo_hi_2585, dataGroup_lo_lo_2585};
  wire [2047:0] dataGroup_hi_2585 = {dataGroup_hi_hi_2585, dataGroup_hi_lo_2585};
  wire [15:0]   dataGroup_25_44 = dataGroup_lo_2585[1647:1632];
  wire [2047:0] dataGroup_lo_2586 = {dataGroup_lo_hi_2586, dataGroup_lo_lo_2586};
  wire [2047:0] dataGroup_hi_2586 = {dataGroup_hi_hi_2586, dataGroup_hi_lo_2586};
  wire [15:0]   dataGroup_26_44 = dataGroup_lo_2586[1711:1696];
  wire [2047:0] dataGroup_lo_2587 = {dataGroup_lo_hi_2587, dataGroup_lo_lo_2587};
  wire [2047:0] dataGroup_hi_2587 = {dataGroup_hi_hi_2587, dataGroup_hi_lo_2587};
  wire [15:0]   dataGroup_27_44 = dataGroup_lo_2587[1775:1760];
  wire [2047:0] dataGroup_lo_2588 = {dataGroup_lo_hi_2588, dataGroup_lo_lo_2588};
  wire [2047:0] dataGroup_hi_2588 = {dataGroup_hi_hi_2588, dataGroup_hi_lo_2588};
  wire [15:0]   dataGroup_28_44 = dataGroup_lo_2588[1839:1824];
  wire [2047:0] dataGroup_lo_2589 = {dataGroup_lo_hi_2589, dataGroup_lo_lo_2589};
  wire [2047:0] dataGroup_hi_2589 = {dataGroup_hi_hi_2589, dataGroup_hi_lo_2589};
  wire [15:0]   dataGroup_29_44 = dataGroup_lo_2589[1903:1888];
  wire [2047:0] dataGroup_lo_2590 = {dataGroup_lo_hi_2590, dataGroup_lo_lo_2590};
  wire [2047:0] dataGroup_hi_2590 = {dataGroup_hi_hi_2590, dataGroup_hi_lo_2590};
  wire [15:0]   dataGroup_30_44 = dataGroup_lo_2590[1967:1952];
  wire [2047:0] dataGroup_lo_2591 = {dataGroup_lo_hi_2591, dataGroup_lo_lo_2591};
  wire [2047:0] dataGroup_hi_2591 = {dataGroup_hi_hi_2591, dataGroup_hi_lo_2591};
  wire [15:0]   dataGroup_31_44 = dataGroup_lo_2591[2031:2016];
  wire [31:0]   res_lo_lo_lo_lo_44 = {dataGroup_1_44, dataGroup_0_44};
  wire [31:0]   res_lo_lo_lo_hi_44 = {dataGroup_3_44, dataGroup_2_44};
  wire [63:0]   res_lo_lo_lo_44 = {res_lo_lo_lo_hi_44, res_lo_lo_lo_lo_44};
  wire [31:0]   res_lo_lo_hi_lo_44 = {dataGroup_5_44, dataGroup_4_44};
  wire [31:0]   res_lo_lo_hi_hi_44 = {dataGroup_7_44, dataGroup_6_44};
  wire [63:0]   res_lo_lo_hi_44 = {res_lo_lo_hi_hi_44, res_lo_lo_hi_lo_44};
  wire [127:0]  res_lo_lo_44 = {res_lo_lo_hi_44, res_lo_lo_lo_44};
  wire [31:0]   res_lo_hi_lo_lo_44 = {dataGroup_9_44, dataGroup_8_44};
  wire [31:0]   res_lo_hi_lo_hi_44 = {dataGroup_11_44, dataGroup_10_44};
  wire [63:0]   res_lo_hi_lo_44 = {res_lo_hi_lo_hi_44, res_lo_hi_lo_lo_44};
  wire [31:0]   res_lo_hi_hi_lo_44 = {dataGroup_13_44, dataGroup_12_44};
  wire [31:0]   res_lo_hi_hi_hi_44 = {dataGroup_15_44, dataGroup_14_44};
  wire [63:0]   res_lo_hi_hi_44 = {res_lo_hi_hi_hi_44, res_lo_hi_hi_lo_44};
  wire [127:0]  res_lo_hi_44 = {res_lo_hi_hi_44, res_lo_hi_lo_44};
  wire [255:0]  res_lo_44 = {res_lo_hi_44, res_lo_lo_44};
  wire [31:0]   res_hi_lo_lo_lo_44 = {dataGroup_17_44, dataGroup_16_44};
  wire [31:0]   res_hi_lo_lo_hi_44 = {dataGroup_19_44, dataGroup_18_44};
  wire [63:0]   res_hi_lo_lo_44 = {res_hi_lo_lo_hi_44, res_hi_lo_lo_lo_44};
  wire [31:0]   res_hi_lo_hi_lo_44 = {dataGroup_21_44, dataGroup_20_44};
  wire [31:0]   res_hi_lo_hi_hi_44 = {dataGroup_23_44, dataGroup_22_44};
  wire [63:0]   res_hi_lo_hi_44 = {res_hi_lo_hi_hi_44, res_hi_lo_hi_lo_44};
  wire [127:0]  res_hi_lo_44 = {res_hi_lo_hi_44, res_hi_lo_lo_44};
  wire [31:0]   res_hi_hi_lo_lo_44 = {dataGroup_25_44, dataGroup_24_44};
  wire [31:0]   res_hi_hi_lo_hi_44 = {dataGroup_27_44, dataGroup_26_44};
  wire [63:0]   res_hi_hi_lo_44 = {res_hi_hi_lo_hi_44, res_hi_hi_lo_lo_44};
  wire [31:0]   res_hi_hi_hi_lo_44 = {dataGroup_29_44, dataGroup_28_44};
  wire [31:0]   res_hi_hi_hi_hi_44 = {dataGroup_31_44, dataGroup_30_44};
  wire [63:0]   res_hi_hi_hi_44 = {res_hi_hi_hi_hi_44, res_hi_hi_hi_lo_44};
  wire [127:0]  res_hi_hi_44 = {res_hi_hi_hi_44, res_hi_hi_lo_44};
  wire [255:0]  res_hi_44 = {res_hi_hi_44, res_hi_lo_44};
  wire [511:0]  res_90 = {res_hi_44, res_lo_44};
  wire [2047:0] dataGroup_lo_2592 = {dataGroup_lo_hi_2592, dataGroup_lo_lo_2592};
  wire [2047:0] dataGroup_hi_2592 = {dataGroup_hi_hi_2592, dataGroup_hi_lo_2592};
  wire [15:0]   dataGroup_0_45 = dataGroup_lo_2592[63:48];
  wire [2047:0] dataGroup_lo_2593 = {dataGroup_lo_hi_2593, dataGroup_lo_lo_2593};
  wire [2047:0] dataGroup_hi_2593 = {dataGroup_hi_hi_2593, dataGroup_hi_lo_2593};
  wire [15:0]   dataGroup_1_45 = dataGroup_lo_2593[127:112];
  wire [2047:0] dataGroup_lo_2594 = {dataGroup_lo_hi_2594, dataGroup_lo_lo_2594};
  wire [2047:0] dataGroup_hi_2594 = {dataGroup_hi_hi_2594, dataGroup_hi_lo_2594};
  wire [15:0]   dataGroup_2_45 = dataGroup_lo_2594[191:176];
  wire [2047:0] dataGroup_lo_2595 = {dataGroup_lo_hi_2595, dataGroup_lo_lo_2595};
  wire [2047:0] dataGroup_hi_2595 = {dataGroup_hi_hi_2595, dataGroup_hi_lo_2595};
  wire [15:0]   dataGroup_3_45 = dataGroup_lo_2595[255:240];
  wire [2047:0] dataGroup_lo_2596 = {dataGroup_lo_hi_2596, dataGroup_lo_lo_2596};
  wire [2047:0] dataGroup_hi_2596 = {dataGroup_hi_hi_2596, dataGroup_hi_lo_2596};
  wire [15:0]   dataGroup_4_45 = dataGroup_lo_2596[319:304];
  wire [2047:0] dataGroup_lo_2597 = {dataGroup_lo_hi_2597, dataGroup_lo_lo_2597};
  wire [2047:0] dataGroup_hi_2597 = {dataGroup_hi_hi_2597, dataGroup_hi_lo_2597};
  wire [15:0]   dataGroup_5_45 = dataGroup_lo_2597[383:368];
  wire [2047:0] dataGroup_lo_2598 = {dataGroup_lo_hi_2598, dataGroup_lo_lo_2598};
  wire [2047:0] dataGroup_hi_2598 = {dataGroup_hi_hi_2598, dataGroup_hi_lo_2598};
  wire [15:0]   dataGroup_6_45 = dataGroup_lo_2598[447:432];
  wire [2047:0] dataGroup_lo_2599 = {dataGroup_lo_hi_2599, dataGroup_lo_lo_2599};
  wire [2047:0] dataGroup_hi_2599 = {dataGroup_hi_hi_2599, dataGroup_hi_lo_2599};
  wire [15:0]   dataGroup_7_45 = dataGroup_lo_2599[511:496];
  wire [2047:0] dataGroup_lo_2600 = {dataGroup_lo_hi_2600, dataGroup_lo_lo_2600};
  wire [2047:0] dataGroup_hi_2600 = {dataGroup_hi_hi_2600, dataGroup_hi_lo_2600};
  wire [15:0]   dataGroup_8_45 = dataGroup_lo_2600[575:560];
  wire [2047:0] dataGroup_lo_2601 = {dataGroup_lo_hi_2601, dataGroup_lo_lo_2601};
  wire [2047:0] dataGroup_hi_2601 = {dataGroup_hi_hi_2601, dataGroup_hi_lo_2601};
  wire [15:0]   dataGroup_9_45 = dataGroup_lo_2601[639:624];
  wire [2047:0] dataGroup_lo_2602 = {dataGroup_lo_hi_2602, dataGroup_lo_lo_2602};
  wire [2047:0] dataGroup_hi_2602 = {dataGroup_hi_hi_2602, dataGroup_hi_lo_2602};
  wire [15:0]   dataGroup_10_45 = dataGroup_lo_2602[703:688];
  wire [2047:0] dataGroup_lo_2603 = {dataGroup_lo_hi_2603, dataGroup_lo_lo_2603};
  wire [2047:0] dataGroup_hi_2603 = {dataGroup_hi_hi_2603, dataGroup_hi_lo_2603};
  wire [15:0]   dataGroup_11_45 = dataGroup_lo_2603[767:752];
  wire [2047:0] dataGroup_lo_2604 = {dataGroup_lo_hi_2604, dataGroup_lo_lo_2604};
  wire [2047:0] dataGroup_hi_2604 = {dataGroup_hi_hi_2604, dataGroup_hi_lo_2604};
  wire [15:0]   dataGroup_12_45 = dataGroup_lo_2604[831:816];
  wire [2047:0] dataGroup_lo_2605 = {dataGroup_lo_hi_2605, dataGroup_lo_lo_2605};
  wire [2047:0] dataGroup_hi_2605 = {dataGroup_hi_hi_2605, dataGroup_hi_lo_2605};
  wire [15:0]   dataGroup_13_45 = dataGroup_lo_2605[895:880];
  wire [2047:0] dataGroup_lo_2606 = {dataGroup_lo_hi_2606, dataGroup_lo_lo_2606};
  wire [2047:0] dataGroup_hi_2606 = {dataGroup_hi_hi_2606, dataGroup_hi_lo_2606};
  wire [15:0]   dataGroup_14_45 = dataGroup_lo_2606[959:944];
  wire [2047:0] dataGroup_lo_2607 = {dataGroup_lo_hi_2607, dataGroup_lo_lo_2607};
  wire [2047:0] dataGroup_hi_2607 = {dataGroup_hi_hi_2607, dataGroup_hi_lo_2607};
  wire [15:0]   dataGroup_15_45 = dataGroup_lo_2607[1023:1008];
  wire [2047:0] dataGroup_lo_2608 = {dataGroup_lo_hi_2608, dataGroup_lo_lo_2608};
  wire [2047:0] dataGroup_hi_2608 = {dataGroup_hi_hi_2608, dataGroup_hi_lo_2608};
  wire [15:0]   dataGroup_16_45 = dataGroup_lo_2608[1087:1072];
  wire [2047:0] dataGroup_lo_2609 = {dataGroup_lo_hi_2609, dataGroup_lo_lo_2609};
  wire [2047:0] dataGroup_hi_2609 = {dataGroup_hi_hi_2609, dataGroup_hi_lo_2609};
  wire [15:0]   dataGroup_17_45 = dataGroup_lo_2609[1151:1136];
  wire [2047:0] dataGroup_lo_2610 = {dataGroup_lo_hi_2610, dataGroup_lo_lo_2610};
  wire [2047:0] dataGroup_hi_2610 = {dataGroup_hi_hi_2610, dataGroup_hi_lo_2610};
  wire [15:0]   dataGroup_18_45 = dataGroup_lo_2610[1215:1200];
  wire [2047:0] dataGroup_lo_2611 = {dataGroup_lo_hi_2611, dataGroup_lo_lo_2611};
  wire [2047:0] dataGroup_hi_2611 = {dataGroup_hi_hi_2611, dataGroup_hi_lo_2611};
  wire [15:0]   dataGroup_19_45 = dataGroup_lo_2611[1279:1264];
  wire [2047:0] dataGroup_lo_2612 = {dataGroup_lo_hi_2612, dataGroup_lo_lo_2612};
  wire [2047:0] dataGroup_hi_2612 = {dataGroup_hi_hi_2612, dataGroup_hi_lo_2612};
  wire [15:0]   dataGroup_20_45 = dataGroup_lo_2612[1343:1328];
  wire [2047:0] dataGroup_lo_2613 = {dataGroup_lo_hi_2613, dataGroup_lo_lo_2613};
  wire [2047:0] dataGroup_hi_2613 = {dataGroup_hi_hi_2613, dataGroup_hi_lo_2613};
  wire [15:0]   dataGroup_21_45 = dataGroup_lo_2613[1407:1392];
  wire [2047:0] dataGroup_lo_2614 = {dataGroup_lo_hi_2614, dataGroup_lo_lo_2614};
  wire [2047:0] dataGroup_hi_2614 = {dataGroup_hi_hi_2614, dataGroup_hi_lo_2614};
  wire [15:0]   dataGroup_22_45 = dataGroup_lo_2614[1471:1456];
  wire [2047:0] dataGroup_lo_2615 = {dataGroup_lo_hi_2615, dataGroup_lo_lo_2615};
  wire [2047:0] dataGroup_hi_2615 = {dataGroup_hi_hi_2615, dataGroup_hi_lo_2615};
  wire [15:0]   dataGroup_23_45 = dataGroup_lo_2615[1535:1520];
  wire [2047:0] dataGroup_lo_2616 = {dataGroup_lo_hi_2616, dataGroup_lo_lo_2616};
  wire [2047:0] dataGroup_hi_2616 = {dataGroup_hi_hi_2616, dataGroup_hi_lo_2616};
  wire [15:0]   dataGroup_24_45 = dataGroup_lo_2616[1599:1584];
  wire [2047:0] dataGroup_lo_2617 = {dataGroup_lo_hi_2617, dataGroup_lo_lo_2617};
  wire [2047:0] dataGroup_hi_2617 = {dataGroup_hi_hi_2617, dataGroup_hi_lo_2617};
  wire [15:0]   dataGroup_25_45 = dataGroup_lo_2617[1663:1648];
  wire [2047:0] dataGroup_lo_2618 = {dataGroup_lo_hi_2618, dataGroup_lo_lo_2618};
  wire [2047:0] dataGroup_hi_2618 = {dataGroup_hi_hi_2618, dataGroup_hi_lo_2618};
  wire [15:0]   dataGroup_26_45 = dataGroup_lo_2618[1727:1712];
  wire [2047:0] dataGroup_lo_2619 = {dataGroup_lo_hi_2619, dataGroup_lo_lo_2619};
  wire [2047:0] dataGroup_hi_2619 = {dataGroup_hi_hi_2619, dataGroup_hi_lo_2619};
  wire [15:0]   dataGroup_27_45 = dataGroup_lo_2619[1791:1776];
  wire [2047:0] dataGroup_lo_2620 = {dataGroup_lo_hi_2620, dataGroup_lo_lo_2620};
  wire [2047:0] dataGroup_hi_2620 = {dataGroup_hi_hi_2620, dataGroup_hi_lo_2620};
  wire [15:0]   dataGroup_28_45 = dataGroup_lo_2620[1855:1840];
  wire [2047:0] dataGroup_lo_2621 = {dataGroup_lo_hi_2621, dataGroup_lo_lo_2621};
  wire [2047:0] dataGroup_hi_2621 = {dataGroup_hi_hi_2621, dataGroup_hi_lo_2621};
  wire [15:0]   dataGroup_29_45 = dataGroup_lo_2621[1919:1904];
  wire [2047:0] dataGroup_lo_2622 = {dataGroup_lo_hi_2622, dataGroup_lo_lo_2622};
  wire [2047:0] dataGroup_hi_2622 = {dataGroup_hi_hi_2622, dataGroup_hi_lo_2622};
  wire [15:0]   dataGroup_30_45 = dataGroup_lo_2622[1983:1968];
  wire [2047:0] dataGroup_lo_2623 = {dataGroup_lo_hi_2623, dataGroup_lo_lo_2623};
  wire [2047:0] dataGroup_hi_2623 = {dataGroup_hi_hi_2623, dataGroup_hi_lo_2623};
  wire [15:0]   dataGroup_31_45 = dataGroup_lo_2623[2047:2032];
  wire [31:0]   res_lo_lo_lo_lo_45 = {dataGroup_1_45, dataGroup_0_45};
  wire [31:0]   res_lo_lo_lo_hi_45 = {dataGroup_3_45, dataGroup_2_45};
  wire [63:0]   res_lo_lo_lo_45 = {res_lo_lo_lo_hi_45, res_lo_lo_lo_lo_45};
  wire [31:0]   res_lo_lo_hi_lo_45 = {dataGroup_5_45, dataGroup_4_45};
  wire [31:0]   res_lo_lo_hi_hi_45 = {dataGroup_7_45, dataGroup_6_45};
  wire [63:0]   res_lo_lo_hi_45 = {res_lo_lo_hi_hi_45, res_lo_lo_hi_lo_45};
  wire [127:0]  res_lo_lo_45 = {res_lo_lo_hi_45, res_lo_lo_lo_45};
  wire [31:0]   res_lo_hi_lo_lo_45 = {dataGroup_9_45, dataGroup_8_45};
  wire [31:0]   res_lo_hi_lo_hi_45 = {dataGroup_11_45, dataGroup_10_45};
  wire [63:0]   res_lo_hi_lo_45 = {res_lo_hi_lo_hi_45, res_lo_hi_lo_lo_45};
  wire [31:0]   res_lo_hi_hi_lo_45 = {dataGroup_13_45, dataGroup_12_45};
  wire [31:0]   res_lo_hi_hi_hi_45 = {dataGroup_15_45, dataGroup_14_45};
  wire [63:0]   res_lo_hi_hi_45 = {res_lo_hi_hi_hi_45, res_lo_hi_hi_lo_45};
  wire [127:0]  res_lo_hi_45 = {res_lo_hi_hi_45, res_lo_hi_lo_45};
  wire [255:0]  res_lo_45 = {res_lo_hi_45, res_lo_lo_45};
  wire [31:0]   res_hi_lo_lo_lo_45 = {dataGroup_17_45, dataGroup_16_45};
  wire [31:0]   res_hi_lo_lo_hi_45 = {dataGroup_19_45, dataGroup_18_45};
  wire [63:0]   res_hi_lo_lo_45 = {res_hi_lo_lo_hi_45, res_hi_lo_lo_lo_45};
  wire [31:0]   res_hi_lo_hi_lo_45 = {dataGroup_21_45, dataGroup_20_45};
  wire [31:0]   res_hi_lo_hi_hi_45 = {dataGroup_23_45, dataGroup_22_45};
  wire [63:0]   res_hi_lo_hi_45 = {res_hi_lo_hi_hi_45, res_hi_lo_hi_lo_45};
  wire [127:0]  res_hi_lo_45 = {res_hi_lo_hi_45, res_hi_lo_lo_45};
  wire [31:0]   res_hi_hi_lo_lo_45 = {dataGroup_25_45, dataGroup_24_45};
  wire [31:0]   res_hi_hi_lo_hi_45 = {dataGroup_27_45, dataGroup_26_45};
  wire [63:0]   res_hi_hi_lo_45 = {res_hi_hi_lo_hi_45, res_hi_hi_lo_lo_45};
  wire [31:0]   res_hi_hi_hi_lo_45 = {dataGroup_29_45, dataGroup_28_45};
  wire [31:0]   res_hi_hi_hi_hi_45 = {dataGroup_31_45, dataGroup_30_45};
  wire [63:0]   res_hi_hi_hi_45 = {res_hi_hi_hi_hi_45, res_hi_hi_hi_lo_45};
  wire [127:0]  res_hi_hi_45 = {res_hi_hi_hi_45, res_hi_hi_lo_45};
  wire [255:0]  res_hi_45 = {res_hi_hi_45, res_hi_lo_45};
  wire [511:0]  res_91 = {res_hi_45, res_lo_45};
  wire [1023:0] lo_lo_11 = {res_89, res_88};
  wire [1023:0] lo_hi_11 = {res_91, res_90};
  wire [2047:0] lo_11 = {lo_hi_11, lo_lo_11};
  wire [4095:0] regroupLoadData_1_3 = {2048'h0, lo_11};
  wire [2047:0] dataGroup_lo_2624 = {dataGroup_lo_hi_2624, dataGroup_lo_lo_2624};
  wire [2047:0] dataGroup_hi_2624 = {dataGroup_hi_hi_2624, dataGroup_hi_lo_2624};
  wire [15:0]   dataGroup_0_46 = dataGroup_lo_2624[15:0];
  wire [2047:0] dataGroup_lo_2625 = {dataGroup_lo_hi_2625, dataGroup_lo_lo_2625};
  wire [2047:0] dataGroup_hi_2625 = {dataGroup_hi_hi_2625, dataGroup_hi_lo_2625};
  wire [15:0]   dataGroup_1_46 = dataGroup_lo_2625[95:80];
  wire [2047:0] dataGroup_lo_2626 = {dataGroup_lo_hi_2626, dataGroup_lo_lo_2626};
  wire [2047:0] dataGroup_hi_2626 = {dataGroup_hi_hi_2626, dataGroup_hi_lo_2626};
  wire [15:0]   dataGroup_2_46 = dataGroup_lo_2626[175:160];
  wire [2047:0] dataGroup_lo_2627 = {dataGroup_lo_hi_2627, dataGroup_lo_lo_2627};
  wire [2047:0] dataGroup_hi_2627 = {dataGroup_hi_hi_2627, dataGroup_hi_lo_2627};
  wire [15:0]   dataGroup_3_46 = dataGroup_lo_2627[255:240];
  wire [2047:0] dataGroup_lo_2628 = {dataGroup_lo_hi_2628, dataGroup_lo_lo_2628};
  wire [2047:0] dataGroup_hi_2628 = {dataGroup_hi_hi_2628, dataGroup_hi_lo_2628};
  wire [15:0]   dataGroup_4_46 = dataGroup_lo_2628[335:320];
  wire [2047:0] dataGroup_lo_2629 = {dataGroup_lo_hi_2629, dataGroup_lo_lo_2629};
  wire [2047:0] dataGroup_hi_2629 = {dataGroup_hi_hi_2629, dataGroup_hi_lo_2629};
  wire [15:0]   dataGroup_5_46 = dataGroup_lo_2629[415:400];
  wire [2047:0] dataGroup_lo_2630 = {dataGroup_lo_hi_2630, dataGroup_lo_lo_2630};
  wire [2047:0] dataGroup_hi_2630 = {dataGroup_hi_hi_2630, dataGroup_hi_lo_2630};
  wire [15:0]   dataGroup_6_46 = dataGroup_lo_2630[495:480];
  wire [2047:0] dataGroup_lo_2631 = {dataGroup_lo_hi_2631, dataGroup_lo_lo_2631};
  wire [2047:0] dataGroup_hi_2631 = {dataGroup_hi_hi_2631, dataGroup_hi_lo_2631};
  wire [15:0]   dataGroup_7_46 = dataGroup_lo_2631[575:560];
  wire [2047:0] dataGroup_lo_2632 = {dataGroup_lo_hi_2632, dataGroup_lo_lo_2632};
  wire [2047:0] dataGroup_hi_2632 = {dataGroup_hi_hi_2632, dataGroup_hi_lo_2632};
  wire [15:0]   dataGroup_8_46 = dataGroup_lo_2632[655:640];
  wire [2047:0] dataGroup_lo_2633 = {dataGroup_lo_hi_2633, dataGroup_lo_lo_2633};
  wire [2047:0] dataGroup_hi_2633 = {dataGroup_hi_hi_2633, dataGroup_hi_lo_2633};
  wire [15:0]   dataGroup_9_46 = dataGroup_lo_2633[735:720];
  wire [2047:0] dataGroup_lo_2634 = {dataGroup_lo_hi_2634, dataGroup_lo_lo_2634};
  wire [2047:0] dataGroup_hi_2634 = {dataGroup_hi_hi_2634, dataGroup_hi_lo_2634};
  wire [15:0]   dataGroup_10_46 = dataGroup_lo_2634[815:800];
  wire [2047:0] dataGroup_lo_2635 = {dataGroup_lo_hi_2635, dataGroup_lo_lo_2635};
  wire [2047:0] dataGroup_hi_2635 = {dataGroup_hi_hi_2635, dataGroup_hi_lo_2635};
  wire [15:0]   dataGroup_11_46 = dataGroup_lo_2635[895:880];
  wire [2047:0] dataGroup_lo_2636 = {dataGroup_lo_hi_2636, dataGroup_lo_lo_2636};
  wire [2047:0] dataGroup_hi_2636 = {dataGroup_hi_hi_2636, dataGroup_hi_lo_2636};
  wire [15:0]   dataGroup_12_46 = dataGroup_lo_2636[975:960];
  wire [2047:0] dataGroup_lo_2637 = {dataGroup_lo_hi_2637, dataGroup_lo_lo_2637};
  wire [2047:0] dataGroup_hi_2637 = {dataGroup_hi_hi_2637, dataGroup_hi_lo_2637};
  wire [15:0]   dataGroup_13_46 = dataGroup_lo_2637[1055:1040];
  wire [2047:0] dataGroup_lo_2638 = {dataGroup_lo_hi_2638, dataGroup_lo_lo_2638};
  wire [2047:0] dataGroup_hi_2638 = {dataGroup_hi_hi_2638, dataGroup_hi_lo_2638};
  wire [15:0]   dataGroup_14_46 = dataGroup_lo_2638[1135:1120];
  wire [2047:0] dataGroup_lo_2639 = {dataGroup_lo_hi_2639, dataGroup_lo_lo_2639};
  wire [2047:0] dataGroup_hi_2639 = {dataGroup_hi_hi_2639, dataGroup_hi_lo_2639};
  wire [15:0]   dataGroup_15_46 = dataGroup_lo_2639[1215:1200];
  wire [2047:0] dataGroup_lo_2640 = {dataGroup_lo_hi_2640, dataGroup_lo_lo_2640};
  wire [2047:0] dataGroup_hi_2640 = {dataGroup_hi_hi_2640, dataGroup_hi_lo_2640};
  wire [15:0]   dataGroup_16_46 = dataGroup_lo_2640[1295:1280];
  wire [2047:0] dataGroup_lo_2641 = {dataGroup_lo_hi_2641, dataGroup_lo_lo_2641};
  wire [2047:0] dataGroup_hi_2641 = {dataGroup_hi_hi_2641, dataGroup_hi_lo_2641};
  wire [15:0]   dataGroup_17_46 = dataGroup_lo_2641[1375:1360];
  wire [2047:0] dataGroup_lo_2642 = {dataGroup_lo_hi_2642, dataGroup_lo_lo_2642};
  wire [2047:0] dataGroup_hi_2642 = {dataGroup_hi_hi_2642, dataGroup_hi_lo_2642};
  wire [15:0]   dataGroup_18_46 = dataGroup_lo_2642[1455:1440];
  wire [2047:0] dataGroup_lo_2643 = {dataGroup_lo_hi_2643, dataGroup_lo_lo_2643};
  wire [2047:0] dataGroup_hi_2643 = {dataGroup_hi_hi_2643, dataGroup_hi_lo_2643};
  wire [15:0]   dataGroup_19_46 = dataGroup_lo_2643[1535:1520];
  wire [2047:0] dataGroup_lo_2644 = {dataGroup_lo_hi_2644, dataGroup_lo_lo_2644};
  wire [2047:0] dataGroup_hi_2644 = {dataGroup_hi_hi_2644, dataGroup_hi_lo_2644};
  wire [15:0]   dataGroup_20_46 = dataGroup_lo_2644[1615:1600];
  wire [2047:0] dataGroup_lo_2645 = {dataGroup_lo_hi_2645, dataGroup_lo_lo_2645};
  wire [2047:0] dataGroup_hi_2645 = {dataGroup_hi_hi_2645, dataGroup_hi_lo_2645};
  wire [15:0]   dataGroup_21_46 = dataGroup_lo_2645[1695:1680];
  wire [2047:0] dataGroup_lo_2646 = {dataGroup_lo_hi_2646, dataGroup_lo_lo_2646};
  wire [2047:0] dataGroup_hi_2646 = {dataGroup_hi_hi_2646, dataGroup_hi_lo_2646};
  wire [15:0]   dataGroup_22_46 = dataGroup_lo_2646[1775:1760];
  wire [2047:0] dataGroup_lo_2647 = {dataGroup_lo_hi_2647, dataGroup_lo_lo_2647};
  wire [2047:0] dataGroup_hi_2647 = {dataGroup_hi_hi_2647, dataGroup_hi_lo_2647};
  wire [15:0]   dataGroup_23_46 = dataGroup_lo_2647[1855:1840];
  wire [2047:0] dataGroup_lo_2648 = {dataGroup_lo_hi_2648, dataGroup_lo_lo_2648};
  wire [2047:0] dataGroup_hi_2648 = {dataGroup_hi_hi_2648, dataGroup_hi_lo_2648};
  wire [15:0]   dataGroup_24_46 = dataGroup_lo_2648[1935:1920];
  wire [2047:0] dataGroup_lo_2649 = {dataGroup_lo_hi_2649, dataGroup_lo_lo_2649};
  wire [2047:0] dataGroup_hi_2649 = {dataGroup_hi_hi_2649, dataGroup_hi_lo_2649};
  wire [15:0]   dataGroup_25_46 = dataGroup_lo_2649[2015:2000];
  wire [2047:0] dataGroup_lo_2650 = {dataGroup_lo_hi_2650, dataGroup_lo_lo_2650};
  wire [2047:0] dataGroup_hi_2650 = {dataGroup_hi_hi_2650, dataGroup_hi_lo_2650};
  wire [15:0]   dataGroup_26_46 = dataGroup_hi_2650[47:32];
  wire [2047:0] dataGroup_lo_2651 = {dataGroup_lo_hi_2651, dataGroup_lo_lo_2651};
  wire [2047:0] dataGroup_hi_2651 = {dataGroup_hi_hi_2651, dataGroup_hi_lo_2651};
  wire [15:0]   dataGroup_27_46 = dataGroup_hi_2651[127:112];
  wire [2047:0] dataGroup_lo_2652 = {dataGroup_lo_hi_2652, dataGroup_lo_lo_2652};
  wire [2047:0] dataGroup_hi_2652 = {dataGroup_hi_hi_2652, dataGroup_hi_lo_2652};
  wire [15:0]   dataGroup_28_46 = dataGroup_hi_2652[207:192];
  wire [2047:0] dataGroup_lo_2653 = {dataGroup_lo_hi_2653, dataGroup_lo_lo_2653};
  wire [2047:0] dataGroup_hi_2653 = {dataGroup_hi_hi_2653, dataGroup_hi_lo_2653};
  wire [15:0]   dataGroup_29_46 = dataGroup_hi_2653[287:272];
  wire [2047:0] dataGroup_lo_2654 = {dataGroup_lo_hi_2654, dataGroup_lo_lo_2654};
  wire [2047:0] dataGroup_hi_2654 = {dataGroup_hi_hi_2654, dataGroup_hi_lo_2654};
  wire [15:0]   dataGroup_30_46 = dataGroup_hi_2654[367:352];
  wire [2047:0] dataGroup_lo_2655 = {dataGroup_lo_hi_2655, dataGroup_lo_lo_2655};
  wire [2047:0] dataGroup_hi_2655 = {dataGroup_hi_hi_2655, dataGroup_hi_lo_2655};
  wire [15:0]   dataGroup_31_46 = dataGroup_hi_2655[447:432];
  wire [31:0]   res_lo_lo_lo_lo_46 = {dataGroup_1_46, dataGroup_0_46};
  wire [31:0]   res_lo_lo_lo_hi_46 = {dataGroup_3_46, dataGroup_2_46};
  wire [63:0]   res_lo_lo_lo_46 = {res_lo_lo_lo_hi_46, res_lo_lo_lo_lo_46};
  wire [31:0]   res_lo_lo_hi_lo_46 = {dataGroup_5_46, dataGroup_4_46};
  wire [31:0]   res_lo_lo_hi_hi_46 = {dataGroup_7_46, dataGroup_6_46};
  wire [63:0]   res_lo_lo_hi_46 = {res_lo_lo_hi_hi_46, res_lo_lo_hi_lo_46};
  wire [127:0]  res_lo_lo_46 = {res_lo_lo_hi_46, res_lo_lo_lo_46};
  wire [31:0]   res_lo_hi_lo_lo_46 = {dataGroup_9_46, dataGroup_8_46};
  wire [31:0]   res_lo_hi_lo_hi_46 = {dataGroup_11_46, dataGroup_10_46};
  wire [63:0]   res_lo_hi_lo_46 = {res_lo_hi_lo_hi_46, res_lo_hi_lo_lo_46};
  wire [31:0]   res_lo_hi_hi_lo_46 = {dataGroup_13_46, dataGroup_12_46};
  wire [31:0]   res_lo_hi_hi_hi_46 = {dataGroup_15_46, dataGroup_14_46};
  wire [63:0]   res_lo_hi_hi_46 = {res_lo_hi_hi_hi_46, res_lo_hi_hi_lo_46};
  wire [127:0]  res_lo_hi_46 = {res_lo_hi_hi_46, res_lo_hi_lo_46};
  wire [255:0]  res_lo_46 = {res_lo_hi_46, res_lo_lo_46};
  wire [31:0]   res_hi_lo_lo_lo_46 = {dataGroup_17_46, dataGroup_16_46};
  wire [31:0]   res_hi_lo_lo_hi_46 = {dataGroup_19_46, dataGroup_18_46};
  wire [63:0]   res_hi_lo_lo_46 = {res_hi_lo_lo_hi_46, res_hi_lo_lo_lo_46};
  wire [31:0]   res_hi_lo_hi_lo_46 = {dataGroup_21_46, dataGroup_20_46};
  wire [31:0]   res_hi_lo_hi_hi_46 = {dataGroup_23_46, dataGroup_22_46};
  wire [63:0]   res_hi_lo_hi_46 = {res_hi_lo_hi_hi_46, res_hi_lo_hi_lo_46};
  wire [127:0]  res_hi_lo_46 = {res_hi_lo_hi_46, res_hi_lo_lo_46};
  wire [31:0]   res_hi_hi_lo_lo_46 = {dataGroup_25_46, dataGroup_24_46};
  wire [31:0]   res_hi_hi_lo_hi_46 = {dataGroup_27_46, dataGroup_26_46};
  wire [63:0]   res_hi_hi_lo_46 = {res_hi_hi_lo_hi_46, res_hi_hi_lo_lo_46};
  wire [31:0]   res_hi_hi_hi_lo_46 = {dataGroup_29_46, dataGroup_28_46};
  wire [31:0]   res_hi_hi_hi_hi_46 = {dataGroup_31_46, dataGroup_30_46};
  wire [63:0]   res_hi_hi_hi_46 = {res_hi_hi_hi_hi_46, res_hi_hi_hi_lo_46};
  wire [127:0]  res_hi_hi_46 = {res_hi_hi_hi_46, res_hi_hi_lo_46};
  wire [255:0]  res_hi_46 = {res_hi_hi_46, res_hi_lo_46};
  wire [511:0]  res_96 = {res_hi_46, res_lo_46};
  wire [2047:0] dataGroup_lo_2656 = {dataGroup_lo_hi_2656, dataGroup_lo_lo_2656};
  wire [2047:0] dataGroup_hi_2656 = {dataGroup_hi_hi_2656, dataGroup_hi_lo_2656};
  wire [15:0]   dataGroup_0_47 = dataGroup_lo_2656[31:16];
  wire [2047:0] dataGroup_lo_2657 = {dataGroup_lo_hi_2657, dataGroup_lo_lo_2657};
  wire [2047:0] dataGroup_hi_2657 = {dataGroup_hi_hi_2657, dataGroup_hi_lo_2657};
  wire [15:0]   dataGroup_1_47 = dataGroup_lo_2657[111:96];
  wire [2047:0] dataGroup_lo_2658 = {dataGroup_lo_hi_2658, dataGroup_lo_lo_2658};
  wire [2047:0] dataGroup_hi_2658 = {dataGroup_hi_hi_2658, dataGroup_hi_lo_2658};
  wire [15:0]   dataGroup_2_47 = dataGroup_lo_2658[191:176];
  wire [2047:0] dataGroup_lo_2659 = {dataGroup_lo_hi_2659, dataGroup_lo_lo_2659};
  wire [2047:0] dataGroup_hi_2659 = {dataGroup_hi_hi_2659, dataGroup_hi_lo_2659};
  wire [15:0]   dataGroup_3_47 = dataGroup_lo_2659[271:256];
  wire [2047:0] dataGroup_lo_2660 = {dataGroup_lo_hi_2660, dataGroup_lo_lo_2660};
  wire [2047:0] dataGroup_hi_2660 = {dataGroup_hi_hi_2660, dataGroup_hi_lo_2660};
  wire [15:0]   dataGroup_4_47 = dataGroup_lo_2660[351:336];
  wire [2047:0] dataGroup_lo_2661 = {dataGroup_lo_hi_2661, dataGroup_lo_lo_2661};
  wire [2047:0] dataGroup_hi_2661 = {dataGroup_hi_hi_2661, dataGroup_hi_lo_2661};
  wire [15:0]   dataGroup_5_47 = dataGroup_lo_2661[431:416];
  wire [2047:0] dataGroup_lo_2662 = {dataGroup_lo_hi_2662, dataGroup_lo_lo_2662};
  wire [2047:0] dataGroup_hi_2662 = {dataGroup_hi_hi_2662, dataGroup_hi_lo_2662};
  wire [15:0]   dataGroup_6_47 = dataGroup_lo_2662[511:496];
  wire [2047:0] dataGroup_lo_2663 = {dataGroup_lo_hi_2663, dataGroup_lo_lo_2663};
  wire [2047:0] dataGroup_hi_2663 = {dataGroup_hi_hi_2663, dataGroup_hi_lo_2663};
  wire [15:0]   dataGroup_7_47 = dataGroup_lo_2663[591:576];
  wire [2047:0] dataGroup_lo_2664 = {dataGroup_lo_hi_2664, dataGroup_lo_lo_2664};
  wire [2047:0] dataGroup_hi_2664 = {dataGroup_hi_hi_2664, dataGroup_hi_lo_2664};
  wire [15:0]   dataGroup_8_47 = dataGroup_lo_2664[671:656];
  wire [2047:0] dataGroup_lo_2665 = {dataGroup_lo_hi_2665, dataGroup_lo_lo_2665};
  wire [2047:0] dataGroup_hi_2665 = {dataGroup_hi_hi_2665, dataGroup_hi_lo_2665};
  wire [15:0]   dataGroup_9_47 = dataGroup_lo_2665[751:736];
  wire [2047:0] dataGroup_lo_2666 = {dataGroup_lo_hi_2666, dataGroup_lo_lo_2666};
  wire [2047:0] dataGroup_hi_2666 = {dataGroup_hi_hi_2666, dataGroup_hi_lo_2666};
  wire [15:0]   dataGroup_10_47 = dataGroup_lo_2666[831:816];
  wire [2047:0] dataGroup_lo_2667 = {dataGroup_lo_hi_2667, dataGroup_lo_lo_2667};
  wire [2047:0] dataGroup_hi_2667 = {dataGroup_hi_hi_2667, dataGroup_hi_lo_2667};
  wire [15:0]   dataGroup_11_47 = dataGroup_lo_2667[911:896];
  wire [2047:0] dataGroup_lo_2668 = {dataGroup_lo_hi_2668, dataGroup_lo_lo_2668};
  wire [2047:0] dataGroup_hi_2668 = {dataGroup_hi_hi_2668, dataGroup_hi_lo_2668};
  wire [15:0]   dataGroup_12_47 = dataGroup_lo_2668[991:976];
  wire [2047:0] dataGroup_lo_2669 = {dataGroup_lo_hi_2669, dataGroup_lo_lo_2669};
  wire [2047:0] dataGroup_hi_2669 = {dataGroup_hi_hi_2669, dataGroup_hi_lo_2669};
  wire [15:0]   dataGroup_13_47 = dataGroup_lo_2669[1071:1056];
  wire [2047:0] dataGroup_lo_2670 = {dataGroup_lo_hi_2670, dataGroup_lo_lo_2670};
  wire [2047:0] dataGroup_hi_2670 = {dataGroup_hi_hi_2670, dataGroup_hi_lo_2670};
  wire [15:0]   dataGroup_14_47 = dataGroup_lo_2670[1151:1136];
  wire [2047:0] dataGroup_lo_2671 = {dataGroup_lo_hi_2671, dataGroup_lo_lo_2671};
  wire [2047:0] dataGroup_hi_2671 = {dataGroup_hi_hi_2671, dataGroup_hi_lo_2671};
  wire [15:0]   dataGroup_15_47 = dataGroup_lo_2671[1231:1216];
  wire [2047:0] dataGroup_lo_2672 = {dataGroup_lo_hi_2672, dataGroup_lo_lo_2672};
  wire [2047:0] dataGroup_hi_2672 = {dataGroup_hi_hi_2672, dataGroup_hi_lo_2672};
  wire [15:0]   dataGroup_16_47 = dataGroup_lo_2672[1311:1296];
  wire [2047:0] dataGroup_lo_2673 = {dataGroup_lo_hi_2673, dataGroup_lo_lo_2673};
  wire [2047:0] dataGroup_hi_2673 = {dataGroup_hi_hi_2673, dataGroup_hi_lo_2673};
  wire [15:0]   dataGroup_17_47 = dataGroup_lo_2673[1391:1376];
  wire [2047:0] dataGroup_lo_2674 = {dataGroup_lo_hi_2674, dataGroup_lo_lo_2674};
  wire [2047:0] dataGroup_hi_2674 = {dataGroup_hi_hi_2674, dataGroup_hi_lo_2674};
  wire [15:0]   dataGroup_18_47 = dataGroup_lo_2674[1471:1456];
  wire [2047:0] dataGroup_lo_2675 = {dataGroup_lo_hi_2675, dataGroup_lo_lo_2675};
  wire [2047:0] dataGroup_hi_2675 = {dataGroup_hi_hi_2675, dataGroup_hi_lo_2675};
  wire [15:0]   dataGroup_19_47 = dataGroup_lo_2675[1551:1536];
  wire [2047:0] dataGroup_lo_2676 = {dataGroup_lo_hi_2676, dataGroup_lo_lo_2676};
  wire [2047:0] dataGroup_hi_2676 = {dataGroup_hi_hi_2676, dataGroup_hi_lo_2676};
  wire [15:0]   dataGroup_20_47 = dataGroup_lo_2676[1631:1616];
  wire [2047:0] dataGroup_lo_2677 = {dataGroup_lo_hi_2677, dataGroup_lo_lo_2677};
  wire [2047:0] dataGroup_hi_2677 = {dataGroup_hi_hi_2677, dataGroup_hi_lo_2677};
  wire [15:0]   dataGroup_21_47 = dataGroup_lo_2677[1711:1696];
  wire [2047:0] dataGroup_lo_2678 = {dataGroup_lo_hi_2678, dataGroup_lo_lo_2678};
  wire [2047:0] dataGroup_hi_2678 = {dataGroup_hi_hi_2678, dataGroup_hi_lo_2678};
  wire [15:0]   dataGroup_22_47 = dataGroup_lo_2678[1791:1776];
  wire [2047:0] dataGroup_lo_2679 = {dataGroup_lo_hi_2679, dataGroup_lo_lo_2679};
  wire [2047:0] dataGroup_hi_2679 = {dataGroup_hi_hi_2679, dataGroup_hi_lo_2679};
  wire [15:0]   dataGroup_23_47 = dataGroup_lo_2679[1871:1856];
  wire [2047:0] dataGroup_lo_2680 = {dataGroup_lo_hi_2680, dataGroup_lo_lo_2680};
  wire [2047:0] dataGroup_hi_2680 = {dataGroup_hi_hi_2680, dataGroup_hi_lo_2680};
  wire [15:0]   dataGroup_24_47 = dataGroup_lo_2680[1951:1936];
  wire [2047:0] dataGroup_lo_2681 = {dataGroup_lo_hi_2681, dataGroup_lo_lo_2681};
  wire [2047:0] dataGroup_hi_2681 = {dataGroup_hi_hi_2681, dataGroup_hi_lo_2681};
  wire [15:0]   dataGroup_25_47 = dataGroup_lo_2681[2031:2016];
  wire [2047:0] dataGroup_lo_2682 = {dataGroup_lo_hi_2682, dataGroup_lo_lo_2682};
  wire [2047:0] dataGroup_hi_2682 = {dataGroup_hi_hi_2682, dataGroup_hi_lo_2682};
  wire [15:0]   dataGroup_26_47 = dataGroup_hi_2682[63:48];
  wire [2047:0] dataGroup_lo_2683 = {dataGroup_lo_hi_2683, dataGroup_lo_lo_2683};
  wire [2047:0] dataGroup_hi_2683 = {dataGroup_hi_hi_2683, dataGroup_hi_lo_2683};
  wire [15:0]   dataGroup_27_47 = dataGroup_hi_2683[143:128];
  wire [2047:0] dataGroup_lo_2684 = {dataGroup_lo_hi_2684, dataGroup_lo_lo_2684};
  wire [2047:0] dataGroup_hi_2684 = {dataGroup_hi_hi_2684, dataGroup_hi_lo_2684};
  wire [15:0]   dataGroup_28_47 = dataGroup_hi_2684[223:208];
  wire [2047:0] dataGroup_lo_2685 = {dataGroup_lo_hi_2685, dataGroup_lo_lo_2685};
  wire [2047:0] dataGroup_hi_2685 = {dataGroup_hi_hi_2685, dataGroup_hi_lo_2685};
  wire [15:0]   dataGroup_29_47 = dataGroup_hi_2685[303:288];
  wire [2047:0] dataGroup_lo_2686 = {dataGroup_lo_hi_2686, dataGroup_lo_lo_2686};
  wire [2047:0] dataGroup_hi_2686 = {dataGroup_hi_hi_2686, dataGroup_hi_lo_2686};
  wire [15:0]   dataGroup_30_47 = dataGroup_hi_2686[383:368];
  wire [2047:0] dataGroup_lo_2687 = {dataGroup_lo_hi_2687, dataGroup_lo_lo_2687};
  wire [2047:0] dataGroup_hi_2687 = {dataGroup_hi_hi_2687, dataGroup_hi_lo_2687};
  wire [15:0]   dataGroup_31_47 = dataGroup_hi_2687[463:448];
  wire [31:0]   res_lo_lo_lo_lo_47 = {dataGroup_1_47, dataGroup_0_47};
  wire [31:0]   res_lo_lo_lo_hi_47 = {dataGroup_3_47, dataGroup_2_47};
  wire [63:0]   res_lo_lo_lo_47 = {res_lo_lo_lo_hi_47, res_lo_lo_lo_lo_47};
  wire [31:0]   res_lo_lo_hi_lo_47 = {dataGroup_5_47, dataGroup_4_47};
  wire [31:0]   res_lo_lo_hi_hi_47 = {dataGroup_7_47, dataGroup_6_47};
  wire [63:0]   res_lo_lo_hi_47 = {res_lo_lo_hi_hi_47, res_lo_lo_hi_lo_47};
  wire [127:0]  res_lo_lo_47 = {res_lo_lo_hi_47, res_lo_lo_lo_47};
  wire [31:0]   res_lo_hi_lo_lo_47 = {dataGroup_9_47, dataGroup_8_47};
  wire [31:0]   res_lo_hi_lo_hi_47 = {dataGroup_11_47, dataGroup_10_47};
  wire [63:0]   res_lo_hi_lo_47 = {res_lo_hi_lo_hi_47, res_lo_hi_lo_lo_47};
  wire [31:0]   res_lo_hi_hi_lo_47 = {dataGroup_13_47, dataGroup_12_47};
  wire [31:0]   res_lo_hi_hi_hi_47 = {dataGroup_15_47, dataGroup_14_47};
  wire [63:0]   res_lo_hi_hi_47 = {res_lo_hi_hi_hi_47, res_lo_hi_hi_lo_47};
  wire [127:0]  res_lo_hi_47 = {res_lo_hi_hi_47, res_lo_hi_lo_47};
  wire [255:0]  res_lo_47 = {res_lo_hi_47, res_lo_lo_47};
  wire [31:0]   res_hi_lo_lo_lo_47 = {dataGroup_17_47, dataGroup_16_47};
  wire [31:0]   res_hi_lo_lo_hi_47 = {dataGroup_19_47, dataGroup_18_47};
  wire [63:0]   res_hi_lo_lo_47 = {res_hi_lo_lo_hi_47, res_hi_lo_lo_lo_47};
  wire [31:0]   res_hi_lo_hi_lo_47 = {dataGroup_21_47, dataGroup_20_47};
  wire [31:0]   res_hi_lo_hi_hi_47 = {dataGroup_23_47, dataGroup_22_47};
  wire [63:0]   res_hi_lo_hi_47 = {res_hi_lo_hi_hi_47, res_hi_lo_hi_lo_47};
  wire [127:0]  res_hi_lo_47 = {res_hi_lo_hi_47, res_hi_lo_lo_47};
  wire [31:0]   res_hi_hi_lo_lo_47 = {dataGroup_25_47, dataGroup_24_47};
  wire [31:0]   res_hi_hi_lo_hi_47 = {dataGroup_27_47, dataGroup_26_47};
  wire [63:0]   res_hi_hi_lo_47 = {res_hi_hi_lo_hi_47, res_hi_hi_lo_lo_47};
  wire [31:0]   res_hi_hi_hi_lo_47 = {dataGroup_29_47, dataGroup_28_47};
  wire [31:0]   res_hi_hi_hi_hi_47 = {dataGroup_31_47, dataGroup_30_47};
  wire [63:0]   res_hi_hi_hi_47 = {res_hi_hi_hi_hi_47, res_hi_hi_hi_lo_47};
  wire [127:0]  res_hi_hi_47 = {res_hi_hi_hi_47, res_hi_hi_lo_47};
  wire [255:0]  res_hi_47 = {res_hi_hi_47, res_hi_lo_47};
  wire [511:0]  res_97 = {res_hi_47, res_lo_47};
  wire [2047:0] dataGroup_lo_2688 = {dataGroup_lo_hi_2688, dataGroup_lo_lo_2688};
  wire [2047:0] dataGroup_hi_2688 = {dataGroup_hi_hi_2688, dataGroup_hi_lo_2688};
  wire [15:0]   dataGroup_0_48 = dataGroup_lo_2688[47:32];
  wire [2047:0] dataGroup_lo_2689 = {dataGroup_lo_hi_2689, dataGroup_lo_lo_2689};
  wire [2047:0] dataGroup_hi_2689 = {dataGroup_hi_hi_2689, dataGroup_hi_lo_2689};
  wire [15:0]   dataGroup_1_48 = dataGroup_lo_2689[127:112];
  wire [2047:0] dataGroup_lo_2690 = {dataGroup_lo_hi_2690, dataGroup_lo_lo_2690};
  wire [2047:0] dataGroup_hi_2690 = {dataGroup_hi_hi_2690, dataGroup_hi_lo_2690};
  wire [15:0]   dataGroup_2_48 = dataGroup_lo_2690[207:192];
  wire [2047:0] dataGroup_lo_2691 = {dataGroup_lo_hi_2691, dataGroup_lo_lo_2691};
  wire [2047:0] dataGroup_hi_2691 = {dataGroup_hi_hi_2691, dataGroup_hi_lo_2691};
  wire [15:0]   dataGroup_3_48 = dataGroup_lo_2691[287:272];
  wire [2047:0] dataGroup_lo_2692 = {dataGroup_lo_hi_2692, dataGroup_lo_lo_2692};
  wire [2047:0] dataGroup_hi_2692 = {dataGroup_hi_hi_2692, dataGroup_hi_lo_2692};
  wire [15:0]   dataGroup_4_48 = dataGroup_lo_2692[367:352];
  wire [2047:0] dataGroup_lo_2693 = {dataGroup_lo_hi_2693, dataGroup_lo_lo_2693};
  wire [2047:0] dataGroup_hi_2693 = {dataGroup_hi_hi_2693, dataGroup_hi_lo_2693};
  wire [15:0]   dataGroup_5_48 = dataGroup_lo_2693[447:432];
  wire [2047:0] dataGroup_lo_2694 = {dataGroup_lo_hi_2694, dataGroup_lo_lo_2694};
  wire [2047:0] dataGroup_hi_2694 = {dataGroup_hi_hi_2694, dataGroup_hi_lo_2694};
  wire [15:0]   dataGroup_6_48 = dataGroup_lo_2694[527:512];
  wire [2047:0] dataGroup_lo_2695 = {dataGroup_lo_hi_2695, dataGroup_lo_lo_2695};
  wire [2047:0] dataGroup_hi_2695 = {dataGroup_hi_hi_2695, dataGroup_hi_lo_2695};
  wire [15:0]   dataGroup_7_48 = dataGroup_lo_2695[607:592];
  wire [2047:0] dataGroup_lo_2696 = {dataGroup_lo_hi_2696, dataGroup_lo_lo_2696};
  wire [2047:0] dataGroup_hi_2696 = {dataGroup_hi_hi_2696, dataGroup_hi_lo_2696};
  wire [15:0]   dataGroup_8_48 = dataGroup_lo_2696[687:672];
  wire [2047:0] dataGroup_lo_2697 = {dataGroup_lo_hi_2697, dataGroup_lo_lo_2697};
  wire [2047:0] dataGroup_hi_2697 = {dataGroup_hi_hi_2697, dataGroup_hi_lo_2697};
  wire [15:0]   dataGroup_9_48 = dataGroup_lo_2697[767:752];
  wire [2047:0] dataGroup_lo_2698 = {dataGroup_lo_hi_2698, dataGroup_lo_lo_2698};
  wire [2047:0] dataGroup_hi_2698 = {dataGroup_hi_hi_2698, dataGroup_hi_lo_2698};
  wire [15:0]   dataGroup_10_48 = dataGroup_lo_2698[847:832];
  wire [2047:0] dataGroup_lo_2699 = {dataGroup_lo_hi_2699, dataGroup_lo_lo_2699};
  wire [2047:0] dataGroup_hi_2699 = {dataGroup_hi_hi_2699, dataGroup_hi_lo_2699};
  wire [15:0]   dataGroup_11_48 = dataGroup_lo_2699[927:912];
  wire [2047:0] dataGroup_lo_2700 = {dataGroup_lo_hi_2700, dataGroup_lo_lo_2700};
  wire [2047:0] dataGroup_hi_2700 = {dataGroup_hi_hi_2700, dataGroup_hi_lo_2700};
  wire [15:0]   dataGroup_12_48 = dataGroup_lo_2700[1007:992];
  wire [2047:0] dataGroup_lo_2701 = {dataGroup_lo_hi_2701, dataGroup_lo_lo_2701};
  wire [2047:0] dataGroup_hi_2701 = {dataGroup_hi_hi_2701, dataGroup_hi_lo_2701};
  wire [15:0]   dataGroup_13_48 = dataGroup_lo_2701[1087:1072];
  wire [2047:0] dataGroup_lo_2702 = {dataGroup_lo_hi_2702, dataGroup_lo_lo_2702};
  wire [2047:0] dataGroup_hi_2702 = {dataGroup_hi_hi_2702, dataGroup_hi_lo_2702};
  wire [15:0]   dataGroup_14_48 = dataGroup_lo_2702[1167:1152];
  wire [2047:0] dataGroup_lo_2703 = {dataGroup_lo_hi_2703, dataGroup_lo_lo_2703};
  wire [2047:0] dataGroup_hi_2703 = {dataGroup_hi_hi_2703, dataGroup_hi_lo_2703};
  wire [15:0]   dataGroup_15_48 = dataGroup_lo_2703[1247:1232];
  wire [2047:0] dataGroup_lo_2704 = {dataGroup_lo_hi_2704, dataGroup_lo_lo_2704};
  wire [2047:0] dataGroup_hi_2704 = {dataGroup_hi_hi_2704, dataGroup_hi_lo_2704};
  wire [15:0]   dataGroup_16_48 = dataGroup_lo_2704[1327:1312];
  wire [2047:0] dataGroup_lo_2705 = {dataGroup_lo_hi_2705, dataGroup_lo_lo_2705};
  wire [2047:0] dataGroup_hi_2705 = {dataGroup_hi_hi_2705, dataGroup_hi_lo_2705};
  wire [15:0]   dataGroup_17_48 = dataGroup_lo_2705[1407:1392];
  wire [2047:0] dataGroup_lo_2706 = {dataGroup_lo_hi_2706, dataGroup_lo_lo_2706};
  wire [2047:0] dataGroup_hi_2706 = {dataGroup_hi_hi_2706, dataGroup_hi_lo_2706};
  wire [15:0]   dataGroup_18_48 = dataGroup_lo_2706[1487:1472];
  wire [2047:0] dataGroup_lo_2707 = {dataGroup_lo_hi_2707, dataGroup_lo_lo_2707};
  wire [2047:0] dataGroup_hi_2707 = {dataGroup_hi_hi_2707, dataGroup_hi_lo_2707};
  wire [15:0]   dataGroup_19_48 = dataGroup_lo_2707[1567:1552];
  wire [2047:0] dataGroup_lo_2708 = {dataGroup_lo_hi_2708, dataGroup_lo_lo_2708};
  wire [2047:0] dataGroup_hi_2708 = {dataGroup_hi_hi_2708, dataGroup_hi_lo_2708};
  wire [15:0]   dataGroup_20_48 = dataGroup_lo_2708[1647:1632];
  wire [2047:0] dataGroup_lo_2709 = {dataGroup_lo_hi_2709, dataGroup_lo_lo_2709};
  wire [2047:0] dataGroup_hi_2709 = {dataGroup_hi_hi_2709, dataGroup_hi_lo_2709};
  wire [15:0]   dataGroup_21_48 = dataGroup_lo_2709[1727:1712];
  wire [2047:0] dataGroup_lo_2710 = {dataGroup_lo_hi_2710, dataGroup_lo_lo_2710};
  wire [2047:0] dataGroup_hi_2710 = {dataGroup_hi_hi_2710, dataGroup_hi_lo_2710};
  wire [15:0]   dataGroup_22_48 = dataGroup_lo_2710[1807:1792];
  wire [2047:0] dataGroup_lo_2711 = {dataGroup_lo_hi_2711, dataGroup_lo_lo_2711};
  wire [2047:0] dataGroup_hi_2711 = {dataGroup_hi_hi_2711, dataGroup_hi_lo_2711};
  wire [15:0]   dataGroup_23_48 = dataGroup_lo_2711[1887:1872];
  wire [2047:0] dataGroup_lo_2712 = {dataGroup_lo_hi_2712, dataGroup_lo_lo_2712};
  wire [2047:0] dataGroup_hi_2712 = {dataGroup_hi_hi_2712, dataGroup_hi_lo_2712};
  wire [15:0]   dataGroup_24_48 = dataGroup_lo_2712[1967:1952];
  wire [2047:0] dataGroup_lo_2713 = {dataGroup_lo_hi_2713, dataGroup_lo_lo_2713};
  wire [2047:0] dataGroup_hi_2713 = {dataGroup_hi_hi_2713, dataGroup_hi_lo_2713};
  wire [15:0]   dataGroup_25_48 = dataGroup_lo_2713[2047:2032];
  wire [2047:0] dataGroup_lo_2714 = {dataGroup_lo_hi_2714, dataGroup_lo_lo_2714};
  wire [2047:0] dataGroup_hi_2714 = {dataGroup_hi_hi_2714, dataGroup_hi_lo_2714};
  wire [15:0]   dataGroup_26_48 = dataGroup_hi_2714[79:64];
  wire [2047:0] dataGroup_lo_2715 = {dataGroup_lo_hi_2715, dataGroup_lo_lo_2715};
  wire [2047:0] dataGroup_hi_2715 = {dataGroup_hi_hi_2715, dataGroup_hi_lo_2715};
  wire [15:0]   dataGroup_27_48 = dataGroup_hi_2715[159:144];
  wire [2047:0] dataGroup_lo_2716 = {dataGroup_lo_hi_2716, dataGroup_lo_lo_2716};
  wire [2047:0] dataGroup_hi_2716 = {dataGroup_hi_hi_2716, dataGroup_hi_lo_2716};
  wire [15:0]   dataGroup_28_48 = dataGroup_hi_2716[239:224];
  wire [2047:0] dataGroup_lo_2717 = {dataGroup_lo_hi_2717, dataGroup_lo_lo_2717};
  wire [2047:0] dataGroup_hi_2717 = {dataGroup_hi_hi_2717, dataGroup_hi_lo_2717};
  wire [15:0]   dataGroup_29_48 = dataGroup_hi_2717[319:304];
  wire [2047:0] dataGroup_lo_2718 = {dataGroup_lo_hi_2718, dataGroup_lo_lo_2718};
  wire [2047:0] dataGroup_hi_2718 = {dataGroup_hi_hi_2718, dataGroup_hi_lo_2718};
  wire [15:0]   dataGroup_30_48 = dataGroup_hi_2718[399:384];
  wire [2047:0] dataGroup_lo_2719 = {dataGroup_lo_hi_2719, dataGroup_lo_lo_2719};
  wire [2047:0] dataGroup_hi_2719 = {dataGroup_hi_hi_2719, dataGroup_hi_lo_2719};
  wire [15:0]   dataGroup_31_48 = dataGroup_hi_2719[479:464];
  wire [31:0]   res_lo_lo_lo_lo_48 = {dataGroup_1_48, dataGroup_0_48};
  wire [31:0]   res_lo_lo_lo_hi_48 = {dataGroup_3_48, dataGroup_2_48};
  wire [63:0]   res_lo_lo_lo_48 = {res_lo_lo_lo_hi_48, res_lo_lo_lo_lo_48};
  wire [31:0]   res_lo_lo_hi_lo_48 = {dataGroup_5_48, dataGroup_4_48};
  wire [31:0]   res_lo_lo_hi_hi_48 = {dataGroup_7_48, dataGroup_6_48};
  wire [63:0]   res_lo_lo_hi_48 = {res_lo_lo_hi_hi_48, res_lo_lo_hi_lo_48};
  wire [127:0]  res_lo_lo_48 = {res_lo_lo_hi_48, res_lo_lo_lo_48};
  wire [31:0]   res_lo_hi_lo_lo_48 = {dataGroup_9_48, dataGroup_8_48};
  wire [31:0]   res_lo_hi_lo_hi_48 = {dataGroup_11_48, dataGroup_10_48};
  wire [63:0]   res_lo_hi_lo_48 = {res_lo_hi_lo_hi_48, res_lo_hi_lo_lo_48};
  wire [31:0]   res_lo_hi_hi_lo_48 = {dataGroup_13_48, dataGroup_12_48};
  wire [31:0]   res_lo_hi_hi_hi_48 = {dataGroup_15_48, dataGroup_14_48};
  wire [63:0]   res_lo_hi_hi_48 = {res_lo_hi_hi_hi_48, res_lo_hi_hi_lo_48};
  wire [127:0]  res_lo_hi_48 = {res_lo_hi_hi_48, res_lo_hi_lo_48};
  wire [255:0]  res_lo_48 = {res_lo_hi_48, res_lo_lo_48};
  wire [31:0]   res_hi_lo_lo_lo_48 = {dataGroup_17_48, dataGroup_16_48};
  wire [31:0]   res_hi_lo_lo_hi_48 = {dataGroup_19_48, dataGroup_18_48};
  wire [63:0]   res_hi_lo_lo_48 = {res_hi_lo_lo_hi_48, res_hi_lo_lo_lo_48};
  wire [31:0]   res_hi_lo_hi_lo_48 = {dataGroup_21_48, dataGroup_20_48};
  wire [31:0]   res_hi_lo_hi_hi_48 = {dataGroup_23_48, dataGroup_22_48};
  wire [63:0]   res_hi_lo_hi_48 = {res_hi_lo_hi_hi_48, res_hi_lo_hi_lo_48};
  wire [127:0]  res_hi_lo_48 = {res_hi_lo_hi_48, res_hi_lo_lo_48};
  wire [31:0]   res_hi_hi_lo_lo_48 = {dataGroup_25_48, dataGroup_24_48};
  wire [31:0]   res_hi_hi_lo_hi_48 = {dataGroup_27_48, dataGroup_26_48};
  wire [63:0]   res_hi_hi_lo_48 = {res_hi_hi_lo_hi_48, res_hi_hi_lo_lo_48};
  wire [31:0]   res_hi_hi_hi_lo_48 = {dataGroup_29_48, dataGroup_28_48};
  wire [31:0]   res_hi_hi_hi_hi_48 = {dataGroup_31_48, dataGroup_30_48};
  wire [63:0]   res_hi_hi_hi_48 = {res_hi_hi_hi_hi_48, res_hi_hi_hi_lo_48};
  wire [127:0]  res_hi_hi_48 = {res_hi_hi_hi_48, res_hi_hi_lo_48};
  wire [255:0]  res_hi_48 = {res_hi_hi_48, res_hi_lo_48};
  wire [511:0]  res_98 = {res_hi_48, res_lo_48};
  wire [2047:0] dataGroup_lo_2720 = {dataGroup_lo_hi_2720, dataGroup_lo_lo_2720};
  wire [2047:0] dataGroup_hi_2720 = {dataGroup_hi_hi_2720, dataGroup_hi_lo_2720};
  wire [15:0]   dataGroup_0_49 = dataGroup_lo_2720[63:48];
  wire [2047:0] dataGroup_lo_2721 = {dataGroup_lo_hi_2721, dataGroup_lo_lo_2721};
  wire [2047:0] dataGroup_hi_2721 = {dataGroup_hi_hi_2721, dataGroup_hi_lo_2721};
  wire [15:0]   dataGroup_1_49 = dataGroup_lo_2721[143:128];
  wire [2047:0] dataGroup_lo_2722 = {dataGroup_lo_hi_2722, dataGroup_lo_lo_2722};
  wire [2047:0] dataGroup_hi_2722 = {dataGroup_hi_hi_2722, dataGroup_hi_lo_2722};
  wire [15:0]   dataGroup_2_49 = dataGroup_lo_2722[223:208];
  wire [2047:0] dataGroup_lo_2723 = {dataGroup_lo_hi_2723, dataGroup_lo_lo_2723};
  wire [2047:0] dataGroup_hi_2723 = {dataGroup_hi_hi_2723, dataGroup_hi_lo_2723};
  wire [15:0]   dataGroup_3_49 = dataGroup_lo_2723[303:288];
  wire [2047:0] dataGroup_lo_2724 = {dataGroup_lo_hi_2724, dataGroup_lo_lo_2724};
  wire [2047:0] dataGroup_hi_2724 = {dataGroup_hi_hi_2724, dataGroup_hi_lo_2724};
  wire [15:0]   dataGroup_4_49 = dataGroup_lo_2724[383:368];
  wire [2047:0] dataGroup_lo_2725 = {dataGroup_lo_hi_2725, dataGroup_lo_lo_2725};
  wire [2047:0] dataGroup_hi_2725 = {dataGroup_hi_hi_2725, dataGroup_hi_lo_2725};
  wire [15:0]   dataGroup_5_49 = dataGroup_lo_2725[463:448];
  wire [2047:0] dataGroup_lo_2726 = {dataGroup_lo_hi_2726, dataGroup_lo_lo_2726};
  wire [2047:0] dataGroup_hi_2726 = {dataGroup_hi_hi_2726, dataGroup_hi_lo_2726};
  wire [15:0]   dataGroup_6_49 = dataGroup_lo_2726[543:528];
  wire [2047:0] dataGroup_lo_2727 = {dataGroup_lo_hi_2727, dataGroup_lo_lo_2727};
  wire [2047:0] dataGroup_hi_2727 = {dataGroup_hi_hi_2727, dataGroup_hi_lo_2727};
  wire [15:0]   dataGroup_7_49 = dataGroup_lo_2727[623:608];
  wire [2047:0] dataGroup_lo_2728 = {dataGroup_lo_hi_2728, dataGroup_lo_lo_2728};
  wire [2047:0] dataGroup_hi_2728 = {dataGroup_hi_hi_2728, dataGroup_hi_lo_2728};
  wire [15:0]   dataGroup_8_49 = dataGroup_lo_2728[703:688];
  wire [2047:0] dataGroup_lo_2729 = {dataGroup_lo_hi_2729, dataGroup_lo_lo_2729};
  wire [2047:0] dataGroup_hi_2729 = {dataGroup_hi_hi_2729, dataGroup_hi_lo_2729};
  wire [15:0]   dataGroup_9_49 = dataGroup_lo_2729[783:768];
  wire [2047:0] dataGroup_lo_2730 = {dataGroup_lo_hi_2730, dataGroup_lo_lo_2730};
  wire [2047:0] dataGroup_hi_2730 = {dataGroup_hi_hi_2730, dataGroup_hi_lo_2730};
  wire [15:0]   dataGroup_10_49 = dataGroup_lo_2730[863:848];
  wire [2047:0] dataGroup_lo_2731 = {dataGroup_lo_hi_2731, dataGroup_lo_lo_2731};
  wire [2047:0] dataGroup_hi_2731 = {dataGroup_hi_hi_2731, dataGroup_hi_lo_2731};
  wire [15:0]   dataGroup_11_49 = dataGroup_lo_2731[943:928];
  wire [2047:0] dataGroup_lo_2732 = {dataGroup_lo_hi_2732, dataGroup_lo_lo_2732};
  wire [2047:0] dataGroup_hi_2732 = {dataGroup_hi_hi_2732, dataGroup_hi_lo_2732};
  wire [15:0]   dataGroup_12_49 = dataGroup_lo_2732[1023:1008];
  wire [2047:0] dataGroup_lo_2733 = {dataGroup_lo_hi_2733, dataGroup_lo_lo_2733};
  wire [2047:0] dataGroup_hi_2733 = {dataGroup_hi_hi_2733, dataGroup_hi_lo_2733};
  wire [15:0]   dataGroup_13_49 = dataGroup_lo_2733[1103:1088];
  wire [2047:0] dataGroup_lo_2734 = {dataGroup_lo_hi_2734, dataGroup_lo_lo_2734};
  wire [2047:0] dataGroup_hi_2734 = {dataGroup_hi_hi_2734, dataGroup_hi_lo_2734};
  wire [15:0]   dataGroup_14_49 = dataGroup_lo_2734[1183:1168];
  wire [2047:0] dataGroup_lo_2735 = {dataGroup_lo_hi_2735, dataGroup_lo_lo_2735};
  wire [2047:0] dataGroup_hi_2735 = {dataGroup_hi_hi_2735, dataGroup_hi_lo_2735};
  wire [15:0]   dataGroup_15_49 = dataGroup_lo_2735[1263:1248];
  wire [2047:0] dataGroup_lo_2736 = {dataGroup_lo_hi_2736, dataGroup_lo_lo_2736};
  wire [2047:0] dataGroup_hi_2736 = {dataGroup_hi_hi_2736, dataGroup_hi_lo_2736};
  wire [15:0]   dataGroup_16_49 = dataGroup_lo_2736[1343:1328];
  wire [2047:0] dataGroup_lo_2737 = {dataGroup_lo_hi_2737, dataGroup_lo_lo_2737};
  wire [2047:0] dataGroup_hi_2737 = {dataGroup_hi_hi_2737, dataGroup_hi_lo_2737};
  wire [15:0]   dataGroup_17_49 = dataGroup_lo_2737[1423:1408];
  wire [2047:0] dataGroup_lo_2738 = {dataGroup_lo_hi_2738, dataGroup_lo_lo_2738};
  wire [2047:0] dataGroup_hi_2738 = {dataGroup_hi_hi_2738, dataGroup_hi_lo_2738};
  wire [15:0]   dataGroup_18_49 = dataGroup_lo_2738[1503:1488];
  wire [2047:0] dataGroup_lo_2739 = {dataGroup_lo_hi_2739, dataGroup_lo_lo_2739};
  wire [2047:0] dataGroup_hi_2739 = {dataGroup_hi_hi_2739, dataGroup_hi_lo_2739};
  wire [15:0]   dataGroup_19_49 = dataGroup_lo_2739[1583:1568];
  wire [2047:0] dataGroup_lo_2740 = {dataGroup_lo_hi_2740, dataGroup_lo_lo_2740};
  wire [2047:0] dataGroup_hi_2740 = {dataGroup_hi_hi_2740, dataGroup_hi_lo_2740};
  wire [15:0]   dataGroup_20_49 = dataGroup_lo_2740[1663:1648];
  wire [2047:0] dataGroup_lo_2741 = {dataGroup_lo_hi_2741, dataGroup_lo_lo_2741};
  wire [2047:0] dataGroup_hi_2741 = {dataGroup_hi_hi_2741, dataGroup_hi_lo_2741};
  wire [15:0]   dataGroup_21_49 = dataGroup_lo_2741[1743:1728];
  wire [2047:0] dataGroup_lo_2742 = {dataGroup_lo_hi_2742, dataGroup_lo_lo_2742};
  wire [2047:0] dataGroup_hi_2742 = {dataGroup_hi_hi_2742, dataGroup_hi_lo_2742};
  wire [15:0]   dataGroup_22_49 = dataGroup_lo_2742[1823:1808];
  wire [2047:0] dataGroup_lo_2743 = {dataGroup_lo_hi_2743, dataGroup_lo_lo_2743};
  wire [2047:0] dataGroup_hi_2743 = {dataGroup_hi_hi_2743, dataGroup_hi_lo_2743};
  wire [15:0]   dataGroup_23_49 = dataGroup_lo_2743[1903:1888];
  wire [2047:0] dataGroup_lo_2744 = {dataGroup_lo_hi_2744, dataGroup_lo_lo_2744};
  wire [2047:0] dataGroup_hi_2744 = {dataGroup_hi_hi_2744, dataGroup_hi_lo_2744};
  wire [15:0]   dataGroup_24_49 = dataGroup_lo_2744[1983:1968];
  wire [2047:0] dataGroup_lo_2745 = {dataGroup_lo_hi_2745, dataGroup_lo_lo_2745};
  wire [2047:0] dataGroup_hi_2745 = {dataGroup_hi_hi_2745, dataGroup_hi_lo_2745};
  wire [15:0]   dataGroup_25_49 = dataGroup_hi_2745[15:0];
  wire [2047:0] dataGroup_lo_2746 = {dataGroup_lo_hi_2746, dataGroup_lo_lo_2746};
  wire [2047:0] dataGroup_hi_2746 = {dataGroup_hi_hi_2746, dataGroup_hi_lo_2746};
  wire [15:0]   dataGroup_26_49 = dataGroup_hi_2746[95:80];
  wire [2047:0] dataGroup_lo_2747 = {dataGroup_lo_hi_2747, dataGroup_lo_lo_2747};
  wire [2047:0] dataGroup_hi_2747 = {dataGroup_hi_hi_2747, dataGroup_hi_lo_2747};
  wire [15:0]   dataGroup_27_49 = dataGroup_hi_2747[175:160];
  wire [2047:0] dataGroup_lo_2748 = {dataGroup_lo_hi_2748, dataGroup_lo_lo_2748};
  wire [2047:0] dataGroup_hi_2748 = {dataGroup_hi_hi_2748, dataGroup_hi_lo_2748};
  wire [15:0]   dataGroup_28_49 = dataGroup_hi_2748[255:240];
  wire [2047:0] dataGroup_lo_2749 = {dataGroup_lo_hi_2749, dataGroup_lo_lo_2749};
  wire [2047:0] dataGroup_hi_2749 = {dataGroup_hi_hi_2749, dataGroup_hi_lo_2749};
  wire [15:0]   dataGroup_29_49 = dataGroup_hi_2749[335:320];
  wire [2047:0] dataGroup_lo_2750 = {dataGroup_lo_hi_2750, dataGroup_lo_lo_2750};
  wire [2047:0] dataGroup_hi_2750 = {dataGroup_hi_hi_2750, dataGroup_hi_lo_2750};
  wire [15:0]   dataGroup_30_49 = dataGroup_hi_2750[415:400];
  wire [2047:0] dataGroup_lo_2751 = {dataGroup_lo_hi_2751, dataGroup_lo_lo_2751};
  wire [2047:0] dataGroup_hi_2751 = {dataGroup_hi_hi_2751, dataGroup_hi_lo_2751};
  wire [15:0]   dataGroup_31_49 = dataGroup_hi_2751[495:480];
  wire [31:0]   res_lo_lo_lo_lo_49 = {dataGroup_1_49, dataGroup_0_49};
  wire [31:0]   res_lo_lo_lo_hi_49 = {dataGroup_3_49, dataGroup_2_49};
  wire [63:0]   res_lo_lo_lo_49 = {res_lo_lo_lo_hi_49, res_lo_lo_lo_lo_49};
  wire [31:0]   res_lo_lo_hi_lo_49 = {dataGroup_5_49, dataGroup_4_49};
  wire [31:0]   res_lo_lo_hi_hi_49 = {dataGroup_7_49, dataGroup_6_49};
  wire [63:0]   res_lo_lo_hi_49 = {res_lo_lo_hi_hi_49, res_lo_lo_hi_lo_49};
  wire [127:0]  res_lo_lo_49 = {res_lo_lo_hi_49, res_lo_lo_lo_49};
  wire [31:0]   res_lo_hi_lo_lo_49 = {dataGroup_9_49, dataGroup_8_49};
  wire [31:0]   res_lo_hi_lo_hi_49 = {dataGroup_11_49, dataGroup_10_49};
  wire [63:0]   res_lo_hi_lo_49 = {res_lo_hi_lo_hi_49, res_lo_hi_lo_lo_49};
  wire [31:0]   res_lo_hi_hi_lo_49 = {dataGroup_13_49, dataGroup_12_49};
  wire [31:0]   res_lo_hi_hi_hi_49 = {dataGroup_15_49, dataGroup_14_49};
  wire [63:0]   res_lo_hi_hi_49 = {res_lo_hi_hi_hi_49, res_lo_hi_hi_lo_49};
  wire [127:0]  res_lo_hi_49 = {res_lo_hi_hi_49, res_lo_hi_lo_49};
  wire [255:0]  res_lo_49 = {res_lo_hi_49, res_lo_lo_49};
  wire [31:0]   res_hi_lo_lo_lo_49 = {dataGroup_17_49, dataGroup_16_49};
  wire [31:0]   res_hi_lo_lo_hi_49 = {dataGroup_19_49, dataGroup_18_49};
  wire [63:0]   res_hi_lo_lo_49 = {res_hi_lo_lo_hi_49, res_hi_lo_lo_lo_49};
  wire [31:0]   res_hi_lo_hi_lo_49 = {dataGroup_21_49, dataGroup_20_49};
  wire [31:0]   res_hi_lo_hi_hi_49 = {dataGroup_23_49, dataGroup_22_49};
  wire [63:0]   res_hi_lo_hi_49 = {res_hi_lo_hi_hi_49, res_hi_lo_hi_lo_49};
  wire [127:0]  res_hi_lo_49 = {res_hi_lo_hi_49, res_hi_lo_lo_49};
  wire [31:0]   res_hi_hi_lo_lo_49 = {dataGroup_25_49, dataGroup_24_49};
  wire [31:0]   res_hi_hi_lo_hi_49 = {dataGroup_27_49, dataGroup_26_49};
  wire [63:0]   res_hi_hi_lo_49 = {res_hi_hi_lo_hi_49, res_hi_hi_lo_lo_49};
  wire [31:0]   res_hi_hi_hi_lo_49 = {dataGroup_29_49, dataGroup_28_49};
  wire [31:0]   res_hi_hi_hi_hi_49 = {dataGroup_31_49, dataGroup_30_49};
  wire [63:0]   res_hi_hi_hi_49 = {res_hi_hi_hi_hi_49, res_hi_hi_hi_lo_49};
  wire [127:0]  res_hi_hi_49 = {res_hi_hi_hi_49, res_hi_hi_lo_49};
  wire [255:0]  res_hi_49 = {res_hi_hi_49, res_hi_lo_49};
  wire [511:0]  res_99 = {res_hi_49, res_lo_49};
  wire [2047:0] dataGroup_lo_2752 = {dataGroup_lo_hi_2752, dataGroup_lo_lo_2752};
  wire [2047:0] dataGroup_hi_2752 = {dataGroup_hi_hi_2752, dataGroup_hi_lo_2752};
  wire [15:0]   dataGroup_0_50 = dataGroup_lo_2752[79:64];
  wire [2047:0] dataGroup_lo_2753 = {dataGroup_lo_hi_2753, dataGroup_lo_lo_2753};
  wire [2047:0] dataGroup_hi_2753 = {dataGroup_hi_hi_2753, dataGroup_hi_lo_2753};
  wire [15:0]   dataGroup_1_50 = dataGroup_lo_2753[159:144];
  wire [2047:0] dataGroup_lo_2754 = {dataGroup_lo_hi_2754, dataGroup_lo_lo_2754};
  wire [2047:0] dataGroup_hi_2754 = {dataGroup_hi_hi_2754, dataGroup_hi_lo_2754};
  wire [15:0]   dataGroup_2_50 = dataGroup_lo_2754[239:224];
  wire [2047:0] dataGroup_lo_2755 = {dataGroup_lo_hi_2755, dataGroup_lo_lo_2755};
  wire [2047:0] dataGroup_hi_2755 = {dataGroup_hi_hi_2755, dataGroup_hi_lo_2755};
  wire [15:0]   dataGroup_3_50 = dataGroup_lo_2755[319:304];
  wire [2047:0] dataGroup_lo_2756 = {dataGroup_lo_hi_2756, dataGroup_lo_lo_2756};
  wire [2047:0] dataGroup_hi_2756 = {dataGroup_hi_hi_2756, dataGroup_hi_lo_2756};
  wire [15:0]   dataGroup_4_50 = dataGroup_lo_2756[399:384];
  wire [2047:0] dataGroup_lo_2757 = {dataGroup_lo_hi_2757, dataGroup_lo_lo_2757};
  wire [2047:0] dataGroup_hi_2757 = {dataGroup_hi_hi_2757, dataGroup_hi_lo_2757};
  wire [15:0]   dataGroup_5_50 = dataGroup_lo_2757[479:464];
  wire [2047:0] dataGroup_lo_2758 = {dataGroup_lo_hi_2758, dataGroup_lo_lo_2758};
  wire [2047:0] dataGroup_hi_2758 = {dataGroup_hi_hi_2758, dataGroup_hi_lo_2758};
  wire [15:0]   dataGroup_6_50 = dataGroup_lo_2758[559:544];
  wire [2047:0] dataGroup_lo_2759 = {dataGroup_lo_hi_2759, dataGroup_lo_lo_2759};
  wire [2047:0] dataGroup_hi_2759 = {dataGroup_hi_hi_2759, dataGroup_hi_lo_2759};
  wire [15:0]   dataGroup_7_50 = dataGroup_lo_2759[639:624];
  wire [2047:0] dataGroup_lo_2760 = {dataGroup_lo_hi_2760, dataGroup_lo_lo_2760};
  wire [2047:0] dataGroup_hi_2760 = {dataGroup_hi_hi_2760, dataGroup_hi_lo_2760};
  wire [15:0]   dataGroup_8_50 = dataGroup_lo_2760[719:704];
  wire [2047:0] dataGroup_lo_2761 = {dataGroup_lo_hi_2761, dataGroup_lo_lo_2761};
  wire [2047:0] dataGroup_hi_2761 = {dataGroup_hi_hi_2761, dataGroup_hi_lo_2761};
  wire [15:0]   dataGroup_9_50 = dataGroup_lo_2761[799:784];
  wire [2047:0] dataGroup_lo_2762 = {dataGroup_lo_hi_2762, dataGroup_lo_lo_2762};
  wire [2047:0] dataGroup_hi_2762 = {dataGroup_hi_hi_2762, dataGroup_hi_lo_2762};
  wire [15:0]   dataGroup_10_50 = dataGroup_lo_2762[879:864];
  wire [2047:0] dataGroup_lo_2763 = {dataGroup_lo_hi_2763, dataGroup_lo_lo_2763};
  wire [2047:0] dataGroup_hi_2763 = {dataGroup_hi_hi_2763, dataGroup_hi_lo_2763};
  wire [15:0]   dataGroup_11_50 = dataGroup_lo_2763[959:944];
  wire [2047:0] dataGroup_lo_2764 = {dataGroup_lo_hi_2764, dataGroup_lo_lo_2764};
  wire [2047:0] dataGroup_hi_2764 = {dataGroup_hi_hi_2764, dataGroup_hi_lo_2764};
  wire [15:0]   dataGroup_12_50 = dataGroup_lo_2764[1039:1024];
  wire [2047:0] dataGroup_lo_2765 = {dataGroup_lo_hi_2765, dataGroup_lo_lo_2765};
  wire [2047:0] dataGroup_hi_2765 = {dataGroup_hi_hi_2765, dataGroup_hi_lo_2765};
  wire [15:0]   dataGroup_13_50 = dataGroup_lo_2765[1119:1104];
  wire [2047:0] dataGroup_lo_2766 = {dataGroup_lo_hi_2766, dataGroup_lo_lo_2766};
  wire [2047:0] dataGroup_hi_2766 = {dataGroup_hi_hi_2766, dataGroup_hi_lo_2766};
  wire [15:0]   dataGroup_14_50 = dataGroup_lo_2766[1199:1184];
  wire [2047:0] dataGroup_lo_2767 = {dataGroup_lo_hi_2767, dataGroup_lo_lo_2767};
  wire [2047:0] dataGroup_hi_2767 = {dataGroup_hi_hi_2767, dataGroup_hi_lo_2767};
  wire [15:0]   dataGroup_15_50 = dataGroup_lo_2767[1279:1264];
  wire [2047:0] dataGroup_lo_2768 = {dataGroup_lo_hi_2768, dataGroup_lo_lo_2768};
  wire [2047:0] dataGroup_hi_2768 = {dataGroup_hi_hi_2768, dataGroup_hi_lo_2768};
  wire [15:0]   dataGroup_16_50 = dataGroup_lo_2768[1359:1344];
  wire [2047:0] dataGroup_lo_2769 = {dataGroup_lo_hi_2769, dataGroup_lo_lo_2769};
  wire [2047:0] dataGroup_hi_2769 = {dataGroup_hi_hi_2769, dataGroup_hi_lo_2769};
  wire [15:0]   dataGroup_17_50 = dataGroup_lo_2769[1439:1424];
  wire [2047:0] dataGroup_lo_2770 = {dataGroup_lo_hi_2770, dataGroup_lo_lo_2770};
  wire [2047:0] dataGroup_hi_2770 = {dataGroup_hi_hi_2770, dataGroup_hi_lo_2770};
  wire [15:0]   dataGroup_18_50 = dataGroup_lo_2770[1519:1504];
  wire [2047:0] dataGroup_lo_2771 = {dataGroup_lo_hi_2771, dataGroup_lo_lo_2771};
  wire [2047:0] dataGroup_hi_2771 = {dataGroup_hi_hi_2771, dataGroup_hi_lo_2771};
  wire [15:0]   dataGroup_19_50 = dataGroup_lo_2771[1599:1584];
  wire [2047:0] dataGroup_lo_2772 = {dataGroup_lo_hi_2772, dataGroup_lo_lo_2772};
  wire [2047:0] dataGroup_hi_2772 = {dataGroup_hi_hi_2772, dataGroup_hi_lo_2772};
  wire [15:0]   dataGroup_20_50 = dataGroup_lo_2772[1679:1664];
  wire [2047:0] dataGroup_lo_2773 = {dataGroup_lo_hi_2773, dataGroup_lo_lo_2773};
  wire [2047:0] dataGroup_hi_2773 = {dataGroup_hi_hi_2773, dataGroup_hi_lo_2773};
  wire [15:0]   dataGroup_21_50 = dataGroup_lo_2773[1759:1744];
  wire [2047:0] dataGroup_lo_2774 = {dataGroup_lo_hi_2774, dataGroup_lo_lo_2774};
  wire [2047:0] dataGroup_hi_2774 = {dataGroup_hi_hi_2774, dataGroup_hi_lo_2774};
  wire [15:0]   dataGroup_22_50 = dataGroup_lo_2774[1839:1824];
  wire [2047:0] dataGroup_lo_2775 = {dataGroup_lo_hi_2775, dataGroup_lo_lo_2775};
  wire [2047:0] dataGroup_hi_2775 = {dataGroup_hi_hi_2775, dataGroup_hi_lo_2775};
  wire [15:0]   dataGroup_23_50 = dataGroup_lo_2775[1919:1904];
  wire [2047:0] dataGroup_lo_2776 = {dataGroup_lo_hi_2776, dataGroup_lo_lo_2776};
  wire [2047:0] dataGroup_hi_2776 = {dataGroup_hi_hi_2776, dataGroup_hi_lo_2776};
  wire [15:0]   dataGroup_24_50 = dataGroup_lo_2776[1999:1984];
  wire [2047:0] dataGroup_lo_2777 = {dataGroup_lo_hi_2777, dataGroup_lo_lo_2777};
  wire [2047:0] dataGroup_hi_2777 = {dataGroup_hi_hi_2777, dataGroup_hi_lo_2777};
  wire [15:0]   dataGroup_25_50 = dataGroup_hi_2777[31:16];
  wire [2047:0] dataGroup_lo_2778 = {dataGroup_lo_hi_2778, dataGroup_lo_lo_2778};
  wire [2047:0] dataGroup_hi_2778 = {dataGroup_hi_hi_2778, dataGroup_hi_lo_2778};
  wire [15:0]   dataGroup_26_50 = dataGroup_hi_2778[111:96];
  wire [2047:0] dataGroup_lo_2779 = {dataGroup_lo_hi_2779, dataGroup_lo_lo_2779};
  wire [2047:0] dataGroup_hi_2779 = {dataGroup_hi_hi_2779, dataGroup_hi_lo_2779};
  wire [15:0]   dataGroup_27_50 = dataGroup_hi_2779[191:176];
  wire [2047:0] dataGroup_lo_2780 = {dataGroup_lo_hi_2780, dataGroup_lo_lo_2780};
  wire [2047:0] dataGroup_hi_2780 = {dataGroup_hi_hi_2780, dataGroup_hi_lo_2780};
  wire [15:0]   dataGroup_28_50 = dataGroup_hi_2780[271:256];
  wire [2047:0] dataGroup_lo_2781 = {dataGroup_lo_hi_2781, dataGroup_lo_lo_2781};
  wire [2047:0] dataGroup_hi_2781 = {dataGroup_hi_hi_2781, dataGroup_hi_lo_2781};
  wire [15:0]   dataGroup_29_50 = dataGroup_hi_2781[351:336];
  wire [2047:0] dataGroup_lo_2782 = {dataGroup_lo_hi_2782, dataGroup_lo_lo_2782};
  wire [2047:0] dataGroup_hi_2782 = {dataGroup_hi_hi_2782, dataGroup_hi_lo_2782};
  wire [15:0]   dataGroup_30_50 = dataGroup_hi_2782[431:416];
  wire [2047:0] dataGroup_lo_2783 = {dataGroup_lo_hi_2783, dataGroup_lo_lo_2783};
  wire [2047:0] dataGroup_hi_2783 = {dataGroup_hi_hi_2783, dataGroup_hi_lo_2783};
  wire [15:0]   dataGroup_31_50 = dataGroup_hi_2783[511:496];
  wire [31:0]   res_lo_lo_lo_lo_50 = {dataGroup_1_50, dataGroup_0_50};
  wire [31:0]   res_lo_lo_lo_hi_50 = {dataGroup_3_50, dataGroup_2_50};
  wire [63:0]   res_lo_lo_lo_50 = {res_lo_lo_lo_hi_50, res_lo_lo_lo_lo_50};
  wire [31:0]   res_lo_lo_hi_lo_50 = {dataGroup_5_50, dataGroup_4_50};
  wire [31:0]   res_lo_lo_hi_hi_50 = {dataGroup_7_50, dataGroup_6_50};
  wire [63:0]   res_lo_lo_hi_50 = {res_lo_lo_hi_hi_50, res_lo_lo_hi_lo_50};
  wire [127:0]  res_lo_lo_50 = {res_lo_lo_hi_50, res_lo_lo_lo_50};
  wire [31:0]   res_lo_hi_lo_lo_50 = {dataGroup_9_50, dataGroup_8_50};
  wire [31:0]   res_lo_hi_lo_hi_50 = {dataGroup_11_50, dataGroup_10_50};
  wire [63:0]   res_lo_hi_lo_50 = {res_lo_hi_lo_hi_50, res_lo_hi_lo_lo_50};
  wire [31:0]   res_lo_hi_hi_lo_50 = {dataGroup_13_50, dataGroup_12_50};
  wire [31:0]   res_lo_hi_hi_hi_50 = {dataGroup_15_50, dataGroup_14_50};
  wire [63:0]   res_lo_hi_hi_50 = {res_lo_hi_hi_hi_50, res_lo_hi_hi_lo_50};
  wire [127:0]  res_lo_hi_50 = {res_lo_hi_hi_50, res_lo_hi_lo_50};
  wire [255:0]  res_lo_50 = {res_lo_hi_50, res_lo_lo_50};
  wire [31:0]   res_hi_lo_lo_lo_50 = {dataGroup_17_50, dataGroup_16_50};
  wire [31:0]   res_hi_lo_lo_hi_50 = {dataGroup_19_50, dataGroup_18_50};
  wire [63:0]   res_hi_lo_lo_50 = {res_hi_lo_lo_hi_50, res_hi_lo_lo_lo_50};
  wire [31:0]   res_hi_lo_hi_lo_50 = {dataGroup_21_50, dataGroup_20_50};
  wire [31:0]   res_hi_lo_hi_hi_50 = {dataGroup_23_50, dataGroup_22_50};
  wire [63:0]   res_hi_lo_hi_50 = {res_hi_lo_hi_hi_50, res_hi_lo_hi_lo_50};
  wire [127:0]  res_hi_lo_50 = {res_hi_lo_hi_50, res_hi_lo_lo_50};
  wire [31:0]   res_hi_hi_lo_lo_50 = {dataGroup_25_50, dataGroup_24_50};
  wire [31:0]   res_hi_hi_lo_hi_50 = {dataGroup_27_50, dataGroup_26_50};
  wire [63:0]   res_hi_hi_lo_50 = {res_hi_hi_lo_hi_50, res_hi_hi_lo_lo_50};
  wire [31:0]   res_hi_hi_hi_lo_50 = {dataGroup_29_50, dataGroup_28_50};
  wire [31:0]   res_hi_hi_hi_hi_50 = {dataGroup_31_50, dataGroup_30_50};
  wire [63:0]   res_hi_hi_hi_50 = {res_hi_hi_hi_hi_50, res_hi_hi_hi_lo_50};
  wire [127:0]  res_hi_hi_50 = {res_hi_hi_hi_50, res_hi_hi_lo_50};
  wire [255:0]  res_hi_50 = {res_hi_hi_50, res_hi_lo_50};
  wire [511:0]  res_100 = {res_hi_50, res_lo_50};
  wire [1023:0] lo_lo_12 = {res_97, res_96};
  wire [1023:0] lo_hi_12 = {res_99, res_98};
  wire [2047:0] lo_12 = {lo_hi_12, lo_lo_12};
  wire [1023:0] hi_lo_12 = {512'h0, res_100};
  wire [2047:0] hi_12 = {1024'h0, hi_lo_12};
  wire [4095:0] regroupLoadData_1_4 = {hi_12, lo_12};
  wire [2047:0] dataGroup_lo_2784 = {dataGroup_lo_hi_2784, dataGroup_lo_lo_2784};
  wire [2047:0] dataGroup_hi_2784 = {dataGroup_hi_hi_2784, dataGroup_hi_lo_2784};
  wire [15:0]   dataGroup_0_51 = dataGroup_lo_2784[15:0];
  wire [2047:0] dataGroup_lo_2785 = {dataGroup_lo_hi_2785, dataGroup_lo_lo_2785};
  wire [2047:0] dataGroup_hi_2785 = {dataGroup_hi_hi_2785, dataGroup_hi_lo_2785};
  wire [15:0]   dataGroup_1_51 = dataGroup_lo_2785[111:96];
  wire [2047:0] dataGroup_lo_2786 = {dataGroup_lo_hi_2786, dataGroup_lo_lo_2786};
  wire [2047:0] dataGroup_hi_2786 = {dataGroup_hi_hi_2786, dataGroup_hi_lo_2786};
  wire [15:0]   dataGroup_2_51 = dataGroup_lo_2786[207:192];
  wire [2047:0] dataGroup_lo_2787 = {dataGroup_lo_hi_2787, dataGroup_lo_lo_2787};
  wire [2047:0] dataGroup_hi_2787 = {dataGroup_hi_hi_2787, dataGroup_hi_lo_2787};
  wire [15:0]   dataGroup_3_51 = dataGroup_lo_2787[303:288];
  wire [2047:0] dataGroup_lo_2788 = {dataGroup_lo_hi_2788, dataGroup_lo_lo_2788};
  wire [2047:0] dataGroup_hi_2788 = {dataGroup_hi_hi_2788, dataGroup_hi_lo_2788};
  wire [15:0]   dataGroup_4_51 = dataGroup_lo_2788[399:384];
  wire [2047:0] dataGroup_lo_2789 = {dataGroup_lo_hi_2789, dataGroup_lo_lo_2789};
  wire [2047:0] dataGroup_hi_2789 = {dataGroup_hi_hi_2789, dataGroup_hi_lo_2789};
  wire [15:0]   dataGroup_5_51 = dataGroup_lo_2789[495:480];
  wire [2047:0] dataGroup_lo_2790 = {dataGroup_lo_hi_2790, dataGroup_lo_lo_2790};
  wire [2047:0] dataGroup_hi_2790 = {dataGroup_hi_hi_2790, dataGroup_hi_lo_2790};
  wire [15:0]   dataGroup_6_51 = dataGroup_lo_2790[591:576];
  wire [2047:0] dataGroup_lo_2791 = {dataGroup_lo_hi_2791, dataGroup_lo_lo_2791};
  wire [2047:0] dataGroup_hi_2791 = {dataGroup_hi_hi_2791, dataGroup_hi_lo_2791};
  wire [15:0]   dataGroup_7_51 = dataGroup_lo_2791[687:672];
  wire [2047:0] dataGroup_lo_2792 = {dataGroup_lo_hi_2792, dataGroup_lo_lo_2792};
  wire [2047:0] dataGroup_hi_2792 = {dataGroup_hi_hi_2792, dataGroup_hi_lo_2792};
  wire [15:0]   dataGroup_8_51 = dataGroup_lo_2792[783:768];
  wire [2047:0] dataGroup_lo_2793 = {dataGroup_lo_hi_2793, dataGroup_lo_lo_2793};
  wire [2047:0] dataGroup_hi_2793 = {dataGroup_hi_hi_2793, dataGroup_hi_lo_2793};
  wire [15:0]   dataGroup_9_51 = dataGroup_lo_2793[879:864];
  wire [2047:0] dataGroup_lo_2794 = {dataGroup_lo_hi_2794, dataGroup_lo_lo_2794};
  wire [2047:0] dataGroup_hi_2794 = {dataGroup_hi_hi_2794, dataGroup_hi_lo_2794};
  wire [15:0]   dataGroup_10_51 = dataGroup_lo_2794[975:960];
  wire [2047:0] dataGroup_lo_2795 = {dataGroup_lo_hi_2795, dataGroup_lo_lo_2795};
  wire [2047:0] dataGroup_hi_2795 = {dataGroup_hi_hi_2795, dataGroup_hi_lo_2795};
  wire [15:0]   dataGroup_11_51 = dataGroup_lo_2795[1071:1056];
  wire [2047:0] dataGroup_lo_2796 = {dataGroup_lo_hi_2796, dataGroup_lo_lo_2796};
  wire [2047:0] dataGroup_hi_2796 = {dataGroup_hi_hi_2796, dataGroup_hi_lo_2796};
  wire [15:0]   dataGroup_12_51 = dataGroup_lo_2796[1167:1152];
  wire [2047:0] dataGroup_lo_2797 = {dataGroup_lo_hi_2797, dataGroup_lo_lo_2797};
  wire [2047:0] dataGroup_hi_2797 = {dataGroup_hi_hi_2797, dataGroup_hi_lo_2797};
  wire [15:0]   dataGroup_13_51 = dataGroup_lo_2797[1263:1248];
  wire [2047:0] dataGroup_lo_2798 = {dataGroup_lo_hi_2798, dataGroup_lo_lo_2798};
  wire [2047:0] dataGroup_hi_2798 = {dataGroup_hi_hi_2798, dataGroup_hi_lo_2798};
  wire [15:0]   dataGroup_14_51 = dataGroup_lo_2798[1359:1344];
  wire [2047:0] dataGroup_lo_2799 = {dataGroup_lo_hi_2799, dataGroup_lo_lo_2799};
  wire [2047:0] dataGroup_hi_2799 = {dataGroup_hi_hi_2799, dataGroup_hi_lo_2799};
  wire [15:0]   dataGroup_15_51 = dataGroup_lo_2799[1455:1440];
  wire [2047:0] dataGroup_lo_2800 = {dataGroup_lo_hi_2800, dataGroup_lo_lo_2800};
  wire [2047:0] dataGroup_hi_2800 = {dataGroup_hi_hi_2800, dataGroup_hi_lo_2800};
  wire [15:0]   dataGroup_16_51 = dataGroup_lo_2800[1551:1536];
  wire [2047:0] dataGroup_lo_2801 = {dataGroup_lo_hi_2801, dataGroup_lo_lo_2801};
  wire [2047:0] dataGroup_hi_2801 = {dataGroup_hi_hi_2801, dataGroup_hi_lo_2801};
  wire [15:0]   dataGroup_17_51 = dataGroup_lo_2801[1647:1632];
  wire [2047:0] dataGroup_lo_2802 = {dataGroup_lo_hi_2802, dataGroup_lo_lo_2802};
  wire [2047:0] dataGroup_hi_2802 = {dataGroup_hi_hi_2802, dataGroup_hi_lo_2802};
  wire [15:0]   dataGroup_18_51 = dataGroup_lo_2802[1743:1728];
  wire [2047:0] dataGroup_lo_2803 = {dataGroup_lo_hi_2803, dataGroup_lo_lo_2803};
  wire [2047:0] dataGroup_hi_2803 = {dataGroup_hi_hi_2803, dataGroup_hi_lo_2803};
  wire [15:0]   dataGroup_19_51 = dataGroup_lo_2803[1839:1824];
  wire [2047:0] dataGroup_lo_2804 = {dataGroup_lo_hi_2804, dataGroup_lo_lo_2804};
  wire [2047:0] dataGroup_hi_2804 = {dataGroup_hi_hi_2804, dataGroup_hi_lo_2804};
  wire [15:0]   dataGroup_20_51 = dataGroup_lo_2804[1935:1920];
  wire [2047:0] dataGroup_lo_2805 = {dataGroup_lo_hi_2805, dataGroup_lo_lo_2805};
  wire [2047:0] dataGroup_hi_2805 = {dataGroup_hi_hi_2805, dataGroup_hi_lo_2805};
  wire [15:0]   dataGroup_21_51 = dataGroup_lo_2805[2031:2016];
  wire [2047:0] dataGroup_lo_2806 = {dataGroup_lo_hi_2806, dataGroup_lo_lo_2806};
  wire [2047:0] dataGroup_hi_2806 = {dataGroup_hi_hi_2806, dataGroup_hi_lo_2806};
  wire [15:0]   dataGroup_22_51 = dataGroup_hi_2806[79:64];
  wire [2047:0] dataGroup_lo_2807 = {dataGroup_lo_hi_2807, dataGroup_lo_lo_2807};
  wire [2047:0] dataGroup_hi_2807 = {dataGroup_hi_hi_2807, dataGroup_hi_lo_2807};
  wire [15:0]   dataGroup_23_51 = dataGroup_hi_2807[175:160];
  wire [2047:0] dataGroup_lo_2808 = {dataGroup_lo_hi_2808, dataGroup_lo_lo_2808};
  wire [2047:0] dataGroup_hi_2808 = {dataGroup_hi_hi_2808, dataGroup_hi_lo_2808};
  wire [15:0]   dataGroup_24_51 = dataGroup_hi_2808[271:256];
  wire [2047:0] dataGroup_lo_2809 = {dataGroup_lo_hi_2809, dataGroup_lo_lo_2809};
  wire [2047:0] dataGroup_hi_2809 = {dataGroup_hi_hi_2809, dataGroup_hi_lo_2809};
  wire [15:0]   dataGroup_25_51 = dataGroup_hi_2809[367:352];
  wire [2047:0] dataGroup_lo_2810 = {dataGroup_lo_hi_2810, dataGroup_lo_lo_2810};
  wire [2047:0] dataGroup_hi_2810 = {dataGroup_hi_hi_2810, dataGroup_hi_lo_2810};
  wire [15:0]   dataGroup_26_51 = dataGroup_hi_2810[463:448];
  wire [2047:0] dataGroup_lo_2811 = {dataGroup_lo_hi_2811, dataGroup_lo_lo_2811};
  wire [2047:0] dataGroup_hi_2811 = {dataGroup_hi_hi_2811, dataGroup_hi_lo_2811};
  wire [15:0]   dataGroup_27_51 = dataGroup_hi_2811[559:544];
  wire [2047:0] dataGroup_lo_2812 = {dataGroup_lo_hi_2812, dataGroup_lo_lo_2812};
  wire [2047:0] dataGroup_hi_2812 = {dataGroup_hi_hi_2812, dataGroup_hi_lo_2812};
  wire [15:0]   dataGroup_28_51 = dataGroup_hi_2812[655:640];
  wire [2047:0] dataGroup_lo_2813 = {dataGroup_lo_hi_2813, dataGroup_lo_lo_2813};
  wire [2047:0] dataGroup_hi_2813 = {dataGroup_hi_hi_2813, dataGroup_hi_lo_2813};
  wire [15:0]   dataGroup_29_51 = dataGroup_hi_2813[751:736];
  wire [2047:0] dataGroup_lo_2814 = {dataGroup_lo_hi_2814, dataGroup_lo_lo_2814};
  wire [2047:0] dataGroup_hi_2814 = {dataGroup_hi_hi_2814, dataGroup_hi_lo_2814};
  wire [15:0]   dataGroup_30_51 = dataGroup_hi_2814[847:832];
  wire [2047:0] dataGroup_lo_2815 = {dataGroup_lo_hi_2815, dataGroup_lo_lo_2815};
  wire [2047:0] dataGroup_hi_2815 = {dataGroup_hi_hi_2815, dataGroup_hi_lo_2815};
  wire [15:0]   dataGroup_31_51 = dataGroup_hi_2815[943:928];
  wire [31:0]   res_lo_lo_lo_lo_51 = {dataGroup_1_51, dataGroup_0_51};
  wire [31:0]   res_lo_lo_lo_hi_51 = {dataGroup_3_51, dataGroup_2_51};
  wire [63:0]   res_lo_lo_lo_51 = {res_lo_lo_lo_hi_51, res_lo_lo_lo_lo_51};
  wire [31:0]   res_lo_lo_hi_lo_51 = {dataGroup_5_51, dataGroup_4_51};
  wire [31:0]   res_lo_lo_hi_hi_51 = {dataGroup_7_51, dataGroup_6_51};
  wire [63:0]   res_lo_lo_hi_51 = {res_lo_lo_hi_hi_51, res_lo_lo_hi_lo_51};
  wire [127:0]  res_lo_lo_51 = {res_lo_lo_hi_51, res_lo_lo_lo_51};
  wire [31:0]   res_lo_hi_lo_lo_51 = {dataGroup_9_51, dataGroup_8_51};
  wire [31:0]   res_lo_hi_lo_hi_51 = {dataGroup_11_51, dataGroup_10_51};
  wire [63:0]   res_lo_hi_lo_51 = {res_lo_hi_lo_hi_51, res_lo_hi_lo_lo_51};
  wire [31:0]   res_lo_hi_hi_lo_51 = {dataGroup_13_51, dataGroup_12_51};
  wire [31:0]   res_lo_hi_hi_hi_51 = {dataGroup_15_51, dataGroup_14_51};
  wire [63:0]   res_lo_hi_hi_51 = {res_lo_hi_hi_hi_51, res_lo_hi_hi_lo_51};
  wire [127:0]  res_lo_hi_51 = {res_lo_hi_hi_51, res_lo_hi_lo_51};
  wire [255:0]  res_lo_51 = {res_lo_hi_51, res_lo_lo_51};
  wire [31:0]   res_hi_lo_lo_lo_51 = {dataGroup_17_51, dataGroup_16_51};
  wire [31:0]   res_hi_lo_lo_hi_51 = {dataGroup_19_51, dataGroup_18_51};
  wire [63:0]   res_hi_lo_lo_51 = {res_hi_lo_lo_hi_51, res_hi_lo_lo_lo_51};
  wire [31:0]   res_hi_lo_hi_lo_51 = {dataGroup_21_51, dataGroup_20_51};
  wire [31:0]   res_hi_lo_hi_hi_51 = {dataGroup_23_51, dataGroup_22_51};
  wire [63:0]   res_hi_lo_hi_51 = {res_hi_lo_hi_hi_51, res_hi_lo_hi_lo_51};
  wire [127:0]  res_hi_lo_51 = {res_hi_lo_hi_51, res_hi_lo_lo_51};
  wire [31:0]   res_hi_hi_lo_lo_51 = {dataGroup_25_51, dataGroup_24_51};
  wire [31:0]   res_hi_hi_lo_hi_51 = {dataGroup_27_51, dataGroup_26_51};
  wire [63:0]   res_hi_hi_lo_51 = {res_hi_hi_lo_hi_51, res_hi_hi_lo_lo_51};
  wire [31:0]   res_hi_hi_hi_lo_51 = {dataGroup_29_51, dataGroup_28_51};
  wire [31:0]   res_hi_hi_hi_hi_51 = {dataGroup_31_51, dataGroup_30_51};
  wire [63:0]   res_hi_hi_hi_51 = {res_hi_hi_hi_hi_51, res_hi_hi_hi_lo_51};
  wire [127:0]  res_hi_hi_51 = {res_hi_hi_hi_51, res_hi_hi_lo_51};
  wire [255:0]  res_hi_51 = {res_hi_hi_51, res_hi_lo_51};
  wire [511:0]  res_104 = {res_hi_51, res_lo_51};
  wire [2047:0] dataGroup_lo_2816 = {dataGroup_lo_hi_2816, dataGroup_lo_lo_2816};
  wire [2047:0] dataGroup_hi_2816 = {dataGroup_hi_hi_2816, dataGroup_hi_lo_2816};
  wire [15:0]   dataGroup_0_52 = dataGroup_lo_2816[31:16];
  wire [2047:0] dataGroup_lo_2817 = {dataGroup_lo_hi_2817, dataGroup_lo_lo_2817};
  wire [2047:0] dataGroup_hi_2817 = {dataGroup_hi_hi_2817, dataGroup_hi_lo_2817};
  wire [15:0]   dataGroup_1_52 = dataGroup_lo_2817[127:112];
  wire [2047:0] dataGroup_lo_2818 = {dataGroup_lo_hi_2818, dataGroup_lo_lo_2818};
  wire [2047:0] dataGroup_hi_2818 = {dataGroup_hi_hi_2818, dataGroup_hi_lo_2818};
  wire [15:0]   dataGroup_2_52 = dataGroup_lo_2818[223:208];
  wire [2047:0] dataGroup_lo_2819 = {dataGroup_lo_hi_2819, dataGroup_lo_lo_2819};
  wire [2047:0] dataGroup_hi_2819 = {dataGroup_hi_hi_2819, dataGroup_hi_lo_2819};
  wire [15:0]   dataGroup_3_52 = dataGroup_lo_2819[319:304];
  wire [2047:0] dataGroup_lo_2820 = {dataGroup_lo_hi_2820, dataGroup_lo_lo_2820};
  wire [2047:0] dataGroup_hi_2820 = {dataGroup_hi_hi_2820, dataGroup_hi_lo_2820};
  wire [15:0]   dataGroup_4_52 = dataGroup_lo_2820[415:400];
  wire [2047:0] dataGroup_lo_2821 = {dataGroup_lo_hi_2821, dataGroup_lo_lo_2821};
  wire [2047:0] dataGroup_hi_2821 = {dataGroup_hi_hi_2821, dataGroup_hi_lo_2821};
  wire [15:0]   dataGroup_5_52 = dataGroup_lo_2821[511:496];
  wire [2047:0] dataGroup_lo_2822 = {dataGroup_lo_hi_2822, dataGroup_lo_lo_2822};
  wire [2047:0] dataGroup_hi_2822 = {dataGroup_hi_hi_2822, dataGroup_hi_lo_2822};
  wire [15:0]   dataGroup_6_52 = dataGroup_lo_2822[607:592];
  wire [2047:0] dataGroup_lo_2823 = {dataGroup_lo_hi_2823, dataGroup_lo_lo_2823};
  wire [2047:0] dataGroup_hi_2823 = {dataGroup_hi_hi_2823, dataGroup_hi_lo_2823};
  wire [15:0]   dataGroup_7_52 = dataGroup_lo_2823[703:688];
  wire [2047:0] dataGroup_lo_2824 = {dataGroup_lo_hi_2824, dataGroup_lo_lo_2824};
  wire [2047:0] dataGroup_hi_2824 = {dataGroup_hi_hi_2824, dataGroup_hi_lo_2824};
  wire [15:0]   dataGroup_8_52 = dataGroup_lo_2824[799:784];
  wire [2047:0] dataGroup_lo_2825 = {dataGroup_lo_hi_2825, dataGroup_lo_lo_2825};
  wire [2047:0] dataGroup_hi_2825 = {dataGroup_hi_hi_2825, dataGroup_hi_lo_2825};
  wire [15:0]   dataGroup_9_52 = dataGroup_lo_2825[895:880];
  wire [2047:0] dataGroup_lo_2826 = {dataGroup_lo_hi_2826, dataGroup_lo_lo_2826};
  wire [2047:0] dataGroup_hi_2826 = {dataGroup_hi_hi_2826, dataGroup_hi_lo_2826};
  wire [15:0]   dataGroup_10_52 = dataGroup_lo_2826[991:976];
  wire [2047:0] dataGroup_lo_2827 = {dataGroup_lo_hi_2827, dataGroup_lo_lo_2827};
  wire [2047:0] dataGroup_hi_2827 = {dataGroup_hi_hi_2827, dataGroup_hi_lo_2827};
  wire [15:0]   dataGroup_11_52 = dataGroup_lo_2827[1087:1072];
  wire [2047:0] dataGroup_lo_2828 = {dataGroup_lo_hi_2828, dataGroup_lo_lo_2828};
  wire [2047:0] dataGroup_hi_2828 = {dataGroup_hi_hi_2828, dataGroup_hi_lo_2828};
  wire [15:0]   dataGroup_12_52 = dataGroup_lo_2828[1183:1168];
  wire [2047:0] dataGroup_lo_2829 = {dataGroup_lo_hi_2829, dataGroup_lo_lo_2829};
  wire [2047:0] dataGroup_hi_2829 = {dataGroup_hi_hi_2829, dataGroup_hi_lo_2829};
  wire [15:0]   dataGroup_13_52 = dataGroup_lo_2829[1279:1264];
  wire [2047:0] dataGroup_lo_2830 = {dataGroup_lo_hi_2830, dataGroup_lo_lo_2830};
  wire [2047:0] dataGroup_hi_2830 = {dataGroup_hi_hi_2830, dataGroup_hi_lo_2830};
  wire [15:0]   dataGroup_14_52 = dataGroup_lo_2830[1375:1360];
  wire [2047:0] dataGroup_lo_2831 = {dataGroup_lo_hi_2831, dataGroup_lo_lo_2831};
  wire [2047:0] dataGroup_hi_2831 = {dataGroup_hi_hi_2831, dataGroup_hi_lo_2831};
  wire [15:0]   dataGroup_15_52 = dataGroup_lo_2831[1471:1456];
  wire [2047:0] dataGroup_lo_2832 = {dataGroup_lo_hi_2832, dataGroup_lo_lo_2832};
  wire [2047:0] dataGroup_hi_2832 = {dataGroup_hi_hi_2832, dataGroup_hi_lo_2832};
  wire [15:0]   dataGroup_16_52 = dataGroup_lo_2832[1567:1552];
  wire [2047:0] dataGroup_lo_2833 = {dataGroup_lo_hi_2833, dataGroup_lo_lo_2833};
  wire [2047:0] dataGroup_hi_2833 = {dataGroup_hi_hi_2833, dataGroup_hi_lo_2833};
  wire [15:0]   dataGroup_17_52 = dataGroup_lo_2833[1663:1648];
  wire [2047:0] dataGroup_lo_2834 = {dataGroup_lo_hi_2834, dataGroup_lo_lo_2834};
  wire [2047:0] dataGroup_hi_2834 = {dataGroup_hi_hi_2834, dataGroup_hi_lo_2834};
  wire [15:0]   dataGroup_18_52 = dataGroup_lo_2834[1759:1744];
  wire [2047:0] dataGroup_lo_2835 = {dataGroup_lo_hi_2835, dataGroup_lo_lo_2835};
  wire [2047:0] dataGroup_hi_2835 = {dataGroup_hi_hi_2835, dataGroup_hi_lo_2835};
  wire [15:0]   dataGroup_19_52 = dataGroup_lo_2835[1855:1840];
  wire [2047:0] dataGroup_lo_2836 = {dataGroup_lo_hi_2836, dataGroup_lo_lo_2836};
  wire [2047:0] dataGroup_hi_2836 = {dataGroup_hi_hi_2836, dataGroup_hi_lo_2836};
  wire [15:0]   dataGroup_20_52 = dataGroup_lo_2836[1951:1936];
  wire [2047:0] dataGroup_lo_2837 = {dataGroup_lo_hi_2837, dataGroup_lo_lo_2837};
  wire [2047:0] dataGroup_hi_2837 = {dataGroup_hi_hi_2837, dataGroup_hi_lo_2837};
  wire [15:0]   dataGroup_21_52 = dataGroup_lo_2837[2047:2032];
  wire [2047:0] dataGroup_lo_2838 = {dataGroup_lo_hi_2838, dataGroup_lo_lo_2838};
  wire [2047:0] dataGroup_hi_2838 = {dataGroup_hi_hi_2838, dataGroup_hi_lo_2838};
  wire [15:0]   dataGroup_22_52 = dataGroup_hi_2838[95:80];
  wire [2047:0] dataGroup_lo_2839 = {dataGroup_lo_hi_2839, dataGroup_lo_lo_2839};
  wire [2047:0] dataGroup_hi_2839 = {dataGroup_hi_hi_2839, dataGroup_hi_lo_2839};
  wire [15:0]   dataGroup_23_52 = dataGroup_hi_2839[191:176];
  wire [2047:0] dataGroup_lo_2840 = {dataGroup_lo_hi_2840, dataGroup_lo_lo_2840};
  wire [2047:0] dataGroup_hi_2840 = {dataGroup_hi_hi_2840, dataGroup_hi_lo_2840};
  wire [15:0]   dataGroup_24_52 = dataGroup_hi_2840[287:272];
  wire [2047:0] dataGroup_lo_2841 = {dataGroup_lo_hi_2841, dataGroup_lo_lo_2841};
  wire [2047:0] dataGroup_hi_2841 = {dataGroup_hi_hi_2841, dataGroup_hi_lo_2841};
  wire [15:0]   dataGroup_25_52 = dataGroup_hi_2841[383:368];
  wire [2047:0] dataGroup_lo_2842 = {dataGroup_lo_hi_2842, dataGroup_lo_lo_2842};
  wire [2047:0] dataGroup_hi_2842 = {dataGroup_hi_hi_2842, dataGroup_hi_lo_2842};
  wire [15:0]   dataGroup_26_52 = dataGroup_hi_2842[479:464];
  wire [2047:0] dataGroup_lo_2843 = {dataGroup_lo_hi_2843, dataGroup_lo_lo_2843};
  wire [2047:0] dataGroup_hi_2843 = {dataGroup_hi_hi_2843, dataGroup_hi_lo_2843};
  wire [15:0]   dataGroup_27_52 = dataGroup_hi_2843[575:560];
  wire [2047:0] dataGroup_lo_2844 = {dataGroup_lo_hi_2844, dataGroup_lo_lo_2844};
  wire [2047:0] dataGroup_hi_2844 = {dataGroup_hi_hi_2844, dataGroup_hi_lo_2844};
  wire [15:0]   dataGroup_28_52 = dataGroup_hi_2844[671:656];
  wire [2047:0] dataGroup_lo_2845 = {dataGroup_lo_hi_2845, dataGroup_lo_lo_2845};
  wire [2047:0] dataGroup_hi_2845 = {dataGroup_hi_hi_2845, dataGroup_hi_lo_2845};
  wire [15:0]   dataGroup_29_52 = dataGroup_hi_2845[767:752];
  wire [2047:0] dataGroup_lo_2846 = {dataGroup_lo_hi_2846, dataGroup_lo_lo_2846};
  wire [2047:0] dataGroup_hi_2846 = {dataGroup_hi_hi_2846, dataGroup_hi_lo_2846};
  wire [15:0]   dataGroup_30_52 = dataGroup_hi_2846[863:848];
  wire [2047:0] dataGroup_lo_2847 = {dataGroup_lo_hi_2847, dataGroup_lo_lo_2847};
  wire [2047:0] dataGroup_hi_2847 = {dataGroup_hi_hi_2847, dataGroup_hi_lo_2847};
  wire [15:0]   dataGroup_31_52 = dataGroup_hi_2847[959:944];
  wire [31:0]   res_lo_lo_lo_lo_52 = {dataGroup_1_52, dataGroup_0_52};
  wire [31:0]   res_lo_lo_lo_hi_52 = {dataGroup_3_52, dataGroup_2_52};
  wire [63:0]   res_lo_lo_lo_52 = {res_lo_lo_lo_hi_52, res_lo_lo_lo_lo_52};
  wire [31:0]   res_lo_lo_hi_lo_52 = {dataGroup_5_52, dataGroup_4_52};
  wire [31:0]   res_lo_lo_hi_hi_52 = {dataGroup_7_52, dataGroup_6_52};
  wire [63:0]   res_lo_lo_hi_52 = {res_lo_lo_hi_hi_52, res_lo_lo_hi_lo_52};
  wire [127:0]  res_lo_lo_52 = {res_lo_lo_hi_52, res_lo_lo_lo_52};
  wire [31:0]   res_lo_hi_lo_lo_52 = {dataGroup_9_52, dataGroup_8_52};
  wire [31:0]   res_lo_hi_lo_hi_52 = {dataGroup_11_52, dataGroup_10_52};
  wire [63:0]   res_lo_hi_lo_52 = {res_lo_hi_lo_hi_52, res_lo_hi_lo_lo_52};
  wire [31:0]   res_lo_hi_hi_lo_52 = {dataGroup_13_52, dataGroup_12_52};
  wire [31:0]   res_lo_hi_hi_hi_52 = {dataGroup_15_52, dataGroup_14_52};
  wire [63:0]   res_lo_hi_hi_52 = {res_lo_hi_hi_hi_52, res_lo_hi_hi_lo_52};
  wire [127:0]  res_lo_hi_52 = {res_lo_hi_hi_52, res_lo_hi_lo_52};
  wire [255:0]  res_lo_52 = {res_lo_hi_52, res_lo_lo_52};
  wire [31:0]   res_hi_lo_lo_lo_52 = {dataGroup_17_52, dataGroup_16_52};
  wire [31:0]   res_hi_lo_lo_hi_52 = {dataGroup_19_52, dataGroup_18_52};
  wire [63:0]   res_hi_lo_lo_52 = {res_hi_lo_lo_hi_52, res_hi_lo_lo_lo_52};
  wire [31:0]   res_hi_lo_hi_lo_52 = {dataGroup_21_52, dataGroup_20_52};
  wire [31:0]   res_hi_lo_hi_hi_52 = {dataGroup_23_52, dataGroup_22_52};
  wire [63:0]   res_hi_lo_hi_52 = {res_hi_lo_hi_hi_52, res_hi_lo_hi_lo_52};
  wire [127:0]  res_hi_lo_52 = {res_hi_lo_hi_52, res_hi_lo_lo_52};
  wire [31:0]   res_hi_hi_lo_lo_52 = {dataGroup_25_52, dataGroup_24_52};
  wire [31:0]   res_hi_hi_lo_hi_52 = {dataGroup_27_52, dataGroup_26_52};
  wire [63:0]   res_hi_hi_lo_52 = {res_hi_hi_lo_hi_52, res_hi_hi_lo_lo_52};
  wire [31:0]   res_hi_hi_hi_lo_52 = {dataGroup_29_52, dataGroup_28_52};
  wire [31:0]   res_hi_hi_hi_hi_52 = {dataGroup_31_52, dataGroup_30_52};
  wire [63:0]   res_hi_hi_hi_52 = {res_hi_hi_hi_hi_52, res_hi_hi_hi_lo_52};
  wire [127:0]  res_hi_hi_52 = {res_hi_hi_hi_52, res_hi_hi_lo_52};
  wire [255:0]  res_hi_52 = {res_hi_hi_52, res_hi_lo_52};
  wire [511:0]  res_105 = {res_hi_52, res_lo_52};
  wire [2047:0] dataGroup_lo_2848 = {dataGroup_lo_hi_2848, dataGroup_lo_lo_2848};
  wire [2047:0] dataGroup_hi_2848 = {dataGroup_hi_hi_2848, dataGroup_hi_lo_2848};
  wire [15:0]   dataGroup_0_53 = dataGroup_lo_2848[47:32];
  wire [2047:0] dataGroup_lo_2849 = {dataGroup_lo_hi_2849, dataGroup_lo_lo_2849};
  wire [2047:0] dataGroup_hi_2849 = {dataGroup_hi_hi_2849, dataGroup_hi_lo_2849};
  wire [15:0]   dataGroup_1_53 = dataGroup_lo_2849[143:128];
  wire [2047:0] dataGroup_lo_2850 = {dataGroup_lo_hi_2850, dataGroup_lo_lo_2850};
  wire [2047:0] dataGroup_hi_2850 = {dataGroup_hi_hi_2850, dataGroup_hi_lo_2850};
  wire [15:0]   dataGroup_2_53 = dataGroup_lo_2850[239:224];
  wire [2047:0] dataGroup_lo_2851 = {dataGroup_lo_hi_2851, dataGroup_lo_lo_2851};
  wire [2047:0] dataGroup_hi_2851 = {dataGroup_hi_hi_2851, dataGroup_hi_lo_2851};
  wire [15:0]   dataGroup_3_53 = dataGroup_lo_2851[335:320];
  wire [2047:0] dataGroup_lo_2852 = {dataGroup_lo_hi_2852, dataGroup_lo_lo_2852};
  wire [2047:0] dataGroup_hi_2852 = {dataGroup_hi_hi_2852, dataGroup_hi_lo_2852};
  wire [15:0]   dataGroup_4_53 = dataGroup_lo_2852[431:416];
  wire [2047:0] dataGroup_lo_2853 = {dataGroup_lo_hi_2853, dataGroup_lo_lo_2853};
  wire [2047:0] dataGroup_hi_2853 = {dataGroup_hi_hi_2853, dataGroup_hi_lo_2853};
  wire [15:0]   dataGroup_5_53 = dataGroup_lo_2853[527:512];
  wire [2047:0] dataGroup_lo_2854 = {dataGroup_lo_hi_2854, dataGroup_lo_lo_2854};
  wire [2047:0] dataGroup_hi_2854 = {dataGroup_hi_hi_2854, dataGroup_hi_lo_2854};
  wire [15:0]   dataGroup_6_53 = dataGroup_lo_2854[623:608];
  wire [2047:0] dataGroup_lo_2855 = {dataGroup_lo_hi_2855, dataGroup_lo_lo_2855};
  wire [2047:0] dataGroup_hi_2855 = {dataGroup_hi_hi_2855, dataGroup_hi_lo_2855};
  wire [15:0]   dataGroup_7_53 = dataGroup_lo_2855[719:704];
  wire [2047:0] dataGroup_lo_2856 = {dataGroup_lo_hi_2856, dataGroup_lo_lo_2856};
  wire [2047:0] dataGroup_hi_2856 = {dataGroup_hi_hi_2856, dataGroup_hi_lo_2856};
  wire [15:0]   dataGroup_8_53 = dataGroup_lo_2856[815:800];
  wire [2047:0] dataGroup_lo_2857 = {dataGroup_lo_hi_2857, dataGroup_lo_lo_2857};
  wire [2047:0] dataGroup_hi_2857 = {dataGroup_hi_hi_2857, dataGroup_hi_lo_2857};
  wire [15:0]   dataGroup_9_53 = dataGroup_lo_2857[911:896];
  wire [2047:0] dataGroup_lo_2858 = {dataGroup_lo_hi_2858, dataGroup_lo_lo_2858};
  wire [2047:0] dataGroup_hi_2858 = {dataGroup_hi_hi_2858, dataGroup_hi_lo_2858};
  wire [15:0]   dataGroup_10_53 = dataGroup_lo_2858[1007:992];
  wire [2047:0] dataGroup_lo_2859 = {dataGroup_lo_hi_2859, dataGroup_lo_lo_2859};
  wire [2047:0] dataGroup_hi_2859 = {dataGroup_hi_hi_2859, dataGroup_hi_lo_2859};
  wire [15:0]   dataGroup_11_53 = dataGroup_lo_2859[1103:1088];
  wire [2047:0] dataGroup_lo_2860 = {dataGroup_lo_hi_2860, dataGroup_lo_lo_2860};
  wire [2047:0] dataGroup_hi_2860 = {dataGroup_hi_hi_2860, dataGroup_hi_lo_2860};
  wire [15:0]   dataGroup_12_53 = dataGroup_lo_2860[1199:1184];
  wire [2047:0] dataGroup_lo_2861 = {dataGroup_lo_hi_2861, dataGroup_lo_lo_2861};
  wire [2047:0] dataGroup_hi_2861 = {dataGroup_hi_hi_2861, dataGroup_hi_lo_2861};
  wire [15:0]   dataGroup_13_53 = dataGroup_lo_2861[1295:1280];
  wire [2047:0] dataGroup_lo_2862 = {dataGroup_lo_hi_2862, dataGroup_lo_lo_2862};
  wire [2047:0] dataGroup_hi_2862 = {dataGroup_hi_hi_2862, dataGroup_hi_lo_2862};
  wire [15:0]   dataGroup_14_53 = dataGroup_lo_2862[1391:1376];
  wire [2047:0] dataGroup_lo_2863 = {dataGroup_lo_hi_2863, dataGroup_lo_lo_2863};
  wire [2047:0] dataGroup_hi_2863 = {dataGroup_hi_hi_2863, dataGroup_hi_lo_2863};
  wire [15:0]   dataGroup_15_53 = dataGroup_lo_2863[1487:1472];
  wire [2047:0] dataGroup_lo_2864 = {dataGroup_lo_hi_2864, dataGroup_lo_lo_2864};
  wire [2047:0] dataGroup_hi_2864 = {dataGroup_hi_hi_2864, dataGroup_hi_lo_2864};
  wire [15:0]   dataGroup_16_53 = dataGroup_lo_2864[1583:1568];
  wire [2047:0] dataGroup_lo_2865 = {dataGroup_lo_hi_2865, dataGroup_lo_lo_2865};
  wire [2047:0] dataGroup_hi_2865 = {dataGroup_hi_hi_2865, dataGroup_hi_lo_2865};
  wire [15:0]   dataGroup_17_53 = dataGroup_lo_2865[1679:1664];
  wire [2047:0] dataGroup_lo_2866 = {dataGroup_lo_hi_2866, dataGroup_lo_lo_2866};
  wire [2047:0] dataGroup_hi_2866 = {dataGroup_hi_hi_2866, dataGroup_hi_lo_2866};
  wire [15:0]   dataGroup_18_53 = dataGroup_lo_2866[1775:1760];
  wire [2047:0] dataGroup_lo_2867 = {dataGroup_lo_hi_2867, dataGroup_lo_lo_2867};
  wire [2047:0] dataGroup_hi_2867 = {dataGroup_hi_hi_2867, dataGroup_hi_lo_2867};
  wire [15:0]   dataGroup_19_53 = dataGroup_lo_2867[1871:1856];
  wire [2047:0] dataGroup_lo_2868 = {dataGroup_lo_hi_2868, dataGroup_lo_lo_2868};
  wire [2047:0] dataGroup_hi_2868 = {dataGroup_hi_hi_2868, dataGroup_hi_lo_2868};
  wire [15:0]   dataGroup_20_53 = dataGroup_lo_2868[1967:1952];
  wire [2047:0] dataGroup_lo_2869 = {dataGroup_lo_hi_2869, dataGroup_lo_lo_2869};
  wire [2047:0] dataGroup_hi_2869 = {dataGroup_hi_hi_2869, dataGroup_hi_lo_2869};
  wire [15:0]   dataGroup_21_53 = dataGroup_hi_2869[15:0];
  wire [2047:0] dataGroup_lo_2870 = {dataGroup_lo_hi_2870, dataGroup_lo_lo_2870};
  wire [2047:0] dataGroup_hi_2870 = {dataGroup_hi_hi_2870, dataGroup_hi_lo_2870};
  wire [15:0]   dataGroup_22_53 = dataGroup_hi_2870[111:96];
  wire [2047:0] dataGroup_lo_2871 = {dataGroup_lo_hi_2871, dataGroup_lo_lo_2871};
  wire [2047:0] dataGroup_hi_2871 = {dataGroup_hi_hi_2871, dataGroup_hi_lo_2871};
  wire [15:0]   dataGroup_23_53 = dataGroup_hi_2871[207:192];
  wire [2047:0] dataGroup_lo_2872 = {dataGroup_lo_hi_2872, dataGroup_lo_lo_2872};
  wire [2047:0] dataGroup_hi_2872 = {dataGroup_hi_hi_2872, dataGroup_hi_lo_2872};
  wire [15:0]   dataGroup_24_53 = dataGroup_hi_2872[303:288];
  wire [2047:0] dataGroup_lo_2873 = {dataGroup_lo_hi_2873, dataGroup_lo_lo_2873};
  wire [2047:0] dataGroup_hi_2873 = {dataGroup_hi_hi_2873, dataGroup_hi_lo_2873};
  wire [15:0]   dataGroup_25_53 = dataGroup_hi_2873[399:384];
  wire [2047:0] dataGroup_lo_2874 = {dataGroup_lo_hi_2874, dataGroup_lo_lo_2874};
  wire [2047:0] dataGroup_hi_2874 = {dataGroup_hi_hi_2874, dataGroup_hi_lo_2874};
  wire [15:0]   dataGroup_26_53 = dataGroup_hi_2874[495:480];
  wire [2047:0] dataGroup_lo_2875 = {dataGroup_lo_hi_2875, dataGroup_lo_lo_2875};
  wire [2047:0] dataGroup_hi_2875 = {dataGroup_hi_hi_2875, dataGroup_hi_lo_2875};
  wire [15:0]   dataGroup_27_53 = dataGroup_hi_2875[591:576];
  wire [2047:0] dataGroup_lo_2876 = {dataGroup_lo_hi_2876, dataGroup_lo_lo_2876};
  wire [2047:0] dataGroup_hi_2876 = {dataGroup_hi_hi_2876, dataGroup_hi_lo_2876};
  wire [15:0]   dataGroup_28_53 = dataGroup_hi_2876[687:672];
  wire [2047:0] dataGroup_lo_2877 = {dataGroup_lo_hi_2877, dataGroup_lo_lo_2877};
  wire [2047:0] dataGroup_hi_2877 = {dataGroup_hi_hi_2877, dataGroup_hi_lo_2877};
  wire [15:0]   dataGroup_29_53 = dataGroup_hi_2877[783:768];
  wire [2047:0] dataGroup_lo_2878 = {dataGroup_lo_hi_2878, dataGroup_lo_lo_2878};
  wire [2047:0] dataGroup_hi_2878 = {dataGroup_hi_hi_2878, dataGroup_hi_lo_2878};
  wire [15:0]   dataGroup_30_53 = dataGroup_hi_2878[879:864];
  wire [2047:0] dataGroup_lo_2879 = {dataGroup_lo_hi_2879, dataGroup_lo_lo_2879};
  wire [2047:0] dataGroup_hi_2879 = {dataGroup_hi_hi_2879, dataGroup_hi_lo_2879};
  wire [15:0]   dataGroup_31_53 = dataGroup_hi_2879[975:960];
  wire [31:0]   res_lo_lo_lo_lo_53 = {dataGroup_1_53, dataGroup_0_53};
  wire [31:0]   res_lo_lo_lo_hi_53 = {dataGroup_3_53, dataGroup_2_53};
  wire [63:0]   res_lo_lo_lo_53 = {res_lo_lo_lo_hi_53, res_lo_lo_lo_lo_53};
  wire [31:0]   res_lo_lo_hi_lo_53 = {dataGroup_5_53, dataGroup_4_53};
  wire [31:0]   res_lo_lo_hi_hi_53 = {dataGroup_7_53, dataGroup_6_53};
  wire [63:0]   res_lo_lo_hi_53 = {res_lo_lo_hi_hi_53, res_lo_lo_hi_lo_53};
  wire [127:0]  res_lo_lo_53 = {res_lo_lo_hi_53, res_lo_lo_lo_53};
  wire [31:0]   res_lo_hi_lo_lo_53 = {dataGroup_9_53, dataGroup_8_53};
  wire [31:0]   res_lo_hi_lo_hi_53 = {dataGroup_11_53, dataGroup_10_53};
  wire [63:0]   res_lo_hi_lo_53 = {res_lo_hi_lo_hi_53, res_lo_hi_lo_lo_53};
  wire [31:0]   res_lo_hi_hi_lo_53 = {dataGroup_13_53, dataGroup_12_53};
  wire [31:0]   res_lo_hi_hi_hi_53 = {dataGroup_15_53, dataGroup_14_53};
  wire [63:0]   res_lo_hi_hi_53 = {res_lo_hi_hi_hi_53, res_lo_hi_hi_lo_53};
  wire [127:0]  res_lo_hi_53 = {res_lo_hi_hi_53, res_lo_hi_lo_53};
  wire [255:0]  res_lo_53 = {res_lo_hi_53, res_lo_lo_53};
  wire [31:0]   res_hi_lo_lo_lo_53 = {dataGroup_17_53, dataGroup_16_53};
  wire [31:0]   res_hi_lo_lo_hi_53 = {dataGroup_19_53, dataGroup_18_53};
  wire [63:0]   res_hi_lo_lo_53 = {res_hi_lo_lo_hi_53, res_hi_lo_lo_lo_53};
  wire [31:0]   res_hi_lo_hi_lo_53 = {dataGroup_21_53, dataGroup_20_53};
  wire [31:0]   res_hi_lo_hi_hi_53 = {dataGroup_23_53, dataGroup_22_53};
  wire [63:0]   res_hi_lo_hi_53 = {res_hi_lo_hi_hi_53, res_hi_lo_hi_lo_53};
  wire [127:0]  res_hi_lo_53 = {res_hi_lo_hi_53, res_hi_lo_lo_53};
  wire [31:0]   res_hi_hi_lo_lo_53 = {dataGroup_25_53, dataGroup_24_53};
  wire [31:0]   res_hi_hi_lo_hi_53 = {dataGroup_27_53, dataGroup_26_53};
  wire [63:0]   res_hi_hi_lo_53 = {res_hi_hi_lo_hi_53, res_hi_hi_lo_lo_53};
  wire [31:0]   res_hi_hi_hi_lo_53 = {dataGroup_29_53, dataGroup_28_53};
  wire [31:0]   res_hi_hi_hi_hi_53 = {dataGroup_31_53, dataGroup_30_53};
  wire [63:0]   res_hi_hi_hi_53 = {res_hi_hi_hi_hi_53, res_hi_hi_hi_lo_53};
  wire [127:0]  res_hi_hi_53 = {res_hi_hi_hi_53, res_hi_hi_lo_53};
  wire [255:0]  res_hi_53 = {res_hi_hi_53, res_hi_lo_53};
  wire [511:0]  res_106 = {res_hi_53, res_lo_53};
  wire [2047:0] dataGroup_lo_2880 = {dataGroup_lo_hi_2880, dataGroup_lo_lo_2880};
  wire [2047:0] dataGroup_hi_2880 = {dataGroup_hi_hi_2880, dataGroup_hi_lo_2880};
  wire [15:0]   dataGroup_0_54 = dataGroup_lo_2880[63:48];
  wire [2047:0] dataGroup_lo_2881 = {dataGroup_lo_hi_2881, dataGroup_lo_lo_2881};
  wire [2047:0] dataGroup_hi_2881 = {dataGroup_hi_hi_2881, dataGroup_hi_lo_2881};
  wire [15:0]   dataGroup_1_54 = dataGroup_lo_2881[159:144];
  wire [2047:0] dataGroup_lo_2882 = {dataGroup_lo_hi_2882, dataGroup_lo_lo_2882};
  wire [2047:0] dataGroup_hi_2882 = {dataGroup_hi_hi_2882, dataGroup_hi_lo_2882};
  wire [15:0]   dataGroup_2_54 = dataGroup_lo_2882[255:240];
  wire [2047:0] dataGroup_lo_2883 = {dataGroup_lo_hi_2883, dataGroup_lo_lo_2883};
  wire [2047:0] dataGroup_hi_2883 = {dataGroup_hi_hi_2883, dataGroup_hi_lo_2883};
  wire [15:0]   dataGroup_3_54 = dataGroup_lo_2883[351:336];
  wire [2047:0] dataGroup_lo_2884 = {dataGroup_lo_hi_2884, dataGroup_lo_lo_2884};
  wire [2047:0] dataGroup_hi_2884 = {dataGroup_hi_hi_2884, dataGroup_hi_lo_2884};
  wire [15:0]   dataGroup_4_54 = dataGroup_lo_2884[447:432];
  wire [2047:0] dataGroup_lo_2885 = {dataGroup_lo_hi_2885, dataGroup_lo_lo_2885};
  wire [2047:0] dataGroup_hi_2885 = {dataGroup_hi_hi_2885, dataGroup_hi_lo_2885};
  wire [15:0]   dataGroup_5_54 = dataGroup_lo_2885[543:528];
  wire [2047:0] dataGroup_lo_2886 = {dataGroup_lo_hi_2886, dataGroup_lo_lo_2886};
  wire [2047:0] dataGroup_hi_2886 = {dataGroup_hi_hi_2886, dataGroup_hi_lo_2886};
  wire [15:0]   dataGroup_6_54 = dataGroup_lo_2886[639:624];
  wire [2047:0] dataGroup_lo_2887 = {dataGroup_lo_hi_2887, dataGroup_lo_lo_2887};
  wire [2047:0] dataGroup_hi_2887 = {dataGroup_hi_hi_2887, dataGroup_hi_lo_2887};
  wire [15:0]   dataGroup_7_54 = dataGroup_lo_2887[735:720];
  wire [2047:0] dataGroup_lo_2888 = {dataGroup_lo_hi_2888, dataGroup_lo_lo_2888};
  wire [2047:0] dataGroup_hi_2888 = {dataGroup_hi_hi_2888, dataGroup_hi_lo_2888};
  wire [15:0]   dataGroup_8_54 = dataGroup_lo_2888[831:816];
  wire [2047:0] dataGroup_lo_2889 = {dataGroup_lo_hi_2889, dataGroup_lo_lo_2889};
  wire [2047:0] dataGroup_hi_2889 = {dataGroup_hi_hi_2889, dataGroup_hi_lo_2889};
  wire [15:0]   dataGroup_9_54 = dataGroup_lo_2889[927:912];
  wire [2047:0] dataGroup_lo_2890 = {dataGroup_lo_hi_2890, dataGroup_lo_lo_2890};
  wire [2047:0] dataGroup_hi_2890 = {dataGroup_hi_hi_2890, dataGroup_hi_lo_2890};
  wire [15:0]   dataGroup_10_54 = dataGroup_lo_2890[1023:1008];
  wire [2047:0] dataGroup_lo_2891 = {dataGroup_lo_hi_2891, dataGroup_lo_lo_2891};
  wire [2047:0] dataGroup_hi_2891 = {dataGroup_hi_hi_2891, dataGroup_hi_lo_2891};
  wire [15:0]   dataGroup_11_54 = dataGroup_lo_2891[1119:1104];
  wire [2047:0] dataGroup_lo_2892 = {dataGroup_lo_hi_2892, dataGroup_lo_lo_2892};
  wire [2047:0] dataGroup_hi_2892 = {dataGroup_hi_hi_2892, dataGroup_hi_lo_2892};
  wire [15:0]   dataGroup_12_54 = dataGroup_lo_2892[1215:1200];
  wire [2047:0] dataGroup_lo_2893 = {dataGroup_lo_hi_2893, dataGroup_lo_lo_2893};
  wire [2047:0] dataGroup_hi_2893 = {dataGroup_hi_hi_2893, dataGroup_hi_lo_2893};
  wire [15:0]   dataGroup_13_54 = dataGroup_lo_2893[1311:1296];
  wire [2047:0] dataGroup_lo_2894 = {dataGroup_lo_hi_2894, dataGroup_lo_lo_2894};
  wire [2047:0] dataGroup_hi_2894 = {dataGroup_hi_hi_2894, dataGroup_hi_lo_2894};
  wire [15:0]   dataGroup_14_54 = dataGroup_lo_2894[1407:1392];
  wire [2047:0] dataGroup_lo_2895 = {dataGroup_lo_hi_2895, dataGroup_lo_lo_2895};
  wire [2047:0] dataGroup_hi_2895 = {dataGroup_hi_hi_2895, dataGroup_hi_lo_2895};
  wire [15:0]   dataGroup_15_54 = dataGroup_lo_2895[1503:1488];
  wire [2047:0] dataGroup_lo_2896 = {dataGroup_lo_hi_2896, dataGroup_lo_lo_2896};
  wire [2047:0] dataGroup_hi_2896 = {dataGroup_hi_hi_2896, dataGroup_hi_lo_2896};
  wire [15:0]   dataGroup_16_54 = dataGroup_lo_2896[1599:1584];
  wire [2047:0] dataGroup_lo_2897 = {dataGroup_lo_hi_2897, dataGroup_lo_lo_2897};
  wire [2047:0] dataGroup_hi_2897 = {dataGroup_hi_hi_2897, dataGroup_hi_lo_2897};
  wire [15:0]   dataGroup_17_54 = dataGroup_lo_2897[1695:1680];
  wire [2047:0] dataGroup_lo_2898 = {dataGroup_lo_hi_2898, dataGroup_lo_lo_2898};
  wire [2047:0] dataGroup_hi_2898 = {dataGroup_hi_hi_2898, dataGroup_hi_lo_2898};
  wire [15:0]   dataGroup_18_54 = dataGroup_lo_2898[1791:1776];
  wire [2047:0] dataGroup_lo_2899 = {dataGroup_lo_hi_2899, dataGroup_lo_lo_2899};
  wire [2047:0] dataGroup_hi_2899 = {dataGroup_hi_hi_2899, dataGroup_hi_lo_2899};
  wire [15:0]   dataGroup_19_54 = dataGroup_lo_2899[1887:1872];
  wire [2047:0] dataGroup_lo_2900 = {dataGroup_lo_hi_2900, dataGroup_lo_lo_2900};
  wire [2047:0] dataGroup_hi_2900 = {dataGroup_hi_hi_2900, dataGroup_hi_lo_2900};
  wire [15:0]   dataGroup_20_54 = dataGroup_lo_2900[1983:1968];
  wire [2047:0] dataGroup_lo_2901 = {dataGroup_lo_hi_2901, dataGroup_lo_lo_2901};
  wire [2047:0] dataGroup_hi_2901 = {dataGroup_hi_hi_2901, dataGroup_hi_lo_2901};
  wire [15:0]   dataGroup_21_54 = dataGroup_hi_2901[31:16];
  wire [2047:0] dataGroup_lo_2902 = {dataGroup_lo_hi_2902, dataGroup_lo_lo_2902};
  wire [2047:0] dataGroup_hi_2902 = {dataGroup_hi_hi_2902, dataGroup_hi_lo_2902};
  wire [15:0]   dataGroup_22_54 = dataGroup_hi_2902[127:112];
  wire [2047:0] dataGroup_lo_2903 = {dataGroup_lo_hi_2903, dataGroup_lo_lo_2903};
  wire [2047:0] dataGroup_hi_2903 = {dataGroup_hi_hi_2903, dataGroup_hi_lo_2903};
  wire [15:0]   dataGroup_23_54 = dataGroup_hi_2903[223:208];
  wire [2047:0] dataGroup_lo_2904 = {dataGroup_lo_hi_2904, dataGroup_lo_lo_2904};
  wire [2047:0] dataGroup_hi_2904 = {dataGroup_hi_hi_2904, dataGroup_hi_lo_2904};
  wire [15:0]   dataGroup_24_54 = dataGroup_hi_2904[319:304];
  wire [2047:0] dataGroup_lo_2905 = {dataGroup_lo_hi_2905, dataGroup_lo_lo_2905};
  wire [2047:0] dataGroup_hi_2905 = {dataGroup_hi_hi_2905, dataGroup_hi_lo_2905};
  wire [15:0]   dataGroup_25_54 = dataGroup_hi_2905[415:400];
  wire [2047:0] dataGroup_lo_2906 = {dataGroup_lo_hi_2906, dataGroup_lo_lo_2906};
  wire [2047:0] dataGroup_hi_2906 = {dataGroup_hi_hi_2906, dataGroup_hi_lo_2906};
  wire [15:0]   dataGroup_26_54 = dataGroup_hi_2906[511:496];
  wire [2047:0] dataGroup_lo_2907 = {dataGroup_lo_hi_2907, dataGroup_lo_lo_2907};
  wire [2047:0] dataGroup_hi_2907 = {dataGroup_hi_hi_2907, dataGroup_hi_lo_2907};
  wire [15:0]   dataGroup_27_54 = dataGroup_hi_2907[607:592];
  wire [2047:0] dataGroup_lo_2908 = {dataGroup_lo_hi_2908, dataGroup_lo_lo_2908};
  wire [2047:0] dataGroup_hi_2908 = {dataGroup_hi_hi_2908, dataGroup_hi_lo_2908};
  wire [15:0]   dataGroup_28_54 = dataGroup_hi_2908[703:688];
  wire [2047:0] dataGroup_lo_2909 = {dataGroup_lo_hi_2909, dataGroup_lo_lo_2909};
  wire [2047:0] dataGroup_hi_2909 = {dataGroup_hi_hi_2909, dataGroup_hi_lo_2909};
  wire [15:0]   dataGroup_29_54 = dataGroup_hi_2909[799:784];
  wire [2047:0] dataGroup_lo_2910 = {dataGroup_lo_hi_2910, dataGroup_lo_lo_2910};
  wire [2047:0] dataGroup_hi_2910 = {dataGroup_hi_hi_2910, dataGroup_hi_lo_2910};
  wire [15:0]   dataGroup_30_54 = dataGroup_hi_2910[895:880];
  wire [2047:0] dataGroup_lo_2911 = {dataGroup_lo_hi_2911, dataGroup_lo_lo_2911};
  wire [2047:0] dataGroup_hi_2911 = {dataGroup_hi_hi_2911, dataGroup_hi_lo_2911};
  wire [15:0]   dataGroup_31_54 = dataGroup_hi_2911[991:976];
  wire [31:0]   res_lo_lo_lo_lo_54 = {dataGroup_1_54, dataGroup_0_54};
  wire [31:0]   res_lo_lo_lo_hi_54 = {dataGroup_3_54, dataGroup_2_54};
  wire [63:0]   res_lo_lo_lo_54 = {res_lo_lo_lo_hi_54, res_lo_lo_lo_lo_54};
  wire [31:0]   res_lo_lo_hi_lo_54 = {dataGroup_5_54, dataGroup_4_54};
  wire [31:0]   res_lo_lo_hi_hi_54 = {dataGroup_7_54, dataGroup_6_54};
  wire [63:0]   res_lo_lo_hi_54 = {res_lo_lo_hi_hi_54, res_lo_lo_hi_lo_54};
  wire [127:0]  res_lo_lo_54 = {res_lo_lo_hi_54, res_lo_lo_lo_54};
  wire [31:0]   res_lo_hi_lo_lo_54 = {dataGroup_9_54, dataGroup_8_54};
  wire [31:0]   res_lo_hi_lo_hi_54 = {dataGroup_11_54, dataGroup_10_54};
  wire [63:0]   res_lo_hi_lo_54 = {res_lo_hi_lo_hi_54, res_lo_hi_lo_lo_54};
  wire [31:0]   res_lo_hi_hi_lo_54 = {dataGroup_13_54, dataGroup_12_54};
  wire [31:0]   res_lo_hi_hi_hi_54 = {dataGroup_15_54, dataGroup_14_54};
  wire [63:0]   res_lo_hi_hi_54 = {res_lo_hi_hi_hi_54, res_lo_hi_hi_lo_54};
  wire [127:0]  res_lo_hi_54 = {res_lo_hi_hi_54, res_lo_hi_lo_54};
  wire [255:0]  res_lo_54 = {res_lo_hi_54, res_lo_lo_54};
  wire [31:0]   res_hi_lo_lo_lo_54 = {dataGroup_17_54, dataGroup_16_54};
  wire [31:0]   res_hi_lo_lo_hi_54 = {dataGroup_19_54, dataGroup_18_54};
  wire [63:0]   res_hi_lo_lo_54 = {res_hi_lo_lo_hi_54, res_hi_lo_lo_lo_54};
  wire [31:0]   res_hi_lo_hi_lo_54 = {dataGroup_21_54, dataGroup_20_54};
  wire [31:0]   res_hi_lo_hi_hi_54 = {dataGroup_23_54, dataGroup_22_54};
  wire [63:0]   res_hi_lo_hi_54 = {res_hi_lo_hi_hi_54, res_hi_lo_hi_lo_54};
  wire [127:0]  res_hi_lo_54 = {res_hi_lo_hi_54, res_hi_lo_lo_54};
  wire [31:0]   res_hi_hi_lo_lo_54 = {dataGroup_25_54, dataGroup_24_54};
  wire [31:0]   res_hi_hi_lo_hi_54 = {dataGroup_27_54, dataGroup_26_54};
  wire [63:0]   res_hi_hi_lo_54 = {res_hi_hi_lo_hi_54, res_hi_hi_lo_lo_54};
  wire [31:0]   res_hi_hi_hi_lo_54 = {dataGroup_29_54, dataGroup_28_54};
  wire [31:0]   res_hi_hi_hi_hi_54 = {dataGroup_31_54, dataGroup_30_54};
  wire [63:0]   res_hi_hi_hi_54 = {res_hi_hi_hi_hi_54, res_hi_hi_hi_lo_54};
  wire [127:0]  res_hi_hi_54 = {res_hi_hi_hi_54, res_hi_hi_lo_54};
  wire [255:0]  res_hi_54 = {res_hi_hi_54, res_hi_lo_54};
  wire [511:0]  res_107 = {res_hi_54, res_lo_54};
  wire [2047:0] dataGroup_lo_2912 = {dataGroup_lo_hi_2912, dataGroup_lo_lo_2912};
  wire [2047:0] dataGroup_hi_2912 = {dataGroup_hi_hi_2912, dataGroup_hi_lo_2912};
  wire [15:0]   dataGroup_0_55 = dataGroup_lo_2912[79:64];
  wire [2047:0] dataGroup_lo_2913 = {dataGroup_lo_hi_2913, dataGroup_lo_lo_2913};
  wire [2047:0] dataGroup_hi_2913 = {dataGroup_hi_hi_2913, dataGroup_hi_lo_2913};
  wire [15:0]   dataGroup_1_55 = dataGroup_lo_2913[175:160];
  wire [2047:0] dataGroup_lo_2914 = {dataGroup_lo_hi_2914, dataGroup_lo_lo_2914};
  wire [2047:0] dataGroup_hi_2914 = {dataGroup_hi_hi_2914, dataGroup_hi_lo_2914};
  wire [15:0]   dataGroup_2_55 = dataGroup_lo_2914[271:256];
  wire [2047:0] dataGroup_lo_2915 = {dataGroup_lo_hi_2915, dataGroup_lo_lo_2915};
  wire [2047:0] dataGroup_hi_2915 = {dataGroup_hi_hi_2915, dataGroup_hi_lo_2915};
  wire [15:0]   dataGroup_3_55 = dataGroup_lo_2915[367:352];
  wire [2047:0] dataGroup_lo_2916 = {dataGroup_lo_hi_2916, dataGroup_lo_lo_2916};
  wire [2047:0] dataGroup_hi_2916 = {dataGroup_hi_hi_2916, dataGroup_hi_lo_2916};
  wire [15:0]   dataGroup_4_55 = dataGroup_lo_2916[463:448];
  wire [2047:0] dataGroup_lo_2917 = {dataGroup_lo_hi_2917, dataGroup_lo_lo_2917};
  wire [2047:0] dataGroup_hi_2917 = {dataGroup_hi_hi_2917, dataGroup_hi_lo_2917};
  wire [15:0]   dataGroup_5_55 = dataGroup_lo_2917[559:544];
  wire [2047:0] dataGroup_lo_2918 = {dataGroup_lo_hi_2918, dataGroup_lo_lo_2918};
  wire [2047:0] dataGroup_hi_2918 = {dataGroup_hi_hi_2918, dataGroup_hi_lo_2918};
  wire [15:0]   dataGroup_6_55 = dataGroup_lo_2918[655:640];
  wire [2047:0] dataGroup_lo_2919 = {dataGroup_lo_hi_2919, dataGroup_lo_lo_2919};
  wire [2047:0] dataGroup_hi_2919 = {dataGroup_hi_hi_2919, dataGroup_hi_lo_2919};
  wire [15:0]   dataGroup_7_55 = dataGroup_lo_2919[751:736];
  wire [2047:0] dataGroup_lo_2920 = {dataGroup_lo_hi_2920, dataGroup_lo_lo_2920};
  wire [2047:0] dataGroup_hi_2920 = {dataGroup_hi_hi_2920, dataGroup_hi_lo_2920};
  wire [15:0]   dataGroup_8_55 = dataGroup_lo_2920[847:832];
  wire [2047:0] dataGroup_lo_2921 = {dataGroup_lo_hi_2921, dataGroup_lo_lo_2921};
  wire [2047:0] dataGroup_hi_2921 = {dataGroup_hi_hi_2921, dataGroup_hi_lo_2921};
  wire [15:0]   dataGroup_9_55 = dataGroup_lo_2921[943:928];
  wire [2047:0] dataGroup_lo_2922 = {dataGroup_lo_hi_2922, dataGroup_lo_lo_2922};
  wire [2047:0] dataGroup_hi_2922 = {dataGroup_hi_hi_2922, dataGroup_hi_lo_2922};
  wire [15:0]   dataGroup_10_55 = dataGroup_lo_2922[1039:1024];
  wire [2047:0] dataGroup_lo_2923 = {dataGroup_lo_hi_2923, dataGroup_lo_lo_2923};
  wire [2047:0] dataGroup_hi_2923 = {dataGroup_hi_hi_2923, dataGroup_hi_lo_2923};
  wire [15:0]   dataGroup_11_55 = dataGroup_lo_2923[1135:1120];
  wire [2047:0] dataGroup_lo_2924 = {dataGroup_lo_hi_2924, dataGroup_lo_lo_2924};
  wire [2047:0] dataGroup_hi_2924 = {dataGroup_hi_hi_2924, dataGroup_hi_lo_2924};
  wire [15:0]   dataGroup_12_55 = dataGroup_lo_2924[1231:1216];
  wire [2047:0] dataGroup_lo_2925 = {dataGroup_lo_hi_2925, dataGroup_lo_lo_2925};
  wire [2047:0] dataGroup_hi_2925 = {dataGroup_hi_hi_2925, dataGroup_hi_lo_2925};
  wire [15:0]   dataGroup_13_55 = dataGroup_lo_2925[1327:1312];
  wire [2047:0] dataGroup_lo_2926 = {dataGroup_lo_hi_2926, dataGroup_lo_lo_2926};
  wire [2047:0] dataGroup_hi_2926 = {dataGroup_hi_hi_2926, dataGroup_hi_lo_2926};
  wire [15:0]   dataGroup_14_55 = dataGroup_lo_2926[1423:1408];
  wire [2047:0] dataGroup_lo_2927 = {dataGroup_lo_hi_2927, dataGroup_lo_lo_2927};
  wire [2047:0] dataGroup_hi_2927 = {dataGroup_hi_hi_2927, dataGroup_hi_lo_2927};
  wire [15:0]   dataGroup_15_55 = dataGroup_lo_2927[1519:1504];
  wire [2047:0] dataGroup_lo_2928 = {dataGroup_lo_hi_2928, dataGroup_lo_lo_2928};
  wire [2047:0] dataGroup_hi_2928 = {dataGroup_hi_hi_2928, dataGroup_hi_lo_2928};
  wire [15:0]   dataGroup_16_55 = dataGroup_lo_2928[1615:1600];
  wire [2047:0] dataGroup_lo_2929 = {dataGroup_lo_hi_2929, dataGroup_lo_lo_2929};
  wire [2047:0] dataGroup_hi_2929 = {dataGroup_hi_hi_2929, dataGroup_hi_lo_2929};
  wire [15:0]   dataGroup_17_55 = dataGroup_lo_2929[1711:1696];
  wire [2047:0] dataGroup_lo_2930 = {dataGroup_lo_hi_2930, dataGroup_lo_lo_2930};
  wire [2047:0] dataGroup_hi_2930 = {dataGroup_hi_hi_2930, dataGroup_hi_lo_2930};
  wire [15:0]   dataGroup_18_55 = dataGroup_lo_2930[1807:1792];
  wire [2047:0] dataGroup_lo_2931 = {dataGroup_lo_hi_2931, dataGroup_lo_lo_2931};
  wire [2047:0] dataGroup_hi_2931 = {dataGroup_hi_hi_2931, dataGroup_hi_lo_2931};
  wire [15:0]   dataGroup_19_55 = dataGroup_lo_2931[1903:1888];
  wire [2047:0] dataGroup_lo_2932 = {dataGroup_lo_hi_2932, dataGroup_lo_lo_2932};
  wire [2047:0] dataGroup_hi_2932 = {dataGroup_hi_hi_2932, dataGroup_hi_lo_2932};
  wire [15:0]   dataGroup_20_55 = dataGroup_lo_2932[1999:1984];
  wire [2047:0] dataGroup_lo_2933 = {dataGroup_lo_hi_2933, dataGroup_lo_lo_2933};
  wire [2047:0] dataGroup_hi_2933 = {dataGroup_hi_hi_2933, dataGroup_hi_lo_2933};
  wire [15:0]   dataGroup_21_55 = dataGroup_hi_2933[47:32];
  wire [2047:0] dataGroup_lo_2934 = {dataGroup_lo_hi_2934, dataGroup_lo_lo_2934};
  wire [2047:0] dataGroup_hi_2934 = {dataGroup_hi_hi_2934, dataGroup_hi_lo_2934};
  wire [15:0]   dataGroup_22_55 = dataGroup_hi_2934[143:128];
  wire [2047:0] dataGroup_lo_2935 = {dataGroup_lo_hi_2935, dataGroup_lo_lo_2935};
  wire [2047:0] dataGroup_hi_2935 = {dataGroup_hi_hi_2935, dataGroup_hi_lo_2935};
  wire [15:0]   dataGroup_23_55 = dataGroup_hi_2935[239:224];
  wire [2047:0] dataGroup_lo_2936 = {dataGroup_lo_hi_2936, dataGroup_lo_lo_2936};
  wire [2047:0] dataGroup_hi_2936 = {dataGroup_hi_hi_2936, dataGroup_hi_lo_2936};
  wire [15:0]   dataGroup_24_55 = dataGroup_hi_2936[335:320];
  wire [2047:0] dataGroup_lo_2937 = {dataGroup_lo_hi_2937, dataGroup_lo_lo_2937};
  wire [2047:0] dataGroup_hi_2937 = {dataGroup_hi_hi_2937, dataGroup_hi_lo_2937};
  wire [15:0]   dataGroup_25_55 = dataGroup_hi_2937[431:416];
  wire [2047:0] dataGroup_lo_2938 = {dataGroup_lo_hi_2938, dataGroup_lo_lo_2938};
  wire [2047:0] dataGroup_hi_2938 = {dataGroup_hi_hi_2938, dataGroup_hi_lo_2938};
  wire [15:0]   dataGroup_26_55 = dataGroup_hi_2938[527:512];
  wire [2047:0] dataGroup_lo_2939 = {dataGroup_lo_hi_2939, dataGroup_lo_lo_2939};
  wire [2047:0] dataGroup_hi_2939 = {dataGroup_hi_hi_2939, dataGroup_hi_lo_2939};
  wire [15:0]   dataGroup_27_55 = dataGroup_hi_2939[623:608];
  wire [2047:0] dataGroup_lo_2940 = {dataGroup_lo_hi_2940, dataGroup_lo_lo_2940};
  wire [2047:0] dataGroup_hi_2940 = {dataGroup_hi_hi_2940, dataGroup_hi_lo_2940};
  wire [15:0]   dataGroup_28_55 = dataGroup_hi_2940[719:704];
  wire [2047:0] dataGroup_lo_2941 = {dataGroup_lo_hi_2941, dataGroup_lo_lo_2941};
  wire [2047:0] dataGroup_hi_2941 = {dataGroup_hi_hi_2941, dataGroup_hi_lo_2941};
  wire [15:0]   dataGroup_29_55 = dataGroup_hi_2941[815:800];
  wire [2047:0] dataGroup_lo_2942 = {dataGroup_lo_hi_2942, dataGroup_lo_lo_2942};
  wire [2047:0] dataGroup_hi_2942 = {dataGroup_hi_hi_2942, dataGroup_hi_lo_2942};
  wire [15:0]   dataGroup_30_55 = dataGroup_hi_2942[911:896];
  wire [2047:0] dataGroup_lo_2943 = {dataGroup_lo_hi_2943, dataGroup_lo_lo_2943};
  wire [2047:0] dataGroup_hi_2943 = {dataGroup_hi_hi_2943, dataGroup_hi_lo_2943};
  wire [15:0]   dataGroup_31_55 = dataGroup_hi_2943[1007:992];
  wire [31:0]   res_lo_lo_lo_lo_55 = {dataGroup_1_55, dataGroup_0_55};
  wire [31:0]   res_lo_lo_lo_hi_55 = {dataGroup_3_55, dataGroup_2_55};
  wire [63:0]   res_lo_lo_lo_55 = {res_lo_lo_lo_hi_55, res_lo_lo_lo_lo_55};
  wire [31:0]   res_lo_lo_hi_lo_55 = {dataGroup_5_55, dataGroup_4_55};
  wire [31:0]   res_lo_lo_hi_hi_55 = {dataGroup_7_55, dataGroup_6_55};
  wire [63:0]   res_lo_lo_hi_55 = {res_lo_lo_hi_hi_55, res_lo_lo_hi_lo_55};
  wire [127:0]  res_lo_lo_55 = {res_lo_lo_hi_55, res_lo_lo_lo_55};
  wire [31:0]   res_lo_hi_lo_lo_55 = {dataGroup_9_55, dataGroup_8_55};
  wire [31:0]   res_lo_hi_lo_hi_55 = {dataGroup_11_55, dataGroup_10_55};
  wire [63:0]   res_lo_hi_lo_55 = {res_lo_hi_lo_hi_55, res_lo_hi_lo_lo_55};
  wire [31:0]   res_lo_hi_hi_lo_55 = {dataGroup_13_55, dataGroup_12_55};
  wire [31:0]   res_lo_hi_hi_hi_55 = {dataGroup_15_55, dataGroup_14_55};
  wire [63:0]   res_lo_hi_hi_55 = {res_lo_hi_hi_hi_55, res_lo_hi_hi_lo_55};
  wire [127:0]  res_lo_hi_55 = {res_lo_hi_hi_55, res_lo_hi_lo_55};
  wire [255:0]  res_lo_55 = {res_lo_hi_55, res_lo_lo_55};
  wire [31:0]   res_hi_lo_lo_lo_55 = {dataGroup_17_55, dataGroup_16_55};
  wire [31:0]   res_hi_lo_lo_hi_55 = {dataGroup_19_55, dataGroup_18_55};
  wire [63:0]   res_hi_lo_lo_55 = {res_hi_lo_lo_hi_55, res_hi_lo_lo_lo_55};
  wire [31:0]   res_hi_lo_hi_lo_55 = {dataGroup_21_55, dataGroup_20_55};
  wire [31:0]   res_hi_lo_hi_hi_55 = {dataGroup_23_55, dataGroup_22_55};
  wire [63:0]   res_hi_lo_hi_55 = {res_hi_lo_hi_hi_55, res_hi_lo_hi_lo_55};
  wire [127:0]  res_hi_lo_55 = {res_hi_lo_hi_55, res_hi_lo_lo_55};
  wire [31:0]   res_hi_hi_lo_lo_55 = {dataGroup_25_55, dataGroup_24_55};
  wire [31:0]   res_hi_hi_lo_hi_55 = {dataGroup_27_55, dataGroup_26_55};
  wire [63:0]   res_hi_hi_lo_55 = {res_hi_hi_lo_hi_55, res_hi_hi_lo_lo_55};
  wire [31:0]   res_hi_hi_hi_lo_55 = {dataGroup_29_55, dataGroup_28_55};
  wire [31:0]   res_hi_hi_hi_hi_55 = {dataGroup_31_55, dataGroup_30_55};
  wire [63:0]   res_hi_hi_hi_55 = {res_hi_hi_hi_hi_55, res_hi_hi_hi_lo_55};
  wire [127:0]  res_hi_hi_55 = {res_hi_hi_hi_55, res_hi_hi_lo_55};
  wire [255:0]  res_hi_55 = {res_hi_hi_55, res_hi_lo_55};
  wire [511:0]  res_108 = {res_hi_55, res_lo_55};
  wire [2047:0] dataGroup_lo_2944 = {dataGroup_lo_hi_2944, dataGroup_lo_lo_2944};
  wire [2047:0] dataGroup_hi_2944 = {dataGroup_hi_hi_2944, dataGroup_hi_lo_2944};
  wire [15:0]   dataGroup_0_56 = dataGroup_lo_2944[95:80];
  wire [2047:0] dataGroup_lo_2945 = {dataGroup_lo_hi_2945, dataGroup_lo_lo_2945};
  wire [2047:0] dataGroup_hi_2945 = {dataGroup_hi_hi_2945, dataGroup_hi_lo_2945};
  wire [15:0]   dataGroup_1_56 = dataGroup_lo_2945[191:176];
  wire [2047:0] dataGroup_lo_2946 = {dataGroup_lo_hi_2946, dataGroup_lo_lo_2946};
  wire [2047:0] dataGroup_hi_2946 = {dataGroup_hi_hi_2946, dataGroup_hi_lo_2946};
  wire [15:0]   dataGroup_2_56 = dataGroup_lo_2946[287:272];
  wire [2047:0] dataGroup_lo_2947 = {dataGroup_lo_hi_2947, dataGroup_lo_lo_2947};
  wire [2047:0] dataGroup_hi_2947 = {dataGroup_hi_hi_2947, dataGroup_hi_lo_2947};
  wire [15:0]   dataGroup_3_56 = dataGroup_lo_2947[383:368];
  wire [2047:0] dataGroup_lo_2948 = {dataGroup_lo_hi_2948, dataGroup_lo_lo_2948};
  wire [2047:0] dataGroup_hi_2948 = {dataGroup_hi_hi_2948, dataGroup_hi_lo_2948};
  wire [15:0]   dataGroup_4_56 = dataGroup_lo_2948[479:464];
  wire [2047:0] dataGroup_lo_2949 = {dataGroup_lo_hi_2949, dataGroup_lo_lo_2949};
  wire [2047:0] dataGroup_hi_2949 = {dataGroup_hi_hi_2949, dataGroup_hi_lo_2949};
  wire [15:0]   dataGroup_5_56 = dataGroup_lo_2949[575:560];
  wire [2047:0] dataGroup_lo_2950 = {dataGroup_lo_hi_2950, dataGroup_lo_lo_2950};
  wire [2047:0] dataGroup_hi_2950 = {dataGroup_hi_hi_2950, dataGroup_hi_lo_2950};
  wire [15:0]   dataGroup_6_56 = dataGroup_lo_2950[671:656];
  wire [2047:0] dataGroup_lo_2951 = {dataGroup_lo_hi_2951, dataGroup_lo_lo_2951};
  wire [2047:0] dataGroup_hi_2951 = {dataGroup_hi_hi_2951, dataGroup_hi_lo_2951};
  wire [15:0]   dataGroup_7_56 = dataGroup_lo_2951[767:752];
  wire [2047:0] dataGroup_lo_2952 = {dataGroup_lo_hi_2952, dataGroup_lo_lo_2952};
  wire [2047:0] dataGroup_hi_2952 = {dataGroup_hi_hi_2952, dataGroup_hi_lo_2952};
  wire [15:0]   dataGroup_8_56 = dataGroup_lo_2952[863:848];
  wire [2047:0] dataGroup_lo_2953 = {dataGroup_lo_hi_2953, dataGroup_lo_lo_2953};
  wire [2047:0] dataGroup_hi_2953 = {dataGroup_hi_hi_2953, dataGroup_hi_lo_2953};
  wire [15:0]   dataGroup_9_56 = dataGroup_lo_2953[959:944];
  wire [2047:0] dataGroup_lo_2954 = {dataGroup_lo_hi_2954, dataGroup_lo_lo_2954};
  wire [2047:0] dataGroup_hi_2954 = {dataGroup_hi_hi_2954, dataGroup_hi_lo_2954};
  wire [15:0]   dataGroup_10_56 = dataGroup_lo_2954[1055:1040];
  wire [2047:0] dataGroup_lo_2955 = {dataGroup_lo_hi_2955, dataGroup_lo_lo_2955};
  wire [2047:0] dataGroup_hi_2955 = {dataGroup_hi_hi_2955, dataGroup_hi_lo_2955};
  wire [15:0]   dataGroup_11_56 = dataGroup_lo_2955[1151:1136];
  wire [2047:0] dataGroup_lo_2956 = {dataGroup_lo_hi_2956, dataGroup_lo_lo_2956};
  wire [2047:0] dataGroup_hi_2956 = {dataGroup_hi_hi_2956, dataGroup_hi_lo_2956};
  wire [15:0]   dataGroup_12_56 = dataGroup_lo_2956[1247:1232];
  wire [2047:0] dataGroup_lo_2957 = {dataGroup_lo_hi_2957, dataGroup_lo_lo_2957};
  wire [2047:0] dataGroup_hi_2957 = {dataGroup_hi_hi_2957, dataGroup_hi_lo_2957};
  wire [15:0]   dataGroup_13_56 = dataGroup_lo_2957[1343:1328];
  wire [2047:0] dataGroup_lo_2958 = {dataGroup_lo_hi_2958, dataGroup_lo_lo_2958};
  wire [2047:0] dataGroup_hi_2958 = {dataGroup_hi_hi_2958, dataGroup_hi_lo_2958};
  wire [15:0]   dataGroup_14_56 = dataGroup_lo_2958[1439:1424];
  wire [2047:0] dataGroup_lo_2959 = {dataGroup_lo_hi_2959, dataGroup_lo_lo_2959};
  wire [2047:0] dataGroup_hi_2959 = {dataGroup_hi_hi_2959, dataGroup_hi_lo_2959};
  wire [15:0]   dataGroup_15_56 = dataGroup_lo_2959[1535:1520];
  wire [2047:0] dataGroup_lo_2960 = {dataGroup_lo_hi_2960, dataGroup_lo_lo_2960};
  wire [2047:0] dataGroup_hi_2960 = {dataGroup_hi_hi_2960, dataGroup_hi_lo_2960};
  wire [15:0]   dataGroup_16_56 = dataGroup_lo_2960[1631:1616];
  wire [2047:0] dataGroup_lo_2961 = {dataGroup_lo_hi_2961, dataGroup_lo_lo_2961};
  wire [2047:0] dataGroup_hi_2961 = {dataGroup_hi_hi_2961, dataGroup_hi_lo_2961};
  wire [15:0]   dataGroup_17_56 = dataGroup_lo_2961[1727:1712];
  wire [2047:0] dataGroup_lo_2962 = {dataGroup_lo_hi_2962, dataGroup_lo_lo_2962};
  wire [2047:0] dataGroup_hi_2962 = {dataGroup_hi_hi_2962, dataGroup_hi_lo_2962};
  wire [15:0]   dataGroup_18_56 = dataGroup_lo_2962[1823:1808];
  wire [2047:0] dataGroup_lo_2963 = {dataGroup_lo_hi_2963, dataGroup_lo_lo_2963};
  wire [2047:0] dataGroup_hi_2963 = {dataGroup_hi_hi_2963, dataGroup_hi_lo_2963};
  wire [15:0]   dataGroup_19_56 = dataGroup_lo_2963[1919:1904];
  wire [2047:0] dataGroup_lo_2964 = {dataGroup_lo_hi_2964, dataGroup_lo_lo_2964};
  wire [2047:0] dataGroup_hi_2964 = {dataGroup_hi_hi_2964, dataGroup_hi_lo_2964};
  wire [15:0]   dataGroup_20_56 = dataGroup_lo_2964[2015:2000];
  wire [2047:0] dataGroup_lo_2965 = {dataGroup_lo_hi_2965, dataGroup_lo_lo_2965};
  wire [2047:0] dataGroup_hi_2965 = {dataGroup_hi_hi_2965, dataGroup_hi_lo_2965};
  wire [15:0]   dataGroup_21_56 = dataGroup_hi_2965[63:48];
  wire [2047:0] dataGroup_lo_2966 = {dataGroup_lo_hi_2966, dataGroup_lo_lo_2966};
  wire [2047:0] dataGroup_hi_2966 = {dataGroup_hi_hi_2966, dataGroup_hi_lo_2966};
  wire [15:0]   dataGroup_22_56 = dataGroup_hi_2966[159:144];
  wire [2047:0] dataGroup_lo_2967 = {dataGroup_lo_hi_2967, dataGroup_lo_lo_2967};
  wire [2047:0] dataGroup_hi_2967 = {dataGroup_hi_hi_2967, dataGroup_hi_lo_2967};
  wire [15:0]   dataGroup_23_56 = dataGroup_hi_2967[255:240];
  wire [2047:0] dataGroup_lo_2968 = {dataGroup_lo_hi_2968, dataGroup_lo_lo_2968};
  wire [2047:0] dataGroup_hi_2968 = {dataGroup_hi_hi_2968, dataGroup_hi_lo_2968};
  wire [15:0]   dataGroup_24_56 = dataGroup_hi_2968[351:336];
  wire [2047:0] dataGroup_lo_2969 = {dataGroup_lo_hi_2969, dataGroup_lo_lo_2969};
  wire [2047:0] dataGroup_hi_2969 = {dataGroup_hi_hi_2969, dataGroup_hi_lo_2969};
  wire [15:0]   dataGroup_25_56 = dataGroup_hi_2969[447:432];
  wire [2047:0] dataGroup_lo_2970 = {dataGroup_lo_hi_2970, dataGroup_lo_lo_2970};
  wire [2047:0] dataGroup_hi_2970 = {dataGroup_hi_hi_2970, dataGroup_hi_lo_2970};
  wire [15:0]   dataGroup_26_56 = dataGroup_hi_2970[543:528];
  wire [2047:0] dataGroup_lo_2971 = {dataGroup_lo_hi_2971, dataGroup_lo_lo_2971};
  wire [2047:0] dataGroup_hi_2971 = {dataGroup_hi_hi_2971, dataGroup_hi_lo_2971};
  wire [15:0]   dataGroup_27_56 = dataGroup_hi_2971[639:624];
  wire [2047:0] dataGroup_lo_2972 = {dataGroup_lo_hi_2972, dataGroup_lo_lo_2972};
  wire [2047:0] dataGroup_hi_2972 = {dataGroup_hi_hi_2972, dataGroup_hi_lo_2972};
  wire [15:0]   dataGroup_28_56 = dataGroup_hi_2972[735:720];
  wire [2047:0] dataGroup_lo_2973 = {dataGroup_lo_hi_2973, dataGroup_lo_lo_2973};
  wire [2047:0] dataGroup_hi_2973 = {dataGroup_hi_hi_2973, dataGroup_hi_lo_2973};
  wire [15:0]   dataGroup_29_56 = dataGroup_hi_2973[831:816];
  wire [2047:0] dataGroup_lo_2974 = {dataGroup_lo_hi_2974, dataGroup_lo_lo_2974};
  wire [2047:0] dataGroup_hi_2974 = {dataGroup_hi_hi_2974, dataGroup_hi_lo_2974};
  wire [15:0]   dataGroup_30_56 = dataGroup_hi_2974[927:912];
  wire [2047:0] dataGroup_lo_2975 = {dataGroup_lo_hi_2975, dataGroup_lo_lo_2975};
  wire [2047:0] dataGroup_hi_2975 = {dataGroup_hi_hi_2975, dataGroup_hi_lo_2975};
  wire [15:0]   dataGroup_31_56 = dataGroup_hi_2975[1023:1008];
  wire [31:0]   res_lo_lo_lo_lo_56 = {dataGroup_1_56, dataGroup_0_56};
  wire [31:0]   res_lo_lo_lo_hi_56 = {dataGroup_3_56, dataGroup_2_56};
  wire [63:0]   res_lo_lo_lo_56 = {res_lo_lo_lo_hi_56, res_lo_lo_lo_lo_56};
  wire [31:0]   res_lo_lo_hi_lo_56 = {dataGroup_5_56, dataGroup_4_56};
  wire [31:0]   res_lo_lo_hi_hi_56 = {dataGroup_7_56, dataGroup_6_56};
  wire [63:0]   res_lo_lo_hi_56 = {res_lo_lo_hi_hi_56, res_lo_lo_hi_lo_56};
  wire [127:0]  res_lo_lo_56 = {res_lo_lo_hi_56, res_lo_lo_lo_56};
  wire [31:0]   res_lo_hi_lo_lo_56 = {dataGroup_9_56, dataGroup_8_56};
  wire [31:0]   res_lo_hi_lo_hi_56 = {dataGroup_11_56, dataGroup_10_56};
  wire [63:0]   res_lo_hi_lo_56 = {res_lo_hi_lo_hi_56, res_lo_hi_lo_lo_56};
  wire [31:0]   res_lo_hi_hi_lo_56 = {dataGroup_13_56, dataGroup_12_56};
  wire [31:0]   res_lo_hi_hi_hi_56 = {dataGroup_15_56, dataGroup_14_56};
  wire [63:0]   res_lo_hi_hi_56 = {res_lo_hi_hi_hi_56, res_lo_hi_hi_lo_56};
  wire [127:0]  res_lo_hi_56 = {res_lo_hi_hi_56, res_lo_hi_lo_56};
  wire [255:0]  res_lo_56 = {res_lo_hi_56, res_lo_lo_56};
  wire [31:0]   res_hi_lo_lo_lo_56 = {dataGroup_17_56, dataGroup_16_56};
  wire [31:0]   res_hi_lo_lo_hi_56 = {dataGroup_19_56, dataGroup_18_56};
  wire [63:0]   res_hi_lo_lo_56 = {res_hi_lo_lo_hi_56, res_hi_lo_lo_lo_56};
  wire [31:0]   res_hi_lo_hi_lo_56 = {dataGroup_21_56, dataGroup_20_56};
  wire [31:0]   res_hi_lo_hi_hi_56 = {dataGroup_23_56, dataGroup_22_56};
  wire [63:0]   res_hi_lo_hi_56 = {res_hi_lo_hi_hi_56, res_hi_lo_hi_lo_56};
  wire [127:0]  res_hi_lo_56 = {res_hi_lo_hi_56, res_hi_lo_lo_56};
  wire [31:0]   res_hi_hi_lo_lo_56 = {dataGroup_25_56, dataGroup_24_56};
  wire [31:0]   res_hi_hi_lo_hi_56 = {dataGroup_27_56, dataGroup_26_56};
  wire [63:0]   res_hi_hi_lo_56 = {res_hi_hi_lo_hi_56, res_hi_hi_lo_lo_56};
  wire [31:0]   res_hi_hi_hi_lo_56 = {dataGroup_29_56, dataGroup_28_56};
  wire [31:0]   res_hi_hi_hi_hi_56 = {dataGroup_31_56, dataGroup_30_56};
  wire [63:0]   res_hi_hi_hi_56 = {res_hi_hi_hi_hi_56, res_hi_hi_hi_lo_56};
  wire [127:0]  res_hi_hi_56 = {res_hi_hi_hi_56, res_hi_hi_lo_56};
  wire [255:0]  res_hi_56 = {res_hi_hi_56, res_hi_lo_56};
  wire [511:0]  res_109 = {res_hi_56, res_lo_56};
  wire [1023:0] lo_lo_13 = {res_105, res_104};
  wire [1023:0] lo_hi_13 = {res_107, res_106};
  wire [2047:0] lo_13 = {lo_hi_13, lo_lo_13};
  wire [1023:0] hi_lo_13 = {res_109, res_108};
  wire [2047:0] hi_13 = {1024'h0, hi_lo_13};
  wire [4095:0] regroupLoadData_1_5 = {hi_13, lo_13};
  wire [2047:0] dataGroup_lo_2976 = {dataGroup_lo_hi_2976, dataGroup_lo_lo_2976};
  wire [2047:0] dataGroup_hi_2976 = {dataGroup_hi_hi_2976, dataGroup_hi_lo_2976};
  wire [15:0]   dataGroup_0_57 = dataGroup_lo_2976[15:0];
  wire [2047:0] dataGroup_lo_2977 = {dataGroup_lo_hi_2977, dataGroup_lo_lo_2977};
  wire [2047:0] dataGroup_hi_2977 = {dataGroup_hi_hi_2977, dataGroup_hi_lo_2977};
  wire [15:0]   dataGroup_1_57 = dataGroup_lo_2977[127:112];
  wire [2047:0] dataGroup_lo_2978 = {dataGroup_lo_hi_2978, dataGroup_lo_lo_2978};
  wire [2047:0] dataGroup_hi_2978 = {dataGroup_hi_hi_2978, dataGroup_hi_lo_2978};
  wire [15:0]   dataGroup_2_57 = dataGroup_lo_2978[239:224];
  wire [2047:0] dataGroup_lo_2979 = {dataGroup_lo_hi_2979, dataGroup_lo_lo_2979};
  wire [2047:0] dataGroup_hi_2979 = {dataGroup_hi_hi_2979, dataGroup_hi_lo_2979};
  wire [15:0]   dataGroup_3_57 = dataGroup_lo_2979[351:336];
  wire [2047:0] dataGroup_lo_2980 = {dataGroup_lo_hi_2980, dataGroup_lo_lo_2980};
  wire [2047:0] dataGroup_hi_2980 = {dataGroup_hi_hi_2980, dataGroup_hi_lo_2980};
  wire [15:0]   dataGroup_4_57 = dataGroup_lo_2980[463:448];
  wire [2047:0] dataGroup_lo_2981 = {dataGroup_lo_hi_2981, dataGroup_lo_lo_2981};
  wire [2047:0] dataGroup_hi_2981 = {dataGroup_hi_hi_2981, dataGroup_hi_lo_2981};
  wire [15:0]   dataGroup_5_57 = dataGroup_lo_2981[575:560];
  wire [2047:0] dataGroup_lo_2982 = {dataGroup_lo_hi_2982, dataGroup_lo_lo_2982};
  wire [2047:0] dataGroup_hi_2982 = {dataGroup_hi_hi_2982, dataGroup_hi_lo_2982};
  wire [15:0]   dataGroup_6_57 = dataGroup_lo_2982[687:672];
  wire [2047:0] dataGroup_lo_2983 = {dataGroup_lo_hi_2983, dataGroup_lo_lo_2983};
  wire [2047:0] dataGroup_hi_2983 = {dataGroup_hi_hi_2983, dataGroup_hi_lo_2983};
  wire [15:0]   dataGroup_7_57 = dataGroup_lo_2983[799:784];
  wire [2047:0] dataGroup_lo_2984 = {dataGroup_lo_hi_2984, dataGroup_lo_lo_2984};
  wire [2047:0] dataGroup_hi_2984 = {dataGroup_hi_hi_2984, dataGroup_hi_lo_2984};
  wire [15:0]   dataGroup_8_57 = dataGroup_lo_2984[911:896];
  wire [2047:0] dataGroup_lo_2985 = {dataGroup_lo_hi_2985, dataGroup_lo_lo_2985};
  wire [2047:0] dataGroup_hi_2985 = {dataGroup_hi_hi_2985, dataGroup_hi_lo_2985};
  wire [15:0]   dataGroup_9_57 = dataGroup_lo_2985[1023:1008];
  wire [2047:0] dataGroup_lo_2986 = {dataGroup_lo_hi_2986, dataGroup_lo_lo_2986};
  wire [2047:0] dataGroup_hi_2986 = {dataGroup_hi_hi_2986, dataGroup_hi_lo_2986};
  wire [15:0]   dataGroup_10_57 = dataGroup_lo_2986[1135:1120];
  wire [2047:0] dataGroup_lo_2987 = {dataGroup_lo_hi_2987, dataGroup_lo_lo_2987};
  wire [2047:0] dataGroup_hi_2987 = {dataGroup_hi_hi_2987, dataGroup_hi_lo_2987};
  wire [15:0]   dataGroup_11_57 = dataGroup_lo_2987[1247:1232];
  wire [2047:0] dataGroup_lo_2988 = {dataGroup_lo_hi_2988, dataGroup_lo_lo_2988};
  wire [2047:0] dataGroup_hi_2988 = {dataGroup_hi_hi_2988, dataGroup_hi_lo_2988};
  wire [15:0]   dataGroup_12_57 = dataGroup_lo_2988[1359:1344];
  wire [2047:0] dataGroup_lo_2989 = {dataGroup_lo_hi_2989, dataGroup_lo_lo_2989};
  wire [2047:0] dataGroup_hi_2989 = {dataGroup_hi_hi_2989, dataGroup_hi_lo_2989};
  wire [15:0]   dataGroup_13_57 = dataGroup_lo_2989[1471:1456];
  wire [2047:0] dataGroup_lo_2990 = {dataGroup_lo_hi_2990, dataGroup_lo_lo_2990};
  wire [2047:0] dataGroup_hi_2990 = {dataGroup_hi_hi_2990, dataGroup_hi_lo_2990};
  wire [15:0]   dataGroup_14_57 = dataGroup_lo_2990[1583:1568];
  wire [2047:0] dataGroup_lo_2991 = {dataGroup_lo_hi_2991, dataGroup_lo_lo_2991};
  wire [2047:0] dataGroup_hi_2991 = {dataGroup_hi_hi_2991, dataGroup_hi_lo_2991};
  wire [15:0]   dataGroup_15_57 = dataGroup_lo_2991[1695:1680];
  wire [2047:0] dataGroup_lo_2992 = {dataGroup_lo_hi_2992, dataGroup_lo_lo_2992};
  wire [2047:0] dataGroup_hi_2992 = {dataGroup_hi_hi_2992, dataGroup_hi_lo_2992};
  wire [15:0]   dataGroup_16_57 = dataGroup_lo_2992[1807:1792];
  wire [2047:0] dataGroup_lo_2993 = {dataGroup_lo_hi_2993, dataGroup_lo_lo_2993};
  wire [2047:0] dataGroup_hi_2993 = {dataGroup_hi_hi_2993, dataGroup_hi_lo_2993};
  wire [15:0]   dataGroup_17_57 = dataGroup_lo_2993[1919:1904];
  wire [2047:0] dataGroup_lo_2994 = {dataGroup_lo_hi_2994, dataGroup_lo_lo_2994};
  wire [2047:0] dataGroup_hi_2994 = {dataGroup_hi_hi_2994, dataGroup_hi_lo_2994};
  wire [15:0]   dataGroup_18_57 = dataGroup_lo_2994[2031:2016];
  wire [2047:0] dataGroup_lo_2995 = {dataGroup_lo_hi_2995, dataGroup_lo_lo_2995};
  wire [2047:0] dataGroup_hi_2995 = {dataGroup_hi_hi_2995, dataGroup_hi_lo_2995};
  wire [15:0]   dataGroup_19_57 = dataGroup_hi_2995[95:80];
  wire [2047:0] dataGroup_lo_2996 = {dataGroup_lo_hi_2996, dataGroup_lo_lo_2996};
  wire [2047:0] dataGroup_hi_2996 = {dataGroup_hi_hi_2996, dataGroup_hi_lo_2996};
  wire [15:0]   dataGroup_20_57 = dataGroup_hi_2996[207:192];
  wire [2047:0] dataGroup_lo_2997 = {dataGroup_lo_hi_2997, dataGroup_lo_lo_2997};
  wire [2047:0] dataGroup_hi_2997 = {dataGroup_hi_hi_2997, dataGroup_hi_lo_2997};
  wire [15:0]   dataGroup_21_57 = dataGroup_hi_2997[319:304];
  wire [2047:0] dataGroup_lo_2998 = {dataGroup_lo_hi_2998, dataGroup_lo_lo_2998};
  wire [2047:0] dataGroup_hi_2998 = {dataGroup_hi_hi_2998, dataGroup_hi_lo_2998};
  wire [15:0]   dataGroup_22_57 = dataGroup_hi_2998[431:416];
  wire [2047:0] dataGroup_lo_2999 = {dataGroup_lo_hi_2999, dataGroup_lo_lo_2999};
  wire [2047:0] dataGroup_hi_2999 = {dataGroup_hi_hi_2999, dataGroup_hi_lo_2999};
  wire [15:0]   dataGroup_23_57 = dataGroup_hi_2999[543:528];
  wire [2047:0] dataGroup_lo_3000 = {dataGroup_lo_hi_3000, dataGroup_lo_lo_3000};
  wire [2047:0] dataGroup_hi_3000 = {dataGroup_hi_hi_3000, dataGroup_hi_lo_3000};
  wire [15:0]   dataGroup_24_57 = dataGroup_hi_3000[655:640];
  wire [2047:0] dataGroup_lo_3001 = {dataGroup_lo_hi_3001, dataGroup_lo_lo_3001};
  wire [2047:0] dataGroup_hi_3001 = {dataGroup_hi_hi_3001, dataGroup_hi_lo_3001};
  wire [15:0]   dataGroup_25_57 = dataGroup_hi_3001[767:752];
  wire [2047:0] dataGroup_lo_3002 = {dataGroup_lo_hi_3002, dataGroup_lo_lo_3002};
  wire [2047:0] dataGroup_hi_3002 = {dataGroup_hi_hi_3002, dataGroup_hi_lo_3002};
  wire [15:0]   dataGroup_26_57 = dataGroup_hi_3002[879:864];
  wire [2047:0] dataGroup_lo_3003 = {dataGroup_lo_hi_3003, dataGroup_lo_lo_3003};
  wire [2047:0] dataGroup_hi_3003 = {dataGroup_hi_hi_3003, dataGroup_hi_lo_3003};
  wire [15:0]   dataGroup_27_57 = dataGroup_hi_3003[991:976];
  wire [2047:0] dataGroup_lo_3004 = {dataGroup_lo_hi_3004, dataGroup_lo_lo_3004};
  wire [2047:0] dataGroup_hi_3004 = {dataGroup_hi_hi_3004, dataGroup_hi_lo_3004};
  wire [15:0]   dataGroup_28_57 = dataGroup_hi_3004[1103:1088];
  wire [2047:0] dataGroup_lo_3005 = {dataGroup_lo_hi_3005, dataGroup_lo_lo_3005};
  wire [2047:0] dataGroup_hi_3005 = {dataGroup_hi_hi_3005, dataGroup_hi_lo_3005};
  wire [15:0]   dataGroup_29_57 = dataGroup_hi_3005[1215:1200];
  wire [2047:0] dataGroup_lo_3006 = {dataGroup_lo_hi_3006, dataGroup_lo_lo_3006};
  wire [2047:0] dataGroup_hi_3006 = {dataGroup_hi_hi_3006, dataGroup_hi_lo_3006};
  wire [15:0]   dataGroup_30_57 = dataGroup_hi_3006[1327:1312];
  wire [2047:0] dataGroup_lo_3007 = {dataGroup_lo_hi_3007, dataGroup_lo_lo_3007};
  wire [2047:0] dataGroup_hi_3007 = {dataGroup_hi_hi_3007, dataGroup_hi_lo_3007};
  wire [15:0]   dataGroup_31_57 = dataGroup_hi_3007[1439:1424];
  wire [31:0]   res_lo_lo_lo_lo_57 = {dataGroup_1_57, dataGroup_0_57};
  wire [31:0]   res_lo_lo_lo_hi_57 = {dataGroup_3_57, dataGroup_2_57};
  wire [63:0]   res_lo_lo_lo_57 = {res_lo_lo_lo_hi_57, res_lo_lo_lo_lo_57};
  wire [31:0]   res_lo_lo_hi_lo_57 = {dataGroup_5_57, dataGroup_4_57};
  wire [31:0]   res_lo_lo_hi_hi_57 = {dataGroup_7_57, dataGroup_6_57};
  wire [63:0]   res_lo_lo_hi_57 = {res_lo_lo_hi_hi_57, res_lo_lo_hi_lo_57};
  wire [127:0]  res_lo_lo_57 = {res_lo_lo_hi_57, res_lo_lo_lo_57};
  wire [31:0]   res_lo_hi_lo_lo_57 = {dataGroup_9_57, dataGroup_8_57};
  wire [31:0]   res_lo_hi_lo_hi_57 = {dataGroup_11_57, dataGroup_10_57};
  wire [63:0]   res_lo_hi_lo_57 = {res_lo_hi_lo_hi_57, res_lo_hi_lo_lo_57};
  wire [31:0]   res_lo_hi_hi_lo_57 = {dataGroup_13_57, dataGroup_12_57};
  wire [31:0]   res_lo_hi_hi_hi_57 = {dataGroup_15_57, dataGroup_14_57};
  wire [63:0]   res_lo_hi_hi_57 = {res_lo_hi_hi_hi_57, res_lo_hi_hi_lo_57};
  wire [127:0]  res_lo_hi_57 = {res_lo_hi_hi_57, res_lo_hi_lo_57};
  wire [255:0]  res_lo_57 = {res_lo_hi_57, res_lo_lo_57};
  wire [31:0]   res_hi_lo_lo_lo_57 = {dataGroup_17_57, dataGroup_16_57};
  wire [31:0]   res_hi_lo_lo_hi_57 = {dataGroup_19_57, dataGroup_18_57};
  wire [63:0]   res_hi_lo_lo_57 = {res_hi_lo_lo_hi_57, res_hi_lo_lo_lo_57};
  wire [31:0]   res_hi_lo_hi_lo_57 = {dataGroup_21_57, dataGroup_20_57};
  wire [31:0]   res_hi_lo_hi_hi_57 = {dataGroup_23_57, dataGroup_22_57};
  wire [63:0]   res_hi_lo_hi_57 = {res_hi_lo_hi_hi_57, res_hi_lo_hi_lo_57};
  wire [127:0]  res_hi_lo_57 = {res_hi_lo_hi_57, res_hi_lo_lo_57};
  wire [31:0]   res_hi_hi_lo_lo_57 = {dataGroup_25_57, dataGroup_24_57};
  wire [31:0]   res_hi_hi_lo_hi_57 = {dataGroup_27_57, dataGroup_26_57};
  wire [63:0]   res_hi_hi_lo_57 = {res_hi_hi_lo_hi_57, res_hi_hi_lo_lo_57};
  wire [31:0]   res_hi_hi_hi_lo_57 = {dataGroup_29_57, dataGroup_28_57};
  wire [31:0]   res_hi_hi_hi_hi_57 = {dataGroup_31_57, dataGroup_30_57};
  wire [63:0]   res_hi_hi_hi_57 = {res_hi_hi_hi_hi_57, res_hi_hi_hi_lo_57};
  wire [127:0]  res_hi_hi_57 = {res_hi_hi_hi_57, res_hi_hi_lo_57};
  wire [255:0]  res_hi_57 = {res_hi_hi_57, res_hi_lo_57};
  wire [511:0]  res_112 = {res_hi_57, res_lo_57};
  wire [2047:0] dataGroup_lo_3008 = {dataGroup_lo_hi_3008, dataGroup_lo_lo_3008};
  wire [2047:0] dataGroup_hi_3008 = {dataGroup_hi_hi_3008, dataGroup_hi_lo_3008};
  wire [15:0]   dataGroup_0_58 = dataGroup_lo_3008[31:16];
  wire [2047:0] dataGroup_lo_3009 = {dataGroup_lo_hi_3009, dataGroup_lo_lo_3009};
  wire [2047:0] dataGroup_hi_3009 = {dataGroup_hi_hi_3009, dataGroup_hi_lo_3009};
  wire [15:0]   dataGroup_1_58 = dataGroup_lo_3009[143:128];
  wire [2047:0] dataGroup_lo_3010 = {dataGroup_lo_hi_3010, dataGroup_lo_lo_3010};
  wire [2047:0] dataGroup_hi_3010 = {dataGroup_hi_hi_3010, dataGroup_hi_lo_3010};
  wire [15:0]   dataGroup_2_58 = dataGroup_lo_3010[255:240];
  wire [2047:0] dataGroup_lo_3011 = {dataGroup_lo_hi_3011, dataGroup_lo_lo_3011};
  wire [2047:0] dataGroup_hi_3011 = {dataGroup_hi_hi_3011, dataGroup_hi_lo_3011};
  wire [15:0]   dataGroup_3_58 = dataGroup_lo_3011[367:352];
  wire [2047:0] dataGroup_lo_3012 = {dataGroup_lo_hi_3012, dataGroup_lo_lo_3012};
  wire [2047:0] dataGroup_hi_3012 = {dataGroup_hi_hi_3012, dataGroup_hi_lo_3012};
  wire [15:0]   dataGroup_4_58 = dataGroup_lo_3012[479:464];
  wire [2047:0] dataGroup_lo_3013 = {dataGroup_lo_hi_3013, dataGroup_lo_lo_3013};
  wire [2047:0] dataGroup_hi_3013 = {dataGroup_hi_hi_3013, dataGroup_hi_lo_3013};
  wire [15:0]   dataGroup_5_58 = dataGroup_lo_3013[591:576];
  wire [2047:0] dataGroup_lo_3014 = {dataGroup_lo_hi_3014, dataGroup_lo_lo_3014};
  wire [2047:0] dataGroup_hi_3014 = {dataGroup_hi_hi_3014, dataGroup_hi_lo_3014};
  wire [15:0]   dataGroup_6_58 = dataGroup_lo_3014[703:688];
  wire [2047:0] dataGroup_lo_3015 = {dataGroup_lo_hi_3015, dataGroup_lo_lo_3015};
  wire [2047:0] dataGroup_hi_3015 = {dataGroup_hi_hi_3015, dataGroup_hi_lo_3015};
  wire [15:0]   dataGroup_7_58 = dataGroup_lo_3015[815:800];
  wire [2047:0] dataGroup_lo_3016 = {dataGroup_lo_hi_3016, dataGroup_lo_lo_3016};
  wire [2047:0] dataGroup_hi_3016 = {dataGroup_hi_hi_3016, dataGroup_hi_lo_3016};
  wire [15:0]   dataGroup_8_58 = dataGroup_lo_3016[927:912];
  wire [2047:0] dataGroup_lo_3017 = {dataGroup_lo_hi_3017, dataGroup_lo_lo_3017};
  wire [2047:0] dataGroup_hi_3017 = {dataGroup_hi_hi_3017, dataGroup_hi_lo_3017};
  wire [15:0]   dataGroup_9_58 = dataGroup_lo_3017[1039:1024];
  wire [2047:0] dataGroup_lo_3018 = {dataGroup_lo_hi_3018, dataGroup_lo_lo_3018};
  wire [2047:0] dataGroup_hi_3018 = {dataGroup_hi_hi_3018, dataGroup_hi_lo_3018};
  wire [15:0]   dataGroup_10_58 = dataGroup_lo_3018[1151:1136];
  wire [2047:0] dataGroup_lo_3019 = {dataGroup_lo_hi_3019, dataGroup_lo_lo_3019};
  wire [2047:0] dataGroup_hi_3019 = {dataGroup_hi_hi_3019, dataGroup_hi_lo_3019};
  wire [15:0]   dataGroup_11_58 = dataGroup_lo_3019[1263:1248];
  wire [2047:0] dataGroup_lo_3020 = {dataGroup_lo_hi_3020, dataGroup_lo_lo_3020};
  wire [2047:0] dataGroup_hi_3020 = {dataGroup_hi_hi_3020, dataGroup_hi_lo_3020};
  wire [15:0]   dataGroup_12_58 = dataGroup_lo_3020[1375:1360];
  wire [2047:0] dataGroup_lo_3021 = {dataGroup_lo_hi_3021, dataGroup_lo_lo_3021};
  wire [2047:0] dataGroup_hi_3021 = {dataGroup_hi_hi_3021, dataGroup_hi_lo_3021};
  wire [15:0]   dataGroup_13_58 = dataGroup_lo_3021[1487:1472];
  wire [2047:0] dataGroup_lo_3022 = {dataGroup_lo_hi_3022, dataGroup_lo_lo_3022};
  wire [2047:0] dataGroup_hi_3022 = {dataGroup_hi_hi_3022, dataGroup_hi_lo_3022};
  wire [15:0]   dataGroup_14_58 = dataGroup_lo_3022[1599:1584];
  wire [2047:0] dataGroup_lo_3023 = {dataGroup_lo_hi_3023, dataGroup_lo_lo_3023};
  wire [2047:0] dataGroup_hi_3023 = {dataGroup_hi_hi_3023, dataGroup_hi_lo_3023};
  wire [15:0]   dataGroup_15_58 = dataGroup_lo_3023[1711:1696];
  wire [2047:0] dataGroup_lo_3024 = {dataGroup_lo_hi_3024, dataGroup_lo_lo_3024};
  wire [2047:0] dataGroup_hi_3024 = {dataGroup_hi_hi_3024, dataGroup_hi_lo_3024};
  wire [15:0]   dataGroup_16_58 = dataGroup_lo_3024[1823:1808];
  wire [2047:0] dataGroup_lo_3025 = {dataGroup_lo_hi_3025, dataGroup_lo_lo_3025};
  wire [2047:0] dataGroup_hi_3025 = {dataGroup_hi_hi_3025, dataGroup_hi_lo_3025};
  wire [15:0]   dataGroup_17_58 = dataGroup_lo_3025[1935:1920];
  wire [2047:0] dataGroup_lo_3026 = {dataGroup_lo_hi_3026, dataGroup_lo_lo_3026};
  wire [2047:0] dataGroup_hi_3026 = {dataGroup_hi_hi_3026, dataGroup_hi_lo_3026};
  wire [15:0]   dataGroup_18_58 = dataGroup_lo_3026[2047:2032];
  wire [2047:0] dataGroup_lo_3027 = {dataGroup_lo_hi_3027, dataGroup_lo_lo_3027};
  wire [2047:0] dataGroup_hi_3027 = {dataGroup_hi_hi_3027, dataGroup_hi_lo_3027};
  wire [15:0]   dataGroup_19_58 = dataGroup_hi_3027[111:96];
  wire [2047:0] dataGroup_lo_3028 = {dataGroup_lo_hi_3028, dataGroup_lo_lo_3028};
  wire [2047:0] dataGroup_hi_3028 = {dataGroup_hi_hi_3028, dataGroup_hi_lo_3028};
  wire [15:0]   dataGroup_20_58 = dataGroup_hi_3028[223:208];
  wire [2047:0] dataGroup_lo_3029 = {dataGroup_lo_hi_3029, dataGroup_lo_lo_3029};
  wire [2047:0] dataGroup_hi_3029 = {dataGroup_hi_hi_3029, dataGroup_hi_lo_3029};
  wire [15:0]   dataGroup_21_58 = dataGroup_hi_3029[335:320];
  wire [2047:0] dataGroup_lo_3030 = {dataGroup_lo_hi_3030, dataGroup_lo_lo_3030};
  wire [2047:0] dataGroup_hi_3030 = {dataGroup_hi_hi_3030, dataGroup_hi_lo_3030};
  wire [15:0]   dataGroup_22_58 = dataGroup_hi_3030[447:432];
  wire [2047:0] dataGroup_lo_3031 = {dataGroup_lo_hi_3031, dataGroup_lo_lo_3031};
  wire [2047:0] dataGroup_hi_3031 = {dataGroup_hi_hi_3031, dataGroup_hi_lo_3031};
  wire [15:0]   dataGroup_23_58 = dataGroup_hi_3031[559:544];
  wire [2047:0] dataGroup_lo_3032 = {dataGroup_lo_hi_3032, dataGroup_lo_lo_3032};
  wire [2047:0] dataGroup_hi_3032 = {dataGroup_hi_hi_3032, dataGroup_hi_lo_3032};
  wire [15:0]   dataGroup_24_58 = dataGroup_hi_3032[671:656];
  wire [2047:0] dataGroup_lo_3033 = {dataGroup_lo_hi_3033, dataGroup_lo_lo_3033};
  wire [2047:0] dataGroup_hi_3033 = {dataGroup_hi_hi_3033, dataGroup_hi_lo_3033};
  wire [15:0]   dataGroup_25_58 = dataGroup_hi_3033[783:768];
  wire [2047:0] dataGroup_lo_3034 = {dataGroup_lo_hi_3034, dataGroup_lo_lo_3034};
  wire [2047:0] dataGroup_hi_3034 = {dataGroup_hi_hi_3034, dataGroup_hi_lo_3034};
  wire [15:0]   dataGroup_26_58 = dataGroup_hi_3034[895:880];
  wire [2047:0] dataGroup_lo_3035 = {dataGroup_lo_hi_3035, dataGroup_lo_lo_3035};
  wire [2047:0] dataGroup_hi_3035 = {dataGroup_hi_hi_3035, dataGroup_hi_lo_3035};
  wire [15:0]   dataGroup_27_58 = dataGroup_hi_3035[1007:992];
  wire [2047:0] dataGroup_lo_3036 = {dataGroup_lo_hi_3036, dataGroup_lo_lo_3036};
  wire [2047:0] dataGroup_hi_3036 = {dataGroup_hi_hi_3036, dataGroup_hi_lo_3036};
  wire [15:0]   dataGroup_28_58 = dataGroup_hi_3036[1119:1104];
  wire [2047:0] dataGroup_lo_3037 = {dataGroup_lo_hi_3037, dataGroup_lo_lo_3037};
  wire [2047:0] dataGroup_hi_3037 = {dataGroup_hi_hi_3037, dataGroup_hi_lo_3037};
  wire [15:0]   dataGroup_29_58 = dataGroup_hi_3037[1231:1216];
  wire [2047:0] dataGroup_lo_3038 = {dataGroup_lo_hi_3038, dataGroup_lo_lo_3038};
  wire [2047:0] dataGroup_hi_3038 = {dataGroup_hi_hi_3038, dataGroup_hi_lo_3038};
  wire [15:0]   dataGroup_30_58 = dataGroup_hi_3038[1343:1328];
  wire [2047:0] dataGroup_lo_3039 = {dataGroup_lo_hi_3039, dataGroup_lo_lo_3039};
  wire [2047:0] dataGroup_hi_3039 = {dataGroup_hi_hi_3039, dataGroup_hi_lo_3039};
  wire [15:0]   dataGroup_31_58 = dataGroup_hi_3039[1455:1440];
  wire [31:0]   res_lo_lo_lo_lo_58 = {dataGroup_1_58, dataGroup_0_58};
  wire [31:0]   res_lo_lo_lo_hi_58 = {dataGroup_3_58, dataGroup_2_58};
  wire [63:0]   res_lo_lo_lo_58 = {res_lo_lo_lo_hi_58, res_lo_lo_lo_lo_58};
  wire [31:0]   res_lo_lo_hi_lo_58 = {dataGroup_5_58, dataGroup_4_58};
  wire [31:0]   res_lo_lo_hi_hi_58 = {dataGroup_7_58, dataGroup_6_58};
  wire [63:0]   res_lo_lo_hi_58 = {res_lo_lo_hi_hi_58, res_lo_lo_hi_lo_58};
  wire [127:0]  res_lo_lo_58 = {res_lo_lo_hi_58, res_lo_lo_lo_58};
  wire [31:0]   res_lo_hi_lo_lo_58 = {dataGroup_9_58, dataGroup_8_58};
  wire [31:0]   res_lo_hi_lo_hi_58 = {dataGroup_11_58, dataGroup_10_58};
  wire [63:0]   res_lo_hi_lo_58 = {res_lo_hi_lo_hi_58, res_lo_hi_lo_lo_58};
  wire [31:0]   res_lo_hi_hi_lo_58 = {dataGroup_13_58, dataGroup_12_58};
  wire [31:0]   res_lo_hi_hi_hi_58 = {dataGroup_15_58, dataGroup_14_58};
  wire [63:0]   res_lo_hi_hi_58 = {res_lo_hi_hi_hi_58, res_lo_hi_hi_lo_58};
  wire [127:0]  res_lo_hi_58 = {res_lo_hi_hi_58, res_lo_hi_lo_58};
  wire [255:0]  res_lo_58 = {res_lo_hi_58, res_lo_lo_58};
  wire [31:0]   res_hi_lo_lo_lo_58 = {dataGroup_17_58, dataGroup_16_58};
  wire [31:0]   res_hi_lo_lo_hi_58 = {dataGroup_19_58, dataGroup_18_58};
  wire [63:0]   res_hi_lo_lo_58 = {res_hi_lo_lo_hi_58, res_hi_lo_lo_lo_58};
  wire [31:0]   res_hi_lo_hi_lo_58 = {dataGroup_21_58, dataGroup_20_58};
  wire [31:0]   res_hi_lo_hi_hi_58 = {dataGroup_23_58, dataGroup_22_58};
  wire [63:0]   res_hi_lo_hi_58 = {res_hi_lo_hi_hi_58, res_hi_lo_hi_lo_58};
  wire [127:0]  res_hi_lo_58 = {res_hi_lo_hi_58, res_hi_lo_lo_58};
  wire [31:0]   res_hi_hi_lo_lo_58 = {dataGroup_25_58, dataGroup_24_58};
  wire [31:0]   res_hi_hi_lo_hi_58 = {dataGroup_27_58, dataGroup_26_58};
  wire [63:0]   res_hi_hi_lo_58 = {res_hi_hi_lo_hi_58, res_hi_hi_lo_lo_58};
  wire [31:0]   res_hi_hi_hi_lo_58 = {dataGroup_29_58, dataGroup_28_58};
  wire [31:0]   res_hi_hi_hi_hi_58 = {dataGroup_31_58, dataGroup_30_58};
  wire [63:0]   res_hi_hi_hi_58 = {res_hi_hi_hi_hi_58, res_hi_hi_hi_lo_58};
  wire [127:0]  res_hi_hi_58 = {res_hi_hi_hi_58, res_hi_hi_lo_58};
  wire [255:0]  res_hi_58 = {res_hi_hi_58, res_hi_lo_58};
  wire [511:0]  res_113 = {res_hi_58, res_lo_58};
  wire [2047:0] dataGroup_lo_3040 = {dataGroup_lo_hi_3040, dataGroup_lo_lo_3040};
  wire [2047:0] dataGroup_hi_3040 = {dataGroup_hi_hi_3040, dataGroup_hi_lo_3040};
  wire [15:0]   dataGroup_0_59 = dataGroup_lo_3040[47:32];
  wire [2047:0] dataGroup_lo_3041 = {dataGroup_lo_hi_3041, dataGroup_lo_lo_3041};
  wire [2047:0] dataGroup_hi_3041 = {dataGroup_hi_hi_3041, dataGroup_hi_lo_3041};
  wire [15:0]   dataGroup_1_59 = dataGroup_lo_3041[159:144];
  wire [2047:0] dataGroup_lo_3042 = {dataGroup_lo_hi_3042, dataGroup_lo_lo_3042};
  wire [2047:0] dataGroup_hi_3042 = {dataGroup_hi_hi_3042, dataGroup_hi_lo_3042};
  wire [15:0]   dataGroup_2_59 = dataGroup_lo_3042[271:256];
  wire [2047:0] dataGroup_lo_3043 = {dataGroup_lo_hi_3043, dataGroup_lo_lo_3043};
  wire [2047:0] dataGroup_hi_3043 = {dataGroup_hi_hi_3043, dataGroup_hi_lo_3043};
  wire [15:0]   dataGroup_3_59 = dataGroup_lo_3043[383:368];
  wire [2047:0] dataGroup_lo_3044 = {dataGroup_lo_hi_3044, dataGroup_lo_lo_3044};
  wire [2047:0] dataGroup_hi_3044 = {dataGroup_hi_hi_3044, dataGroup_hi_lo_3044};
  wire [15:0]   dataGroup_4_59 = dataGroup_lo_3044[495:480];
  wire [2047:0] dataGroup_lo_3045 = {dataGroup_lo_hi_3045, dataGroup_lo_lo_3045};
  wire [2047:0] dataGroup_hi_3045 = {dataGroup_hi_hi_3045, dataGroup_hi_lo_3045};
  wire [15:0]   dataGroup_5_59 = dataGroup_lo_3045[607:592];
  wire [2047:0] dataGroup_lo_3046 = {dataGroup_lo_hi_3046, dataGroup_lo_lo_3046};
  wire [2047:0] dataGroup_hi_3046 = {dataGroup_hi_hi_3046, dataGroup_hi_lo_3046};
  wire [15:0]   dataGroup_6_59 = dataGroup_lo_3046[719:704];
  wire [2047:0] dataGroup_lo_3047 = {dataGroup_lo_hi_3047, dataGroup_lo_lo_3047};
  wire [2047:0] dataGroup_hi_3047 = {dataGroup_hi_hi_3047, dataGroup_hi_lo_3047};
  wire [15:0]   dataGroup_7_59 = dataGroup_lo_3047[831:816];
  wire [2047:0] dataGroup_lo_3048 = {dataGroup_lo_hi_3048, dataGroup_lo_lo_3048};
  wire [2047:0] dataGroup_hi_3048 = {dataGroup_hi_hi_3048, dataGroup_hi_lo_3048};
  wire [15:0]   dataGroup_8_59 = dataGroup_lo_3048[943:928];
  wire [2047:0] dataGroup_lo_3049 = {dataGroup_lo_hi_3049, dataGroup_lo_lo_3049};
  wire [2047:0] dataGroup_hi_3049 = {dataGroup_hi_hi_3049, dataGroup_hi_lo_3049};
  wire [15:0]   dataGroup_9_59 = dataGroup_lo_3049[1055:1040];
  wire [2047:0] dataGroup_lo_3050 = {dataGroup_lo_hi_3050, dataGroup_lo_lo_3050};
  wire [2047:0] dataGroup_hi_3050 = {dataGroup_hi_hi_3050, dataGroup_hi_lo_3050};
  wire [15:0]   dataGroup_10_59 = dataGroup_lo_3050[1167:1152];
  wire [2047:0] dataGroup_lo_3051 = {dataGroup_lo_hi_3051, dataGroup_lo_lo_3051};
  wire [2047:0] dataGroup_hi_3051 = {dataGroup_hi_hi_3051, dataGroup_hi_lo_3051};
  wire [15:0]   dataGroup_11_59 = dataGroup_lo_3051[1279:1264];
  wire [2047:0] dataGroup_lo_3052 = {dataGroup_lo_hi_3052, dataGroup_lo_lo_3052};
  wire [2047:0] dataGroup_hi_3052 = {dataGroup_hi_hi_3052, dataGroup_hi_lo_3052};
  wire [15:0]   dataGroup_12_59 = dataGroup_lo_3052[1391:1376];
  wire [2047:0] dataGroup_lo_3053 = {dataGroup_lo_hi_3053, dataGroup_lo_lo_3053};
  wire [2047:0] dataGroup_hi_3053 = {dataGroup_hi_hi_3053, dataGroup_hi_lo_3053};
  wire [15:0]   dataGroup_13_59 = dataGroup_lo_3053[1503:1488];
  wire [2047:0] dataGroup_lo_3054 = {dataGroup_lo_hi_3054, dataGroup_lo_lo_3054};
  wire [2047:0] dataGroup_hi_3054 = {dataGroup_hi_hi_3054, dataGroup_hi_lo_3054};
  wire [15:0]   dataGroup_14_59 = dataGroup_lo_3054[1615:1600];
  wire [2047:0] dataGroup_lo_3055 = {dataGroup_lo_hi_3055, dataGroup_lo_lo_3055};
  wire [2047:0] dataGroup_hi_3055 = {dataGroup_hi_hi_3055, dataGroup_hi_lo_3055};
  wire [15:0]   dataGroup_15_59 = dataGroup_lo_3055[1727:1712];
  wire [2047:0] dataGroup_lo_3056 = {dataGroup_lo_hi_3056, dataGroup_lo_lo_3056};
  wire [2047:0] dataGroup_hi_3056 = {dataGroup_hi_hi_3056, dataGroup_hi_lo_3056};
  wire [15:0]   dataGroup_16_59 = dataGroup_lo_3056[1839:1824];
  wire [2047:0] dataGroup_lo_3057 = {dataGroup_lo_hi_3057, dataGroup_lo_lo_3057};
  wire [2047:0] dataGroup_hi_3057 = {dataGroup_hi_hi_3057, dataGroup_hi_lo_3057};
  wire [15:0]   dataGroup_17_59 = dataGroup_lo_3057[1951:1936];
  wire [2047:0] dataGroup_lo_3058 = {dataGroup_lo_hi_3058, dataGroup_lo_lo_3058};
  wire [2047:0] dataGroup_hi_3058 = {dataGroup_hi_hi_3058, dataGroup_hi_lo_3058};
  wire [15:0]   dataGroup_18_59 = dataGroup_hi_3058[15:0];
  wire [2047:0] dataGroup_lo_3059 = {dataGroup_lo_hi_3059, dataGroup_lo_lo_3059};
  wire [2047:0] dataGroup_hi_3059 = {dataGroup_hi_hi_3059, dataGroup_hi_lo_3059};
  wire [15:0]   dataGroup_19_59 = dataGroup_hi_3059[127:112];
  wire [2047:0] dataGroup_lo_3060 = {dataGroup_lo_hi_3060, dataGroup_lo_lo_3060};
  wire [2047:0] dataGroup_hi_3060 = {dataGroup_hi_hi_3060, dataGroup_hi_lo_3060};
  wire [15:0]   dataGroup_20_59 = dataGroup_hi_3060[239:224];
  wire [2047:0] dataGroup_lo_3061 = {dataGroup_lo_hi_3061, dataGroup_lo_lo_3061};
  wire [2047:0] dataGroup_hi_3061 = {dataGroup_hi_hi_3061, dataGroup_hi_lo_3061};
  wire [15:0]   dataGroup_21_59 = dataGroup_hi_3061[351:336];
  wire [2047:0] dataGroup_lo_3062 = {dataGroup_lo_hi_3062, dataGroup_lo_lo_3062};
  wire [2047:0] dataGroup_hi_3062 = {dataGroup_hi_hi_3062, dataGroup_hi_lo_3062};
  wire [15:0]   dataGroup_22_59 = dataGroup_hi_3062[463:448];
  wire [2047:0] dataGroup_lo_3063 = {dataGroup_lo_hi_3063, dataGroup_lo_lo_3063};
  wire [2047:0] dataGroup_hi_3063 = {dataGroup_hi_hi_3063, dataGroup_hi_lo_3063};
  wire [15:0]   dataGroup_23_59 = dataGroup_hi_3063[575:560];
  wire [2047:0] dataGroup_lo_3064 = {dataGroup_lo_hi_3064, dataGroup_lo_lo_3064};
  wire [2047:0] dataGroup_hi_3064 = {dataGroup_hi_hi_3064, dataGroup_hi_lo_3064};
  wire [15:0]   dataGroup_24_59 = dataGroup_hi_3064[687:672];
  wire [2047:0] dataGroup_lo_3065 = {dataGroup_lo_hi_3065, dataGroup_lo_lo_3065};
  wire [2047:0] dataGroup_hi_3065 = {dataGroup_hi_hi_3065, dataGroup_hi_lo_3065};
  wire [15:0]   dataGroup_25_59 = dataGroup_hi_3065[799:784];
  wire [2047:0] dataGroup_lo_3066 = {dataGroup_lo_hi_3066, dataGroup_lo_lo_3066};
  wire [2047:0] dataGroup_hi_3066 = {dataGroup_hi_hi_3066, dataGroup_hi_lo_3066};
  wire [15:0]   dataGroup_26_59 = dataGroup_hi_3066[911:896];
  wire [2047:0] dataGroup_lo_3067 = {dataGroup_lo_hi_3067, dataGroup_lo_lo_3067};
  wire [2047:0] dataGroup_hi_3067 = {dataGroup_hi_hi_3067, dataGroup_hi_lo_3067};
  wire [15:0]   dataGroup_27_59 = dataGroup_hi_3067[1023:1008];
  wire [2047:0] dataGroup_lo_3068 = {dataGroup_lo_hi_3068, dataGroup_lo_lo_3068};
  wire [2047:0] dataGroup_hi_3068 = {dataGroup_hi_hi_3068, dataGroup_hi_lo_3068};
  wire [15:0]   dataGroup_28_59 = dataGroup_hi_3068[1135:1120];
  wire [2047:0] dataGroup_lo_3069 = {dataGroup_lo_hi_3069, dataGroup_lo_lo_3069};
  wire [2047:0] dataGroup_hi_3069 = {dataGroup_hi_hi_3069, dataGroup_hi_lo_3069};
  wire [15:0]   dataGroup_29_59 = dataGroup_hi_3069[1247:1232];
  wire [2047:0] dataGroup_lo_3070 = {dataGroup_lo_hi_3070, dataGroup_lo_lo_3070};
  wire [2047:0] dataGroup_hi_3070 = {dataGroup_hi_hi_3070, dataGroup_hi_lo_3070};
  wire [15:0]   dataGroup_30_59 = dataGroup_hi_3070[1359:1344];
  wire [2047:0] dataGroup_lo_3071 = {dataGroup_lo_hi_3071, dataGroup_lo_lo_3071};
  wire [2047:0] dataGroup_hi_3071 = {dataGroup_hi_hi_3071, dataGroup_hi_lo_3071};
  wire [15:0]   dataGroup_31_59 = dataGroup_hi_3071[1471:1456];
  wire [31:0]   res_lo_lo_lo_lo_59 = {dataGroup_1_59, dataGroup_0_59};
  wire [31:0]   res_lo_lo_lo_hi_59 = {dataGroup_3_59, dataGroup_2_59};
  wire [63:0]   res_lo_lo_lo_59 = {res_lo_lo_lo_hi_59, res_lo_lo_lo_lo_59};
  wire [31:0]   res_lo_lo_hi_lo_59 = {dataGroup_5_59, dataGroup_4_59};
  wire [31:0]   res_lo_lo_hi_hi_59 = {dataGroup_7_59, dataGroup_6_59};
  wire [63:0]   res_lo_lo_hi_59 = {res_lo_lo_hi_hi_59, res_lo_lo_hi_lo_59};
  wire [127:0]  res_lo_lo_59 = {res_lo_lo_hi_59, res_lo_lo_lo_59};
  wire [31:0]   res_lo_hi_lo_lo_59 = {dataGroup_9_59, dataGroup_8_59};
  wire [31:0]   res_lo_hi_lo_hi_59 = {dataGroup_11_59, dataGroup_10_59};
  wire [63:0]   res_lo_hi_lo_59 = {res_lo_hi_lo_hi_59, res_lo_hi_lo_lo_59};
  wire [31:0]   res_lo_hi_hi_lo_59 = {dataGroup_13_59, dataGroup_12_59};
  wire [31:0]   res_lo_hi_hi_hi_59 = {dataGroup_15_59, dataGroup_14_59};
  wire [63:0]   res_lo_hi_hi_59 = {res_lo_hi_hi_hi_59, res_lo_hi_hi_lo_59};
  wire [127:0]  res_lo_hi_59 = {res_lo_hi_hi_59, res_lo_hi_lo_59};
  wire [255:0]  res_lo_59 = {res_lo_hi_59, res_lo_lo_59};
  wire [31:0]   res_hi_lo_lo_lo_59 = {dataGroup_17_59, dataGroup_16_59};
  wire [31:0]   res_hi_lo_lo_hi_59 = {dataGroup_19_59, dataGroup_18_59};
  wire [63:0]   res_hi_lo_lo_59 = {res_hi_lo_lo_hi_59, res_hi_lo_lo_lo_59};
  wire [31:0]   res_hi_lo_hi_lo_59 = {dataGroup_21_59, dataGroup_20_59};
  wire [31:0]   res_hi_lo_hi_hi_59 = {dataGroup_23_59, dataGroup_22_59};
  wire [63:0]   res_hi_lo_hi_59 = {res_hi_lo_hi_hi_59, res_hi_lo_hi_lo_59};
  wire [127:0]  res_hi_lo_59 = {res_hi_lo_hi_59, res_hi_lo_lo_59};
  wire [31:0]   res_hi_hi_lo_lo_59 = {dataGroup_25_59, dataGroup_24_59};
  wire [31:0]   res_hi_hi_lo_hi_59 = {dataGroup_27_59, dataGroup_26_59};
  wire [63:0]   res_hi_hi_lo_59 = {res_hi_hi_lo_hi_59, res_hi_hi_lo_lo_59};
  wire [31:0]   res_hi_hi_hi_lo_59 = {dataGroup_29_59, dataGroup_28_59};
  wire [31:0]   res_hi_hi_hi_hi_59 = {dataGroup_31_59, dataGroup_30_59};
  wire [63:0]   res_hi_hi_hi_59 = {res_hi_hi_hi_hi_59, res_hi_hi_hi_lo_59};
  wire [127:0]  res_hi_hi_59 = {res_hi_hi_hi_59, res_hi_hi_lo_59};
  wire [255:0]  res_hi_59 = {res_hi_hi_59, res_hi_lo_59};
  wire [511:0]  res_114 = {res_hi_59, res_lo_59};
  wire [2047:0] dataGroup_lo_3072 = {dataGroup_lo_hi_3072, dataGroup_lo_lo_3072};
  wire [2047:0] dataGroup_hi_3072 = {dataGroup_hi_hi_3072, dataGroup_hi_lo_3072};
  wire [15:0]   dataGroup_0_60 = dataGroup_lo_3072[63:48];
  wire [2047:0] dataGroup_lo_3073 = {dataGroup_lo_hi_3073, dataGroup_lo_lo_3073};
  wire [2047:0] dataGroup_hi_3073 = {dataGroup_hi_hi_3073, dataGroup_hi_lo_3073};
  wire [15:0]   dataGroup_1_60 = dataGroup_lo_3073[175:160];
  wire [2047:0] dataGroup_lo_3074 = {dataGroup_lo_hi_3074, dataGroup_lo_lo_3074};
  wire [2047:0] dataGroup_hi_3074 = {dataGroup_hi_hi_3074, dataGroup_hi_lo_3074};
  wire [15:0]   dataGroup_2_60 = dataGroup_lo_3074[287:272];
  wire [2047:0] dataGroup_lo_3075 = {dataGroup_lo_hi_3075, dataGroup_lo_lo_3075};
  wire [2047:0] dataGroup_hi_3075 = {dataGroup_hi_hi_3075, dataGroup_hi_lo_3075};
  wire [15:0]   dataGroup_3_60 = dataGroup_lo_3075[399:384];
  wire [2047:0] dataGroup_lo_3076 = {dataGroup_lo_hi_3076, dataGroup_lo_lo_3076};
  wire [2047:0] dataGroup_hi_3076 = {dataGroup_hi_hi_3076, dataGroup_hi_lo_3076};
  wire [15:0]   dataGroup_4_60 = dataGroup_lo_3076[511:496];
  wire [2047:0] dataGroup_lo_3077 = {dataGroup_lo_hi_3077, dataGroup_lo_lo_3077};
  wire [2047:0] dataGroup_hi_3077 = {dataGroup_hi_hi_3077, dataGroup_hi_lo_3077};
  wire [15:0]   dataGroup_5_60 = dataGroup_lo_3077[623:608];
  wire [2047:0] dataGroup_lo_3078 = {dataGroup_lo_hi_3078, dataGroup_lo_lo_3078};
  wire [2047:0] dataGroup_hi_3078 = {dataGroup_hi_hi_3078, dataGroup_hi_lo_3078};
  wire [15:0]   dataGroup_6_60 = dataGroup_lo_3078[735:720];
  wire [2047:0] dataGroup_lo_3079 = {dataGroup_lo_hi_3079, dataGroup_lo_lo_3079};
  wire [2047:0] dataGroup_hi_3079 = {dataGroup_hi_hi_3079, dataGroup_hi_lo_3079};
  wire [15:0]   dataGroup_7_60 = dataGroup_lo_3079[847:832];
  wire [2047:0] dataGroup_lo_3080 = {dataGroup_lo_hi_3080, dataGroup_lo_lo_3080};
  wire [2047:0] dataGroup_hi_3080 = {dataGroup_hi_hi_3080, dataGroup_hi_lo_3080};
  wire [15:0]   dataGroup_8_60 = dataGroup_lo_3080[959:944];
  wire [2047:0] dataGroup_lo_3081 = {dataGroup_lo_hi_3081, dataGroup_lo_lo_3081};
  wire [2047:0] dataGroup_hi_3081 = {dataGroup_hi_hi_3081, dataGroup_hi_lo_3081};
  wire [15:0]   dataGroup_9_60 = dataGroup_lo_3081[1071:1056];
  wire [2047:0] dataGroup_lo_3082 = {dataGroup_lo_hi_3082, dataGroup_lo_lo_3082};
  wire [2047:0] dataGroup_hi_3082 = {dataGroup_hi_hi_3082, dataGroup_hi_lo_3082};
  wire [15:0]   dataGroup_10_60 = dataGroup_lo_3082[1183:1168];
  wire [2047:0] dataGroup_lo_3083 = {dataGroup_lo_hi_3083, dataGroup_lo_lo_3083};
  wire [2047:0] dataGroup_hi_3083 = {dataGroup_hi_hi_3083, dataGroup_hi_lo_3083};
  wire [15:0]   dataGroup_11_60 = dataGroup_lo_3083[1295:1280];
  wire [2047:0] dataGroup_lo_3084 = {dataGroup_lo_hi_3084, dataGroup_lo_lo_3084};
  wire [2047:0] dataGroup_hi_3084 = {dataGroup_hi_hi_3084, dataGroup_hi_lo_3084};
  wire [15:0]   dataGroup_12_60 = dataGroup_lo_3084[1407:1392];
  wire [2047:0] dataGroup_lo_3085 = {dataGroup_lo_hi_3085, dataGroup_lo_lo_3085};
  wire [2047:0] dataGroup_hi_3085 = {dataGroup_hi_hi_3085, dataGroup_hi_lo_3085};
  wire [15:0]   dataGroup_13_60 = dataGroup_lo_3085[1519:1504];
  wire [2047:0] dataGroup_lo_3086 = {dataGroup_lo_hi_3086, dataGroup_lo_lo_3086};
  wire [2047:0] dataGroup_hi_3086 = {dataGroup_hi_hi_3086, dataGroup_hi_lo_3086};
  wire [15:0]   dataGroup_14_60 = dataGroup_lo_3086[1631:1616];
  wire [2047:0] dataGroup_lo_3087 = {dataGroup_lo_hi_3087, dataGroup_lo_lo_3087};
  wire [2047:0] dataGroup_hi_3087 = {dataGroup_hi_hi_3087, dataGroup_hi_lo_3087};
  wire [15:0]   dataGroup_15_60 = dataGroup_lo_3087[1743:1728];
  wire [2047:0] dataGroup_lo_3088 = {dataGroup_lo_hi_3088, dataGroup_lo_lo_3088};
  wire [2047:0] dataGroup_hi_3088 = {dataGroup_hi_hi_3088, dataGroup_hi_lo_3088};
  wire [15:0]   dataGroup_16_60 = dataGroup_lo_3088[1855:1840];
  wire [2047:0] dataGroup_lo_3089 = {dataGroup_lo_hi_3089, dataGroup_lo_lo_3089};
  wire [2047:0] dataGroup_hi_3089 = {dataGroup_hi_hi_3089, dataGroup_hi_lo_3089};
  wire [15:0]   dataGroup_17_60 = dataGroup_lo_3089[1967:1952];
  wire [2047:0] dataGroup_lo_3090 = {dataGroup_lo_hi_3090, dataGroup_lo_lo_3090};
  wire [2047:0] dataGroup_hi_3090 = {dataGroup_hi_hi_3090, dataGroup_hi_lo_3090};
  wire [15:0]   dataGroup_18_60 = dataGroup_hi_3090[31:16];
  wire [2047:0] dataGroup_lo_3091 = {dataGroup_lo_hi_3091, dataGroup_lo_lo_3091};
  wire [2047:0] dataGroup_hi_3091 = {dataGroup_hi_hi_3091, dataGroup_hi_lo_3091};
  wire [15:0]   dataGroup_19_60 = dataGroup_hi_3091[143:128];
  wire [2047:0] dataGroup_lo_3092 = {dataGroup_lo_hi_3092, dataGroup_lo_lo_3092};
  wire [2047:0] dataGroup_hi_3092 = {dataGroup_hi_hi_3092, dataGroup_hi_lo_3092};
  wire [15:0]   dataGroup_20_60 = dataGroup_hi_3092[255:240];
  wire [2047:0] dataGroup_lo_3093 = {dataGroup_lo_hi_3093, dataGroup_lo_lo_3093};
  wire [2047:0] dataGroup_hi_3093 = {dataGroup_hi_hi_3093, dataGroup_hi_lo_3093};
  wire [15:0]   dataGroup_21_60 = dataGroup_hi_3093[367:352];
  wire [2047:0] dataGroup_lo_3094 = {dataGroup_lo_hi_3094, dataGroup_lo_lo_3094};
  wire [2047:0] dataGroup_hi_3094 = {dataGroup_hi_hi_3094, dataGroup_hi_lo_3094};
  wire [15:0]   dataGroup_22_60 = dataGroup_hi_3094[479:464];
  wire [2047:0] dataGroup_lo_3095 = {dataGroup_lo_hi_3095, dataGroup_lo_lo_3095};
  wire [2047:0] dataGroup_hi_3095 = {dataGroup_hi_hi_3095, dataGroup_hi_lo_3095};
  wire [15:0]   dataGroup_23_60 = dataGroup_hi_3095[591:576];
  wire [2047:0] dataGroup_lo_3096 = {dataGroup_lo_hi_3096, dataGroup_lo_lo_3096};
  wire [2047:0] dataGroup_hi_3096 = {dataGroup_hi_hi_3096, dataGroup_hi_lo_3096};
  wire [15:0]   dataGroup_24_60 = dataGroup_hi_3096[703:688];
  wire [2047:0] dataGroup_lo_3097 = {dataGroup_lo_hi_3097, dataGroup_lo_lo_3097};
  wire [2047:0] dataGroup_hi_3097 = {dataGroup_hi_hi_3097, dataGroup_hi_lo_3097};
  wire [15:0]   dataGroup_25_60 = dataGroup_hi_3097[815:800];
  wire [2047:0] dataGroup_lo_3098 = {dataGroup_lo_hi_3098, dataGroup_lo_lo_3098};
  wire [2047:0] dataGroup_hi_3098 = {dataGroup_hi_hi_3098, dataGroup_hi_lo_3098};
  wire [15:0]   dataGroup_26_60 = dataGroup_hi_3098[927:912];
  wire [2047:0] dataGroup_lo_3099 = {dataGroup_lo_hi_3099, dataGroup_lo_lo_3099};
  wire [2047:0] dataGroup_hi_3099 = {dataGroup_hi_hi_3099, dataGroup_hi_lo_3099};
  wire [15:0]   dataGroup_27_60 = dataGroup_hi_3099[1039:1024];
  wire [2047:0] dataGroup_lo_3100 = {dataGroup_lo_hi_3100, dataGroup_lo_lo_3100};
  wire [2047:0] dataGroup_hi_3100 = {dataGroup_hi_hi_3100, dataGroup_hi_lo_3100};
  wire [15:0]   dataGroup_28_60 = dataGroup_hi_3100[1151:1136];
  wire [2047:0] dataGroup_lo_3101 = {dataGroup_lo_hi_3101, dataGroup_lo_lo_3101};
  wire [2047:0] dataGroup_hi_3101 = {dataGroup_hi_hi_3101, dataGroup_hi_lo_3101};
  wire [15:0]   dataGroup_29_60 = dataGroup_hi_3101[1263:1248];
  wire [2047:0] dataGroup_lo_3102 = {dataGroup_lo_hi_3102, dataGroup_lo_lo_3102};
  wire [2047:0] dataGroup_hi_3102 = {dataGroup_hi_hi_3102, dataGroup_hi_lo_3102};
  wire [15:0]   dataGroup_30_60 = dataGroup_hi_3102[1375:1360];
  wire [2047:0] dataGroup_lo_3103 = {dataGroup_lo_hi_3103, dataGroup_lo_lo_3103};
  wire [2047:0] dataGroup_hi_3103 = {dataGroup_hi_hi_3103, dataGroup_hi_lo_3103};
  wire [15:0]   dataGroup_31_60 = dataGroup_hi_3103[1487:1472];
  wire [31:0]   res_lo_lo_lo_lo_60 = {dataGroup_1_60, dataGroup_0_60};
  wire [31:0]   res_lo_lo_lo_hi_60 = {dataGroup_3_60, dataGroup_2_60};
  wire [63:0]   res_lo_lo_lo_60 = {res_lo_lo_lo_hi_60, res_lo_lo_lo_lo_60};
  wire [31:0]   res_lo_lo_hi_lo_60 = {dataGroup_5_60, dataGroup_4_60};
  wire [31:0]   res_lo_lo_hi_hi_60 = {dataGroup_7_60, dataGroup_6_60};
  wire [63:0]   res_lo_lo_hi_60 = {res_lo_lo_hi_hi_60, res_lo_lo_hi_lo_60};
  wire [127:0]  res_lo_lo_60 = {res_lo_lo_hi_60, res_lo_lo_lo_60};
  wire [31:0]   res_lo_hi_lo_lo_60 = {dataGroup_9_60, dataGroup_8_60};
  wire [31:0]   res_lo_hi_lo_hi_60 = {dataGroup_11_60, dataGroup_10_60};
  wire [63:0]   res_lo_hi_lo_60 = {res_lo_hi_lo_hi_60, res_lo_hi_lo_lo_60};
  wire [31:0]   res_lo_hi_hi_lo_60 = {dataGroup_13_60, dataGroup_12_60};
  wire [31:0]   res_lo_hi_hi_hi_60 = {dataGroup_15_60, dataGroup_14_60};
  wire [63:0]   res_lo_hi_hi_60 = {res_lo_hi_hi_hi_60, res_lo_hi_hi_lo_60};
  wire [127:0]  res_lo_hi_60 = {res_lo_hi_hi_60, res_lo_hi_lo_60};
  wire [255:0]  res_lo_60 = {res_lo_hi_60, res_lo_lo_60};
  wire [31:0]   res_hi_lo_lo_lo_60 = {dataGroup_17_60, dataGroup_16_60};
  wire [31:0]   res_hi_lo_lo_hi_60 = {dataGroup_19_60, dataGroup_18_60};
  wire [63:0]   res_hi_lo_lo_60 = {res_hi_lo_lo_hi_60, res_hi_lo_lo_lo_60};
  wire [31:0]   res_hi_lo_hi_lo_60 = {dataGroup_21_60, dataGroup_20_60};
  wire [31:0]   res_hi_lo_hi_hi_60 = {dataGroup_23_60, dataGroup_22_60};
  wire [63:0]   res_hi_lo_hi_60 = {res_hi_lo_hi_hi_60, res_hi_lo_hi_lo_60};
  wire [127:0]  res_hi_lo_60 = {res_hi_lo_hi_60, res_hi_lo_lo_60};
  wire [31:0]   res_hi_hi_lo_lo_60 = {dataGroup_25_60, dataGroup_24_60};
  wire [31:0]   res_hi_hi_lo_hi_60 = {dataGroup_27_60, dataGroup_26_60};
  wire [63:0]   res_hi_hi_lo_60 = {res_hi_hi_lo_hi_60, res_hi_hi_lo_lo_60};
  wire [31:0]   res_hi_hi_hi_lo_60 = {dataGroup_29_60, dataGroup_28_60};
  wire [31:0]   res_hi_hi_hi_hi_60 = {dataGroup_31_60, dataGroup_30_60};
  wire [63:0]   res_hi_hi_hi_60 = {res_hi_hi_hi_hi_60, res_hi_hi_hi_lo_60};
  wire [127:0]  res_hi_hi_60 = {res_hi_hi_hi_60, res_hi_hi_lo_60};
  wire [255:0]  res_hi_60 = {res_hi_hi_60, res_hi_lo_60};
  wire [511:0]  res_115 = {res_hi_60, res_lo_60};
  wire [2047:0] dataGroup_lo_3104 = {dataGroup_lo_hi_3104, dataGroup_lo_lo_3104};
  wire [2047:0] dataGroup_hi_3104 = {dataGroup_hi_hi_3104, dataGroup_hi_lo_3104};
  wire [15:0]   dataGroup_0_61 = dataGroup_lo_3104[79:64];
  wire [2047:0] dataGroup_lo_3105 = {dataGroup_lo_hi_3105, dataGroup_lo_lo_3105};
  wire [2047:0] dataGroup_hi_3105 = {dataGroup_hi_hi_3105, dataGroup_hi_lo_3105};
  wire [15:0]   dataGroup_1_61 = dataGroup_lo_3105[191:176];
  wire [2047:0] dataGroup_lo_3106 = {dataGroup_lo_hi_3106, dataGroup_lo_lo_3106};
  wire [2047:0] dataGroup_hi_3106 = {dataGroup_hi_hi_3106, dataGroup_hi_lo_3106};
  wire [15:0]   dataGroup_2_61 = dataGroup_lo_3106[303:288];
  wire [2047:0] dataGroup_lo_3107 = {dataGroup_lo_hi_3107, dataGroup_lo_lo_3107};
  wire [2047:0] dataGroup_hi_3107 = {dataGroup_hi_hi_3107, dataGroup_hi_lo_3107};
  wire [15:0]   dataGroup_3_61 = dataGroup_lo_3107[415:400];
  wire [2047:0] dataGroup_lo_3108 = {dataGroup_lo_hi_3108, dataGroup_lo_lo_3108};
  wire [2047:0] dataGroup_hi_3108 = {dataGroup_hi_hi_3108, dataGroup_hi_lo_3108};
  wire [15:0]   dataGroup_4_61 = dataGroup_lo_3108[527:512];
  wire [2047:0] dataGroup_lo_3109 = {dataGroup_lo_hi_3109, dataGroup_lo_lo_3109};
  wire [2047:0] dataGroup_hi_3109 = {dataGroup_hi_hi_3109, dataGroup_hi_lo_3109};
  wire [15:0]   dataGroup_5_61 = dataGroup_lo_3109[639:624];
  wire [2047:0] dataGroup_lo_3110 = {dataGroup_lo_hi_3110, dataGroup_lo_lo_3110};
  wire [2047:0] dataGroup_hi_3110 = {dataGroup_hi_hi_3110, dataGroup_hi_lo_3110};
  wire [15:0]   dataGroup_6_61 = dataGroup_lo_3110[751:736];
  wire [2047:0] dataGroup_lo_3111 = {dataGroup_lo_hi_3111, dataGroup_lo_lo_3111};
  wire [2047:0] dataGroup_hi_3111 = {dataGroup_hi_hi_3111, dataGroup_hi_lo_3111};
  wire [15:0]   dataGroup_7_61 = dataGroup_lo_3111[863:848];
  wire [2047:0] dataGroup_lo_3112 = {dataGroup_lo_hi_3112, dataGroup_lo_lo_3112};
  wire [2047:0] dataGroup_hi_3112 = {dataGroup_hi_hi_3112, dataGroup_hi_lo_3112};
  wire [15:0]   dataGroup_8_61 = dataGroup_lo_3112[975:960];
  wire [2047:0] dataGroup_lo_3113 = {dataGroup_lo_hi_3113, dataGroup_lo_lo_3113};
  wire [2047:0] dataGroup_hi_3113 = {dataGroup_hi_hi_3113, dataGroup_hi_lo_3113};
  wire [15:0]   dataGroup_9_61 = dataGroup_lo_3113[1087:1072];
  wire [2047:0] dataGroup_lo_3114 = {dataGroup_lo_hi_3114, dataGroup_lo_lo_3114};
  wire [2047:0] dataGroup_hi_3114 = {dataGroup_hi_hi_3114, dataGroup_hi_lo_3114};
  wire [15:0]   dataGroup_10_61 = dataGroup_lo_3114[1199:1184];
  wire [2047:0] dataGroup_lo_3115 = {dataGroup_lo_hi_3115, dataGroup_lo_lo_3115};
  wire [2047:0] dataGroup_hi_3115 = {dataGroup_hi_hi_3115, dataGroup_hi_lo_3115};
  wire [15:0]   dataGroup_11_61 = dataGroup_lo_3115[1311:1296];
  wire [2047:0] dataGroup_lo_3116 = {dataGroup_lo_hi_3116, dataGroup_lo_lo_3116};
  wire [2047:0] dataGroup_hi_3116 = {dataGroup_hi_hi_3116, dataGroup_hi_lo_3116};
  wire [15:0]   dataGroup_12_61 = dataGroup_lo_3116[1423:1408];
  wire [2047:0] dataGroup_lo_3117 = {dataGroup_lo_hi_3117, dataGroup_lo_lo_3117};
  wire [2047:0] dataGroup_hi_3117 = {dataGroup_hi_hi_3117, dataGroup_hi_lo_3117};
  wire [15:0]   dataGroup_13_61 = dataGroup_lo_3117[1535:1520];
  wire [2047:0] dataGroup_lo_3118 = {dataGroup_lo_hi_3118, dataGroup_lo_lo_3118};
  wire [2047:0] dataGroup_hi_3118 = {dataGroup_hi_hi_3118, dataGroup_hi_lo_3118};
  wire [15:0]   dataGroup_14_61 = dataGroup_lo_3118[1647:1632];
  wire [2047:0] dataGroup_lo_3119 = {dataGroup_lo_hi_3119, dataGroup_lo_lo_3119};
  wire [2047:0] dataGroup_hi_3119 = {dataGroup_hi_hi_3119, dataGroup_hi_lo_3119};
  wire [15:0]   dataGroup_15_61 = dataGroup_lo_3119[1759:1744];
  wire [2047:0] dataGroup_lo_3120 = {dataGroup_lo_hi_3120, dataGroup_lo_lo_3120};
  wire [2047:0] dataGroup_hi_3120 = {dataGroup_hi_hi_3120, dataGroup_hi_lo_3120};
  wire [15:0]   dataGroup_16_61 = dataGroup_lo_3120[1871:1856];
  wire [2047:0] dataGroup_lo_3121 = {dataGroup_lo_hi_3121, dataGroup_lo_lo_3121};
  wire [2047:0] dataGroup_hi_3121 = {dataGroup_hi_hi_3121, dataGroup_hi_lo_3121};
  wire [15:0]   dataGroup_17_61 = dataGroup_lo_3121[1983:1968];
  wire [2047:0] dataGroup_lo_3122 = {dataGroup_lo_hi_3122, dataGroup_lo_lo_3122};
  wire [2047:0] dataGroup_hi_3122 = {dataGroup_hi_hi_3122, dataGroup_hi_lo_3122};
  wire [15:0]   dataGroup_18_61 = dataGroup_hi_3122[47:32];
  wire [2047:0] dataGroup_lo_3123 = {dataGroup_lo_hi_3123, dataGroup_lo_lo_3123};
  wire [2047:0] dataGroup_hi_3123 = {dataGroup_hi_hi_3123, dataGroup_hi_lo_3123};
  wire [15:0]   dataGroup_19_61 = dataGroup_hi_3123[159:144];
  wire [2047:0] dataGroup_lo_3124 = {dataGroup_lo_hi_3124, dataGroup_lo_lo_3124};
  wire [2047:0] dataGroup_hi_3124 = {dataGroup_hi_hi_3124, dataGroup_hi_lo_3124};
  wire [15:0]   dataGroup_20_61 = dataGroup_hi_3124[271:256];
  wire [2047:0] dataGroup_lo_3125 = {dataGroup_lo_hi_3125, dataGroup_lo_lo_3125};
  wire [2047:0] dataGroup_hi_3125 = {dataGroup_hi_hi_3125, dataGroup_hi_lo_3125};
  wire [15:0]   dataGroup_21_61 = dataGroup_hi_3125[383:368];
  wire [2047:0] dataGroup_lo_3126 = {dataGroup_lo_hi_3126, dataGroup_lo_lo_3126};
  wire [2047:0] dataGroup_hi_3126 = {dataGroup_hi_hi_3126, dataGroup_hi_lo_3126};
  wire [15:0]   dataGroup_22_61 = dataGroup_hi_3126[495:480];
  wire [2047:0] dataGroup_lo_3127 = {dataGroup_lo_hi_3127, dataGroup_lo_lo_3127};
  wire [2047:0] dataGroup_hi_3127 = {dataGroup_hi_hi_3127, dataGroup_hi_lo_3127};
  wire [15:0]   dataGroup_23_61 = dataGroup_hi_3127[607:592];
  wire [2047:0] dataGroup_lo_3128 = {dataGroup_lo_hi_3128, dataGroup_lo_lo_3128};
  wire [2047:0] dataGroup_hi_3128 = {dataGroup_hi_hi_3128, dataGroup_hi_lo_3128};
  wire [15:0]   dataGroup_24_61 = dataGroup_hi_3128[719:704];
  wire [2047:0] dataGroup_lo_3129 = {dataGroup_lo_hi_3129, dataGroup_lo_lo_3129};
  wire [2047:0] dataGroup_hi_3129 = {dataGroup_hi_hi_3129, dataGroup_hi_lo_3129};
  wire [15:0]   dataGroup_25_61 = dataGroup_hi_3129[831:816];
  wire [2047:0] dataGroup_lo_3130 = {dataGroup_lo_hi_3130, dataGroup_lo_lo_3130};
  wire [2047:0] dataGroup_hi_3130 = {dataGroup_hi_hi_3130, dataGroup_hi_lo_3130};
  wire [15:0]   dataGroup_26_61 = dataGroup_hi_3130[943:928];
  wire [2047:0] dataGroup_lo_3131 = {dataGroup_lo_hi_3131, dataGroup_lo_lo_3131};
  wire [2047:0] dataGroup_hi_3131 = {dataGroup_hi_hi_3131, dataGroup_hi_lo_3131};
  wire [15:0]   dataGroup_27_61 = dataGroup_hi_3131[1055:1040];
  wire [2047:0] dataGroup_lo_3132 = {dataGroup_lo_hi_3132, dataGroup_lo_lo_3132};
  wire [2047:0] dataGroup_hi_3132 = {dataGroup_hi_hi_3132, dataGroup_hi_lo_3132};
  wire [15:0]   dataGroup_28_61 = dataGroup_hi_3132[1167:1152];
  wire [2047:0] dataGroup_lo_3133 = {dataGroup_lo_hi_3133, dataGroup_lo_lo_3133};
  wire [2047:0] dataGroup_hi_3133 = {dataGroup_hi_hi_3133, dataGroup_hi_lo_3133};
  wire [15:0]   dataGroup_29_61 = dataGroup_hi_3133[1279:1264];
  wire [2047:0] dataGroup_lo_3134 = {dataGroup_lo_hi_3134, dataGroup_lo_lo_3134};
  wire [2047:0] dataGroup_hi_3134 = {dataGroup_hi_hi_3134, dataGroup_hi_lo_3134};
  wire [15:0]   dataGroup_30_61 = dataGroup_hi_3134[1391:1376];
  wire [2047:0] dataGroup_lo_3135 = {dataGroup_lo_hi_3135, dataGroup_lo_lo_3135};
  wire [2047:0] dataGroup_hi_3135 = {dataGroup_hi_hi_3135, dataGroup_hi_lo_3135};
  wire [15:0]   dataGroup_31_61 = dataGroup_hi_3135[1503:1488];
  wire [31:0]   res_lo_lo_lo_lo_61 = {dataGroup_1_61, dataGroup_0_61};
  wire [31:0]   res_lo_lo_lo_hi_61 = {dataGroup_3_61, dataGroup_2_61};
  wire [63:0]   res_lo_lo_lo_61 = {res_lo_lo_lo_hi_61, res_lo_lo_lo_lo_61};
  wire [31:0]   res_lo_lo_hi_lo_61 = {dataGroup_5_61, dataGroup_4_61};
  wire [31:0]   res_lo_lo_hi_hi_61 = {dataGroup_7_61, dataGroup_6_61};
  wire [63:0]   res_lo_lo_hi_61 = {res_lo_lo_hi_hi_61, res_lo_lo_hi_lo_61};
  wire [127:0]  res_lo_lo_61 = {res_lo_lo_hi_61, res_lo_lo_lo_61};
  wire [31:0]   res_lo_hi_lo_lo_61 = {dataGroup_9_61, dataGroup_8_61};
  wire [31:0]   res_lo_hi_lo_hi_61 = {dataGroup_11_61, dataGroup_10_61};
  wire [63:0]   res_lo_hi_lo_61 = {res_lo_hi_lo_hi_61, res_lo_hi_lo_lo_61};
  wire [31:0]   res_lo_hi_hi_lo_61 = {dataGroup_13_61, dataGroup_12_61};
  wire [31:0]   res_lo_hi_hi_hi_61 = {dataGroup_15_61, dataGroup_14_61};
  wire [63:0]   res_lo_hi_hi_61 = {res_lo_hi_hi_hi_61, res_lo_hi_hi_lo_61};
  wire [127:0]  res_lo_hi_61 = {res_lo_hi_hi_61, res_lo_hi_lo_61};
  wire [255:0]  res_lo_61 = {res_lo_hi_61, res_lo_lo_61};
  wire [31:0]   res_hi_lo_lo_lo_61 = {dataGroup_17_61, dataGroup_16_61};
  wire [31:0]   res_hi_lo_lo_hi_61 = {dataGroup_19_61, dataGroup_18_61};
  wire [63:0]   res_hi_lo_lo_61 = {res_hi_lo_lo_hi_61, res_hi_lo_lo_lo_61};
  wire [31:0]   res_hi_lo_hi_lo_61 = {dataGroup_21_61, dataGroup_20_61};
  wire [31:0]   res_hi_lo_hi_hi_61 = {dataGroup_23_61, dataGroup_22_61};
  wire [63:0]   res_hi_lo_hi_61 = {res_hi_lo_hi_hi_61, res_hi_lo_hi_lo_61};
  wire [127:0]  res_hi_lo_61 = {res_hi_lo_hi_61, res_hi_lo_lo_61};
  wire [31:0]   res_hi_hi_lo_lo_61 = {dataGroup_25_61, dataGroup_24_61};
  wire [31:0]   res_hi_hi_lo_hi_61 = {dataGroup_27_61, dataGroup_26_61};
  wire [63:0]   res_hi_hi_lo_61 = {res_hi_hi_lo_hi_61, res_hi_hi_lo_lo_61};
  wire [31:0]   res_hi_hi_hi_lo_61 = {dataGroup_29_61, dataGroup_28_61};
  wire [31:0]   res_hi_hi_hi_hi_61 = {dataGroup_31_61, dataGroup_30_61};
  wire [63:0]   res_hi_hi_hi_61 = {res_hi_hi_hi_hi_61, res_hi_hi_hi_lo_61};
  wire [127:0]  res_hi_hi_61 = {res_hi_hi_hi_61, res_hi_hi_lo_61};
  wire [255:0]  res_hi_61 = {res_hi_hi_61, res_hi_lo_61};
  wire [511:0]  res_116 = {res_hi_61, res_lo_61};
  wire [2047:0] dataGroup_lo_3136 = {dataGroup_lo_hi_3136, dataGroup_lo_lo_3136};
  wire [2047:0] dataGroup_hi_3136 = {dataGroup_hi_hi_3136, dataGroup_hi_lo_3136};
  wire [15:0]   dataGroup_0_62 = dataGroup_lo_3136[95:80];
  wire [2047:0] dataGroup_lo_3137 = {dataGroup_lo_hi_3137, dataGroup_lo_lo_3137};
  wire [2047:0] dataGroup_hi_3137 = {dataGroup_hi_hi_3137, dataGroup_hi_lo_3137};
  wire [15:0]   dataGroup_1_62 = dataGroup_lo_3137[207:192];
  wire [2047:0] dataGroup_lo_3138 = {dataGroup_lo_hi_3138, dataGroup_lo_lo_3138};
  wire [2047:0] dataGroup_hi_3138 = {dataGroup_hi_hi_3138, dataGroup_hi_lo_3138};
  wire [15:0]   dataGroup_2_62 = dataGroup_lo_3138[319:304];
  wire [2047:0] dataGroup_lo_3139 = {dataGroup_lo_hi_3139, dataGroup_lo_lo_3139};
  wire [2047:0] dataGroup_hi_3139 = {dataGroup_hi_hi_3139, dataGroup_hi_lo_3139};
  wire [15:0]   dataGroup_3_62 = dataGroup_lo_3139[431:416];
  wire [2047:0] dataGroup_lo_3140 = {dataGroup_lo_hi_3140, dataGroup_lo_lo_3140};
  wire [2047:0] dataGroup_hi_3140 = {dataGroup_hi_hi_3140, dataGroup_hi_lo_3140};
  wire [15:0]   dataGroup_4_62 = dataGroup_lo_3140[543:528];
  wire [2047:0] dataGroup_lo_3141 = {dataGroup_lo_hi_3141, dataGroup_lo_lo_3141};
  wire [2047:0] dataGroup_hi_3141 = {dataGroup_hi_hi_3141, dataGroup_hi_lo_3141};
  wire [15:0]   dataGroup_5_62 = dataGroup_lo_3141[655:640];
  wire [2047:0] dataGroup_lo_3142 = {dataGroup_lo_hi_3142, dataGroup_lo_lo_3142};
  wire [2047:0] dataGroup_hi_3142 = {dataGroup_hi_hi_3142, dataGroup_hi_lo_3142};
  wire [15:0]   dataGroup_6_62 = dataGroup_lo_3142[767:752];
  wire [2047:0] dataGroup_lo_3143 = {dataGroup_lo_hi_3143, dataGroup_lo_lo_3143};
  wire [2047:0] dataGroup_hi_3143 = {dataGroup_hi_hi_3143, dataGroup_hi_lo_3143};
  wire [15:0]   dataGroup_7_62 = dataGroup_lo_3143[879:864];
  wire [2047:0] dataGroup_lo_3144 = {dataGroup_lo_hi_3144, dataGroup_lo_lo_3144};
  wire [2047:0] dataGroup_hi_3144 = {dataGroup_hi_hi_3144, dataGroup_hi_lo_3144};
  wire [15:0]   dataGroup_8_62 = dataGroup_lo_3144[991:976];
  wire [2047:0] dataGroup_lo_3145 = {dataGroup_lo_hi_3145, dataGroup_lo_lo_3145};
  wire [2047:0] dataGroup_hi_3145 = {dataGroup_hi_hi_3145, dataGroup_hi_lo_3145};
  wire [15:0]   dataGroup_9_62 = dataGroup_lo_3145[1103:1088];
  wire [2047:0] dataGroup_lo_3146 = {dataGroup_lo_hi_3146, dataGroup_lo_lo_3146};
  wire [2047:0] dataGroup_hi_3146 = {dataGroup_hi_hi_3146, dataGroup_hi_lo_3146};
  wire [15:0]   dataGroup_10_62 = dataGroup_lo_3146[1215:1200];
  wire [2047:0] dataGroup_lo_3147 = {dataGroup_lo_hi_3147, dataGroup_lo_lo_3147};
  wire [2047:0] dataGroup_hi_3147 = {dataGroup_hi_hi_3147, dataGroup_hi_lo_3147};
  wire [15:0]   dataGroup_11_62 = dataGroup_lo_3147[1327:1312];
  wire [2047:0] dataGroup_lo_3148 = {dataGroup_lo_hi_3148, dataGroup_lo_lo_3148};
  wire [2047:0] dataGroup_hi_3148 = {dataGroup_hi_hi_3148, dataGroup_hi_lo_3148};
  wire [15:0]   dataGroup_12_62 = dataGroup_lo_3148[1439:1424];
  wire [2047:0] dataGroup_lo_3149 = {dataGroup_lo_hi_3149, dataGroup_lo_lo_3149};
  wire [2047:0] dataGroup_hi_3149 = {dataGroup_hi_hi_3149, dataGroup_hi_lo_3149};
  wire [15:0]   dataGroup_13_62 = dataGroup_lo_3149[1551:1536];
  wire [2047:0] dataGroup_lo_3150 = {dataGroup_lo_hi_3150, dataGroup_lo_lo_3150};
  wire [2047:0] dataGroup_hi_3150 = {dataGroup_hi_hi_3150, dataGroup_hi_lo_3150};
  wire [15:0]   dataGroup_14_62 = dataGroup_lo_3150[1663:1648];
  wire [2047:0] dataGroup_lo_3151 = {dataGroup_lo_hi_3151, dataGroup_lo_lo_3151};
  wire [2047:0] dataGroup_hi_3151 = {dataGroup_hi_hi_3151, dataGroup_hi_lo_3151};
  wire [15:0]   dataGroup_15_62 = dataGroup_lo_3151[1775:1760];
  wire [2047:0] dataGroup_lo_3152 = {dataGroup_lo_hi_3152, dataGroup_lo_lo_3152};
  wire [2047:0] dataGroup_hi_3152 = {dataGroup_hi_hi_3152, dataGroup_hi_lo_3152};
  wire [15:0]   dataGroup_16_62 = dataGroup_lo_3152[1887:1872];
  wire [2047:0] dataGroup_lo_3153 = {dataGroup_lo_hi_3153, dataGroup_lo_lo_3153};
  wire [2047:0] dataGroup_hi_3153 = {dataGroup_hi_hi_3153, dataGroup_hi_lo_3153};
  wire [15:0]   dataGroup_17_62 = dataGroup_lo_3153[1999:1984];
  wire [2047:0] dataGroup_lo_3154 = {dataGroup_lo_hi_3154, dataGroup_lo_lo_3154};
  wire [2047:0] dataGroup_hi_3154 = {dataGroup_hi_hi_3154, dataGroup_hi_lo_3154};
  wire [15:0]   dataGroup_18_62 = dataGroup_hi_3154[63:48];
  wire [2047:0] dataGroup_lo_3155 = {dataGroup_lo_hi_3155, dataGroup_lo_lo_3155};
  wire [2047:0] dataGroup_hi_3155 = {dataGroup_hi_hi_3155, dataGroup_hi_lo_3155};
  wire [15:0]   dataGroup_19_62 = dataGroup_hi_3155[175:160];
  wire [2047:0] dataGroup_lo_3156 = {dataGroup_lo_hi_3156, dataGroup_lo_lo_3156};
  wire [2047:0] dataGroup_hi_3156 = {dataGroup_hi_hi_3156, dataGroup_hi_lo_3156};
  wire [15:0]   dataGroup_20_62 = dataGroup_hi_3156[287:272];
  wire [2047:0] dataGroup_lo_3157 = {dataGroup_lo_hi_3157, dataGroup_lo_lo_3157};
  wire [2047:0] dataGroup_hi_3157 = {dataGroup_hi_hi_3157, dataGroup_hi_lo_3157};
  wire [15:0]   dataGroup_21_62 = dataGroup_hi_3157[399:384];
  wire [2047:0] dataGroup_lo_3158 = {dataGroup_lo_hi_3158, dataGroup_lo_lo_3158};
  wire [2047:0] dataGroup_hi_3158 = {dataGroup_hi_hi_3158, dataGroup_hi_lo_3158};
  wire [15:0]   dataGroup_22_62 = dataGroup_hi_3158[511:496];
  wire [2047:0] dataGroup_lo_3159 = {dataGroup_lo_hi_3159, dataGroup_lo_lo_3159};
  wire [2047:0] dataGroup_hi_3159 = {dataGroup_hi_hi_3159, dataGroup_hi_lo_3159};
  wire [15:0]   dataGroup_23_62 = dataGroup_hi_3159[623:608];
  wire [2047:0] dataGroup_lo_3160 = {dataGroup_lo_hi_3160, dataGroup_lo_lo_3160};
  wire [2047:0] dataGroup_hi_3160 = {dataGroup_hi_hi_3160, dataGroup_hi_lo_3160};
  wire [15:0]   dataGroup_24_62 = dataGroup_hi_3160[735:720];
  wire [2047:0] dataGroup_lo_3161 = {dataGroup_lo_hi_3161, dataGroup_lo_lo_3161};
  wire [2047:0] dataGroup_hi_3161 = {dataGroup_hi_hi_3161, dataGroup_hi_lo_3161};
  wire [15:0]   dataGroup_25_62 = dataGroup_hi_3161[847:832];
  wire [2047:0] dataGroup_lo_3162 = {dataGroup_lo_hi_3162, dataGroup_lo_lo_3162};
  wire [2047:0] dataGroup_hi_3162 = {dataGroup_hi_hi_3162, dataGroup_hi_lo_3162};
  wire [15:0]   dataGroup_26_62 = dataGroup_hi_3162[959:944];
  wire [2047:0] dataGroup_lo_3163 = {dataGroup_lo_hi_3163, dataGroup_lo_lo_3163};
  wire [2047:0] dataGroup_hi_3163 = {dataGroup_hi_hi_3163, dataGroup_hi_lo_3163};
  wire [15:0]   dataGroup_27_62 = dataGroup_hi_3163[1071:1056];
  wire [2047:0] dataGroup_lo_3164 = {dataGroup_lo_hi_3164, dataGroup_lo_lo_3164};
  wire [2047:0] dataGroup_hi_3164 = {dataGroup_hi_hi_3164, dataGroup_hi_lo_3164};
  wire [15:0]   dataGroup_28_62 = dataGroup_hi_3164[1183:1168];
  wire [2047:0] dataGroup_lo_3165 = {dataGroup_lo_hi_3165, dataGroup_lo_lo_3165};
  wire [2047:0] dataGroup_hi_3165 = {dataGroup_hi_hi_3165, dataGroup_hi_lo_3165};
  wire [15:0]   dataGroup_29_62 = dataGroup_hi_3165[1295:1280];
  wire [2047:0] dataGroup_lo_3166 = {dataGroup_lo_hi_3166, dataGroup_lo_lo_3166};
  wire [2047:0] dataGroup_hi_3166 = {dataGroup_hi_hi_3166, dataGroup_hi_lo_3166};
  wire [15:0]   dataGroup_30_62 = dataGroup_hi_3166[1407:1392];
  wire [2047:0] dataGroup_lo_3167 = {dataGroup_lo_hi_3167, dataGroup_lo_lo_3167};
  wire [2047:0] dataGroup_hi_3167 = {dataGroup_hi_hi_3167, dataGroup_hi_lo_3167};
  wire [15:0]   dataGroup_31_62 = dataGroup_hi_3167[1519:1504];
  wire [31:0]   res_lo_lo_lo_lo_62 = {dataGroup_1_62, dataGroup_0_62};
  wire [31:0]   res_lo_lo_lo_hi_62 = {dataGroup_3_62, dataGroup_2_62};
  wire [63:0]   res_lo_lo_lo_62 = {res_lo_lo_lo_hi_62, res_lo_lo_lo_lo_62};
  wire [31:0]   res_lo_lo_hi_lo_62 = {dataGroup_5_62, dataGroup_4_62};
  wire [31:0]   res_lo_lo_hi_hi_62 = {dataGroup_7_62, dataGroup_6_62};
  wire [63:0]   res_lo_lo_hi_62 = {res_lo_lo_hi_hi_62, res_lo_lo_hi_lo_62};
  wire [127:0]  res_lo_lo_62 = {res_lo_lo_hi_62, res_lo_lo_lo_62};
  wire [31:0]   res_lo_hi_lo_lo_62 = {dataGroup_9_62, dataGroup_8_62};
  wire [31:0]   res_lo_hi_lo_hi_62 = {dataGroup_11_62, dataGroup_10_62};
  wire [63:0]   res_lo_hi_lo_62 = {res_lo_hi_lo_hi_62, res_lo_hi_lo_lo_62};
  wire [31:0]   res_lo_hi_hi_lo_62 = {dataGroup_13_62, dataGroup_12_62};
  wire [31:0]   res_lo_hi_hi_hi_62 = {dataGroup_15_62, dataGroup_14_62};
  wire [63:0]   res_lo_hi_hi_62 = {res_lo_hi_hi_hi_62, res_lo_hi_hi_lo_62};
  wire [127:0]  res_lo_hi_62 = {res_lo_hi_hi_62, res_lo_hi_lo_62};
  wire [255:0]  res_lo_62 = {res_lo_hi_62, res_lo_lo_62};
  wire [31:0]   res_hi_lo_lo_lo_62 = {dataGroup_17_62, dataGroup_16_62};
  wire [31:0]   res_hi_lo_lo_hi_62 = {dataGroup_19_62, dataGroup_18_62};
  wire [63:0]   res_hi_lo_lo_62 = {res_hi_lo_lo_hi_62, res_hi_lo_lo_lo_62};
  wire [31:0]   res_hi_lo_hi_lo_62 = {dataGroup_21_62, dataGroup_20_62};
  wire [31:0]   res_hi_lo_hi_hi_62 = {dataGroup_23_62, dataGroup_22_62};
  wire [63:0]   res_hi_lo_hi_62 = {res_hi_lo_hi_hi_62, res_hi_lo_hi_lo_62};
  wire [127:0]  res_hi_lo_62 = {res_hi_lo_hi_62, res_hi_lo_lo_62};
  wire [31:0]   res_hi_hi_lo_lo_62 = {dataGroup_25_62, dataGroup_24_62};
  wire [31:0]   res_hi_hi_lo_hi_62 = {dataGroup_27_62, dataGroup_26_62};
  wire [63:0]   res_hi_hi_lo_62 = {res_hi_hi_lo_hi_62, res_hi_hi_lo_lo_62};
  wire [31:0]   res_hi_hi_hi_lo_62 = {dataGroup_29_62, dataGroup_28_62};
  wire [31:0]   res_hi_hi_hi_hi_62 = {dataGroup_31_62, dataGroup_30_62};
  wire [63:0]   res_hi_hi_hi_62 = {res_hi_hi_hi_hi_62, res_hi_hi_hi_lo_62};
  wire [127:0]  res_hi_hi_62 = {res_hi_hi_hi_62, res_hi_hi_lo_62};
  wire [255:0]  res_hi_62 = {res_hi_hi_62, res_hi_lo_62};
  wire [511:0]  res_117 = {res_hi_62, res_lo_62};
  wire [2047:0] dataGroup_lo_3168 = {dataGroup_lo_hi_3168, dataGroup_lo_lo_3168};
  wire [2047:0] dataGroup_hi_3168 = {dataGroup_hi_hi_3168, dataGroup_hi_lo_3168};
  wire [15:0]   dataGroup_0_63 = dataGroup_lo_3168[111:96];
  wire [2047:0] dataGroup_lo_3169 = {dataGroup_lo_hi_3169, dataGroup_lo_lo_3169};
  wire [2047:0] dataGroup_hi_3169 = {dataGroup_hi_hi_3169, dataGroup_hi_lo_3169};
  wire [15:0]   dataGroup_1_63 = dataGroup_lo_3169[223:208];
  wire [2047:0] dataGroup_lo_3170 = {dataGroup_lo_hi_3170, dataGroup_lo_lo_3170};
  wire [2047:0] dataGroup_hi_3170 = {dataGroup_hi_hi_3170, dataGroup_hi_lo_3170};
  wire [15:0]   dataGroup_2_63 = dataGroup_lo_3170[335:320];
  wire [2047:0] dataGroup_lo_3171 = {dataGroup_lo_hi_3171, dataGroup_lo_lo_3171};
  wire [2047:0] dataGroup_hi_3171 = {dataGroup_hi_hi_3171, dataGroup_hi_lo_3171};
  wire [15:0]   dataGroup_3_63 = dataGroup_lo_3171[447:432];
  wire [2047:0] dataGroup_lo_3172 = {dataGroup_lo_hi_3172, dataGroup_lo_lo_3172};
  wire [2047:0] dataGroup_hi_3172 = {dataGroup_hi_hi_3172, dataGroup_hi_lo_3172};
  wire [15:0]   dataGroup_4_63 = dataGroup_lo_3172[559:544];
  wire [2047:0] dataGroup_lo_3173 = {dataGroup_lo_hi_3173, dataGroup_lo_lo_3173};
  wire [2047:0] dataGroup_hi_3173 = {dataGroup_hi_hi_3173, dataGroup_hi_lo_3173};
  wire [15:0]   dataGroup_5_63 = dataGroup_lo_3173[671:656];
  wire [2047:0] dataGroup_lo_3174 = {dataGroup_lo_hi_3174, dataGroup_lo_lo_3174};
  wire [2047:0] dataGroup_hi_3174 = {dataGroup_hi_hi_3174, dataGroup_hi_lo_3174};
  wire [15:0]   dataGroup_6_63 = dataGroup_lo_3174[783:768];
  wire [2047:0] dataGroup_lo_3175 = {dataGroup_lo_hi_3175, dataGroup_lo_lo_3175};
  wire [2047:0] dataGroup_hi_3175 = {dataGroup_hi_hi_3175, dataGroup_hi_lo_3175};
  wire [15:0]   dataGroup_7_63 = dataGroup_lo_3175[895:880];
  wire [2047:0] dataGroup_lo_3176 = {dataGroup_lo_hi_3176, dataGroup_lo_lo_3176};
  wire [2047:0] dataGroup_hi_3176 = {dataGroup_hi_hi_3176, dataGroup_hi_lo_3176};
  wire [15:0]   dataGroup_8_63 = dataGroup_lo_3176[1007:992];
  wire [2047:0] dataGroup_lo_3177 = {dataGroup_lo_hi_3177, dataGroup_lo_lo_3177};
  wire [2047:0] dataGroup_hi_3177 = {dataGroup_hi_hi_3177, dataGroup_hi_lo_3177};
  wire [15:0]   dataGroup_9_63 = dataGroup_lo_3177[1119:1104];
  wire [2047:0] dataGroup_lo_3178 = {dataGroup_lo_hi_3178, dataGroup_lo_lo_3178};
  wire [2047:0] dataGroup_hi_3178 = {dataGroup_hi_hi_3178, dataGroup_hi_lo_3178};
  wire [15:0]   dataGroup_10_63 = dataGroup_lo_3178[1231:1216];
  wire [2047:0] dataGroup_lo_3179 = {dataGroup_lo_hi_3179, dataGroup_lo_lo_3179};
  wire [2047:0] dataGroup_hi_3179 = {dataGroup_hi_hi_3179, dataGroup_hi_lo_3179};
  wire [15:0]   dataGroup_11_63 = dataGroup_lo_3179[1343:1328];
  wire [2047:0] dataGroup_lo_3180 = {dataGroup_lo_hi_3180, dataGroup_lo_lo_3180};
  wire [2047:0] dataGroup_hi_3180 = {dataGroup_hi_hi_3180, dataGroup_hi_lo_3180};
  wire [15:0]   dataGroup_12_63 = dataGroup_lo_3180[1455:1440];
  wire [2047:0] dataGroup_lo_3181 = {dataGroup_lo_hi_3181, dataGroup_lo_lo_3181};
  wire [2047:0] dataGroup_hi_3181 = {dataGroup_hi_hi_3181, dataGroup_hi_lo_3181};
  wire [15:0]   dataGroup_13_63 = dataGroup_lo_3181[1567:1552];
  wire [2047:0] dataGroup_lo_3182 = {dataGroup_lo_hi_3182, dataGroup_lo_lo_3182};
  wire [2047:0] dataGroup_hi_3182 = {dataGroup_hi_hi_3182, dataGroup_hi_lo_3182};
  wire [15:0]   dataGroup_14_63 = dataGroup_lo_3182[1679:1664];
  wire [2047:0] dataGroup_lo_3183 = {dataGroup_lo_hi_3183, dataGroup_lo_lo_3183};
  wire [2047:0] dataGroup_hi_3183 = {dataGroup_hi_hi_3183, dataGroup_hi_lo_3183};
  wire [15:0]   dataGroup_15_63 = dataGroup_lo_3183[1791:1776];
  wire [2047:0] dataGroup_lo_3184 = {dataGroup_lo_hi_3184, dataGroup_lo_lo_3184};
  wire [2047:0] dataGroup_hi_3184 = {dataGroup_hi_hi_3184, dataGroup_hi_lo_3184};
  wire [15:0]   dataGroup_16_63 = dataGroup_lo_3184[1903:1888];
  wire [2047:0] dataGroup_lo_3185 = {dataGroup_lo_hi_3185, dataGroup_lo_lo_3185};
  wire [2047:0] dataGroup_hi_3185 = {dataGroup_hi_hi_3185, dataGroup_hi_lo_3185};
  wire [15:0]   dataGroup_17_63 = dataGroup_lo_3185[2015:2000];
  wire [2047:0] dataGroup_lo_3186 = {dataGroup_lo_hi_3186, dataGroup_lo_lo_3186};
  wire [2047:0] dataGroup_hi_3186 = {dataGroup_hi_hi_3186, dataGroup_hi_lo_3186};
  wire [15:0]   dataGroup_18_63 = dataGroup_hi_3186[79:64];
  wire [2047:0] dataGroup_lo_3187 = {dataGroup_lo_hi_3187, dataGroup_lo_lo_3187};
  wire [2047:0] dataGroup_hi_3187 = {dataGroup_hi_hi_3187, dataGroup_hi_lo_3187};
  wire [15:0]   dataGroup_19_63 = dataGroup_hi_3187[191:176];
  wire [2047:0] dataGroup_lo_3188 = {dataGroup_lo_hi_3188, dataGroup_lo_lo_3188};
  wire [2047:0] dataGroup_hi_3188 = {dataGroup_hi_hi_3188, dataGroup_hi_lo_3188};
  wire [15:0]   dataGroup_20_63 = dataGroup_hi_3188[303:288];
  wire [2047:0] dataGroup_lo_3189 = {dataGroup_lo_hi_3189, dataGroup_lo_lo_3189};
  wire [2047:0] dataGroup_hi_3189 = {dataGroup_hi_hi_3189, dataGroup_hi_lo_3189};
  wire [15:0]   dataGroup_21_63 = dataGroup_hi_3189[415:400];
  wire [2047:0] dataGroup_lo_3190 = {dataGroup_lo_hi_3190, dataGroup_lo_lo_3190};
  wire [2047:0] dataGroup_hi_3190 = {dataGroup_hi_hi_3190, dataGroup_hi_lo_3190};
  wire [15:0]   dataGroup_22_63 = dataGroup_hi_3190[527:512];
  wire [2047:0] dataGroup_lo_3191 = {dataGroup_lo_hi_3191, dataGroup_lo_lo_3191};
  wire [2047:0] dataGroup_hi_3191 = {dataGroup_hi_hi_3191, dataGroup_hi_lo_3191};
  wire [15:0]   dataGroup_23_63 = dataGroup_hi_3191[639:624];
  wire [2047:0] dataGroup_lo_3192 = {dataGroup_lo_hi_3192, dataGroup_lo_lo_3192};
  wire [2047:0] dataGroup_hi_3192 = {dataGroup_hi_hi_3192, dataGroup_hi_lo_3192};
  wire [15:0]   dataGroup_24_63 = dataGroup_hi_3192[751:736];
  wire [2047:0] dataGroup_lo_3193 = {dataGroup_lo_hi_3193, dataGroup_lo_lo_3193};
  wire [2047:0] dataGroup_hi_3193 = {dataGroup_hi_hi_3193, dataGroup_hi_lo_3193};
  wire [15:0]   dataGroup_25_63 = dataGroup_hi_3193[863:848];
  wire [2047:0] dataGroup_lo_3194 = {dataGroup_lo_hi_3194, dataGroup_lo_lo_3194};
  wire [2047:0] dataGroup_hi_3194 = {dataGroup_hi_hi_3194, dataGroup_hi_lo_3194};
  wire [15:0]   dataGroup_26_63 = dataGroup_hi_3194[975:960];
  wire [2047:0] dataGroup_lo_3195 = {dataGroup_lo_hi_3195, dataGroup_lo_lo_3195};
  wire [2047:0] dataGroup_hi_3195 = {dataGroup_hi_hi_3195, dataGroup_hi_lo_3195};
  wire [15:0]   dataGroup_27_63 = dataGroup_hi_3195[1087:1072];
  wire [2047:0] dataGroup_lo_3196 = {dataGroup_lo_hi_3196, dataGroup_lo_lo_3196};
  wire [2047:0] dataGroup_hi_3196 = {dataGroup_hi_hi_3196, dataGroup_hi_lo_3196};
  wire [15:0]   dataGroup_28_63 = dataGroup_hi_3196[1199:1184];
  wire [2047:0] dataGroup_lo_3197 = {dataGroup_lo_hi_3197, dataGroup_lo_lo_3197};
  wire [2047:0] dataGroup_hi_3197 = {dataGroup_hi_hi_3197, dataGroup_hi_lo_3197};
  wire [15:0]   dataGroup_29_63 = dataGroup_hi_3197[1311:1296];
  wire [2047:0] dataGroup_lo_3198 = {dataGroup_lo_hi_3198, dataGroup_lo_lo_3198};
  wire [2047:0] dataGroup_hi_3198 = {dataGroup_hi_hi_3198, dataGroup_hi_lo_3198};
  wire [15:0]   dataGroup_30_63 = dataGroup_hi_3198[1423:1408];
  wire [2047:0] dataGroup_lo_3199 = {dataGroup_lo_hi_3199, dataGroup_lo_lo_3199};
  wire [2047:0] dataGroup_hi_3199 = {dataGroup_hi_hi_3199, dataGroup_hi_lo_3199};
  wire [15:0]   dataGroup_31_63 = dataGroup_hi_3199[1535:1520];
  wire [31:0]   res_lo_lo_lo_lo_63 = {dataGroup_1_63, dataGroup_0_63};
  wire [31:0]   res_lo_lo_lo_hi_63 = {dataGroup_3_63, dataGroup_2_63};
  wire [63:0]   res_lo_lo_lo_63 = {res_lo_lo_lo_hi_63, res_lo_lo_lo_lo_63};
  wire [31:0]   res_lo_lo_hi_lo_63 = {dataGroup_5_63, dataGroup_4_63};
  wire [31:0]   res_lo_lo_hi_hi_63 = {dataGroup_7_63, dataGroup_6_63};
  wire [63:0]   res_lo_lo_hi_63 = {res_lo_lo_hi_hi_63, res_lo_lo_hi_lo_63};
  wire [127:0]  res_lo_lo_63 = {res_lo_lo_hi_63, res_lo_lo_lo_63};
  wire [31:0]   res_lo_hi_lo_lo_63 = {dataGroup_9_63, dataGroup_8_63};
  wire [31:0]   res_lo_hi_lo_hi_63 = {dataGroup_11_63, dataGroup_10_63};
  wire [63:0]   res_lo_hi_lo_63 = {res_lo_hi_lo_hi_63, res_lo_hi_lo_lo_63};
  wire [31:0]   res_lo_hi_hi_lo_63 = {dataGroup_13_63, dataGroup_12_63};
  wire [31:0]   res_lo_hi_hi_hi_63 = {dataGroup_15_63, dataGroup_14_63};
  wire [63:0]   res_lo_hi_hi_63 = {res_lo_hi_hi_hi_63, res_lo_hi_hi_lo_63};
  wire [127:0]  res_lo_hi_63 = {res_lo_hi_hi_63, res_lo_hi_lo_63};
  wire [255:0]  res_lo_63 = {res_lo_hi_63, res_lo_lo_63};
  wire [31:0]   res_hi_lo_lo_lo_63 = {dataGroup_17_63, dataGroup_16_63};
  wire [31:0]   res_hi_lo_lo_hi_63 = {dataGroup_19_63, dataGroup_18_63};
  wire [63:0]   res_hi_lo_lo_63 = {res_hi_lo_lo_hi_63, res_hi_lo_lo_lo_63};
  wire [31:0]   res_hi_lo_hi_lo_63 = {dataGroup_21_63, dataGroup_20_63};
  wire [31:0]   res_hi_lo_hi_hi_63 = {dataGroup_23_63, dataGroup_22_63};
  wire [63:0]   res_hi_lo_hi_63 = {res_hi_lo_hi_hi_63, res_hi_lo_hi_lo_63};
  wire [127:0]  res_hi_lo_63 = {res_hi_lo_hi_63, res_hi_lo_lo_63};
  wire [31:0]   res_hi_hi_lo_lo_63 = {dataGroup_25_63, dataGroup_24_63};
  wire [31:0]   res_hi_hi_lo_hi_63 = {dataGroup_27_63, dataGroup_26_63};
  wire [63:0]   res_hi_hi_lo_63 = {res_hi_hi_lo_hi_63, res_hi_hi_lo_lo_63};
  wire [31:0]   res_hi_hi_hi_lo_63 = {dataGroup_29_63, dataGroup_28_63};
  wire [31:0]   res_hi_hi_hi_hi_63 = {dataGroup_31_63, dataGroup_30_63};
  wire [63:0]   res_hi_hi_hi_63 = {res_hi_hi_hi_hi_63, res_hi_hi_hi_lo_63};
  wire [127:0]  res_hi_hi_63 = {res_hi_hi_hi_63, res_hi_hi_lo_63};
  wire [255:0]  res_hi_63 = {res_hi_hi_63, res_hi_lo_63};
  wire [511:0]  res_118 = {res_hi_63, res_lo_63};
  wire [1023:0] lo_lo_14 = {res_113, res_112};
  wire [1023:0] lo_hi_14 = {res_115, res_114};
  wire [2047:0] lo_14 = {lo_hi_14, lo_lo_14};
  wire [1023:0] hi_lo_14 = {res_117, res_116};
  wire [1023:0] hi_hi_14 = {512'h0, res_118};
  wire [2047:0] hi_14 = {hi_hi_14, hi_lo_14};
  wire [4095:0] regroupLoadData_1_6 = {hi_14, lo_14};
  wire [2047:0] dataGroup_lo_3200 = {dataGroup_lo_hi_3200, dataGroup_lo_lo_3200};
  wire [2047:0] dataGroup_hi_3200 = {dataGroup_hi_hi_3200, dataGroup_hi_lo_3200};
  wire [15:0]   dataGroup_0_64 = dataGroup_lo_3200[15:0];
  wire [2047:0] dataGroup_lo_3201 = {dataGroup_lo_hi_3201, dataGroup_lo_lo_3201};
  wire [2047:0] dataGroup_hi_3201 = {dataGroup_hi_hi_3201, dataGroup_hi_lo_3201};
  wire [15:0]   dataGroup_1_64 = dataGroup_lo_3201[143:128];
  wire [2047:0] dataGroup_lo_3202 = {dataGroup_lo_hi_3202, dataGroup_lo_lo_3202};
  wire [2047:0] dataGroup_hi_3202 = {dataGroup_hi_hi_3202, dataGroup_hi_lo_3202};
  wire [15:0]   dataGroup_2_64 = dataGroup_lo_3202[271:256];
  wire [2047:0] dataGroup_lo_3203 = {dataGroup_lo_hi_3203, dataGroup_lo_lo_3203};
  wire [2047:0] dataGroup_hi_3203 = {dataGroup_hi_hi_3203, dataGroup_hi_lo_3203};
  wire [15:0]   dataGroup_3_64 = dataGroup_lo_3203[399:384];
  wire [2047:0] dataGroup_lo_3204 = {dataGroup_lo_hi_3204, dataGroup_lo_lo_3204};
  wire [2047:0] dataGroup_hi_3204 = {dataGroup_hi_hi_3204, dataGroup_hi_lo_3204};
  wire [15:0]   dataGroup_4_64 = dataGroup_lo_3204[527:512];
  wire [2047:0] dataGroup_lo_3205 = {dataGroup_lo_hi_3205, dataGroup_lo_lo_3205};
  wire [2047:0] dataGroup_hi_3205 = {dataGroup_hi_hi_3205, dataGroup_hi_lo_3205};
  wire [15:0]   dataGroup_5_64 = dataGroup_lo_3205[655:640];
  wire [2047:0] dataGroup_lo_3206 = {dataGroup_lo_hi_3206, dataGroup_lo_lo_3206};
  wire [2047:0] dataGroup_hi_3206 = {dataGroup_hi_hi_3206, dataGroup_hi_lo_3206};
  wire [15:0]   dataGroup_6_64 = dataGroup_lo_3206[783:768];
  wire [2047:0] dataGroup_lo_3207 = {dataGroup_lo_hi_3207, dataGroup_lo_lo_3207};
  wire [2047:0] dataGroup_hi_3207 = {dataGroup_hi_hi_3207, dataGroup_hi_lo_3207};
  wire [15:0]   dataGroup_7_64 = dataGroup_lo_3207[911:896];
  wire [2047:0] dataGroup_lo_3208 = {dataGroup_lo_hi_3208, dataGroup_lo_lo_3208};
  wire [2047:0] dataGroup_hi_3208 = {dataGroup_hi_hi_3208, dataGroup_hi_lo_3208};
  wire [15:0]   dataGroup_8_64 = dataGroup_lo_3208[1039:1024];
  wire [2047:0] dataGroup_lo_3209 = {dataGroup_lo_hi_3209, dataGroup_lo_lo_3209};
  wire [2047:0] dataGroup_hi_3209 = {dataGroup_hi_hi_3209, dataGroup_hi_lo_3209};
  wire [15:0]   dataGroup_9_64 = dataGroup_lo_3209[1167:1152];
  wire [2047:0] dataGroup_lo_3210 = {dataGroup_lo_hi_3210, dataGroup_lo_lo_3210};
  wire [2047:0] dataGroup_hi_3210 = {dataGroup_hi_hi_3210, dataGroup_hi_lo_3210};
  wire [15:0]   dataGroup_10_64 = dataGroup_lo_3210[1295:1280];
  wire [2047:0] dataGroup_lo_3211 = {dataGroup_lo_hi_3211, dataGroup_lo_lo_3211};
  wire [2047:0] dataGroup_hi_3211 = {dataGroup_hi_hi_3211, dataGroup_hi_lo_3211};
  wire [15:0]   dataGroup_11_64 = dataGroup_lo_3211[1423:1408];
  wire [2047:0] dataGroup_lo_3212 = {dataGroup_lo_hi_3212, dataGroup_lo_lo_3212};
  wire [2047:0] dataGroup_hi_3212 = {dataGroup_hi_hi_3212, dataGroup_hi_lo_3212};
  wire [15:0]   dataGroup_12_64 = dataGroup_lo_3212[1551:1536];
  wire [2047:0] dataGroup_lo_3213 = {dataGroup_lo_hi_3213, dataGroup_lo_lo_3213};
  wire [2047:0] dataGroup_hi_3213 = {dataGroup_hi_hi_3213, dataGroup_hi_lo_3213};
  wire [15:0]   dataGroup_13_64 = dataGroup_lo_3213[1679:1664];
  wire [2047:0] dataGroup_lo_3214 = {dataGroup_lo_hi_3214, dataGroup_lo_lo_3214};
  wire [2047:0] dataGroup_hi_3214 = {dataGroup_hi_hi_3214, dataGroup_hi_lo_3214};
  wire [15:0]   dataGroup_14_64 = dataGroup_lo_3214[1807:1792];
  wire [2047:0] dataGroup_lo_3215 = {dataGroup_lo_hi_3215, dataGroup_lo_lo_3215};
  wire [2047:0] dataGroup_hi_3215 = {dataGroup_hi_hi_3215, dataGroup_hi_lo_3215};
  wire [15:0]   dataGroup_15_64 = dataGroup_lo_3215[1935:1920];
  wire [2047:0] dataGroup_lo_3216 = {dataGroup_lo_hi_3216, dataGroup_lo_lo_3216};
  wire [2047:0] dataGroup_hi_3216 = {dataGroup_hi_hi_3216, dataGroup_hi_lo_3216};
  wire [15:0]   dataGroup_16_64 = dataGroup_hi_3216[15:0];
  wire [2047:0] dataGroup_lo_3217 = {dataGroup_lo_hi_3217, dataGroup_lo_lo_3217};
  wire [2047:0] dataGroup_hi_3217 = {dataGroup_hi_hi_3217, dataGroup_hi_lo_3217};
  wire [15:0]   dataGroup_17_64 = dataGroup_hi_3217[143:128];
  wire [2047:0] dataGroup_lo_3218 = {dataGroup_lo_hi_3218, dataGroup_lo_lo_3218};
  wire [2047:0] dataGroup_hi_3218 = {dataGroup_hi_hi_3218, dataGroup_hi_lo_3218};
  wire [15:0]   dataGroup_18_64 = dataGroup_hi_3218[271:256];
  wire [2047:0] dataGroup_lo_3219 = {dataGroup_lo_hi_3219, dataGroup_lo_lo_3219};
  wire [2047:0] dataGroup_hi_3219 = {dataGroup_hi_hi_3219, dataGroup_hi_lo_3219};
  wire [15:0]   dataGroup_19_64 = dataGroup_hi_3219[399:384];
  wire [2047:0] dataGroup_lo_3220 = {dataGroup_lo_hi_3220, dataGroup_lo_lo_3220};
  wire [2047:0] dataGroup_hi_3220 = {dataGroup_hi_hi_3220, dataGroup_hi_lo_3220};
  wire [15:0]   dataGroup_20_64 = dataGroup_hi_3220[527:512];
  wire [2047:0] dataGroup_lo_3221 = {dataGroup_lo_hi_3221, dataGroup_lo_lo_3221};
  wire [2047:0] dataGroup_hi_3221 = {dataGroup_hi_hi_3221, dataGroup_hi_lo_3221};
  wire [15:0]   dataGroup_21_64 = dataGroup_hi_3221[655:640];
  wire [2047:0] dataGroup_lo_3222 = {dataGroup_lo_hi_3222, dataGroup_lo_lo_3222};
  wire [2047:0] dataGroup_hi_3222 = {dataGroup_hi_hi_3222, dataGroup_hi_lo_3222};
  wire [15:0]   dataGroup_22_64 = dataGroup_hi_3222[783:768];
  wire [2047:0] dataGroup_lo_3223 = {dataGroup_lo_hi_3223, dataGroup_lo_lo_3223};
  wire [2047:0] dataGroup_hi_3223 = {dataGroup_hi_hi_3223, dataGroup_hi_lo_3223};
  wire [15:0]   dataGroup_23_64 = dataGroup_hi_3223[911:896];
  wire [2047:0] dataGroup_lo_3224 = {dataGroup_lo_hi_3224, dataGroup_lo_lo_3224};
  wire [2047:0] dataGroup_hi_3224 = {dataGroup_hi_hi_3224, dataGroup_hi_lo_3224};
  wire [15:0]   dataGroup_24_64 = dataGroup_hi_3224[1039:1024];
  wire [2047:0] dataGroup_lo_3225 = {dataGroup_lo_hi_3225, dataGroup_lo_lo_3225};
  wire [2047:0] dataGroup_hi_3225 = {dataGroup_hi_hi_3225, dataGroup_hi_lo_3225};
  wire [15:0]   dataGroup_25_64 = dataGroup_hi_3225[1167:1152];
  wire [2047:0] dataGroup_lo_3226 = {dataGroup_lo_hi_3226, dataGroup_lo_lo_3226};
  wire [2047:0] dataGroup_hi_3226 = {dataGroup_hi_hi_3226, dataGroup_hi_lo_3226};
  wire [15:0]   dataGroup_26_64 = dataGroup_hi_3226[1295:1280];
  wire [2047:0] dataGroup_lo_3227 = {dataGroup_lo_hi_3227, dataGroup_lo_lo_3227};
  wire [2047:0] dataGroup_hi_3227 = {dataGroup_hi_hi_3227, dataGroup_hi_lo_3227};
  wire [15:0]   dataGroup_27_64 = dataGroup_hi_3227[1423:1408];
  wire [2047:0] dataGroup_lo_3228 = {dataGroup_lo_hi_3228, dataGroup_lo_lo_3228};
  wire [2047:0] dataGroup_hi_3228 = {dataGroup_hi_hi_3228, dataGroup_hi_lo_3228};
  wire [15:0]   dataGroup_28_64 = dataGroup_hi_3228[1551:1536];
  wire [2047:0] dataGroup_lo_3229 = {dataGroup_lo_hi_3229, dataGroup_lo_lo_3229};
  wire [2047:0] dataGroup_hi_3229 = {dataGroup_hi_hi_3229, dataGroup_hi_lo_3229};
  wire [15:0]   dataGroup_29_64 = dataGroup_hi_3229[1679:1664];
  wire [2047:0] dataGroup_lo_3230 = {dataGroup_lo_hi_3230, dataGroup_lo_lo_3230};
  wire [2047:0] dataGroup_hi_3230 = {dataGroup_hi_hi_3230, dataGroup_hi_lo_3230};
  wire [15:0]   dataGroup_30_64 = dataGroup_hi_3230[1807:1792];
  wire [2047:0] dataGroup_lo_3231 = {dataGroup_lo_hi_3231, dataGroup_lo_lo_3231};
  wire [2047:0] dataGroup_hi_3231 = {dataGroup_hi_hi_3231, dataGroup_hi_lo_3231};
  wire [15:0]   dataGroup_31_64 = dataGroup_hi_3231[1935:1920];
  wire [31:0]   res_lo_lo_lo_lo_64 = {dataGroup_1_64, dataGroup_0_64};
  wire [31:0]   res_lo_lo_lo_hi_64 = {dataGroup_3_64, dataGroup_2_64};
  wire [63:0]   res_lo_lo_lo_64 = {res_lo_lo_lo_hi_64, res_lo_lo_lo_lo_64};
  wire [31:0]   res_lo_lo_hi_lo_64 = {dataGroup_5_64, dataGroup_4_64};
  wire [31:0]   res_lo_lo_hi_hi_64 = {dataGroup_7_64, dataGroup_6_64};
  wire [63:0]   res_lo_lo_hi_64 = {res_lo_lo_hi_hi_64, res_lo_lo_hi_lo_64};
  wire [127:0]  res_lo_lo_64 = {res_lo_lo_hi_64, res_lo_lo_lo_64};
  wire [31:0]   res_lo_hi_lo_lo_64 = {dataGroup_9_64, dataGroup_8_64};
  wire [31:0]   res_lo_hi_lo_hi_64 = {dataGroup_11_64, dataGroup_10_64};
  wire [63:0]   res_lo_hi_lo_64 = {res_lo_hi_lo_hi_64, res_lo_hi_lo_lo_64};
  wire [31:0]   res_lo_hi_hi_lo_64 = {dataGroup_13_64, dataGroup_12_64};
  wire [31:0]   res_lo_hi_hi_hi_64 = {dataGroup_15_64, dataGroup_14_64};
  wire [63:0]   res_lo_hi_hi_64 = {res_lo_hi_hi_hi_64, res_lo_hi_hi_lo_64};
  wire [127:0]  res_lo_hi_64 = {res_lo_hi_hi_64, res_lo_hi_lo_64};
  wire [255:0]  res_lo_64 = {res_lo_hi_64, res_lo_lo_64};
  wire [31:0]   res_hi_lo_lo_lo_64 = {dataGroup_17_64, dataGroup_16_64};
  wire [31:0]   res_hi_lo_lo_hi_64 = {dataGroup_19_64, dataGroup_18_64};
  wire [63:0]   res_hi_lo_lo_64 = {res_hi_lo_lo_hi_64, res_hi_lo_lo_lo_64};
  wire [31:0]   res_hi_lo_hi_lo_64 = {dataGroup_21_64, dataGroup_20_64};
  wire [31:0]   res_hi_lo_hi_hi_64 = {dataGroup_23_64, dataGroup_22_64};
  wire [63:0]   res_hi_lo_hi_64 = {res_hi_lo_hi_hi_64, res_hi_lo_hi_lo_64};
  wire [127:0]  res_hi_lo_64 = {res_hi_lo_hi_64, res_hi_lo_lo_64};
  wire [31:0]   res_hi_hi_lo_lo_64 = {dataGroup_25_64, dataGroup_24_64};
  wire [31:0]   res_hi_hi_lo_hi_64 = {dataGroup_27_64, dataGroup_26_64};
  wire [63:0]   res_hi_hi_lo_64 = {res_hi_hi_lo_hi_64, res_hi_hi_lo_lo_64};
  wire [31:0]   res_hi_hi_hi_lo_64 = {dataGroup_29_64, dataGroup_28_64};
  wire [31:0]   res_hi_hi_hi_hi_64 = {dataGroup_31_64, dataGroup_30_64};
  wire [63:0]   res_hi_hi_hi_64 = {res_hi_hi_hi_hi_64, res_hi_hi_hi_lo_64};
  wire [127:0]  res_hi_hi_64 = {res_hi_hi_hi_64, res_hi_hi_lo_64};
  wire [255:0]  res_hi_64 = {res_hi_hi_64, res_hi_lo_64};
  wire [511:0]  res_120 = {res_hi_64, res_lo_64};
  wire [2047:0] dataGroup_lo_3232 = {dataGroup_lo_hi_3232, dataGroup_lo_lo_3232};
  wire [2047:0] dataGroup_hi_3232 = {dataGroup_hi_hi_3232, dataGroup_hi_lo_3232};
  wire [15:0]   dataGroup_0_65 = dataGroup_lo_3232[31:16];
  wire [2047:0] dataGroup_lo_3233 = {dataGroup_lo_hi_3233, dataGroup_lo_lo_3233};
  wire [2047:0] dataGroup_hi_3233 = {dataGroup_hi_hi_3233, dataGroup_hi_lo_3233};
  wire [15:0]   dataGroup_1_65 = dataGroup_lo_3233[159:144];
  wire [2047:0] dataGroup_lo_3234 = {dataGroup_lo_hi_3234, dataGroup_lo_lo_3234};
  wire [2047:0] dataGroup_hi_3234 = {dataGroup_hi_hi_3234, dataGroup_hi_lo_3234};
  wire [15:0]   dataGroup_2_65 = dataGroup_lo_3234[287:272];
  wire [2047:0] dataGroup_lo_3235 = {dataGroup_lo_hi_3235, dataGroup_lo_lo_3235};
  wire [2047:0] dataGroup_hi_3235 = {dataGroup_hi_hi_3235, dataGroup_hi_lo_3235};
  wire [15:0]   dataGroup_3_65 = dataGroup_lo_3235[415:400];
  wire [2047:0] dataGroup_lo_3236 = {dataGroup_lo_hi_3236, dataGroup_lo_lo_3236};
  wire [2047:0] dataGroup_hi_3236 = {dataGroup_hi_hi_3236, dataGroup_hi_lo_3236};
  wire [15:0]   dataGroup_4_65 = dataGroup_lo_3236[543:528];
  wire [2047:0] dataGroup_lo_3237 = {dataGroup_lo_hi_3237, dataGroup_lo_lo_3237};
  wire [2047:0] dataGroup_hi_3237 = {dataGroup_hi_hi_3237, dataGroup_hi_lo_3237};
  wire [15:0]   dataGroup_5_65 = dataGroup_lo_3237[671:656];
  wire [2047:0] dataGroup_lo_3238 = {dataGroup_lo_hi_3238, dataGroup_lo_lo_3238};
  wire [2047:0] dataGroup_hi_3238 = {dataGroup_hi_hi_3238, dataGroup_hi_lo_3238};
  wire [15:0]   dataGroup_6_65 = dataGroup_lo_3238[799:784];
  wire [2047:0] dataGroup_lo_3239 = {dataGroup_lo_hi_3239, dataGroup_lo_lo_3239};
  wire [2047:0] dataGroup_hi_3239 = {dataGroup_hi_hi_3239, dataGroup_hi_lo_3239};
  wire [15:0]   dataGroup_7_65 = dataGroup_lo_3239[927:912];
  wire [2047:0] dataGroup_lo_3240 = {dataGroup_lo_hi_3240, dataGroup_lo_lo_3240};
  wire [2047:0] dataGroup_hi_3240 = {dataGroup_hi_hi_3240, dataGroup_hi_lo_3240};
  wire [15:0]   dataGroup_8_65 = dataGroup_lo_3240[1055:1040];
  wire [2047:0] dataGroup_lo_3241 = {dataGroup_lo_hi_3241, dataGroup_lo_lo_3241};
  wire [2047:0] dataGroup_hi_3241 = {dataGroup_hi_hi_3241, dataGroup_hi_lo_3241};
  wire [15:0]   dataGroup_9_65 = dataGroup_lo_3241[1183:1168];
  wire [2047:0] dataGroup_lo_3242 = {dataGroup_lo_hi_3242, dataGroup_lo_lo_3242};
  wire [2047:0] dataGroup_hi_3242 = {dataGroup_hi_hi_3242, dataGroup_hi_lo_3242};
  wire [15:0]   dataGroup_10_65 = dataGroup_lo_3242[1311:1296];
  wire [2047:0] dataGroup_lo_3243 = {dataGroup_lo_hi_3243, dataGroup_lo_lo_3243};
  wire [2047:0] dataGroup_hi_3243 = {dataGroup_hi_hi_3243, dataGroup_hi_lo_3243};
  wire [15:0]   dataGroup_11_65 = dataGroup_lo_3243[1439:1424];
  wire [2047:0] dataGroup_lo_3244 = {dataGroup_lo_hi_3244, dataGroup_lo_lo_3244};
  wire [2047:0] dataGroup_hi_3244 = {dataGroup_hi_hi_3244, dataGroup_hi_lo_3244};
  wire [15:0]   dataGroup_12_65 = dataGroup_lo_3244[1567:1552];
  wire [2047:0] dataGroup_lo_3245 = {dataGroup_lo_hi_3245, dataGroup_lo_lo_3245};
  wire [2047:0] dataGroup_hi_3245 = {dataGroup_hi_hi_3245, dataGroup_hi_lo_3245};
  wire [15:0]   dataGroup_13_65 = dataGroup_lo_3245[1695:1680];
  wire [2047:0] dataGroup_lo_3246 = {dataGroup_lo_hi_3246, dataGroup_lo_lo_3246};
  wire [2047:0] dataGroup_hi_3246 = {dataGroup_hi_hi_3246, dataGroup_hi_lo_3246};
  wire [15:0]   dataGroup_14_65 = dataGroup_lo_3246[1823:1808];
  wire [2047:0] dataGroup_lo_3247 = {dataGroup_lo_hi_3247, dataGroup_lo_lo_3247};
  wire [2047:0] dataGroup_hi_3247 = {dataGroup_hi_hi_3247, dataGroup_hi_lo_3247};
  wire [15:0]   dataGroup_15_65 = dataGroup_lo_3247[1951:1936];
  wire [2047:0] dataGroup_lo_3248 = {dataGroup_lo_hi_3248, dataGroup_lo_lo_3248};
  wire [2047:0] dataGroup_hi_3248 = {dataGroup_hi_hi_3248, dataGroup_hi_lo_3248};
  wire [15:0]   dataGroup_16_65 = dataGroup_hi_3248[31:16];
  wire [2047:0] dataGroup_lo_3249 = {dataGroup_lo_hi_3249, dataGroup_lo_lo_3249};
  wire [2047:0] dataGroup_hi_3249 = {dataGroup_hi_hi_3249, dataGroup_hi_lo_3249};
  wire [15:0]   dataGroup_17_65 = dataGroup_hi_3249[159:144];
  wire [2047:0] dataGroup_lo_3250 = {dataGroup_lo_hi_3250, dataGroup_lo_lo_3250};
  wire [2047:0] dataGroup_hi_3250 = {dataGroup_hi_hi_3250, dataGroup_hi_lo_3250};
  wire [15:0]   dataGroup_18_65 = dataGroup_hi_3250[287:272];
  wire [2047:0] dataGroup_lo_3251 = {dataGroup_lo_hi_3251, dataGroup_lo_lo_3251};
  wire [2047:0] dataGroup_hi_3251 = {dataGroup_hi_hi_3251, dataGroup_hi_lo_3251};
  wire [15:0]   dataGroup_19_65 = dataGroup_hi_3251[415:400];
  wire [2047:0] dataGroup_lo_3252 = {dataGroup_lo_hi_3252, dataGroup_lo_lo_3252};
  wire [2047:0] dataGroup_hi_3252 = {dataGroup_hi_hi_3252, dataGroup_hi_lo_3252};
  wire [15:0]   dataGroup_20_65 = dataGroup_hi_3252[543:528];
  wire [2047:0] dataGroup_lo_3253 = {dataGroup_lo_hi_3253, dataGroup_lo_lo_3253};
  wire [2047:0] dataGroup_hi_3253 = {dataGroup_hi_hi_3253, dataGroup_hi_lo_3253};
  wire [15:0]   dataGroup_21_65 = dataGroup_hi_3253[671:656];
  wire [2047:0] dataGroup_lo_3254 = {dataGroup_lo_hi_3254, dataGroup_lo_lo_3254};
  wire [2047:0] dataGroup_hi_3254 = {dataGroup_hi_hi_3254, dataGroup_hi_lo_3254};
  wire [15:0]   dataGroup_22_65 = dataGroup_hi_3254[799:784];
  wire [2047:0] dataGroup_lo_3255 = {dataGroup_lo_hi_3255, dataGroup_lo_lo_3255};
  wire [2047:0] dataGroup_hi_3255 = {dataGroup_hi_hi_3255, dataGroup_hi_lo_3255};
  wire [15:0]   dataGroup_23_65 = dataGroup_hi_3255[927:912];
  wire [2047:0] dataGroup_lo_3256 = {dataGroup_lo_hi_3256, dataGroup_lo_lo_3256};
  wire [2047:0] dataGroup_hi_3256 = {dataGroup_hi_hi_3256, dataGroup_hi_lo_3256};
  wire [15:0]   dataGroup_24_65 = dataGroup_hi_3256[1055:1040];
  wire [2047:0] dataGroup_lo_3257 = {dataGroup_lo_hi_3257, dataGroup_lo_lo_3257};
  wire [2047:0] dataGroup_hi_3257 = {dataGroup_hi_hi_3257, dataGroup_hi_lo_3257};
  wire [15:0]   dataGroup_25_65 = dataGroup_hi_3257[1183:1168];
  wire [2047:0] dataGroup_lo_3258 = {dataGroup_lo_hi_3258, dataGroup_lo_lo_3258};
  wire [2047:0] dataGroup_hi_3258 = {dataGroup_hi_hi_3258, dataGroup_hi_lo_3258};
  wire [15:0]   dataGroup_26_65 = dataGroup_hi_3258[1311:1296];
  wire [2047:0] dataGroup_lo_3259 = {dataGroup_lo_hi_3259, dataGroup_lo_lo_3259};
  wire [2047:0] dataGroup_hi_3259 = {dataGroup_hi_hi_3259, dataGroup_hi_lo_3259};
  wire [15:0]   dataGroup_27_65 = dataGroup_hi_3259[1439:1424];
  wire [2047:0] dataGroup_lo_3260 = {dataGroup_lo_hi_3260, dataGroup_lo_lo_3260};
  wire [2047:0] dataGroup_hi_3260 = {dataGroup_hi_hi_3260, dataGroup_hi_lo_3260};
  wire [15:0]   dataGroup_28_65 = dataGroup_hi_3260[1567:1552];
  wire [2047:0] dataGroup_lo_3261 = {dataGroup_lo_hi_3261, dataGroup_lo_lo_3261};
  wire [2047:0] dataGroup_hi_3261 = {dataGroup_hi_hi_3261, dataGroup_hi_lo_3261};
  wire [15:0]   dataGroup_29_65 = dataGroup_hi_3261[1695:1680];
  wire [2047:0] dataGroup_lo_3262 = {dataGroup_lo_hi_3262, dataGroup_lo_lo_3262};
  wire [2047:0] dataGroup_hi_3262 = {dataGroup_hi_hi_3262, dataGroup_hi_lo_3262};
  wire [15:0]   dataGroup_30_65 = dataGroup_hi_3262[1823:1808];
  wire [2047:0] dataGroup_lo_3263 = {dataGroup_lo_hi_3263, dataGroup_lo_lo_3263};
  wire [2047:0] dataGroup_hi_3263 = {dataGroup_hi_hi_3263, dataGroup_hi_lo_3263};
  wire [15:0]   dataGroup_31_65 = dataGroup_hi_3263[1951:1936];
  wire [31:0]   res_lo_lo_lo_lo_65 = {dataGroup_1_65, dataGroup_0_65};
  wire [31:0]   res_lo_lo_lo_hi_65 = {dataGroup_3_65, dataGroup_2_65};
  wire [63:0]   res_lo_lo_lo_65 = {res_lo_lo_lo_hi_65, res_lo_lo_lo_lo_65};
  wire [31:0]   res_lo_lo_hi_lo_65 = {dataGroup_5_65, dataGroup_4_65};
  wire [31:0]   res_lo_lo_hi_hi_65 = {dataGroup_7_65, dataGroup_6_65};
  wire [63:0]   res_lo_lo_hi_65 = {res_lo_lo_hi_hi_65, res_lo_lo_hi_lo_65};
  wire [127:0]  res_lo_lo_65 = {res_lo_lo_hi_65, res_lo_lo_lo_65};
  wire [31:0]   res_lo_hi_lo_lo_65 = {dataGroup_9_65, dataGroup_8_65};
  wire [31:0]   res_lo_hi_lo_hi_65 = {dataGroup_11_65, dataGroup_10_65};
  wire [63:0]   res_lo_hi_lo_65 = {res_lo_hi_lo_hi_65, res_lo_hi_lo_lo_65};
  wire [31:0]   res_lo_hi_hi_lo_65 = {dataGroup_13_65, dataGroup_12_65};
  wire [31:0]   res_lo_hi_hi_hi_65 = {dataGroup_15_65, dataGroup_14_65};
  wire [63:0]   res_lo_hi_hi_65 = {res_lo_hi_hi_hi_65, res_lo_hi_hi_lo_65};
  wire [127:0]  res_lo_hi_65 = {res_lo_hi_hi_65, res_lo_hi_lo_65};
  wire [255:0]  res_lo_65 = {res_lo_hi_65, res_lo_lo_65};
  wire [31:0]   res_hi_lo_lo_lo_65 = {dataGroup_17_65, dataGroup_16_65};
  wire [31:0]   res_hi_lo_lo_hi_65 = {dataGroup_19_65, dataGroup_18_65};
  wire [63:0]   res_hi_lo_lo_65 = {res_hi_lo_lo_hi_65, res_hi_lo_lo_lo_65};
  wire [31:0]   res_hi_lo_hi_lo_65 = {dataGroup_21_65, dataGroup_20_65};
  wire [31:0]   res_hi_lo_hi_hi_65 = {dataGroup_23_65, dataGroup_22_65};
  wire [63:0]   res_hi_lo_hi_65 = {res_hi_lo_hi_hi_65, res_hi_lo_hi_lo_65};
  wire [127:0]  res_hi_lo_65 = {res_hi_lo_hi_65, res_hi_lo_lo_65};
  wire [31:0]   res_hi_hi_lo_lo_65 = {dataGroup_25_65, dataGroup_24_65};
  wire [31:0]   res_hi_hi_lo_hi_65 = {dataGroup_27_65, dataGroup_26_65};
  wire [63:0]   res_hi_hi_lo_65 = {res_hi_hi_lo_hi_65, res_hi_hi_lo_lo_65};
  wire [31:0]   res_hi_hi_hi_lo_65 = {dataGroup_29_65, dataGroup_28_65};
  wire [31:0]   res_hi_hi_hi_hi_65 = {dataGroup_31_65, dataGroup_30_65};
  wire [63:0]   res_hi_hi_hi_65 = {res_hi_hi_hi_hi_65, res_hi_hi_hi_lo_65};
  wire [127:0]  res_hi_hi_65 = {res_hi_hi_hi_65, res_hi_hi_lo_65};
  wire [255:0]  res_hi_65 = {res_hi_hi_65, res_hi_lo_65};
  wire [511:0]  res_121 = {res_hi_65, res_lo_65};
  wire [2047:0] dataGroup_lo_3264 = {dataGroup_lo_hi_3264, dataGroup_lo_lo_3264};
  wire [2047:0] dataGroup_hi_3264 = {dataGroup_hi_hi_3264, dataGroup_hi_lo_3264};
  wire [15:0]   dataGroup_0_66 = dataGroup_lo_3264[47:32];
  wire [2047:0] dataGroup_lo_3265 = {dataGroup_lo_hi_3265, dataGroup_lo_lo_3265};
  wire [2047:0] dataGroup_hi_3265 = {dataGroup_hi_hi_3265, dataGroup_hi_lo_3265};
  wire [15:0]   dataGroup_1_66 = dataGroup_lo_3265[175:160];
  wire [2047:0] dataGroup_lo_3266 = {dataGroup_lo_hi_3266, dataGroup_lo_lo_3266};
  wire [2047:0] dataGroup_hi_3266 = {dataGroup_hi_hi_3266, dataGroup_hi_lo_3266};
  wire [15:0]   dataGroup_2_66 = dataGroup_lo_3266[303:288];
  wire [2047:0] dataGroup_lo_3267 = {dataGroup_lo_hi_3267, dataGroup_lo_lo_3267};
  wire [2047:0] dataGroup_hi_3267 = {dataGroup_hi_hi_3267, dataGroup_hi_lo_3267};
  wire [15:0]   dataGroup_3_66 = dataGroup_lo_3267[431:416];
  wire [2047:0] dataGroup_lo_3268 = {dataGroup_lo_hi_3268, dataGroup_lo_lo_3268};
  wire [2047:0] dataGroup_hi_3268 = {dataGroup_hi_hi_3268, dataGroup_hi_lo_3268};
  wire [15:0]   dataGroup_4_66 = dataGroup_lo_3268[559:544];
  wire [2047:0] dataGroup_lo_3269 = {dataGroup_lo_hi_3269, dataGroup_lo_lo_3269};
  wire [2047:0] dataGroup_hi_3269 = {dataGroup_hi_hi_3269, dataGroup_hi_lo_3269};
  wire [15:0]   dataGroup_5_66 = dataGroup_lo_3269[687:672];
  wire [2047:0] dataGroup_lo_3270 = {dataGroup_lo_hi_3270, dataGroup_lo_lo_3270};
  wire [2047:0] dataGroup_hi_3270 = {dataGroup_hi_hi_3270, dataGroup_hi_lo_3270};
  wire [15:0]   dataGroup_6_66 = dataGroup_lo_3270[815:800];
  wire [2047:0] dataGroup_lo_3271 = {dataGroup_lo_hi_3271, dataGroup_lo_lo_3271};
  wire [2047:0] dataGroup_hi_3271 = {dataGroup_hi_hi_3271, dataGroup_hi_lo_3271};
  wire [15:0]   dataGroup_7_66 = dataGroup_lo_3271[943:928];
  wire [2047:0] dataGroup_lo_3272 = {dataGroup_lo_hi_3272, dataGroup_lo_lo_3272};
  wire [2047:0] dataGroup_hi_3272 = {dataGroup_hi_hi_3272, dataGroup_hi_lo_3272};
  wire [15:0]   dataGroup_8_66 = dataGroup_lo_3272[1071:1056];
  wire [2047:0] dataGroup_lo_3273 = {dataGroup_lo_hi_3273, dataGroup_lo_lo_3273};
  wire [2047:0] dataGroup_hi_3273 = {dataGroup_hi_hi_3273, dataGroup_hi_lo_3273};
  wire [15:0]   dataGroup_9_66 = dataGroup_lo_3273[1199:1184];
  wire [2047:0] dataGroup_lo_3274 = {dataGroup_lo_hi_3274, dataGroup_lo_lo_3274};
  wire [2047:0] dataGroup_hi_3274 = {dataGroup_hi_hi_3274, dataGroup_hi_lo_3274};
  wire [15:0]   dataGroup_10_66 = dataGroup_lo_3274[1327:1312];
  wire [2047:0] dataGroup_lo_3275 = {dataGroup_lo_hi_3275, dataGroup_lo_lo_3275};
  wire [2047:0] dataGroup_hi_3275 = {dataGroup_hi_hi_3275, dataGroup_hi_lo_3275};
  wire [15:0]   dataGroup_11_66 = dataGroup_lo_3275[1455:1440];
  wire [2047:0] dataGroup_lo_3276 = {dataGroup_lo_hi_3276, dataGroup_lo_lo_3276};
  wire [2047:0] dataGroup_hi_3276 = {dataGroup_hi_hi_3276, dataGroup_hi_lo_3276};
  wire [15:0]   dataGroup_12_66 = dataGroup_lo_3276[1583:1568];
  wire [2047:0] dataGroup_lo_3277 = {dataGroup_lo_hi_3277, dataGroup_lo_lo_3277};
  wire [2047:0] dataGroup_hi_3277 = {dataGroup_hi_hi_3277, dataGroup_hi_lo_3277};
  wire [15:0]   dataGroup_13_66 = dataGroup_lo_3277[1711:1696];
  wire [2047:0] dataGroup_lo_3278 = {dataGroup_lo_hi_3278, dataGroup_lo_lo_3278};
  wire [2047:0] dataGroup_hi_3278 = {dataGroup_hi_hi_3278, dataGroup_hi_lo_3278};
  wire [15:0]   dataGroup_14_66 = dataGroup_lo_3278[1839:1824];
  wire [2047:0] dataGroup_lo_3279 = {dataGroup_lo_hi_3279, dataGroup_lo_lo_3279};
  wire [2047:0] dataGroup_hi_3279 = {dataGroup_hi_hi_3279, dataGroup_hi_lo_3279};
  wire [15:0]   dataGroup_15_66 = dataGroup_lo_3279[1967:1952];
  wire [2047:0] dataGroup_lo_3280 = {dataGroup_lo_hi_3280, dataGroup_lo_lo_3280};
  wire [2047:0] dataGroup_hi_3280 = {dataGroup_hi_hi_3280, dataGroup_hi_lo_3280};
  wire [15:0]   dataGroup_16_66 = dataGroup_hi_3280[47:32];
  wire [2047:0] dataGroup_lo_3281 = {dataGroup_lo_hi_3281, dataGroup_lo_lo_3281};
  wire [2047:0] dataGroup_hi_3281 = {dataGroup_hi_hi_3281, dataGroup_hi_lo_3281};
  wire [15:0]   dataGroup_17_66 = dataGroup_hi_3281[175:160];
  wire [2047:0] dataGroup_lo_3282 = {dataGroup_lo_hi_3282, dataGroup_lo_lo_3282};
  wire [2047:0] dataGroup_hi_3282 = {dataGroup_hi_hi_3282, dataGroup_hi_lo_3282};
  wire [15:0]   dataGroup_18_66 = dataGroup_hi_3282[303:288];
  wire [2047:0] dataGroup_lo_3283 = {dataGroup_lo_hi_3283, dataGroup_lo_lo_3283};
  wire [2047:0] dataGroup_hi_3283 = {dataGroup_hi_hi_3283, dataGroup_hi_lo_3283};
  wire [15:0]   dataGroup_19_66 = dataGroup_hi_3283[431:416];
  wire [2047:0] dataGroup_lo_3284 = {dataGroup_lo_hi_3284, dataGroup_lo_lo_3284};
  wire [2047:0] dataGroup_hi_3284 = {dataGroup_hi_hi_3284, dataGroup_hi_lo_3284};
  wire [15:0]   dataGroup_20_66 = dataGroup_hi_3284[559:544];
  wire [2047:0] dataGroup_lo_3285 = {dataGroup_lo_hi_3285, dataGroup_lo_lo_3285};
  wire [2047:0] dataGroup_hi_3285 = {dataGroup_hi_hi_3285, dataGroup_hi_lo_3285};
  wire [15:0]   dataGroup_21_66 = dataGroup_hi_3285[687:672];
  wire [2047:0] dataGroup_lo_3286 = {dataGroup_lo_hi_3286, dataGroup_lo_lo_3286};
  wire [2047:0] dataGroup_hi_3286 = {dataGroup_hi_hi_3286, dataGroup_hi_lo_3286};
  wire [15:0]   dataGroup_22_66 = dataGroup_hi_3286[815:800];
  wire [2047:0] dataGroup_lo_3287 = {dataGroup_lo_hi_3287, dataGroup_lo_lo_3287};
  wire [2047:0] dataGroup_hi_3287 = {dataGroup_hi_hi_3287, dataGroup_hi_lo_3287};
  wire [15:0]   dataGroup_23_66 = dataGroup_hi_3287[943:928];
  wire [2047:0] dataGroup_lo_3288 = {dataGroup_lo_hi_3288, dataGroup_lo_lo_3288};
  wire [2047:0] dataGroup_hi_3288 = {dataGroup_hi_hi_3288, dataGroup_hi_lo_3288};
  wire [15:0]   dataGroup_24_66 = dataGroup_hi_3288[1071:1056];
  wire [2047:0] dataGroup_lo_3289 = {dataGroup_lo_hi_3289, dataGroup_lo_lo_3289};
  wire [2047:0] dataGroup_hi_3289 = {dataGroup_hi_hi_3289, dataGroup_hi_lo_3289};
  wire [15:0]   dataGroup_25_66 = dataGroup_hi_3289[1199:1184];
  wire [2047:0] dataGroup_lo_3290 = {dataGroup_lo_hi_3290, dataGroup_lo_lo_3290};
  wire [2047:0] dataGroup_hi_3290 = {dataGroup_hi_hi_3290, dataGroup_hi_lo_3290};
  wire [15:0]   dataGroup_26_66 = dataGroup_hi_3290[1327:1312];
  wire [2047:0] dataGroup_lo_3291 = {dataGroup_lo_hi_3291, dataGroup_lo_lo_3291};
  wire [2047:0] dataGroup_hi_3291 = {dataGroup_hi_hi_3291, dataGroup_hi_lo_3291};
  wire [15:0]   dataGroup_27_66 = dataGroup_hi_3291[1455:1440];
  wire [2047:0] dataGroup_lo_3292 = {dataGroup_lo_hi_3292, dataGroup_lo_lo_3292};
  wire [2047:0] dataGroup_hi_3292 = {dataGroup_hi_hi_3292, dataGroup_hi_lo_3292};
  wire [15:0]   dataGroup_28_66 = dataGroup_hi_3292[1583:1568];
  wire [2047:0] dataGroup_lo_3293 = {dataGroup_lo_hi_3293, dataGroup_lo_lo_3293};
  wire [2047:0] dataGroup_hi_3293 = {dataGroup_hi_hi_3293, dataGroup_hi_lo_3293};
  wire [15:0]   dataGroup_29_66 = dataGroup_hi_3293[1711:1696];
  wire [2047:0] dataGroup_lo_3294 = {dataGroup_lo_hi_3294, dataGroup_lo_lo_3294};
  wire [2047:0] dataGroup_hi_3294 = {dataGroup_hi_hi_3294, dataGroup_hi_lo_3294};
  wire [15:0]   dataGroup_30_66 = dataGroup_hi_3294[1839:1824];
  wire [2047:0] dataGroup_lo_3295 = {dataGroup_lo_hi_3295, dataGroup_lo_lo_3295};
  wire [2047:0] dataGroup_hi_3295 = {dataGroup_hi_hi_3295, dataGroup_hi_lo_3295};
  wire [15:0]   dataGroup_31_66 = dataGroup_hi_3295[1967:1952];
  wire [31:0]   res_lo_lo_lo_lo_66 = {dataGroup_1_66, dataGroup_0_66};
  wire [31:0]   res_lo_lo_lo_hi_66 = {dataGroup_3_66, dataGroup_2_66};
  wire [63:0]   res_lo_lo_lo_66 = {res_lo_lo_lo_hi_66, res_lo_lo_lo_lo_66};
  wire [31:0]   res_lo_lo_hi_lo_66 = {dataGroup_5_66, dataGroup_4_66};
  wire [31:0]   res_lo_lo_hi_hi_66 = {dataGroup_7_66, dataGroup_6_66};
  wire [63:0]   res_lo_lo_hi_66 = {res_lo_lo_hi_hi_66, res_lo_lo_hi_lo_66};
  wire [127:0]  res_lo_lo_66 = {res_lo_lo_hi_66, res_lo_lo_lo_66};
  wire [31:0]   res_lo_hi_lo_lo_66 = {dataGroup_9_66, dataGroup_8_66};
  wire [31:0]   res_lo_hi_lo_hi_66 = {dataGroup_11_66, dataGroup_10_66};
  wire [63:0]   res_lo_hi_lo_66 = {res_lo_hi_lo_hi_66, res_lo_hi_lo_lo_66};
  wire [31:0]   res_lo_hi_hi_lo_66 = {dataGroup_13_66, dataGroup_12_66};
  wire [31:0]   res_lo_hi_hi_hi_66 = {dataGroup_15_66, dataGroup_14_66};
  wire [63:0]   res_lo_hi_hi_66 = {res_lo_hi_hi_hi_66, res_lo_hi_hi_lo_66};
  wire [127:0]  res_lo_hi_66 = {res_lo_hi_hi_66, res_lo_hi_lo_66};
  wire [255:0]  res_lo_66 = {res_lo_hi_66, res_lo_lo_66};
  wire [31:0]   res_hi_lo_lo_lo_66 = {dataGroup_17_66, dataGroup_16_66};
  wire [31:0]   res_hi_lo_lo_hi_66 = {dataGroup_19_66, dataGroup_18_66};
  wire [63:0]   res_hi_lo_lo_66 = {res_hi_lo_lo_hi_66, res_hi_lo_lo_lo_66};
  wire [31:0]   res_hi_lo_hi_lo_66 = {dataGroup_21_66, dataGroup_20_66};
  wire [31:0]   res_hi_lo_hi_hi_66 = {dataGroup_23_66, dataGroup_22_66};
  wire [63:0]   res_hi_lo_hi_66 = {res_hi_lo_hi_hi_66, res_hi_lo_hi_lo_66};
  wire [127:0]  res_hi_lo_66 = {res_hi_lo_hi_66, res_hi_lo_lo_66};
  wire [31:0]   res_hi_hi_lo_lo_66 = {dataGroup_25_66, dataGroup_24_66};
  wire [31:0]   res_hi_hi_lo_hi_66 = {dataGroup_27_66, dataGroup_26_66};
  wire [63:0]   res_hi_hi_lo_66 = {res_hi_hi_lo_hi_66, res_hi_hi_lo_lo_66};
  wire [31:0]   res_hi_hi_hi_lo_66 = {dataGroup_29_66, dataGroup_28_66};
  wire [31:0]   res_hi_hi_hi_hi_66 = {dataGroup_31_66, dataGroup_30_66};
  wire [63:0]   res_hi_hi_hi_66 = {res_hi_hi_hi_hi_66, res_hi_hi_hi_lo_66};
  wire [127:0]  res_hi_hi_66 = {res_hi_hi_hi_66, res_hi_hi_lo_66};
  wire [255:0]  res_hi_66 = {res_hi_hi_66, res_hi_lo_66};
  wire [511:0]  res_122 = {res_hi_66, res_lo_66};
  wire [2047:0] dataGroup_lo_3296 = {dataGroup_lo_hi_3296, dataGroup_lo_lo_3296};
  wire [2047:0] dataGroup_hi_3296 = {dataGroup_hi_hi_3296, dataGroup_hi_lo_3296};
  wire [15:0]   dataGroup_0_67 = dataGroup_lo_3296[63:48];
  wire [2047:0] dataGroup_lo_3297 = {dataGroup_lo_hi_3297, dataGroup_lo_lo_3297};
  wire [2047:0] dataGroup_hi_3297 = {dataGroup_hi_hi_3297, dataGroup_hi_lo_3297};
  wire [15:0]   dataGroup_1_67 = dataGroup_lo_3297[191:176];
  wire [2047:0] dataGroup_lo_3298 = {dataGroup_lo_hi_3298, dataGroup_lo_lo_3298};
  wire [2047:0] dataGroup_hi_3298 = {dataGroup_hi_hi_3298, dataGroup_hi_lo_3298};
  wire [15:0]   dataGroup_2_67 = dataGroup_lo_3298[319:304];
  wire [2047:0] dataGroup_lo_3299 = {dataGroup_lo_hi_3299, dataGroup_lo_lo_3299};
  wire [2047:0] dataGroup_hi_3299 = {dataGroup_hi_hi_3299, dataGroup_hi_lo_3299};
  wire [15:0]   dataGroup_3_67 = dataGroup_lo_3299[447:432];
  wire [2047:0] dataGroup_lo_3300 = {dataGroup_lo_hi_3300, dataGroup_lo_lo_3300};
  wire [2047:0] dataGroup_hi_3300 = {dataGroup_hi_hi_3300, dataGroup_hi_lo_3300};
  wire [15:0]   dataGroup_4_67 = dataGroup_lo_3300[575:560];
  wire [2047:0] dataGroup_lo_3301 = {dataGroup_lo_hi_3301, dataGroup_lo_lo_3301};
  wire [2047:0] dataGroup_hi_3301 = {dataGroup_hi_hi_3301, dataGroup_hi_lo_3301};
  wire [15:0]   dataGroup_5_67 = dataGroup_lo_3301[703:688];
  wire [2047:0] dataGroup_lo_3302 = {dataGroup_lo_hi_3302, dataGroup_lo_lo_3302};
  wire [2047:0] dataGroup_hi_3302 = {dataGroup_hi_hi_3302, dataGroup_hi_lo_3302};
  wire [15:0]   dataGroup_6_67 = dataGroup_lo_3302[831:816];
  wire [2047:0] dataGroup_lo_3303 = {dataGroup_lo_hi_3303, dataGroup_lo_lo_3303};
  wire [2047:0] dataGroup_hi_3303 = {dataGroup_hi_hi_3303, dataGroup_hi_lo_3303};
  wire [15:0]   dataGroup_7_67 = dataGroup_lo_3303[959:944];
  wire [2047:0] dataGroup_lo_3304 = {dataGroup_lo_hi_3304, dataGroup_lo_lo_3304};
  wire [2047:0] dataGroup_hi_3304 = {dataGroup_hi_hi_3304, dataGroup_hi_lo_3304};
  wire [15:0]   dataGroup_8_67 = dataGroup_lo_3304[1087:1072];
  wire [2047:0] dataGroup_lo_3305 = {dataGroup_lo_hi_3305, dataGroup_lo_lo_3305};
  wire [2047:0] dataGroup_hi_3305 = {dataGroup_hi_hi_3305, dataGroup_hi_lo_3305};
  wire [15:0]   dataGroup_9_67 = dataGroup_lo_3305[1215:1200];
  wire [2047:0] dataGroup_lo_3306 = {dataGroup_lo_hi_3306, dataGroup_lo_lo_3306};
  wire [2047:0] dataGroup_hi_3306 = {dataGroup_hi_hi_3306, dataGroup_hi_lo_3306};
  wire [15:0]   dataGroup_10_67 = dataGroup_lo_3306[1343:1328];
  wire [2047:0] dataGroup_lo_3307 = {dataGroup_lo_hi_3307, dataGroup_lo_lo_3307};
  wire [2047:0] dataGroup_hi_3307 = {dataGroup_hi_hi_3307, dataGroup_hi_lo_3307};
  wire [15:0]   dataGroup_11_67 = dataGroup_lo_3307[1471:1456];
  wire [2047:0] dataGroup_lo_3308 = {dataGroup_lo_hi_3308, dataGroup_lo_lo_3308};
  wire [2047:0] dataGroup_hi_3308 = {dataGroup_hi_hi_3308, dataGroup_hi_lo_3308};
  wire [15:0]   dataGroup_12_67 = dataGroup_lo_3308[1599:1584];
  wire [2047:0] dataGroup_lo_3309 = {dataGroup_lo_hi_3309, dataGroup_lo_lo_3309};
  wire [2047:0] dataGroup_hi_3309 = {dataGroup_hi_hi_3309, dataGroup_hi_lo_3309};
  wire [15:0]   dataGroup_13_67 = dataGroup_lo_3309[1727:1712];
  wire [2047:0] dataGroup_lo_3310 = {dataGroup_lo_hi_3310, dataGroup_lo_lo_3310};
  wire [2047:0] dataGroup_hi_3310 = {dataGroup_hi_hi_3310, dataGroup_hi_lo_3310};
  wire [15:0]   dataGroup_14_67 = dataGroup_lo_3310[1855:1840];
  wire [2047:0] dataGroup_lo_3311 = {dataGroup_lo_hi_3311, dataGroup_lo_lo_3311};
  wire [2047:0] dataGroup_hi_3311 = {dataGroup_hi_hi_3311, dataGroup_hi_lo_3311};
  wire [15:0]   dataGroup_15_67 = dataGroup_lo_3311[1983:1968];
  wire [2047:0] dataGroup_lo_3312 = {dataGroup_lo_hi_3312, dataGroup_lo_lo_3312};
  wire [2047:0] dataGroup_hi_3312 = {dataGroup_hi_hi_3312, dataGroup_hi_lo_3312};
  wire [15:0]   dataGroup_16_67 = dataGroup_hi_3312[63:48];
  wire [2047:0] dataGroup_lo_3313 = {dataGroup_lo_hi_3313, dataGroup_lo_lo_3313};
  wire [2047:0] dataGroup_hi_3313 = {dataGroup_hi_hi_3313, dataGroup_hi_lo_3313};
  wire [15:0]   dataGroup_17_67 = dataGroup_hi_3313[191:176];
  wire [2047:0] dataGroup_lo_3314 = {dataGroup_lo_hi_3314, dataGroup_lo_lo_3314};
  wire [2047:0] dataGroup_hi_3314 = {dataGroup_hi_hi_3314, dataGroup_hi_lo_3314};
  wire [15:0]   dataGroup_18_67 = dataGroup_hi_3314[319:304];
  wire [2047:0] dataGroup_lo_3315 = {dataGroup_lo_hi_3315, dataGroup_lo_lo_3315};
  wire [2047:0] dataGroup_hi_3315 = {dataGroup_hi_hi_3315, dataGroup_hi_lo_3315};
  wire [15:0]   dataGroup_19_67 = dataGroup_hi_3315[447:432];
  wire [2047:0] dataGroup_lo_3316 = {dataGroup_lo_hi_3316, dataGroup_lo_lo_3316};
  wire [2047:0] dataGroup_hi_3316 = {dataGroup_hi_hi_3316, dataGroup_hi_lo_3316};
  wire [15:0]   dataGroup_20_67 = dataGroup_hi_3316[575:560];
  wire [2047:0] dataGroup_lo_3317 = {dataGroup_lo_hi_3317, dataGroup_lo_lo_3317};
  wire [2047:0] dataGroup_hi_3317 = {dataGroup_hi_hi_3317, dataGroup_hi_lo_3317};
  wire [15:0]   dataGroup_21_67 = dataGroup_hi_3317[703:688];
  wire [2047:0] dataGroup_lo_3318 = {dataGroup_lo_hi_3318, dataGroup_lo_lo_3318};
  wire [2047:0] dataGroup_hi_3318 = {dataGroup_hi_hi_3318, dataGroup_hi_lo_3318};
  wire [15:0]   dataGroup_22_67 = dataGroup_hi_3318[831:816];
  wire [2047:0] dataGroup_lo_3319 = {dataGroup_lo_hi_3319, dataGroup_lo_lo_3319};
  wire [2047:0] dataGroup_hi_3319 = {dataGroup_hi_hi_3319, dataGroup_hi_lo_3319};
  wire [15:0]   dataGroup_23_67 = dataGroup_hi_3319[959:944];
  wire [2047:0] dataGroup_lo_3320 = {dataGroup_lo_hi_3320, dataGroup_lo_lo_3320};
  wire [2047:0] dataGroup_hi_3320 = {dataGroup_hi_hi_3320, dataGroup_hi_lo_3320};
  wire [15:0]   dataGroup_24_67 = dataGroup_hi_3320[1087:1072];
  wire [2047:0] dataGroup_lo_3321 = {dataGroup_lo_hi_3321, dataGroup_lo_lo_3321};
  wire [2047:0] dataGroup_hi_3321 = {dataGroup_hi_hi_3321, dataGroup_hi_lo_3321};
  wire [15:0]   dataGroup_25_67 = dataGroup_hi_3321[1215:1200];
  wire [2047:0] dataGroup_lo_3322 = {dataGroup_lo_hi_3322, dataGroup_lo_lo_3322};
  wire [2047:0] dataGroup_hi_3322 = {dataGroup_hi_hi_3322, dataGroup_hi_lo_3322};
  wire [15:0]   dataGroup_26_67 = dataGroup_hi_3322[1343:1328];
  wire [2047:0] dataGroup_lo_3323 = {dataGroup_lo_hi_3323, dataGroup_lo_lo_3323};
  wire [2047:0] dataGroup_hi_3323 = {dataGroup_hi_hi_3323, dataGroup_hi_lo_3323};
  wire [15:0]   dataGroup_27_67 = dataGroup_hi_3323[1471:1456];
  wire [2047:0] dataGroup_lo_3324 = {dataGroup_lo_hi_3324, dataGroup_lo_lo_3324};
  wire [2047:0] dataGroup_hi_3324 = {dataGroup_hi_hi_3324, dataGroup_hi_lo_3324};
  wire [15:0]   dataGroup_28_67 = dataGroup_hi_3324[1599:1584];
  wire [2047:0] dataGroup_lo_3325 = {dataGroup_lo_hi_3325, dataGroup_lo_lo_3325};
  wire [2047:0] dataGroup_hi_3325 = {dataGroup_hi_hi_3325, dataGroup_hi_lo_3325};
  wire [15:0]   dataGroup_29_67 = dataGroup_hi_3325[1727:1712];
  wire [2047:0] dataGroup_lo_3326 = {dataGroup_lo_hi_3326, dataGroup_lo_lo_3326};
  wire [2047:0] dataGroup_hi_3326 = {dataGroup_hi_hi_3326, dataGroup_hi_lo_3326};
  wire [15:0]   dataGroup_30_67 = dataGroup_hi_3326[1855:1840];
  wire [2047:0] dataGroup_lo_3327 = {dataGroup_lo_hi_3327, dataGroup_lo_lo_3327};
  wire [2047:0] dataGroup_hi_3327 = {dataGroup_hi_hi_3327, dataGroup_hi_lo_3327};
  wire [15:0]   dataGroup_31_67 = dataGroup_hi_3327[1983:1968];
  wire [31:0]   res_lo_lo_lo_lo_67 = {dataGroup_1_67, dataGroup_0_67};
  wire [31:0]   res_lo_lo_lo_hi_67 = {dataGroup_3_67, dataGroup_2_67};
  wire [63:0]   res_lo_lo_lo_67 = {res_lo_lo_lo_hi_67, res_lo_lo_lo_lo_67};
  wire [31:0]   res_lo_lo_hi_lo_67 = {dataGroup_5_67, dataGroup_4_67};
  wire [31:0]   res_lo_lo_hi_hi_67 = {dataGroup_7_67, dataGroup_6_67};
  wire [63:0]   res_lo_lo_hi_67 = {res_lo_lo_hi_hi_67, res_lo_lo_hi_lo_67};
  wire [127:0]  res_lo_lo_67 = {res_lo_lo_hi_67, res_lo_lo_lo_67};
  wire [31:0]   res_lo_hi_lo_lo_67 = {dataGroup_9_67, dataGroup_8_67};
  wire [31:0]   res_lo_hi_lo_hi_67 = {dataGroup_11_67, dataGroup_10_67};
  wire [63:0]   res_lo_hi_lo_67 = {res_lo_hi_lo_hi_67, res_lo_hi_lo_lo_67};
  wire [31:0]   res_lo_hi_hi_lo_67 = {dataGroup_13_67, dataGroup_12_67};
  wire [31:0]   res_lo_hi_hi_hi_67 = {dataGroup_15_67, dataGroup_14_67};
  wire [63:0]   res_lo_hi_hi_67 = {res_lo_hi_hi_hi_67, res_lo_hi_hi_lo_67};
  wire [127:0]  res_lo_hi_67 = {res_lo_hi_hi_67, res_lo_hi_lo_67};
  wire [255:0]  res_lo_67 = {res_lo_hi_67, res_lo_lo_67};
  wire [31:0]   res_hi_lo_lo_lo_67 = {dataGroup_17_67, dataGroup_16_67};
  wire [31:0]   res_hi_lo_lo_hi_67 = {dataGroup_19_67, dataGroup_18_67};
  wire [63:0]   res_hi_lo_lo_67 = {res_hi_lo_lo_hi_67, res_hi_lo_lo_lo_67};
  wire [31:0]   res_hi_lo_hi_lo_67 = {dataGroup_21_67, dataGroup_20_67};
  wire [31:0]   res_hi_lo_hi_hi_67 = {dataGroup_23_67, dataGroup_22_67};
  wire [63:0]   res_hi_lo_hi_67 = {res_hi_lo_hi_hi_67, res_hi_lo_hi_lo_67};
  wire [127:0]  res_hi_lo_67 = {res_hi_lo_hi_67, res_hi_lo_lo_67};
  wire [31:0]   res_hi_hi_lo_lo_67 = {dataGroup_25_67, dataGroup_24_67};
  wire [31:0]   res_hi_hi_lo_hi_67 = {dataGroup_27_67, dataGroup_26_67};
  wire [63:0]   res_hi_hi_lo_67 = {res_hi_hi_lo_hi_67, res_hi_hi_lo_lo_67};
  wire [31:0]   res_hi_hi_hi_lo_67 = {dataGroup_29_67, dataGroup_28_67};
  wire [31:0]   res_hi_hi_hi_hi_67 = {dataGroup_31_67, dataGroup_30_67};
  wire [63:0]   res_hi_hi_hi_67 = {res_hi_hi_hi_hi_67, res_hi_hi_hi_lo_67};
  wire [127:0]  res_hi_hi_67 = {res_hi_hi_hi_67, res_hi_hi_lo_67};
  wire [255:0]  res_hi_67 = {res_hi_hi_67, res_hi_lo_67};
  wire [511:0]  res_123 = {res_hi_67, res_lo_67};
  wire [2047:0] dataGroup_lo_3328 = {dataGroup_lo_hi_3328, dataGroup_lo_lo_3328};
  wire [2047:0] dataGroup_hi_3328 = {dataGroup_hi_hi_3328, dataGroup_hi_lo_3328};
  wire [15:0]   dataGroup_0_68 = dataGroup_lo_3328[79:64];
  wire [2047:0] dataGroup_lo_3329 = {dataGroup_lo_hi_3329, dataGroup_lo_lo_3329};
  wire [2047:0] dataGroup_hi_3329 = {dataGroup_hi_hi_3329, dataGroup_hi_lo_3329};
  wire [15:0]   dataGroup_1_68 = dataGroup_lo_3329[207:192];
  wire [2047:0] dataGroup_lo_3330 = {dataGroup_lo_hi_3330, dataGroup_lo_lo_3330};
  wire [2047:0] dataGroup_hi_3330 = {dataGroup_hi_hi_3330, dataGroup_hi_lo_3330};
  wire [15:0]   dataGroup_2_68 = dataGroup_lo_3330[335:320];
  wire [2047:0] dataGroup_lo_3331 = {dataGroup_lo_hi_3331, dataGroup_lo_lo_3331};
  wire [2047:0] dataGroup_hi_3331 = {dataGroup_hi_hi_3331, dataGroup_hi_lo_3331};
  wire [15:0]   dataGroup_3_68 = dataGroup_lo_3331[463:448];
  wire [2047:0] dataGroup_lo_3332 = {dataGroup_lo_hi_3332, dataGroup_lo_lo_3332};
  wire [2047:0] dataGroup_hi_3332 = {dataGroup_hi_hi_3332, dataGroup_hi_lo_3332};
  wire [15:0]   dataGroup_4_68 = dataGroup_lo_3332[591:576];
  wire [2047:0] dataGroup_lo_3333 = {dataGroup_lo_hi_3333, dataGroup_lo_lo_3333};
  wire [2047:0] dataGroup_hi_3333 = {dataGroup_hi_hi_3333, dataGroup_hi_lo_3333};
  wire [15:0]   dataGroup_5_68 = dataGroup_lo_3333[719:704];
  wire [2047:0] dataGroup_lo_3334 = {dataGroup_lo_hi_3334, dataGroup_lo_lo_3334};
  wire [2047:0] dataGroup_hi_3334 = {dataGroup_hi_hi_3334, dataGroup_hi_lo_3334};
  wire [15:0]   dataGroup_6_68 = dataGroup_lo_3334[847:832];
  wire [2047:0] dataGroup_lo_3335 = {dataGroup_lo_hi_3335, dataGroup_lo_lo_3335};
  wire [2047:0] dataGroup_hi_3335 = {dataGroup_hi_hi_3335, dataGroup_hi_lo_3335};
  wire [15:0]   dataGroup_7_68 = dataGroup_lo_3335[975:960];
  wire [2047:0] dataGroup_lo_3336 = {dataGroup_lo_hi_3336, dataGroup_lo_lo_3336};
  wire [2047:0] dataGroup_hi_3336 = {dataGroup_hi_hi_3336, dataGroup_hi_lo_3336};
  wire [15:0]   dataGroup_8_68 = dataGroup_lo_3336[1103:1088];
  wire [2047:0] dataGroup_lo_3337 = {dataGroup_lo_hi_3337, dataGroup_lo_lo_3337};
  wire [2047:0] dataGroup_hi_3337 = {dataGroup_hi_hi_3337, dataGroup_hi_lo_3337};
  wire [15:0]   dataGroup_9_68 = dataGroup_lo_3337[1231:1216];
  wire [2047:0] dataGroup_lo_3338 = {dataGroup_lo_hi_3338, dataGroup_lo_lo_3338};
  wire [2047:0] dataGroup_hi_3338 = {dataGroup_hi_hi_3338, dataGroup_hi_lo_3338};
  wire [15:0]   dataGroup_10_68 = dataGroup_lo_3338[1359:1344];
  wire [2047:0] dataGroup_lo_3339 = {dataGroup_lo_hi_3339, dataGroup_lo_lo_3339};
  wire [2047:0] dataGroup_hi_3339 = {dataGroup_hi_hi_3339, dataGroup_hi_lo_3339};
  wire [15:0]   dataGroup_11_68 = dataGroup_lo_3339[1487:1472];
  wire [2047:0] dataGroup_lo_3340 = {dataGroup_lo_hi_3340, dataGroup_lo_lo_3340};
  wire [2047:0] dataGroup_hi_3340 = {dataGroup_hi_hi_3340, dataGroup_hi_lo_3340};
  wire [15:0]   dataGroup_12_68 = dataGroup_lo_3340[1615:1600];
  wire [2047:0] dataGroup_lo_3341 = {dataGroup_lo_hi_3341, dataGroup_lo_lo_3341};
  wire [2047:0] dataGroup_hi_3341 = {dataGroup_hi_hi_3341, dataGroup_hi_lo_3341};
  wire [15:0]   dataGroup_13_68 = dataGroup_lo_3341[1743:1728];
  wire [2047:0] dataGroup_lo_3342 = {dataGroup_lo_hi_3342, dataGroup_lo_lo_3342};
  wire [2047:0] dataGroup_hi_3342 = {dataGroup_hi_hi_3342, dataGroup_hi_lo_3342};
  wire [15:0]   dataGroup_14_68 = dataGroup_lo_3342[1871:1856];
  wire [2047:0] dataGroup_lo_3343 = {dataGroup_lo_hi_3343, dataGroup_lo_lo_3343};
  wire [2047:0] dataGroup_hi_3343 = {dataGroup_hi_hi_3343, dataGroup_hi_lo_3343};
  wire [15:0]   dataGroup_15_68 = dataGroup_lo_3343[1999:1984];
  wire [2047:0] dataGroup_lo_3344 = {dataGroup_lo_hi_3344, dataGroup_lo_lo_3344};
  wire [2047:0] dataGroup_hi_3344 = {dataGroup_hi_hi_3344, dataGroup_hi_lo_3344};
  wire [15:0]   dataGroup_16_68 = dataGroup_hi_3344[79:64];
  wire [2047:0] dataGroup_lo_3345 = {dataGroup_lo_hi_3345, dataGroup_lo_lo_3345};
  wire [2047:0] dataGroup_hi_3345 = {dataGroup_hi_hi_3345, dataGroup_hi_lo_3345};
  wire [15:0]   dataGroup_17_68 = dataGroup_hi_3345[207:192];
  wire [2047:0] dataGroup_lo_3346 = {dataGroup_lo_hi_3346, dataGroup_lo_lo_3346};
  wire [2047:0] dataGroup_hi_3346 = {dataGroup_hi_hi_3346, dataGroup_hi_lo_3346};
  wire [15:0]   dataGroup_18_68 = dataGroup_hi_3346[335:320];
  wire [2047:0] dataGroup_lo_3347 = {dataGroup_lo_hi_3347, dataGroup_lo_lo_3347};
  wire [2047:0] dataGroup_hi_3347 = {dataGroup_hi_hi_3347, dataGroup_hi_lo_3347};
  wire [15:0]   dataGroup_19_68 = dataGroup_hi_3347[463:448];
  wire [2047:0] dataGroup_lo_3348 = {dataGroup_lo_hi_3348, dataGroup_lo_lo_3348};
  wire [2047:0] dataGroup_hi_3348 = {dataGroup_hi_hi_3348, dataGroup_hi_lo_3348};
  wire [15:0]   dataGroup_20_68 = dataGroup_hi_3348[591:576];
  wire [2047:0] dataGroup_lo_3349 = {dataGroup_lo_hi_3349, dataGroup_lo_lo_3349};
  wire [2047:0] dataGroup_hi_3349 = {dataGroup_hi_hi_3349, dataGroup_hi_lo_3349};
  wire [15:0]   dataGroup_21_68 = dataGroup_hi_3349[719:704];
  wire [2047:0] dataGroup_lo_3350 = {dataGroup_lo_hi_3350, dataGroup_lo_lo_3350};
  wire [2047:0] dataGroup_hi_3350 = {dataGroup_hi_hi_3350, dataGroup_hi_lo_3350};
  wire [15:0]   dataGroup_22_68 = dataGroup_hi_3350[847:832];
  wire [2047:0] dataGroup_lo_3351 = {dataGroup_lo_hi_3351, dataGroup_lo_lo_3351};
  wire [2047:0] dataGroup_hi_3351 = {dataGroup_hi_hi_3351, dataGroup_hi_lo_3351};
  wire [15:0]   dataGroup_23_68 = dataGroup_hi_3351[975:960];
  wire [2047:0] dataGroup_lo_3352 = {dataGroup_lo_hi_3352, dataGroup_lo_lo_3352};
  wire [2047:0] dataGroup_hi_3352 = {dataGroup_hi_hi_3352, dataGroup_hi_lo_3352};
  wire [15:0]   dataGroup_24_68 = dataGroup_hi_3352[1103:1088];
  wire [2047:0] dataGroup_lo_3353 = {dataGroup_lo_hi_3353, dataGroup_lo_lo_3353};
  wire [2047:0] dataGroup_hi_3353 = {dataGroup_hi_hi_3353, dataGroup_hi_lo_3353};
  wire [15:0]   dataGroup_25_68 = dataGroup_hi_3353[1231:1216];
  wire [2047:0] dataGroup_lo_3354 = {dataGroup_lo_hi_3354, dataGroup_lo_lo_3354};
  wire [2047:0] dataGroup_hi_3354 = {dataGroup_hi_hi_3354, dataGroup_hi_lo_3354};
  wire [15:0]   dataGroup_26_68 = dataGroup_hi_3354[1359:1344];
  wire [2047:0] dataGroup_lo_3355 = {dataGroup_lo_hi_3355, dataGroup_lo_lo_3355};
  wire [2047:0] dataGroup_hi_3355 = {dataGroup_hi_hi_3355, dataGroup_hi_lo_3355};
  wire [15:0]   dataGroup_27_68 = dataGroup_hi_3355[1487:1472];
  wire [2047:0] dataGroup_lo_3356 = {dataGroup_lo_hi_3356, dataGroup_lo_lo_3356};
  wire [2047:0] dataGroup_hi_3356 = {dataGroup_hi_hi_3356, dataGroup_hi_lo_3356};
  wire [15:0]   dataGroup_28_68 = dataGroup_hi_3356[1615:1600];
  wire [2047:0] dataGroup_lo_3357 = {dataGroup_lo_hi_3357, dataGroup_lo_lo_3357};
  wire [2047:0] dataGroup_hi_3357 = {dataGroup_hi_hi_3357, dataGroup_hi_lo_3357};
  wire [15:0]   dataGroup_29_68 = dataGroup_hi_3357[1743:1728];
  wire [2047:0] dataGroup_lo_3358 = {dataGroup_lo_hi_3358, dataGroup_lo_lo_3358};
  wire [2047:0] dataGroup_hi_3358 = {dataGroup_hi_hi_3358, dataGroup_hi_lo_3358};
  wire [15:0]   dataGroup_30_68 = dataGroup_hi_3358[1871:1856];
  wire [2047:0] dataGroup_lo_3359 = {dataGroup_lo_hi_3359, dataGroup_lo_lo_3359};
  wire [2047:0] dataGroup_hi_3359 = {dataGroup_hi_hi_3359, dataGroup_hi_lo_3359};
  wire [15:0]   dataGroup_31_68 = dataGroup_hi_3359[1999:1984];
  wire [31:0]   res_lo_lo_lo_lo_68 = {dataGroup_1_68, dataGroup_0_68};
  wire [31:0]   res_lo_lo_lo_hi_68 = {dataGroup_3_68, dataGroup_2_68};
  wire [63:0]   res_lo_lo_lo_68 = {res_lo_lo_lo_hi_68, res_lo_lo_lo_lo_68};
  wire [31:0]   res_lo_lo_hi_lo_68 = {dataGroup_5_68, dataGroup_4_68};
  wire [31:0]   res_lo_lo_hi_hi_68 = {dataGroup_7_68, dataGroup_6_68};
  wire [63:0]   res_lo_lo_hi_68 = {res_lo_lo_hi_hi_68, res_lo_lo_hi_lo_68};
  wire [127:0]  res_lo_lo_68 = {res_lo_lo_hi_68, res_lo_lo_lo_68};
  wire [31:0]   res_lo_hi_lo_lo_68 = {dataGroup_9_68, dataGroup_8_68};
  wire [31:0]   res_lo_hi_lo_hi_68 = {dataGroup_11_68, dataGroup_10_68};
  wire [63:0]   res_lo_hi_lo_68 = {res_lo_hi_lo_hi_68, res_lo_hi_lo_lo_68};
  wire [31:0]   res_lo_hi_hi_lo_68 = {dataGroup_13_68, dataGroup_12_68};
  wire [31:0]   res_lo_hi_hi_hi_68 = {dataGroup_15_68, dataGroup_14_68};
  wire [63:0]   res_lo_hi_hi_68 = {res_lo_hi_hi_hi_68, res_lo_hi_hi_lo_68};
  wire [127:0]  res_lo_hi_68 = {res_lo_hi_hi_68, res_lo_hi_lo_68};
  wire [255:0]  res_lo_68 = {res_lo_hi_68, res_lo_lo_68};
  wire [31:0]   res_hi_lo_lo_lo_68 = {dataGroup_17_68, dataGroup_16_68};
  wire [31:0]   res_hi_lo_lo_hi_68 = {dataGroup_19_68, dataGroup_18_68};
  wire [63:0]   res_hi_lo_lo_68 = {res_hi_lo_lo_hi_68, res_hi_lo_lo_lo_68};
  wire [31:0]   res_hi_lo_hi_lo_68 = {dataGroup_21_68, dataGroup_20_68};
  wire [31:0]   res_hi_lo_hi_hi_68 = {dataGroup_23_68, dataGroup_22_68};
  wire [63:0]   res_hi_lo_hi_68 = {res_hi_lo_hi_hi_68, res_hi_lo_hi_lo_68};
  wire [127:0]  res_hi_lo_68 = {res_hi_lo_hi_68, res_hi_lo_lo_68};
  wire [31:0]   res_hi_hi_lo_lo_68 = {dataGroup_25_68, dataGroup_24_68};
  wire [31:0]   res_hi_hi_lo_hi_68 = {dataGroup_27_68, dataGroup_26_68};
  wire [63:0]   res_hi_hi_lo_68 = {res_hi_hi_lo_hi_68, res_hi_hi_lo_lo_68};
  wire [31:0]   res_hi_hi_hi_lo_68 = {dataGroup_29_68, dataGroup_28_68};
  wire [31:0]   res_hi_hi_hi_hi_68 = {dataGroup_31_68, dataGroup_30_68};
  wire [63:0]   res_hi_hi_hi_68 = {res_hi_hi_hi_hi_68, res_hi_hi_hi_lo_68};
  wire [127:0]  res_hi_hi_68 = {res_hi_hi_hi_68, res_hi_hi_lo_68};
  wire [255:0]  res_hi_68 = {res_hi_hi_68, res_hi_lo_68};
  wire [511:0]  res_124 = {res_hi_68, res_lo_68};
  wire [2047:0] dataGroup_lo_3360 = {dataGroup_lo_hi_3360, dataGroup_lo_lo_3360};
  wire [2047:0] dataGroup_hi_3360 = {dataGroup_hi_hi_3360, dataGroup_hi_lo_3360};
  wire [15:0]   dataGroup_0_69 = dataGroup_lo_3360[95:80];
  wire [2047:0] dataGroup_lo_3361 = {dataGroup_lo_hi_3361, dataGroup_lo_lo_3361};
  wire [2047:0] dataGroup_hi_3361 = {dataGroup_hi_hi_3361, dataGroup_hi_lo_3361};
  wire [15:0]   dataGroup_1_69 = dataGroup_lo_3361[223:208];
  wire [2047:0] dataGroup_lo_3362 = {dataGroup_lo_hi_3362, dataGroup_lo_lo_3362};
  wire [2047:0] dataGroup_hi_3362 = {dataGroup_hi_hi_3362, dataGroup_hi_lo_3362};
  wire [15:0]   dataGroup_2_69 = dataGroup_lo_3362[351:336];
  wire [2047:0] dataGroup_lo_3363 = {dataGroup_lo_hi_3363, dataGroup_lo_lo_3363};
  wire [2047:0] dataGroup_hi_3363 = {dataGroup_hi_hi_3363, dataGroup_hi_lo_3363};
  wire [15:0]   dataGroup_3_69 = dataGroup_lo_3363[479:464];
  wire [2047:0] dataGroup_lo_3364 = {dataGroup_lo_hi_3364, dataGroup_lo_lo_3364};
  wire [2047:0] dataGroup_hi_3364 = {dataGroup_hi_hi_3364, dataGroup_hi_lo_3364};
  wire [15:0]   dataGroup_4_69 = dataGroup_lo_3364[607:592];
  wire [2047:0] dataGroup_lo_3365 = {dataGroup_lo_hi_3365, dataGroup_lo_lo_3365};
  wire [2047:0] dataGroup_hi_3365 = {dataGroup_hi_hi_3365, dataGroup_hi_lo_3365};
  wire [15:0]   dataGroup_5_69 = dataGroup_lo_3365[735:720];
  wire [2047:0] dataGroup_lo_3366 = {dataGroup_lo_hi_3366, dataGroup_lo_lo_3366};
  wire [2047:0] dataGroup_hi_3366 = {dataGroup_hi_hi_3366, dataGroup_hi_lo_3366};
  wire [15:0]   dataGroup_6_69 = dataGroup_lo_3366[863:848];
  wire [2047:0] dataGroup_lo_3367 = {dataGroup_lo_hi_3367, dataGroup_lo_lo_3367};
  wire [2047:0] dataGroup_hi_3367 = {dataGroup_hi_hi_3367, dataGroup_hi_lo_3367};
  wire [15:0]   dataGroup_7_69 = dataGroup_lo_3367[991:976];
  wire [2047:0] dataGroup_lo_3368 = {dataGroup_lo_hi_3368, dataGroup_lo_lo_3368};
  wire [2047:0] dataGroup_hi_3368 = {dataGroup_hi_hi_3368, dataGroup_hi_lo_3368};
  wire [15:0]   dataGroup_8_69 = dataGroup_lo_3368[1119:1104];
  wire [2047:0] dataGroup_lo_3369 = {dataGroup_lo_hi_3369, dataGroup_lo_lo_3369};
  wire [2047:0] dataGroup_hi_3369 = {dataGroup_hi_hi_3369, dataGroup_hi_lo_3369};
  wire [15:0]   dataGroup_9_69 = dataGroup_lo_3369[1247:1232];
  wire [2047:0] dataGroup_lo_3370 = {dataGroup_lo_hi_3370, dataGroup_lo_lo_3370};
  wire [2047:0] dataGroup_hi_3370 = {dataGroup_hi_hi_3370, dataGroup_hi_lo_3370};
  wire [15:0]   dataGroup_10_69 = dataGroup_lo_3370[1375:1360];
  wire [2047:0] dataGroup_lo_3371 = {dataGroup_lo_hi_3371, dataGroup_lo_lo_3371};
  wire [2047:0] dataGroup_hi_3371 = {dataGroup_hi_hi_3371, dataGroup_hi_lo_3371};
  wire [15:0]   dataGroup_11_69 = dataGroup_lo_3371[1503:1488];
  wire [2047:0] dataGroup_lo_3372 = {dataGroup_lo_hi_3372, dataGroup_lo_lo_3372};
  wire [2047:0] dataGroup_hi_3372 = {dataGroup_hi_hi_3372, dataGroup_hi_lo_3372};
  wire [15:0]   dataGroup_12_69 = dataGroup_lo_3372[1631:1616];
  wire [2047:0] dataGroup_lo_3373 = {dataGroup_lo_hi_3373, dataGroup_lo_lo_3373};
  wire [2047:0] dataGroup_hi_3373 = {dataGroup_hi_hi_3373, dataGroup_hi_lo_3373};
  wire [15:0]   dataGroup_13_69 = dataGroup_lo_3373[1759:1744];
  wire [2047:0] dataGroup_lo_3374 = {dataGroup_lo_hi_3374, dataGroup_lo_lo_3374};
  wire [2047:0] dataGroup_hi_3374 = {dataGroup_hi_hi_3374, dataGroup_hi_lo_3374};
  wire [15:0]   dataGroup_14_69 = dataGroup_lo_3374[1887:1872];
  wire [2047:0] dataGroup_lo_3375 = {dataGroup_lo_hi_3375, dataGroup_lo_lo_3375};
  wire [2047:0] dataGroup_hi_3375 = {dataGroup_hi_hi_3375, dataGroup_hi_lo_3375};
  wire [15:0]   dataGroup_15_69 = dataGroup_lo_3375[2015:2000];
  wire [2047:0] dataGroup_lo_3376 = {dataGroup_lo_hi_3376, dataGroup_lo_lo_3376};
  wire [2047:0] dataGroup_hi_3376 = {dataGroup_hi_hi_3376, dataGroup_hi_lo_3376};
  wire [15:0]   dataGroup_16_69 = dataGroup_hi_3376[95:80];
  wire [2047:0] dataGroup_lo_3377 = {dataGroup_lo_hi_3377, dataGroup_lo_lo_3377};
  wire [2047:0] dataGroup_hi_3377 = {dataGroup_hi_hi_3377, dataGroup_hi_lo_3377};
  wire [15:0]   dataGroup_17_69 = dataGroup_hi_3377[223:208];
  wire [2047:0] dataGroup_lo_3378 = {dataGroup_lo_hi_3378, dataGroup_lo_lo_3378};
  wire [2047:0] dataGroup_hi_3378 = {dataGroup_hi_hi_3378, dataGroup_hi_lo_3378};
  wire [15:0]   dataGroup_18_69 = dataGroup_hi_3378[351:336];
  wire [2047:0] dataGroup_lo_3379 = {dataGroup_lo_hi_3379, dataGroup_lo_lo_3379};
  wire [2047:0] dataGroup_hi_3379 = {dataGroup_hi_hi_3379, dataGroup_hi_lo_3379};
  wire [15:0]   dataGroup_19_69 = dataGroup_hi_3379[479:464];
  wire [2047:0] dataGroup_lo_3380 = {dataGroup_lo_hi_3380, dataGroup_lo_lo_3380};
  wire [2047:0] dataGroup_hi_3380 = {dataGroup_hi_hi_3380, dataGroup_hi_lo_3380};
  wire [15:0]   dataGroup_20_69 = dataGroup_hi_3380[607:592];
  wire [2047:0] dataGroup_lo_3381 = {dataGroup_lo_hi_3381, dataGroup_lo_lo_3381};
  wire [2047:0] dataGroup_hi_3381 = {dataGroup_hi_hi_3381, dataGroup_hi_lo_3381};
  wire [15:0]   dataGroup_21_69 = dataGroup_hi_3381[735:720];
  wire [2047:0] dataGroup_lo_3382 = {dataGroup_lo_hi_3382, dataGroup_lo_lo_3382};
  wire [2047:0] dataGroup_hi_3382 = {dataGroup_hi_hi_3382, dataGroup_hi_lo_3382};
  wire [15:0]   dataGroup_22_69 = dataGroup_hi_3382[863:848];
  wire [2047:0] dataGroup_lo_3383 = {dataGroup_lo_hi_3383, dataGroup_lo_lo_3383};
  wire [2047:0] dataGroup_hi_3383 = {dataGroup_hi_hi_3383, dataGroup_hi_lo_3383};
  wire [15:0]   dataGroup_23_69 = dataGroup_hi_3383[991:976];
  wire [2047:0] dataGroup_lo_3384 = {dataGroup_lo_hi_3384, dataGroup_lo_lo_3384};
  wire [2047:0] dataGroup_hi_3384 = {dataGroup_hi_hi_3384, dataGroup_hi_lo_3384};
  wire [15:0]   dataGroup_24_69 = dataGroup_hi_3384[1119:1104];
  wire [2047:0] dataGroup_lo_3385 = {dataGroup_lo_hi_3385, dataGroup_lo_lo_3385};
  wire [2047:0] dataGroup_hi_3385 = {dataGroup_hi_hi_3385, dataGroup_hi_lo_3385};
  wire [15:0]   dataGroup_25_69 = dataGroup_hi_3385[1247:1232];
  wire [2047:0] dataGroup_lo_3386 = {dataGroup_lo_hi_3386, dataGroup_lo_lo_3386};
  wire [2047:0] dataGroup_hi_3386 = {dataGroup_hi_hi_3386, dataGroup_hi_lo_3386};
  wire [15:0]   dataGroup_26_69 = dataGroup_hi_3386[1375:1360];
  wire [2047:0] dataGroup_lo_3387 = {dataGroup_lo_hi_3387, dataGroup_lo_lo_3387};
  wire [2047:0] dataGroup_hi_3387 = {dataGroup_hi_hi_3387, dataGroup_hi_lo_3387};
  wire [15:0]   dataGroup_27_69 = dataGroup_hi_3387[1503:1488];
  wire [2047:0] dataGroup_lo_3388 = {dataGroup_lo_hi_3388, dataGroup_lo_lo_3388};
  wire [2047:0] dataGroup_hi_3388 = {dataGroup_hi_hi_3388, dataGroup_hi_lo_3388};
  wire [15:0]   dataGroup_28_69 = dataGroup_hi_3388[1631:1616];
  wire [2047:0] dataGroup_lo_3389 = {dataGroup_lo_hi_3389, dataGroup_lo_lo_3389};
  wire [2047:0] dataGroup_hi_3389 = {dataGroup_hi_hi_3389, dataGroup_hi_lo_3389};
  wire [15:0]   dataGroup_29_69 = dataGroup_hi_3389[1759:1744];
  wire [2047:0] dataGroup_lo_3390 = {dataGroup_lo_hi_3390, dataGroup_lo_lo_3390};
  wire [2047:0] dataGroup_hi_3390 = {dataGroup_hi_hi_3390, dataGroup_hi_lo_3390};
  wire [15:0]   dataGroup_30_69 = dataGroup_hi_3390[1887:1872];
  wire [2047:0] dataGroup_lo_3391 = {dataGroup_lo_hi_3391, dataGroup_lo_lo_3391};
  wire [2047:0] dataGroup_hi_3391 = {dataGroup_hi_hi_3391, dataGroup_hi_lo_3391};
  wire [15:0]   dataGroup_31_69 = dataGroup_hi_3391[2015:2000];
  wire [31:0]   res_lo_lo_lo_lo_69 = {dataGroup_1_69, dataGroup_0_69};
  wire [31:0]   res_lo_lo_lo_hi_69 = {dataGroup_3_69, dataGroup_2_69};
  wire [63:0]   res_lo_lo_lo_69 = {res_lo_lo_lo_hi_69, res_lo_lo_lo_lo_69};
  wire [31:0]   res_lo_lo_hi_lo_69 = {dataGroup_5_69, dataGroup_4_69};
  wire [31:0]   res_lo_lo_hi_hi_69 = {dataGroup_7_69, dataGroup_6_69};
  wire [63:0]   res_lo_lo_hi_69 = {res_lo_lo_hi_hi_69, res_lo_lo_hi_lo_69};
  wire [127:0]  res_lo_lo_69 = {res_lo_lo_hi_69, res_lo_lo_lo_69};
  wire [31:0]   res_lo_hi_lo_lo_69 = {dataGroup_9_69, dataGroup_8_69};
  wire [31:0]   res_lo_hi_lo_hi_69 = {dataGroup_11_69, dataGroup_10_69};
  wire [63:0]   res_lo_hi_lo_69 = {res_lo_hi_lo_hi_69, res_lo_hi_lo_lo_69};
  wire [31:0]   res_lo_hi_hi_lo_69 = {dataGroup_13_69, dataGroup_12_69};
  wire [31:0]   res_lo_hi_hi_hi_69 = {dataGroup_15_69, dataGroup_14_69};
  wire [63:0]   res_lo_hi_hi_69 = {res_lo_hi_hi_hi_69, res_lo_hi_hi_lo_69};
  wire [127:0]  res_lo_hi_69 = {res_lo_hi_hi_69, res_lo_hi_lo_69};
  wire [255:0]  res_lo_69 = {res_lo_hi_69, res_lo_lo_69};
  wire [31:0]   res_hi_lo_lo_lo_69 = {dataGroup_17_69, dataGroup_16_69};
  wire [31:0]   res_hi_lo_lo_hi_69 = {dataGroup_19_69, dataGroup_18_69};
  wire [63:0]   res_hi_lo_lo_69 = {res_hi_lo_lo_hi_69, res_hi_lo_lo_lo_69};
  wire [31:0]   res_hi_lo_hi_lo_69 = {dataGroup_21_69, dataGroup_20_69};
  wire [31:0]   res_hi_lo_hi_hi_69 = {dataGroup_23_69, dataGroup_22_69};
  wire [63:0]   res_hi_lo_hi_69 = {res_hi_lo_hi_hi_69, res_hi_lo_hi_lo_69};
  wire [127:0]  res_hi_lo_69 = {res_hi_lo_hi_69, res_hi_lo_lo_69};
  wire [31:0]   res_hi_hi_lo_lo_69 = {dataGroup_25_69, dataGroup_24_69};
  wire [31:0]   res_hi_hi_lo_hi_69 = {dataGroup_27_69, dataGroup_26_69};
  wire [63:0]   res_hi_hi_lo_69 = {res_hi_hi_lo_hi_69, res_hi_hi_lo_lo_69};
  wire [31:0]   res_hi_hi_hi_lo_69 = {dataGroup_29_69, dataGroup_28_69};
  wire [31:0]   res_hi_hi_hi_hi_69 = {dataGroup_31_69, dataGroup_30_69};
  wire [63:0]   res_hi_hi_hi_69 = {res_hi_hi_hi_hi_69, res_hi_hi_hi_lo_69};
  wire [127:0]  res_hi_hi_69 = {res_hi_hi_hi_69, res_hi_hi_lo_69};
  wire [255:0]  res_hi_69 = {res_hi_hi_69, res_hi_lo_69};
  wire [511:0]  res_125 = {res_hi_69, res_lo_69};
  wire [2047:0] dataGroup_lo_3392 = {dataGroup_lo_hi_3392, dataGroup_lo_lo_3392};
  wire [2047:0] dataGroup_hi_3392 = {dataGroup_hi_hi_3392, dataGroup_hi_lo_3392};
  wire [15:0]   dataGroup_0_70 = dataGroup_lo_3392[111:96];
  wire [2047:0] dataGroup_lo_3393 = {dataGroup_lo_hi_3393, dataGroup_lo_lo_3393};
  wire [2047:0] dataGroup_hi_3393 = {dataGroup_hi_hi_3393, dataGroup_hi_lo_3393};
  wire [15:0]   dataGroup_1_70 = dataGroup_lo_3393[239:224];
  wire [2047:0] dataGroup_lo_3394 = {dataGroup_lo_hi_3394, dataGroup_lo_lo_3394};
  wire [2047:0] dataGroup_hi_3394 = {dataGroup_hi_hi_3394, dataGroup_hi_lo_3394};
  wire [15:0]   dataGroup_2_70 = dataGroup_lo_3394[367:352];
  wire [2047:0] dataGroup_lo_3395 = {dataGroup_lo_hi_3395, dataGroup_lo_lo_3395};
  wire [2047:0] dataGroup_hi_3395 = {dataGroup_hi_hi_3395, dataGroup_hi_lo_3395};
  wire [15:0]   dataGroup_3_70 = dataGroup_lo_3395[495:480];
  wire [2047:0] dataGroup_lo_3396 = {dataGroup_lo_hi_3396, dataGroup_lo_lo_3396};
  wire [2047:0] dataGroup_hi_3396 = {dataGroup_hi_hi_3396, dataGroup_hi_lo_3396};
  wire [15:0]   dataGroup_4_70 = dataGroup_lo_3396[623:608];
  wire [2047:0] dataGroup_lo_3397 = {dataGroup_lo_hi_3397, dataGroup_lo_lo_3397};
  wire [2047:0] dataGroup_hi_3397 = {dataGroup_hi_hi_3397, dataGroup_hi_lo_3397};
  wire [15:0]   dataGroup_5_70 = dataGroup_lo_3397[751:736];
  wire [2047:0] dataGroup_lo_3398 = {dataGroup_lo_hi_3398, dataGroup_lo_lo_3398};
  wire [2047:0] dataGroup_hi_3398 = {dataGroup_hi_hi_3398, dataGroup_hi_lo_3398};
  wire [15:0]   dataGroup_6_70 = dataGroup_lo_3398[879:864];
  wire [2047:0] dataGroup_lo_3399 = {dataGroup_lo_hi_3399, dataGroup_lo_lo_3399};
  wire [2047:0] dataGroup_hi_3399 = {dataGroup_hi_hi_3399, dataGroup_hi_lo_3399};
  wire [15:0]   dataGroup_7_70 = dataGroup_lo_3399[1007:992];
  wire [2047:0] dataGroup_lo_3400 = {dataGroup_lo_hi_3400, dataGroup_lo_lo_3400};
  wire [2047:0] dataGroup_hi_3400 = {dataGroup_hi_hi_3400, dataGroup_hi_lo_3400};
  wire [15:0]   dataGroup_8_70 = dataGroup_lo_3400[1135:1120];
  wire [2047:0] dataGroup_lo_3401 = {dataGroup_lo_hi_3401, dataGroup_lo_lo_3401};
  wire [2047:0] dataGroup_hi_3401 = {dataGroup_hi_hi_3401, dataGroup_hi_lo_3401};
  wire [15:0]   dataGroup_9_70 = dataGroup_lo_3401[1263:1248];
  wire [2047:0] dataGroup_lo_3402 = {dataGroup_lo_hi_3402, dataGroup_lo_lo_3402};
  wire [2047:0] dataGroup_hi_3402 = {dataGroup_hi_hi_3402, dataGroup_hi_lo_3402};
  wire [15:0]   dataGroup_10_70 = dataGroup_lo_3402[1391:1376];
  wire [2047:0] dataGroup_lo_3403 = {dataGroup_lo_hi_3403, dataGroup_lo_lo_3403};
  wire [2047:0] dataGroup_hi_3403 = {dataGroup_hi_hi_3403, dataGroup_hi_lo_3403};
  wire [15:0]   dataGroup_11_70 = dataGroup_lo_3403[1519:1504];
  wire [2047:0] dataGroup_lo_3404 = {dataGroup_lo_hi_3404, dataGroup_lo_lo_3404};
  wire [2047:0] dataGroup_hi_3404 = {dataGroup_hi_hi_3404, dataGroup_hi_lo_3404};
  wire [15:0]   dataGroup_12_70 = dataGroup_lo_3404[1647:1632];
  wire [2047:0] dataGroup_lo_3405 = {dataGroup_lo_hi_3405, dataGroup_lo_lo_3405};
  wire [2047:0] dataGroup_hi_3405 = {dataGroup_hi_hi_3405, dataGroup_hi_lo_3405};
  wire [15:0]   dataGroup_13_70 = dataGroup_lo_3405[1775:1760];
  wire [2047:0] dataGroup_lo_3406 = {dataGroup_lo_hi_3406, dataGroup_lo_lo_3406};
  wire [2047:0] dataGroup_hi_3406 = {dataGroup_hi_hi_3406, dataGroup_hi_lo_3406};
  wire [15:0]   dataGroup_14_70 = dataGroup_lo_3406[1903:1888];
  wire [2047:0] dataGroup_lo_3407 = {dataGroup_lo_hi_3407, dataGroup_lo_lo_3407};
  wire [2047:0] dataGroup_hi_3407 = {dataGroup_hi_hi_3407, dataGroup_hi_lo_3407};
  wire [15:0]   dataGroup_15_70 = dataGroup_lo_3407[2031:2016];
  wire [2047:0] dataGroup_lo_3408 = {dataGroup_lo_hi_3408, dataGroup_lo_lo_3408};
  wire [2047:0] dataGroup_hi_3408 = {dataGroup_hi_hi_3408, dataGroup_hi_lo_3408};
  wire [15:0]   dataGroup_16_70 = dataGroup_hi_3408[111:96];
  wire [2047:0] dataGroup_lo_3409 = {dataGroup_lo_hi_3409, dataGroup_lo_lo_3409};
  wire [2047:0] dataGroup_hi_3409 = {dataGroup_hi_hi_3409, dataGroup_hi_lo_3409};
  wire [15:0]   dataGroup_17_70 = dataGroup_hi_3409[239:224];
  wire [2047:0] dataGroup_lo_3410 = {dataGroup_lo_hi_3410, dataGroup_lo_lo_3410};
  wire [2047:0] dataGroup_hi_3410 = {dataGroup_hi_hi_3410, dataGroup_hi_lo_3410};
  wire [15:0]   dataGroup_18_70 = dataGroup_hi_3410[367:352];
  wire [2047:0] dataGroup_lo_3411 = {dataGroup_lo_hi_3411, dataGroup_lo_lo_3411};
  wire [2047:0] dataGroup_hi_3411 = {dataGroup_hi_hi_3411, dataGroup_hi_lo_3411};
  wire [15:0]   dataGroup_19_70 = dataGroup_hi_3411[495:480];
  wire [2047:0] dataGroup_lo_3412 = {dataGroup_lo_hi_3412, dataGroup_lo_lo_3412};
  wire [2047:0] dataGroup_hi_3412 = {dataGroup_hi_hi_3412, dataGroup_hi_lo_3412};
  wire [15:0]   dataGroup_20_70 = dataGroup_hi_3412[623:608];
  wire [2047:0] dataGroup_lo_3413 = {dataGroup_lo_hi_3413, dataGroup_lo_lo_3413};
  wire [2047:0] dataGroup_hi_3413 = {dataGroup_hi_hi_3413, dataGroup_hi_lo_3413};
  wire [15:0]   dataGroup_21_70 = dataGroup_hi_3413[751:736];
  wire [2047:0] dataGroup_lo_3414 = {dataGroup_lo_hi_3414, dataGroup_lo_lo_3414};
  wire [2047:0] dataGroup_hi_3414 = {dataGroup_hi_hi_3414, dataGroup_hi_lo_3414};
  wire [15:0]   dataGroup_22_70 = dataGroup_hi_3414[879:864];
  wire [2047:0] dataGroup_lo_3415 = {dataGroup_lo_hi_3415, dataGroup_lo_lo_3415};
  wire [2047:0] dataGroup_hi_3415 = {dataGroup_hi_hi_3415, dataGroup_hi_lo_3415};
  wire [15:0]   dataGroup_23_70 = dataGroup_hi_3415[1007:992];
  wire [2047:0] dataGroup_lo_3416 = {dataGroup_lo_hi_3416, dataGroup_lo_lo_3416};
  wire [2047:0] dataGroup_hi_3416 = {dataGroup_hi_hi_3416, dataGroup_hi_lo_3416};
  wire [15:0]   dataGroup_24_70 = dataGroup_hi_3416[1135:1120];
  wire [2047:0] dataGroup_lo_3417 = {dataGroup_lo_hi_3417, dataGroup_lo_lo_3417};
  wire [2047:0] dataGroup_hi_3417 = {dataGroup_hi_hi_3417, dataGroup_hi_lo_3417};
  wire [15:0]   dataGroup_25_70 = dataGroup_hi_3417[1263:1248];
  wire [2047:0] dataGroup_lo_3418 = {dataGroup_lo_hi_3418, dataGroup_lo_lo_3418};
  wire [2047:0] dataGroup_hi_3418 = {dataGroup_hi_hi_3418, dataGroup_hi_lo_3418};
  wire [15:0]   dataGroup_26_70 = dataGroup_hi_3418[1391:1376];
  wire [2047:0] dataGroup_lo_3419 = {dataGroup_lo_hi_3419, dataGroup_lo_lo_3419};
  wire [2047:0] dataGroup_hi_3419 = {dataGroup_hi_hi_3419, dataGroup_hi_lo_3419};
  wire [15:0]   dataGroup_27_70 = dataGroup_hi_3419[1519:1504];
  wire [2047:0] dataGroup_lo_3420 = {dataGroup_lo_hi_3420, dataGroup_lo_lo_3420};
  wire [2047:0] dataGroup_hi_3420 = {dataGroup_hi_hi_3420, dataGroup_hi_lo_3420};
  wire [15:0]   dataGroup_28_70 = dataGroup_hi_3420[1647:1632];
  wire [2047:0] dataGroup_lo_3421 = {dataGroup_lo_hi_3421, dataGroup_lo_lo_3421};
  wire [2047:0] dataGroup_hi_3421 = {dataGroup_hi_hi_3421, dataGroup_hi_lo_3421};
  wire [15:0]   dataGroup_29_70 = dataGroup_hi_3421[1775:1760];
  wire [2047:0] dataGroup_lo_3422 = {dataGroup_lo_hi_3422, dataGroup_lo_lo_3422};
  wire [2047:0] dataGroup_hi_3422 = {dataGroup_hi_hi_3422, dataGroup_hi_lo_3422};
  wire [15:0]   dataGroup_30_70 = dataGroup_hi_3422[1903:1888];
  wire [2047:0] dataGroup_lo_3423 = {dataGroup_lo_hi_3423, dataGroup_lo_lo_3423};
  wire [2047:0] dataGroup_hi_3423 = {dataGroup_hi_hi_3423, dataGroup_hi_lo_3423};
  wire [15:0]   dataGroup_31_70 = dataGroup_hi_3423[2031:2016];
  wire [31:0]   res_lo_lo_lo_lo_70 = {dataGroup_1_70, dataGroup_0_70};
  wire [31:0]   res_lo_lo_lo_hi_70 = {dataGroup_3_70, dataGroup_2_70};
  wire [63:0]   res_lo_lo_lo_70 = {res_lo_lo_lo_hi_70, res_lo_lo_lo_lo_70};
  wire [31:0]   res_lo_lo_hi_lo_70 = {dataGroup_5_70, dataGroup_4_70};
  wire [31:0]   res_lo_lo_hi_hi_70 = {dataGroup_7_70, dataGroup_6_70};
  wire [63:0]   res_lo_lo_hi_70 = {res_lo_lo_hi_hi_70, res_lo_lo_hi_lo_70};
  wire [127:0]  res_lo_lo_70 = {res_lo_lo_hi_70, res_lo_lo_lo_70};
  wire [31:0]   res_lo_hi_lo_lo_70 = {dataGroup_9_70, dataGroup_8_70};
  wire [31:0]   res_lo_hi_lo_hi_70 = {dataGroup_11_70, dataGroup_10_70};
  wire [63:0]   res_lo_hi_lo_70 = {res_lo_hi_lo_hi_70, res_lo_hi_lo_lo_70};
  wire [31:0]   res_lo_hi_hi_lo_70 = {dataGroup_13_70, dataGroup_12_70};
  wire [31:0]   res_lo_hi_hi_hi_70 = {dataGroup_15_70, dataGroup_14_70};
  wire [63:0]   res_lo_hi_hi_70 = {res_lo_hi_hi_hi_70, res_lo_hi_hi_lo_70};
  wire [127:0]  res_lo_hi_70 = {res_lo_hi_hi_70, res_lo_hi_lo_70};
  wire [255:0]  res_lo_70 = {res_lo_hi_70, res_lo_lo_70};
  wire [31:0]   res_hi_lo_lo_lo_70 = {dataGroup_17_70, dataGroup_16_70};
  wire [31:0]   res_hi_lo_lo_hi_70 = {dataGroup_19_70, dataGroup_18_70};
  wire [63:0]   res_hi_lo_lo_70 = {res_hi_lo_lo_hi_70, res_hi_lo_lo_lo_70};
  wire [31:0]   res_hi_lo_hi_lo_70 = {dataGroup_21_70, dataGroup_20_70};
  wire [31:0]   res_hi_lo_hi_hi_70 = {dataGroup_23_70, dataGroup_22_70};
  wire [63:0]   res_hi_lo_hi_70 = {res_hi_lo_hi_hi_70, res_hi_lo_hi_lo_70};
  wire [127:0]  res_hi_lo_70 = {res_hi_lo_hi_70, res_hi_lo_lo_70};
  wire [31:0]   res_hi_hi_lo_lo_70 = {dataGroup_25_70, dataGroup_24_70};
  wire [31:0]   res_hi_hi_lo_hi_70 = {dataGroup_27_70, dataGroup_26_70};
  wire [63:0]   res_hi_hi_lo_70 = {res_hi_hi_lo_hi_70, res_hi_hi_lo_lo_70};
  wire [31:0]   res_hi_hi_hi_lo_70 = {dataGroup_29_70, dataGroup_28_70};
  wire [31:0]   res_hi_hi_hi_hi_70 = {dataGroup_31_70, dataGroup_30_70};
  wire [63:0]   res_hi_hi_hi_70 = {res_hi_hi_hi_hi_70, res_hi_hi_hi_lo_70};
  wire [127:0]  res_hi_hi_70 = {res_hi_hi_hi_70, res_hi_hi_lo_70};
  wire [255:0]  res_hi_70 = {res_hi_hi_70, res_hi_lo_70};
  wire [511:0]  res_126 = {res_hi_70, res_lo_70};
  wire [2047:0] dataGroup_lo_3424 = {dataGroup_lo_hi_3424, dataGroup_lo_lo_3424};
  wire [2047:0] dataGroup_hi_3424 = {dataGroup_hi_hi_3424, dataGroup_hi_lo_3424};
  wire [15:0]   dataGroup_0_71 = dataGroup_lo_3424[127:112];
  wire [2047:0] dataGroup_lo_3425 = {dataGroup_lo_hi_3425, dataGroup_lo_lo_3425};
  wire [2047:0] dataGroup_hi_3425 = {dataGroup_hi_hi_3425, dataGroup_hi_lo_3425};
  wire [15:0]   dataGroup_1_71 = dataGroup_lo_3425[255:240];
  wire [2047:0] dataGroup_lo_3426 = {dataGroup_lo_hi_3426, dataGroup_lo_lo_3426};
  wire [2047:0] dataGroup_hi_3426 = {dataGroup_hi_hi_3426, dataGroup_hi_lo_3426};
  wire [15:0]   dataGroup_2_71 = dataGroup_lo_3426[383:368];
  wire [2047:0] dataGroup_lo_3427 = {dataGroup_lo_hi_3427, dataGroup_lo_lo_3427};
  wire [2047:0] dataGroup_hi_3427 = {dataGroup_hi_hi_3427, dataGroup_hi_lo_3427};
  wire [15:0]   dataGroup_3_71 = dataGroup_lo_3427[511:496];
  wire [2047:0] dataGroup_lo_3428 = {dataGroup_lo_hi_3428, dataGroup_lo_lo_3428};
  wire [2047:0] dataGroup_hi_3428 = {dataGroup_hi_hi_3428, dataGroup_hi_lo_3428};
  wire [15:0]   dataGroup_4_71 = dataGroup_lo_3428[639:624];
  wire [2047:0] dataGroup_lo_3429 = {dataGroup_lo_hi_3429, dataGroup_lo_lo_3429};
  wire [2047:0] dataGroup_hi_3429 = {dataGroup_hi_hi_3429, dataGroup_hi_lo_3429};
  wire [15:0]   dataGroup_5_71 = dataGroup_lo_3429[767:752];
  wire [2047:0] dataGroup_lo_3430 = {dataGroup_lo_hi_3430, dataGroup_lo_lo_3430};
  wire [2047:0] dataGroup_hi_3430 = {dataGroup_hi_hi_3430, dataGroup_hi_lo_3430};
  wire [15:0]   dataGroup_6_71 = dataGroup_lo_3430[895:880];
  wire [2047:0] dataGroup_lo_3431 = {dataGroup_lo_hi_3431, dataGroup_lo_lo_3431};
  wire [2047:0] dataGroup_hi_3431 = {dataGroup_hi_hi_3431, dataGroup_hi_lo_3431};
  wire [15:0]   dataGroup_7_71 = dataGroup_lo_3431[1023:1008];
  wire [2047:0] dataGroup_lo_3432 = {dataGroup_lo_hi_3432, dataGroup_lo_lo_3432};
  wire [2047:0] dataGroup_hi_3432 = {dataGroup_hi_hi_3432, dataGroup_hi_lo_3432};
  wire [15:0]   dataGroup_8_71 = dataGroup_lo_3432[1151:1136];
  wire [2047:0] dataGroup_lo_3433 = {dataGroup_lo_hi_3433, dataGroup_lo_lo_3433};
  wire [2047:0] dataGroup_hi_3433 = {dataGroup_hi_hi_3433, dataGroup_hi_lo_3433};
  wire [15:0]   dataGroup_9_71 = dataGroup_lo_3433[1279:1264];
  wire [2047:0] dataGroup_lo_3434 = {dataGroup_lo_hi_3434, dataGroup_lo_lo_3434};
  wire [2047:0] dataGroup_hi_3434 = {dataGroup_hi_hi_3434, dataGroup_hi_lo_3434};
  wire [15:0]   dataGroup_10_71 = dataGroup_lo_3434[1407:1392];
  wire [2047:0] dataGroup_lo_3435 = {dataGroup_lo_hi_3435, dataGroup_lo_lo_3435};
  wire [2047:0] dataGroup_hi_3435 = {dataGroup_hi_hi_3435, dataGroup_hi_lo_3435};
  wire [15:0]   dataGroup_11_71 = dataGroup_lo_3435[1535:1520];
  wire [2047:0] dataGroup_lo_3436 = {dataGroup_lo_hi_3436, dataGroup_lo_lo_3436};
  wire [2047:0] dataGroup_hi_3436 = {dataGroup_hi_hi_3436, dataGroup_hi_lo_3436};
  wire [15:0]   dataGroup_12_71 = dataGroup_lo_3436[1663:1648];
  wire [2047:0] dataGroup_lo_3437 = {dataGroup_lo_hi_3437, dataGroup_lo_lo_3437};
  wire [2047:0] dataGroup_hi_3437 = {dataGroup_hi_hi_3437, dataGroup_hi_lo_3437};
  wire [15:0]   dataGroup_13_71 = dataGroup_lo_3437[1791:1776];
  wire [2047:0] dataGroup_lo_3438 = {dataGroup_lo_hi_3438, dataGroup_lo_lo_3438};
  wire [2047:0] dataGroup_hi_3438 = {dataGroup_hi_hi_3438, dataGroup_hi_lo_3438};
  wire [15:0]   dataGroup_14_71 = dataGroup_lo_3438[1919:1904];
  wire [2047:0] dataGroup_lo_3439 = {dataGroup_lo_hi_3439, dataGroup_lo_lo_3439};
  wire [2047:0] dataGroup_hi_3439 = {dataGroup_hi_hi_3439, dataGroup_hi_lo_3439};
  wire [15:0]   dataGroup_15_71 = dataGroup_lo_3439[2047:2032];
  wire [2047:0] dataGroup_lo_3440 = {dataGroup_lo_hi_3440, dataGroup_lo_lo_3440};
  wire [2047:0] dataGroup_hi_3440 = {dataGroup_hi_hi_3440, dataGroup_hi_lo_3440};
  wire [15:0]   dataGroup_16_71 = dataGroup_hi_3440[127:112];
  wire [2047:0] dataGroup_lo_3441 = {dataGroup_lo_hi_3441, dataGroup_lo_lo_3441};
  wire [2047:0] dataGroup_hi_3441 = {dataGroup_hi_hi_3441, dataGroup_hi_lo_3441};
  wire [15:0]   dataGroup_17_71 = dataGroup_hi_3441[255:240];
  wire [2047:0] dataGroup_lo_3442 = {dataGroup_lo_hi_3442, dataGroup_lo_lo_3442};
  wire [2047:0] dataGroup_hi_3442 = {dataGroup_hi_hi_3442, dataGroup_hi_lo_3442};
  wire [15:0]   dataGroup_18_71 = dataGroup_hi_3442[383:368];
  wire [2047:0] dataGroup_lo_3443 = {dataGroup_lo_hi_3443, dataGroup_lo_lo_3443};
  wire [2047:0] dataGroup_hi_3443 = {dataGroup_hi_hi_3443, dataGroup_hi_lo_3443};
  wire [15:0]   dataGroup_19_71 = dataGroup_hi_3443[511:496];
  wire [2047:0] dataGroup_lo_3444 = {dataGroup_lo_hi_3444, dataGroup_lo_lo_3444};
  wire [2047:0] dataGroup_hi_3444 = {dataGroup_hi_hi_3444, dataGroup_hi_lo_3444};
  wire [15:0]   dataGroup_20_71 = dataGroup_hi_3444[639:624];
  wire [2047:0] dataGroup_lo_3445 = {dataGroup_lo_hi_3445, dataGroup_lo_lo_3445};
  wire [2047:0] dataGroup_hi_3445 = {dataGroup_hi_hi_3445, dataGroup_hi_lo_3445};
  wire [15:0]   dataGroup_21_71 = dataGroup_hi_3445[767:752];
  wire [2047:0] dataGroup_lo_3446 = {dataGroup_lo_hi_3446, dataGroup_lo_lo_3446};
  wire [2047:0] dataGroup_hi_3446 = {dataGroup_hi_hi_3446, dataGroup_hi_lo_3446};
  wire [15:0]   dataGroup_22_71 = dataGroup_hi_3446[895:880];
  wire [2047:0] dataGroup_lo_3447 = {dataGroup_lo_hi_3447, dataGroup_lo_lo_3447};
  wire [2047:0] dataGroup_hi_3447 = {dataGroup_hi_hi_3447, dataGroup_hi_lo_3447};
  wire [15:0]   dataGroup_23_71 = dataGroup_hi_3447[1023:1008];
  wire [2047:0] dataGroup_lo_3448 = {dataGroup_lo_hi_3448, dataGroup_lo_lo_3448};
  wire [2047:0] dataGroup_hi_3448 = {dataGroup_hi_hi_3448, dataGroup_hi_lo_3448};
  wire [15:0]   dataGroup_24_71 = dataGroup_hi_3448[1151:1136];
  wire [2047:0] dataGroup_lo_3449 = {dataGroup_lo_hi_3449, dataGroup_lo_lo_3449};
  wire [2047:0] dataGroup_hi_3449 = {dataGroup_hi_hi_3449, dataGroup_hi_lo_3449};
  wire [15:0]   dataGroup_25_71 = dataGroup_hi_3449[1279:1264];
  wire [2047:0] dataGroup_lo_3450 = {dataGroup_lo_hi_3450, dataGroup_lo_lo_3450};
  wire [2047:0] dataGroup_hi_3450 = {dataGroup_hi_hi_3450, dataGroup_hi_lo_3450};
  wire [15:0]   dataGroup_26_71 = dataGroup_hi_3450[1407:1392];
  wire [2047:0] dataGroup_lo_3451 = {dataGroup_lo_hi_3451, dataGroup_lo_lo_3451};
  wire [2047:0] dataGroup_hi_3451 = {dataGroup_hi_hi_3451, dataGroup_hi_lo_3451};
  wire [15:0]   dataGroup_27_71 = dataGroup_hi_3451[1535:1520];
  wire [2047:0] dataGroup_lo_3452 = {dataGroup_lo_hi_3452, dataGroup_lo_lo_3452};
  wire [2047:0] dataGroup_hi_3452 = {dataGroup_hi_hi_3452, dataGroup_hi_lo_3452};
  wire [15:0]   dataGroup_28_71 = dataGroup_hi_3452[1663:1648];
  wire [2047:0] dataGroup_lo_3453 = {dataGroup_lo_hi_3453, dataGroup_lo_lo_3453};
  wire [2047:0] dataGroup_hi_3453 = {dataGroup_hi_hi_3453, dataGroup_hi_lo_3453};
  wire [15:0]   dataGroup_29_71 = dataGroup_hi_3453[1791:1776];
  wire [2047:0] dataGroup_lo_3454 = {dataGroup_lo_hi_3454, dataGroup_lo_lo_3454};
  wire [2047:0] dataGroup_hi_3454 = {dataGroup_hi_hi_3454, dataGroup_hi_lo_3454};
  wire [15:0]   dataGroup_30_71 = dataGroup_hi_3454[1919:1904];
  wire [2047:0] dataGroup_lo_3455 = {dataGroup_lo_hi_3455, dataGroup_lo_lo_3455};
  wire [2047:0] dataGroup_hi_3455 = {dataGroup_hi_hi_3455, dataGroup_hi_lo_3455};
  wire [15:0]   dataGroup_31_71 = dataGroup_hi_3455[2047:2032];
  wire [31:0]   res_lo_lo_lo_lo_71 = {dataGroup_1_71, dataGroup_0_71};
  wire [31:0]   res_lo_lo_lo_hi_71 = {dataGroup_3_71, dataGroup_2_71};
  wire [63:0]   res_lo_lo_lo_71 = {res_lo_lo_lo_hi_71, res_lo_lo_lo_lo_71};
  wire [31:0]   res_lo_lo_hi_lo_71 = {dataGroup_5_71, dataGroup_4_71};
  wire [31:0]   res_lo_lo_hi_hi_71 = {dataGroup_7_71, dataGroup_6_71};
  wire [63:0]   res_lo_lo_hi_71 = {res_lo_lo_hi_hi_71, res_lo_lo_hi_lo_71};
  wire [127:0]  res_lo_lo_71 = {res_lo_lo_hi_71, res_lo_lo_lo_71};
  wire [31:0]   res_lo_hi_lo_lo_71 = {dataGroup_9_71, dataGroup_8_71};
  wire [31:0]   res_lo_hi_lo_hi_71 = {dataGroup_11_71, dataGroup_10_71};
  wire [63:0]   res_lo_hi_lo_71 = {res_lo_hi_lo_hi_71, res_lo_hi_lo_lo_71};
  wire [31:0]   res_lo_hi_hi_lo_71 = {dataGroup_13_71, dataGroup_12_71};
  wire [31:0]   res_lo_hi_hi_hi_71 = {dataGroup_15_71, dataGroup_14_71};
  wire [63:0]   res_lo_hi_hi_71 = {res_lo_hi_hi_hi_71, res_lo_hi_hi_lo_71};
  wire [127:0]  res_lo_hi_71 = {res_lo_hi_hi_71, res_lo_hi_lo_71};
  wire [255:0]  res_lo_71 = {res_lo_hi_71, res_lo_lo_71};
  wire [31:0]   res_hi_lo_lo_lo_71 = {dataGroup_17_71, dataGroup_16_71};
  wire [31:0]   res_hi_lo_lo_hi_71 = {dataGroup_19_71, dataGroup_18_71};
  wire [63:0]   res_hi_lo_lo_71 = {res_hi_lo_lo_hi_71, res_hi_lo_lo_lo_71};
  wire [31:0]   res_hi_lo_hi_lo_71 = {dataGroup_21_71, dataGroup_20_71};
  wire [31:0]   res_hi_lo_hi_hi_71 = {dataGroup_23_71, dataGroup_22_71};
  wire [63:0]   res_hi_lo_hi_71 = {res_hi_lo_hi_hi_71, res_hi_lo_hi_lo_71};
  wire [127:0]  res_hi_lo_71 = {res_hi_lo_hi_71, res_hi_lo_lo_71};
  wire [31:0]   res_hi_hi_lo_lo_71 = {dataGroup_25_71, dataGroup_24_71};
  wire [31:0]   res_hi_hi_lo_hi_71 = {dataGroup_27_71, dataGroup_26_71};
  wire [63:0]   res_hi_hi_lo_71 = {res_hi_hi_lo_hi_71, res_hi_hi_lo_lo_71};
  wire [31:0]   res_hi_hi_hi_lo_71 = {dataGroup_29_71, dataGroup_28_71};
  wire [31:0]   res_hi_hi_hi_hi_71 = {dataGroup_31_71, dataGroup_30_71};
  wire [63:0]   res_hi_hi_hi_71 = {res_hi_hi_hi_hi_71, res_hi_hi_hi_lo_71};
  wire [127:0]  res_hi_hi_71 = {res_hi_hi_hi_71, res_hi_hi_lo_71};
  wire [255:0]  res_hi_71 = {res_hi_hi_71, res_hi_lo_71};
  wire [511:0]  res_127 = {res_hi_71, res_lo_71};
  wire [1023:0] lo_lo_15 = {res_121, res_120};
  wire [1023:0] lo_hi_15 = {res_123, res_122};
  wire [2047:0] lo_15 = {lo_hi_15, lo_lo_15};
  wire [1023:0] hi_lo_15 = {res_125, res_124};
  wire [1023:0] hi_hi_15 = {res_127, res_126};
  wire [2047:0] hi_15 = {hi_hi_15, hi_lo_15};
  wire [4095:0] regroupLoadData_1_7 = {hi_15, lo_15};
  wire [2047:0] dataGroup_lo_3456 = {dataGroup_lo_hi_3456, dataGroup_lo_lo_3456};
  wire [2047:0] dataGroup_hi_3456 = {dataGroup_hi_hi_3456, dataGroup_hi_lo_3456};
  wire [31:0]   dataGroup_0_72 = dataGroup_lo_3456[31:0];
  wire [2047:0] dataGroup_lo_3457 = {dataGroup_lo_hi_3457, dataGroup_lo_lo_3457};
  wire [2047:0] dataGroup_hi_3457 = {dataGroup_hi_hi_3457, dataGroup_hi_lo_3457};
  wire [31:0]   dataGroup_1_72 = dataGroup_lo_3457[63:32];
  wire [2047:0] dataGroup_lo_3458 = {dataGroup_lo_hi_3458, dataGroup_lo_lo_3458};
  wire [2047:0] dataGroup_hi_3458 = {dataGroup_hi_hi_3458, dataGroup_hi_lo_3458};
  wire [31:0]   dataGroup_2_72 = dataGroup_lo_3458[95:64];
  wire [2047:0] dataGroup_lo_3459 = {dataGroup_lo_hi_3459, dataGroup_lo_lo_3459};
  wire [2047:0] dataGroup_hi_3459 = {dataGroup_hi_hi_3459, dataGroup_hi_lo_3459};
  wire [31:0]   dataGroup_3_72 = dataGroup_lo_3459[127:96];
  wire [2047:0] dataGroup_lo_3460 = {dataGroup_lo_hi_3460, dataGroup_lo_lo_3460};
  wire [2047:0] dataGroup_hi_3460 = {dataGroup_hi_hi_3460, dataGroup_hi_lo_3460};
  wire [31:0]   dataGroup_4_72 = dataGroup_lo_3460[159:128];
  wire [2047:0] dataGroup_lo_3461 = {dataGroup_lo_hi_3461, dataGroup_lo_lo_3461};
  wire [2047:0] dataGroup_hi_3461 = {dataGroup_hi_hi_3461, dataGroup_hi_lo_3461};
  wire [31:0]   dataGroup_5_72 = dataGroup_lo_3461[191:160];
  wire [2047:0] dataGroup_lo_3462 = {dataGroup_lo_hi_3462, dataGroup_lo_lo_3462};
  wire [2047:0] dataGroup_hi_3462 = {dataGroup_hi_hi_3462, dataGroup_hi_lo_3462};
  wire [31:0]   dataGroup_6_72 = dataGroup_lo_3462[223:192];
  wire [2047:0] dataGroup_lo_3463 = {dataGroup_lo_hi_3463, dataGroup_lo_lo_3463};
  wire [2047:0] dataGroup_hi_3463 = {dataGroup_hi_hi_3463, dataGroup_hi_lo_3463};
  wire [31:0]   dataGroup_7_72 = dataGroup_lo_3463[255:224];
  wire [2047:0] dataGroup_lo_3464 = {dataGroup_lo_hi_3464, dataGroup_lo_lo_3464};
  wire [2047:0] dataGroup_hi_3464 = {dataGroup_hi_hi_3464, dataGroup_hi_lo_3464};
  wire [31:0]   dataGroup_8_72 = dataGroup_lo_3464[287:256];
  wire [2047:0] dataGroup_lo_3465 = {dataGroup_lo_hi_3465, dataGroup_lo_lo_3465};
  wire [2047:0] dataGroup_hi_3465 = {dataGroup_hi_hi_3465, dataGroup_hi_lo_3465};
  wire [31:0]   dataGroup_9_72 = dataGroup_lo_3465[319:288];
  wire [2047:0] dataGroup_lo_3466 = {dataGroup_lo_hi_3466, dataGroup_lo_lo_3466};
  wire [2047:0] dataGroup_hi_3466 = {dataGroup_hi_hi_3466, dataGroup_hi_lo_3466};
  wire [31:0]   dataGroup_10_72 = dataGroup_lo_3466[351:320];
  wire [2047:0] dataGroup_lo_3467 = {dataGroup_lo_hi_3467, dataGroup_lo_lo_3467};
  wire [2047:0] dataGroup_hi_3467 = {dataGroup_hi_hi_3467, dataGroup_hi_lo_3467};
  wire [31:0]   dataGroup_11_72 = dataGroup_lo_3467[383:352];
  wire [2047:0] dataGroup_lo_3468 = {dataGroup_lo_hi_3468, dataGroup_lo_lo_3468};
  wire [2047:0] dataGroup_hi_3468 = {dataGroup_hi_hi_3468, dataGroup_hi_lo_3468};
  wire [31:0]   dataGroup_12_72 = dataGroup_lo_3468[415:384];
  wire [2047:0] dataGroup_lo_3469 = {dataGroup_lo_hi_3469, dataGroup_lo_lo_3469};
  wire [2047:0] dataGroup_hi_3469 = {dataGroup_hi_hi_3469, dataGroup_hi_lo_3469};
  wire [31:0]   dataGroup_13_72 = dataGroup_lo_3469[447:416];
  wire [2047:0] dataGroup_lo_3470 = {dataGroup_lo_hi_3470, dataGroup_lo_lo_3470};
  wire [2047:0] dataGroup_hi_3470 = {dataGroup_hi_hi_3470, dataGroup_hi_lo_3470};
  wire [31:0]   dataGroup_14_72 = dataGroup_lo_3470[479:448];
  wire [2047:0] dataGroup_lo_3471 = {dataGroup_lo_hi_3471, dataGroup_lo_lo_3471};
  wire [2047:0] dataGroup_hi_3471 = {dataGroup_hi_hi_3471, dataGroup_hi_lo_3471};
  wire [31:0]   dataGroup_15_72 = dataGroup_lo_3471[511:480];
  wire [63:0]   res_lo_lo_lo_72 = {dataGroup_1_72, dataGroup_0_72};
  wire [63:0]   res_lo_lo_hi_72 = {dataGroup_3_72, dataGroup_2_72};
  wire [127:0]  res_lo_lo_72 = {res_lo_lo_hi_72, res_lo_lo_lo_72};
  wire [63:0]   res_lo_hi_lo_72 = {dataGroup_5_72, dataGroup_4_72};
  wire [63:0]   res_lo_hi_hi_72 = {dataGroup_7_72, dataGroup_6_72};
  wire [127:0]  res_lo_hi_72 = {res_lo_hi_hi_72, res_lo_hi_lo_72};
  wire [255:0]  res_lo_72 = {res_lo_hi_72, res_lo_lo_72};
  wire [63:0]   res_hi_lo_lo_72 = {dataGroup_9_72, dataGroup_8_72};
  wire [63:0]   res_hi_lo_hi_72 = {dataGroup_11_72, dataGroup_10_72};
  wire [127:0]  res_hi_lo_72 = {res_hi_lo_hi_72, res_hi_lo_lo_72};
  wire [63:0]   res_hi_hi_lo_72 = {dataGroup_13_72, dataGroup_12_72};
  wire [63:0]   res_hi_hi_hi_72 = {dataGroup_15_72, dataGroup_14_72};
  wire [127:0]  res_hi_hi_72 = {res_hi_hi_hi_72, res_hi_hi_lo_72};
  wire [255:0]  res_hi_72 = {res_hi_hi_72, res_hi_lo_72};
  wire [511:0]  res_128 = {res_hi_72, res_lo_72};
  wire [1023:0] lo_lo_16 = {512'h0, res_128};
  wire [2047:0] lo_16 = {1024'h0, lo_lo_16};
  wire [4095:0] regroupLoadData_2_0 = {2048'h0, lo_16};
  wire [2047:0] dataGroup_lo_3472 = {dataGroup_lo_hi_3472, dataGroup_lo_lo_3472};
  wire [2047:0] dataGroup_hi_3472 = {dataGroup_hi_hi_3472, dataGroup_hi_lo_3472};
  wire [31:0]   dataGroup_0_73 = dataGroup_lo_3472[31:0];
  wire [2047:0] dataGroup_lo_3473 = {dataGroup_lo_hi_3473, dataGroup_lo_lo_3473};
  wire [2047:0] dataGroup_hi_3473 = {dataGroup_hi_hi_3473, dataGroup_hi_lo_3473};
  wire [31:0]   dataGroup_1_73 = dataGroup_lo_3473[95:64];
  wire [2047:0] dataGroup_lo_3474 = {dataGroup_lo_hi_3474, dataGroup_lo_lo_3474};
  wire [2047:0] dataGroup_hi_3474 = {dataGroup_hi_hi_3474, dataGroup_hi_lo_3474};
  wire [31:0]   dataGroup_2_73 = dataGroup_lo_3474[159:128];
  wire [2047:0] dataGroup_lo_3475 = {dataGroup_lo_hi_3475, dataGroup_lo_lo_3475};
  wire [2047:0] dataGroup_hi_3475 = {dataGroup_hi_hi_3475, dataGroup_hi_lo_3475};
  wire [31:0]   dataGroup_3_73 = dataGroup_lo_3475[223:192];
  wire [2047:0] dataGroup_lo_3476 = {dataGroup_lo_hi_3476, dataGroup_lo_lo_3476};
  wire [2047:0] dataGroup_hi_3476 = {dataGroup_hi_hi_3476, dataGroup_hi_lo_3476};
  wire [31:0]   dataGroup_4_73 = dataGroup_lo_3476[287:256];
  wire [2047:0] dataGroup_lo_3477 = {dataGroup_lo_hi_3477, dataGroup_lo_lo_3477};
  wire [2047:0] dataGroup_hi_3477 = {dataGroup_hi_hi_3477, dataGroup_hi_lo_3477};
  wire [31:0]   dataGroup_5_73 = dataGroup_lo_3477[351:320];
  wire [2047:0] dataGroup_lo_3478 = {dataGroup_lo_hi_3478, dataGroup_lo_lo_3478};
  wire [2047:0] dataGroup_hi_3478 = {dataGroup_hi_hi_3478, dataGroup_hi_lo_3478};
  wire [31:0]   dataGroup_6_73 = dataGroup_lo_3478[415:384];
  wire [2047:0] dataGroup_lo_3479 = {dataGroup_lo_hi_3479, dataGroup_lo_lo_3479};
  wire [2047:0] dataGroup_hi_3479 = {dataGroup_hi_hi_3479, dataGroup_hi_lo_3479};
  wire [31:0]   dataGroup_7_73 = dataGroup_lo_3479[479:448];
  wire [2047:0] dataGroup_lo_3480 = {dataGroup_lo_hi_3480, dataGroup_lo_lo_3480};
  wire [2047:0] dataGroup_hi_3480 = {dataGroup_hi_hi_3480, dataGroup_hi_lo_3480};
  wire [31:0]   dataGroup_8_73 = dataGroup_lo_3480[543:512];
  wire [2047:0] dataGroup_lo_3481 = {dataGroup_lo_hi_3481, dataGroup_lo_lo_3481};
  wire [2047:0] dataGroup_hi_3481 = {dataGroup_hi_hi_3481, dataGroup_hi_lo_3481};
  wire [31:0]   dataGroup_9_73 = dataGroup_lo_3481[607:576];
  wire [2047:0] dataGroup_lo_3482 = {dataGroup_lo_hi_3482, dataGroup_lo_lo_3482};
  wire [2047:0] dataGroup_hi_3482 = {dataGroup_hi_hi_3482, dataGroup_hi_lo_3482};
  wire [31:0]   dataGroup_10_73 = dataGroup_lo_3482[671:640];
  wire [2047:0] dataGroup_lo_3483 = {dataGroup_lo_hi_3483, dataGroup_lo_lo_3483};
  wire [2047:0] dataGroup_hi_3483 = {dataGroup_hi_hi_3483, dataGroup_hi_lo_3483};
  wire [31:0]   dataGroup_11_73 = dataGroup_lo_3483[735:704];
  wire [2047:0] dataGroup_lo_3484 = {dataGroup_lo_hi_3484, dataGroup_lo_lo_3484};
  wire [2047:0] dataGroup_hi_3484 = {dataGroup_hi_hi_3484, dataGroup_hi_lo_3484};
  wire [31:0]   dataGroup_12_73 = dataGroup_lo_3484[799:768];
  wire [2047:0] dataGroup_lo_3485 = {dataGroup_lo_hi_3485, dataGroup_lo_lo_3485};
  wire [2047:0] dataGroup_hi_3485 = {dataGroup_hi_hi_3485, dataGroup_hi_lo_3485};
  wire [31:0]   dataGroup_13_73 = dataGroup_lo_3485[863:832];
  wire [2047:0] dataGroup_lo_3486 = {dataGroup_lo_hi_3486, dataGroup_lo_lo_3486};
  wire [2047:0] dataGroup_hi_3486 = {dataGroup_hi_hi_3486, dataGroup_hi_lo_3486};
  wire [31:0]   dataGroup_14_73 = dataGroup_lo_3486[927:896];
  wire [2047:0] dataGroup_lo_3487 = {dataGroup_lo_hi_3487, dataGroup_lo_lo_3487};
  wire [2047:0] dataGroup_hi_3487 = {dataGroup_hi_hi_3487, dataGroup_hi_lo_3487};
  wire [31:0]   dataGroup_15_73 = dataGroup_lo_3487[991:960];
  wire [63:0]   res_lo_lo_lo_73 = {dataGroup_1_73, dataGroup_0_73};
  wire [63:0]   res_lo_lo_hi_73 = {dataGroup_3_73, dataGroup_2_73};
  wire [127:0]  res_lo_lo_73 = {res_lo_lo_hi_73, res_lo_lo_lo_73};
  wire [63:0]   res_lo_hi_lo_73 = {dataGroup_5_73, dataGroup_4_73};
  wire [63:0]   res_lo_hi_hi_73 = {dataGroup_7_73, dataGroup_6_73};
  wire [127:0]  res_lo_hi_73 = {res_lo_hi_hi_73, res_lo_hi_lo_73};
  wire [255:0]  res_lo_73 = {res_lo_hi_73, res_lo_lo_73};
  wire [63:0]   res_hi_lo_lo_73 = {dataGroup_9_73, dataGroup_8_73};
  wire [63:0]   res_hi_lo_hi_73 = {dataGroup_11_73, dataGroup_10_73};
  wire [127:0]  res_hi_lo_73 = {res_hi_lo_hi_73, res_hi_lo_lo_73};
  wire [63:0]   res_hi_hi_lo_73 = {dataGroup_13_73, dataGroup_12_73};
  wire [63:0]   res_hi_hi_hi_73 = {dataGroup_15_73, dataGroup_14_73};
  wire [127:0]  res_hi_hi_73 = {res_hi_hi_hi_73, res_hi_hi_lo_73};
  wire [255:0]  res_hi_73 = {res_hi_hi_73, res_hi_lo_73};
  wire [511:0]  res_136 = {res_hi_73, res_lo_73};
  wire [2047:0] dataGroup_lo_3488 = {dataGroup_lo_hi_3488, dataGroup_lo_lo_3488};
  wire [2047:0] dataGroup_hi_3488 = {dataGroup_hi_hi_3488, dataGroup_hi_lo_3488};
  wire [31:0]   dataGroup_0_74 = dataGroup_lo_3488[63:32];
  wire [2047:0] dataGroup_lo_3489 = {dataGroup_lo_hi_3489, dataGroup_lo_lo_3489};
  wire [2047:0] dataGroup_hi_3489 = {dataGroup_hi_hi_3489, dataGroup_hi_lo_3489};
  wire [31:0]   dataGroup_1_74 = dataGroup_lo_3489[127:96];
  wire [2047:0] dataGroup_lo_3490 = {dataGroup_lo_hi_3490, dataGroup_lo_lo_3490};
  wire [2047:0] dataGroup_hi_3490 = {dataGroup_hi_hi_3490, dataGroup_hi_lo_3490};
  wire [31:0]   dataGroup_2_74 = dataGroup_lo_3490[191:160];
  wire [2047:0] dataGroup_lo_3491 = {dataGroup_lo_hi_3491, dataGroup_lo_lo_3491};
  wire [2047:0] dataGroup_hi_3491 = {dataGroup_hi_hi_3491, dataGroup_hi_lo_3491};
  wire [31:0]   dataGroup_3_74 = dataGroup_lo_3491[255:224];
  wire [2047:0] dataGroup_lo_3492 = {dataGroup_lo_hi_3492, dataGroup_lo_lo_3492};
  wire [2047:0] dataGroup_hi_3492 = {dataGroup_hi_hi_3492, dataGroup_hi_lo_3492};
  wire [31:0]   dataGroup_4_74 = dataGroup_lo_3492[319:288];
  wire [2047:0] dataGroup_lo_3493 = {dataGroup_lo_hi_3493, dataGroup_lo_lo_3493};
  wire [2047:0] dataGroup_hi_3493 = {dataGroup_hi_hi_3493, dataGroup_hi_lo_3493};
  wire [31:0]   dataGroup_5_74 = dataGroup_lo_3493[383:352];
  wire [2047:0] dataGroup_lo_3494 = {dataGroup_lo_hi_3494, dataGroup_lo_lo_3494};
  wire [2047:0] dataGroup_hi_3494 = {dataGroup_hi_hi_3494, dataGroup_hi_lo_3494};
  wire [31:0]   dataGroup_6_74 = dataGroup_lo_3494[447:416];
  wire [2047:0] dataGroup_lo_3495 = {dataGroup_lo_hi_3495, dataGroup_lo_lo_3495};
  wire [2047:0] dataGroup_hi_3495 = {dataGroup_hi_hi_3495, dataGroup_hi_lo_3495};
  wire [31:0]   dataGroup_7_74 = dataGroup_lo_3495[511:480];
  wire [2047:0] dataGroup_lo_3496 = {dataGroup_lo_hi_3496, dataGroup_lo_lo_3496};
  wire [2047:0] dataGroup_hi_3496 = {dataGroup_hi_hi_3496, dataGroup_hi_lo_3496};
  wire [31:0]   dataGroup_8_74 = dataGroup_lo_3496[575:544];
  wire [2047:0] dataGroup_lo_3497 = {dataGroup_lo_hi_3497, dataGroup_lo_lo_3497};
  wire [2047:0] dataGroup_hi_3497 = {dataGroup_hi_hi_3497, dataGroup_hi_lo_3497};
  wire [31:0]   dataGroup_9_74 = dataGroup_lo_3497[639:608];
  wire [2047:0] dataGroup_lo_3498 = {dataGroup_lo_hi_3498, dataGroup_lo_lo_3498};
  wire [2047:0] dataGroup_hi_3498 = {dataGroup_hi_hi_3498, dataGroup_hi_lo_3498};
  wire [31:0]   dataGroup_10_74 = dataGroup_lo_3498[703:672];
  wire [2047:0] dataGroup_lo_3499 = {dataGroup_lo_hi_3499, dataGroup_lo_lo_3499};
  wire [2047:0] dataGroup_hi_3499 = {dataGroup_hi_hi_3499, dataGroup_hi_lo_3499};
  wire [31:0]   dataGroup_11_74 = dataGroup_lo_3499[767:736];
  wire [2047:0] dataGroup_lo_3500 = {dataGroup_lo_hi_3500, dataGroup_lo_lo_3500};
  wire [2047:0] dataGroup_hi_3500 = {dataGroup_hi_hi_3500, dataGroup_hi_lo_3500};
  wire [31:0]   dataGroup_12_74 = dataGroup_lo_3500[831:800];
  wire [2047:0] dataGroup_lo_3501 = {dataGroup_lo_hi_3501, dataGroup_lo_lo_3501};
  wire [2047:0] dataGroup_hi_3501 = {dataGroup_hi_hi_3501, dataGroup_hi_lo_3501};
  wire [31:0]   dataGroup_13_74 = dataGroup_lo_3501[895:864];
  wire [2047:0] dataGroup_lo_3502 = {dataGroup_lo_hi_3502, dataGroup_lo_lo_3502};
  wire [2047:0] dataGroup_hi_3502 = {dataGroup_hi_hi_3502, dataGroup_hi_lo_3502};
  wire [31:0]   dataGroup_14_74 = dataGroup_lo_3502[959:928];
  wire [2047:0] dataGroup_lo_3503 = {dataGroup_lo_hi_3503, dataGroup_lo_lo_3503};
  wire [2047:0] dataGroup_hi_3503 = {dataGroup_hi_hi_3503, dataGroup_hi_lo_3503};
  wire [31:0]   dataGroup_15_74 = dataGroup_lo_3503[1023:992];
  wire [63:0]   res_lo_lo_lo_74 = {dataGroup_1_74, dataGroup_0_74};
  wire [63:0]   res_lo_lo_hi_74 = {dataGroup_3_74, dataGroup_2_74};
  wire [127:0]  res_lo_lo_74 = {res_lo_lo_hi_74, res_lo_lo_lo_74};
  wire [63:0]   res_lo_hi_lo_74 = {dataGroup_5_74, dataGroup_4_74};
  wire [63:0]   res_lo_hi_hi_74 = {dataGroup_7_74, dataGroup_6_74};
  wire [127:0]  res_lo_hi_74 = {res_lo_hi_hi_74, res_lo_hi_lo_74};
  wire [255:0]  res_lo_74 = {res_lo_hi_74, res_lo_lo_74};
  wire [63:0]   res_hi_lo_lo_74 = {dataGroup_9_74, dataGroup_8_74};
  wire [63:0]   res_hi_lo_hi_74 = {dataGroup_11_74, dataGroup_10_74};
  wire [127:0]  res_hi_lo_74 = {res_hi_lo_hi_74, res_hi_lo_lo_74};
  wire [63:0]   res_hi_hi_lo_74 = {dataGroup_13_74, dataGroup_12_74};
  wire [63:0]   res_hi_hi_hi_74 = {dataGroup_15_74, dataGroup_14_74};
  wire [127:0]  res_hi_hi_74 = {res_hi_hi_hi_74, res_hi_hi_lo_74};
  wire [255:0]  res_hi_74 = {res_hi_hi_74, res_hi_lo_74};
  wire [511:0]  res_137 = {res_hi_74, res_lo_74};
  wire [1023:0] lo_lo_17 = {res_137, res_136};
  wire [2047:0] lo_17 = {1024'h0, lo_lo_17};
  wire [4095:0] regroupLoadData_2_1 = {2048'h0, lo_17};
  wire [2047:0] dataGroup_lo_3504 = {dataGroup_lo_hi_3504, dataGroup_lo_lo_3504};
  wire [2047:0] dataGroup_hi_3504 = {dataGroup_hi_hi_3504, dataGroup_hi_lo_3504};
  wire [31:0]   dataGroup_0_75 = dataGroup_lo_3504[31:0];
  wire [2047:0] dataGroup_lo_3505 = {dataGroup_lo_hi_3505, dataGroup_lo_lo_3505};
  wire [2047:0] dataGroup_hi_3505 = {dataGroup_hi_hi_3505, dataGroup_hi_lo_3505};
  wire [31:0]   dataGroup_1_75 = dataGroup_lo_3505[127:96];
  wire [2047:0] dataGroup_lo_3506 = {dataGroup_lo_hi_3506, dataGroup_lo_lo_3506};
  wire [2047:0] dataGroup_hi_3506 = {dataGroup_hi_hi_3506, dataGroup_hi_lo_3506};
  wire [31:0]   dataGroup_2_75 = dataGroup_lo_3506[223:192];
  wire [2047:0] dataGroup_lo_3507 = {dataGroup_lo_hi_3507, dataGroup_lo_lo_3507};
  wire [2047:0] dataGroup_hi_3507 = {dataGroup_hi_hi_3507, dataGroup_hi_lo_3507};
  wire [31:0]   dataGroup_3_75 = dataGroup_lo_3507[319:288];
  wire [2047:0] dataGroup_lo_3508 = {dataGroup_lo_hi_3508, dataGroup_lo_lo_3508};
  wire [2047:0] dataGroup_hi_3508 = {dataGroup_hi_hi_3508, dataGroup_hi_lo_3508};
  wire [31:0]   dataGroup_4_75 = dataGroup_lo_3508[415:384];
  wire [2047:0] dataGroup_lo_3509 = {dataGroup_lo_hi_3509, dataGroup_lo_lo_3509};
  wire [2047:0] dataGroup_hi_3509 = {dataGroup_hi_hi_3509, dataGroup_hi_lo_3509};
  wire [31:0]   dataGroup_5_75 = dataGroup_lo_3509[511:480];
  wire [2047:0] dataGroup_lo_3510 = {dataGroup_lo_hi_3510, dataGroup_lo_lo_3510};
  wire [2047:0] dataGroup_hi_3510 = {dataGroup_hi_hi_3510, dataGroup_hi_lo_3510};
  wire [31:0]   dataGroup_6_75 = dataGroup_lo_3510[607:576];
  wire [2047:0] dataGroup_lo_3511 = {dataGroup_lo_hi_3511, dataGroup_lo_lo_3511};
  wire [2047:0] dataGroup_hi_3511 = {dataGroup_hi_hi_3511, dataGroup_hi_lo_3511};
  wire [31:0]   dataGroup_7_75 = dataGroup_lo_3511[703:672];
  wire [2047:0] dataGroup_lo_3512 = {dataGroup_lo_hi_3512, dataGroup_lo_lo_3512};
  wire [2047:0] dataGroup_hi_3512 = {dataGroup_hi_hi_3512, dataGroup_hi_lo_3512};
  wire [31:0]   dataGroup_8_75 = dataGroup_lo_3512[799:768];
  wire [2047:0] dataGroup_lo_3513 = {dataGroup_lo_hi_3513, dataGroup_lo_lo_3513};
  wire [2047:0] dataGroup_hi_3513 = {dataGroup_hi_hi_3513, dataGroup_hi_lo_3513};
  wire [31:0]   dataGroup_9_75 = dataGroup_lo_3513[895:864];
  wire [2047:0] dataGroup_lo_3514 = {dataGroup_lo_hi_3514, dataGroup_lo_lo_3514};
  wire [2047:0] dataGroup_hi_3514 = {dataGroup_hi_hi_3514, dataGroup_hi_lo_3514};
  wire [31:0]   dataGroup_10_75 = dataGroup_lo_3514[991:960];
  wire [2047:0] dataGroup_lo_3515 = {dataGroup_lo_hi_3515, dataGroup_lo_lo_3515};
  wire [2047:0] dataGroup_hi_3515 = {dataGroup_hi_hi_3515, dataGroup_hi_lo_3515};
  wire [31:0]   dataGroup_11_75 = dataGroup_lo_3515[1087:1056];
  wire [2047:0] dataGroup_lo_3516 = {dataGroup_lo_hi_3516, dataGroup_lo_lo_3516};
  wire [2047:0] dataGroup_hi_3516 = {dataGroup_hi_hi_3516, dataGroup_hi_lo_3516};
  wire [31:0]   dataGroup_12_75 = dataGroup_lo_3516[1183:1152];
  wire [2047:0] dataGroup_lo_3517 = {dataGroup_lo_hi_3517, dataGroup_lo_lo_3517};
  wire [2047:0] dataGroup_hi_3517 = {dataGroup_hi_hi_3517, dataGroup_hi_lo_3517};
  wire [31:0]   dataGroup_13_75 = dataGroup_lo_3517[1279:1248];
  wire [2047:0] dataGroup_lo_3518 = {dataGroup_lo_hi_3518, dataGroup_lo_lo_3518};
  wire [2047:0] dataGroup_hi_3518 = {dataGroup_hi_hi_3518, dataGroup_hi_lo_3518};
  wire [31:0]   dataGroup_14_75 = dataGroup_lo_3518[1375:1344];
  wire [2047:0] dataGroup_lo_3519 = {dataGroup_lo_hi_3519, dataGroup_lo_lo_3519};
  wire [2047:0] dataGroup_hi_3519 = {dataGroup_hi_hi_3519, dataGroup_hi_lo_3519};
  wire [31:0]   dataGroup_15_75 = dataGroup_lo_3519[1471:1440];
  wire [63:0]   res_lo_lo_lo_75 = {dataGroup_1_75, dataGroup_0_75};
  wire [63:0]   res_lo_lo_hi_75 = {dataGroup_3_75, dataGroup_2_75};
  wire [127:0]  res_lo_lo_75 = {res_lo_lo_hi_75, res_lo_lo_lo_75};
  wire [63:0]   res_lo_hi_lo_75 = {dataGroup_5_75, dataGroup_4_75};
  wire [63:0]   res_lo_hi_hi_75 = {dataGroup_7_75, dataGroup_6_75};
  wire [127:0]  res_lo_hi_75 = {res_lo_hi_hi_75, res_lo_hi_lo_75};
  wire [255:0]  res_lo_75 = {res_lo_hi_75, res_lo_lo_75};
  wire [63:0]   res_hi_lo_lo_75 = {dataGroup_9_75, dataGroup_8_75};
  wire [63:0]   res_hi_lo_hi_75 = {dataGroup_11_75, dataGroup_10_75};
  wire [127:0]  res_hi_lo_75 = {res_hi_lo_hi_75, res_hi_lo_lo_75};
  wire [63:0]   res_hi_hi_lo_75 = {dataGroup_13_75, dataGroup_12_75};
  wire [63:0]   res_hi_hi_hi_75 = {dataGroup_15_75, dataGroup_14_75};
  wire [127:0]  res_hi_hi_75 = {res_hi_hi_hi_75, res_hi_hi_lo_75};
  wire [255:0]  res_hi_75 = {res_hi_hi_75, res_hi_lo_75};
  wire [511:0]  res_144 = {res_hi_75, res_lo_75};
  wire [2047:0] dataGroup_lo_3520 = {dataGroup_lo_hi_3520, dataGroup_lo_lo_3520};
  wire [2047:0] dataGroup_hi_3520 = {dataGroup_hi_hi_3520, dataGroup_hi_lo_3520};
  wire [31:0]   dataGroup_0_76 = dataGroup_lo_3520[63:32];
  wire [2047:0] dataGroup_lo_3521 = {dataGroup_lo_hi_3521, dataGroup_lo_lo_3521};
  wire [2047:0] dataGroup_hi_3521 = {dataGroup_hi_hi_3521, dataGroup_hi_lo_3521};
  wire [31:0]   dataGroup_1_76 = dataGroup_lo_3521[159:128];
  wire [2047:0] dataGroup_lo_3522 = {dataGroup_lo_hi_3522, dataGroup_lo_lo_3522};
  wire [2047:0] dataGroup_hi_3522 = {dataGroup_hi_hi_3522, dataGroup_hi_lo_3522};
  wire [31:0]   dataGroup_2_76 = dataGroup_lo_3522[255:224];
  wire [2047:0] dataGroup_lo_3523 = {dataGroup_lo_hi_3523, dataGroup_lo_lo_3523};
  wire [2047:0] dataGroup_hi_3523 = {dataGroup_hi_hi_3523, dataGroup_hi_lo_3523};
  wire [31:0]   dataGroup_3_76 = dataGroup_lo_3523[351:320];
  wire [2047:0] dataGroup_lo_3524 = {dataGroup_lo_hi_3524, dataGroup_lo_lo_3524};
  wire [2047:0] dataGroup_hi_3524 = {dataGroup_hi_hi_3524, dataGroup_hi_lo_3524};
  wire [31:0]   dataGroup_4_76 = dataGroup_lo_3524[447:416];
  wire [2047:0] dataGroup_lo_3525 = {dataGroup_lo_hi_3525, dataGroup_lo_lo_3525};
  wire [2047:0] dataGroup_hi_3525 = {dataGroup_hi_hi_3525, dataGroup_hi_lo_3525};
  wire [31:0]   dataGroup_5_76 = dataGroup_lo_3525[543:512];
  wire [2047:0] dataGroup_lo_3526 = {dataGroup_lo_hi_3526, dataGroup_lo_lo_3526};
  wire [2047:0] dataGroup_hi_3526 = {dataGroup_hi_hi_3526, dataGroup_hi_lo_3526};
  wire [31:0]   dataGroup_6_76 = dataGroup_lo_3526[639:608];
  wire [2047:0] dataGroup_lo_3527 = {dataGroup_lo_hi_3527, dataGroup_lo_lo_3527};
  wire [2047:0] dataGroup_hi_3527 = {dataGroup_hi_hi_3527, dataGroup_hi_lo_3527};
  wire [31:0]   dataGroup_7_76 = dataGroup_lo_3527[735:704];
  wire [2047:0] dataGroup_lo_3528 = {dataGroup_lo_hi_3528, dataGroup_lo_lo_3528};
  wire [2047:0] dataGroup_hi_3528 = {dataGroup_hi_hi_3528, dataGroup_hi_lo_3528};
  wire [31:0]   dataGroup_8_76 = dataGroup_lo_3528[831:800];
  wire [2047:0] dataGroup_lo_3529 = {dataGroup_lo_hi_3529, dataGroup_lo_lo_3529};
  wire [2047:0] dataGroup_hi_3529 = {dataGroup_hi_hi_3529, dataGroup_hi_lo_3529};
  wire [31:0]   dataGroup_9_76 = dataGroup_lo_3529[927:896];
  wire [2047:0] dataGroup_lo_3530 = {dataGroup_lo_hi_3530, dataGroup_lo_lo_3530};
  wire [2047:0] dataGroup_hi_3530 = {dataGroup_hi_hi_3530, dataGroup_hi_lo_3530};
  wire [31:0]   dataGroup_10_76 = dataGroup_lo_3530[1023:992];
  wire [2047:0] dataGroup_lo_3531 = {dataGroup_lo_hi_3531, dataGroup_lo_lo_3531};
  wire [2047:0] dataGroup_hi_3531 = {dataGroup_hi_hi_3531, dataGroup_hi_lo_3531};
  wire [31:0]   dataGroup_11_76 = dataGroup_lo_3531[1119:1088];
  wire [2047:0] dataGroup_lo_3532 = {dataGroup_lo_hi_3532, dataGroup_lo_lo_3532};
  wire [2047:0] dataGroup_hi_3532 = {dataGroup_hi_hi_3532, dataGroup_hi_lo_3532};
  wire [31:0]   dataGroup_12_76 = dataGroup_lo_3532[1215:1184];
  wire [2047:0] dataGroup_lo_3533 = {dataGroup_lo_hi_3533, dataGroup_lo_lo_3533};
  wire [2047:0] dataGroup_hi_3533 = {dataGroup_hi_hi_3533, dataGroup_hi_lo_3533};
  wire [31:0]   dataGroup_13_76 = dataGroup_lo_3533[1311:1280];
  wire [2047:0] dataGroup_lo_3534 = {dataGroup_lo_hi_3534, dataGroup_lo_lo_3534};
  wire [2047:0] dataGroup_hi_3534 = {dataGroup_hi_hi_3534, dataGroup_hi_lo_3534};
  wire [31:0]   dataGroup_14_76 = dataGroup_lo_3534[1407:1376];
  wire [2047:0] dataGroup_lo_3535 = {dataGroup_lo_hi_3535, dataGroup_lo_lo_3535};
  wire [2047:0] dataGroup_hi_3535 = {dataGroup_hi_hi_3535, dataGroup_hi_lo_3535};
  wire [31:0]   dataGroup_15_76 = dataGroup_lo_3535[1503:1472];
  wire [63:0]   res_lo_lo_lo_76 = {dataGroup_1_76, dataGroup_0_76};
  wire [63:0]   res_lo_lo_hi_76 = {dataGroup_3_76, dataGroup_2_76};
  wire [127:0]  res_lo_lo_76 = {res_lo_lo_hi_76, res_lo_lo_lo_76};
  wire [63:0]   res_lo_hi_lo_76 = {dataGroup_5_76, dataGroup_4_76};
  wire [63:0]   res_lo_hi_hi_76 = {dataGroup_7_76, dataGroup_6_76};
  wire [127:0]  res_lo_hi_76 = {res_lo_hi_hi_76, res_lo_hi_lo_76};
  wire [255:0]  res_lo_76 = {res_lo_hi_76, res_lo_lo_76};
  wire [63:0]   res_hi_lo_lo_76 = {dataGroup_9_76, dataGroup_8_76};
  wire [63:0]   res_hi_lo_hi_76 = {dataGroup_11_76, dataGroup_10_76};
  wire [127:0]  res_hi_lo_76 = {res_hi_lo_hi_76, res_hi_lo_lo_76};
  wire [63:0]   res_hi_hi_lo_76 = {dataGroup_13_76, dataGroup_12_76};
  wire [63:0]   res_hi_hi_hi_76 = {dataGroup_15_76, dataGroup_14_76};
  wire [127:0]  res_hi_hi_76 = {res_hi_hi_hi_76, res_hi_hi_lo_76};
  wire [255:0]  res_hi_76 = {res_hi_hi_76, res_hi_lo_76};
  wire [511:0]  res_145 = {res_hi_76, res_lo_76};
  wire [2047:0] dataGroup_lo_3536 = {dataGroup_lo_hi_3536, dataGroup_lo_lo_3536};
  wire [2047:0] dataGroup_hi_3536 = {dataGroup_hi_hi_3536, dataGroup_hi_lo_3536};
  wire [31:0]   dataGroup_0_77 = dataGroup_lo_3536[95:64];
  wire [2047:0] dataGroup_lo_3537 = {dataGroup_lo_hi_3537, dataGroup_lo_lo_3537};
  wire [2047:0] dataGroup_hi_3537 = {dataGroup_hi_hi_3537, dataGroup_hi_lo_3537};
  wire [31:0]   dataGroup_1_77 = dataGroup_lo_3537[191:160];
  wire [2047:0] dataGroup_lo_3538 = {dataGroup_lo_hi_3538, dataGroup_lo_lo_3538};
  wire [2047:0] dataGroup_hi_3538 = {dataGroup_hi_hi_3538, dataGroup_hi_lo_3538};
  wire [31:0]   dataGroup_2_77 = dataGroup_lo_3538[287:256];
  wire [2047:0] dataGroup_lo_3539 = {dataGroup_lo_hi_3539, dataGroup_lo_lo_3539};
  wire [2047:0] dataGroup_hi_3539 = {dataGroup_hi_hi_3539, dataGroup_hi_lo_3539};
  wire [31:0]   dataGroup_3_77 = dataGroup_lo_3539[383:352];
  wire [2047:0] dataGroup_lo_3540 = {dataGroup_lo_hi_3540, dataGroup_lo_lo_3540};
  wire [2047:0] dataGroup_hi_3540 = {dataGroup_hi_hi_3540, dataGroup_hi_lo_3540};
  wire [31:0]   dataGroup_4_77 = dataGroup_lo_3540[479:448];
  wire [2047:0] dataGroup_lo_3541 = {dataGroup_lo_hi_3541, dataGroup_lo_lo_3541};
  wire [2047:0] dataGroup_hi_3541 = {dataGroup_hi_hi_3541, dataGroup_hi_lo_3541};
  wire [31:0]   dataGroup_5_77 = dataGroup_lo_3541[575:544];
  wire [2047:0] dataGroup_lo_3542 = {dataGroup_lo_hi_3542, dataGroup_lo_lo_3542};
  wire [2047:0] dataGroup_hi_3542 = {dataGroup_hi_hi_3542, dataGroup_hi_lo_3542};
  wire [31:0]   dataGroup_6_77 = dataGroup_lo_3542[671:640];
  wire [2047:0] dataGroup_lo_3543 = {dataGroup_lo_hi_3543, dataGroup_lo_lo_3543};
  wire [2047:0] dataGroup_hi_3543 = {dataGroup_hi_hi_3543, dataGroup_hi_lo_3543};
  wire [31:0]   dataGroup_7_77 = dataGroup_lo_3543[767:736];
  wire [2047:0] dataGroup_lo_3544 = {dataGroup_lo_hi_3544, dataGroup_lo_lo_3544};
  wire [2047:0] dataGroup_hi_3544 = {dataGroup_hi_hi_3544, dataGroup_hi_lo_3544};
  wire [31:0]   dataGroup_8_77 = dataGroup_lo_3544[863:832];
  wire [2047:0] dataGroup_lo_3545 = {dataGroup_lo_hi_3545, dataGroup_lo_lo_3545};
  wire [2047:0] dataGroup_hi_3545 = {dataGroup_hi_hi_3545, dataGroup_hi_lo_3545};
  wire [31:0]   dataGroup_9_77 = dataGroup_lo_3545[959:928];
  wire [2047:0] dataGroup_lo_3546 = {dataGroup_lo_hi_3546, dataGroup_lo_lo_3546};
  wire [2047:0] dataGroup_hi_3546 = {dataGroup_hi_hi_3546, dataGroup_hi_lo_3546};
  wire [31:0]   dataGroup_10_77 = dataGroup_lo_3546[1055:1024];
  wire [2047:0] dataGroup_lo_3547 = {dataGroup_lo_hi_3547, dataGroup_lo_lo_3547};
  wire [2047:0] dataGroup_hi_3547 = {dataGroup_hi_hi_3547, dataGroup_hi_lo_3547};
  wire [31:0]   dataGroup_11_77 = dataGroup_lo_3547[1151:1120];
  wire [2047:0] dataGroup_lo_3548 = {dataGroup_lo_hi_3548, dataGroup_lo_lo_3548};
  wire [2047:0] dataGroup_hi_3548 = {dataGroup_hi_hi_3548, dataGroup_hi_lo_3548};
  wire [31:0]   dataGroup_12_77 = dataGroup_lo_3548[1247:1216];
  wire [2047:0] dataGroup_lo_3549 = {dataGroup_lo_hi_3549, dataGroup_lo_lo_3549};
  wire [2047:0] dataGroup_hi_3549 = {dataGroup_hi_hi_3549, dataGroup_hi_lo_3549};
  wire [31:0]   dataGroup_13_77 = dataGroup_lo_3549[1343:1312];
  wire [2047:0] dataGroup_lo_3550 = {dataGroup_lo_hi_3550, dataGroup_lo_lo_3550};
  wire [2047:0] dataGroup_hi_3550 = {dataGroup_hi_hi_3550, dataGroup_hi_lo_3550};
  wire [31:0]   dataGroup_14_77 = dataGroup_lo_3550[1439:1408];
  wire [2047:0] dataGroup_lo_3551 = {dataGroup_lo_hi_3551, dataGroup_lo_lo_3551};
  wire [2047:0] dataGroup_hi_3551 = {dataGroup_hi_hi_3551, dataGroup_hi_lo_3551};
  wire [31:0]   dataGroup_15_77 = dataGroup_lo_3551[1535:1504];
  wire [63:0]   res_lo_lo_lo_77 = {dataGroup_1_77, dataGroup_0_77};
  wire [63:0]   res_lo_lo_hi_77 = {dataGroup_3_77, dataGroup_2_77};
  wire [127:0]  res_lo_lo_77 = {res_lo_lo_hi_77, res_lo_lo_lo_77};
  wire [63:0]   res_lo_hi_lo_77 = {dataGroup_5_77, dataGroup_4_77};
  wire [63:0]   res_lo_hi_hi_77 = {dataGroup_7_77, dataGroup_6_77};
  wire [127:0]  res_lo_hi_77 = {res_lo_hi_hi_77, res_lo_hi_lo_77};
  wire [255:0]  res_lo_77 = {res_lo_hi_77, res_lo_lo_77};
  wire [63:0]   res_hi_lo_lo_77 = {dataGroup_9_77, dataGroup_8_77};
  wire [63:0]   res_hi_lo_hi_77 = {dataGroup_11_77, dataGroup_10_77};
  wire [127:0]  res_hi_lo_77 = {res_hi_lo_hi_77, res_hi_lo_lo_77};
  wire [63:0]   res_hi_hi_lo_77 = {dataGroup_13_77, dataGroup_12_77};
  wire [63:0]   res_hi_hi_hi_77 = {dataGroup_15_77, dataGroup_14_77};
  wire [127:0]  res_hi_hi_77 = {res_hi_hi_hi_77, res_hi_hi_lo_77};
  wire [255:0]  res_hi_77 = {res_hi_hi_77, res_hi_lo_77};
  wire [511:0]  res_146 = {res_hi_77, res_lo_77};
  wire [1023:0] lo_lo_18 = {res_145, res_144};
  wire [1023:0] lo_hi_18 = {512'h0, res_146};
  wire [2047:0] lo_18 = {lo_hi_18, lo_lo_18};
  wire [4095:0] regroupLoadData_2_2 = {2048'h0, lo_18};
  wire [2047:0] dataGroup_lo_3552 = {dataGroup_lo_hi_3552, dataGroup_lo_lo_3552};
  wire [2047:0] dataGroup_hi_3552 = {dataGroup_hi_hi_3552, dataGroup_hi_lo_3552};
  wire [31:0]   dataGroup_0_78 = dataGroup_lo_3552[31:0];
  wire [2047:0] dataGroup_lo_3553 = {dataGroup_lo_hi_3553, dataGroup_lo_lo_3553};
  wire [2047:0] dataGroup_hi_3553 = {dataGroup_hi_hi_3553, dataGroup_hi_lo_3553};
  wire [31:0]   dataGroup_1_78 = dataGroup_lo_3553[159:128];
  wire [2047:0] dataGroup_lo_3554 = {dataGroup_lo_hi_3554, dataGroup_lo_lo_3554};
  wire [2047:0] dataGroup_hi_3554 = {dataGroup_hi_hi_3554, dataGroup_hi_lo_3554};
  wire [31:0]   dataGroup_2_78 = dataGroup_lo_3554[287:256];
  wire [2047:0] dataGroup_lo_3555 = {dataGroup_lo_hi_3555, dataGroup_lo_lo_3555};
  wire [2047:0] dataGroup_hi_3555 = {dataGroup_hi_hi_3555, dataGroup_hi_lo_3555};
  wire [31:0]   dataGroup_3_78 = dataGroup_lo_3555[415:384];
  wire [2047:0] dataGroup_lo_3556 = {dataGroup_lo_hi_3556, dataGroup_lo_lo_3556};
  wire [2047:0] dataGroup_hi_3556 = {dataGroup_hi_hi_3556, dataGroup_hi_lo_3556};
  wire [31:0]   dataGroup_4_78 = dataGroup_lo_3556[543:512];
  wire [2047:0] dataGroup_lo_3557 = {dataGroup_lo_hi_3557, dataGroup_lo_lo_3557};
  wire [2047:0] dataGroup_hi_3557 = {dataGroup_hi_hi_3557, dataGroup_hi_lo_3557};
  wire [31:0]   dataGroup_5_78 = dataGroup_lo_3557[671:640];
  wire [2047:0] dataGroup_lo_3558 = {dataGroup_lo_hi_3558, dataGroup_lo_lo_3558};
  wire [2047:0] dataGroup_hi_3558 = {dataGroup_hi_hi_3558, dataGroup_hi_lo_3558};
  wire [31:0]   dataGroup_6_78 = dataGroup_lo_3558[799:768];
  wire [2047:0] dataGroup_lo_3559 = {dataGroup_lo_hi_3559, dataGroup_lo_lo_3559};
  wire [2047:0] dataGroup_hi_3559 = {dataGroup_hi_hi_3559, dataGroup_hi_lo_3559};
  wire [31:0]   dataGroup_7_78 = dataGroup_lo_3559[927:896];
  wire [2047:0] dataGroup_lo_3560 = {dataGroup_lo_hi_3560, dataGroup_lo_lo_3560};
  wire [2047:0] dataGroup_hi_3560 = {dataGroup_hi_hi_3560, dataGroup_hi_lo_3560};
  wire [31:0]   dataGroup_8_78 = dataGroup_lo_3560[1055:1024];
  wire [2047:0] dataGroup_lo_3561 = {dataGroup_lo_hi_3561, dataGroup_lo_lo_3561};
  wire [2047:0] dataGroup_hi_3561 = {dataGroup_hi_hi_3561, dataGroup_hi_lo_3561};
  wire [31:0]   dataGroup_9_78 = dataGroup_lo_3561[1183:1152];
  wire [2047:0] dataGroup_lo_3562 = {dataGroup_lo_hi_3562, dataGroup_lo_lo_3562};
  wire [2047:0] dataGroup_hi_3562 = {dataGroup_hi_hi_3562, dataGroup_hi_lo_3562};
  wire [31:0]   dataGroup_10_78 = dataGroup_lo_3562[1311:1280];
  wire [2047:0] dataGroup_lo_3563 = {dataGroup_lo_hi_3563, dataGroup_lo_lo_3563};
  wire [2047:0] dataGroup_hi_3563 = {dataGroup_hi_hi_3563, dataGroup_hi_lo_3563};
  wire [31:0]   dataGroup_11_78 = dataGroup_lo_3563[1439:1408];
  wire [2047:0] dataGroup_lo_3564 = {dataGroup_lo_hi_3564, dataGroup_lo_lo_3564};
  wire [2047:0] dataGroup_hi_3564 = {dataGroup_hi_hi_3564, dataGroup_hi_lo_3564};
  wire [31:0]   dataGroup_12_78 = dataGroup_lo_3564[1567:1536];
  wire [2047:0] dataGroup_lo_3565 = {dataGroup_lo_hi_3565, dataGroup_lo_lo_3565};
  wire [2047:0] dataGroup_hi_3565 = {dataGroup_hi_hi_3565, dataGroup_hi_lo_3565};
  wire [31:0]   dataGroup_13_78 = dataGroup_lo_3565[1695:1664];
  wire [2047:0] dataGroup_lo_3566 = {dataGroup_lo_hi_3566, dataGroup_lo_lo_3566};
  wire [2047:0] dataGroup_hi_3566 = {dataGroup_hi_hi_3566, dataGroup_hi_lo_3566};
  wire [31:0]   dataGroup_14_78 = dataGroup_lo_3566[1823:1792];
  wire [2047:0] dataGroup_lo_3567 = {dataGroup_lo_hi_3567, dataGroup_lo_lo_3567};
  wire [2047:0] dataGroup_hi_3567 = {dataGroup_hi_hi_3567, dataGroup_hi_lo_3567};
  wire [31:0]   dataGroup_15_78 = dataGroup_lo_3567[1951:1920];
  wire [63:0]   res_lo_lo_lo_78 = {dataGroup_1_78, dataGroup_0_78};
  wire [63:0]   res_lo_lo_hi_78 = {dataGroup_3_78, dataGroup_2_78};
  wire [127:0]  res_lo_lo_78 = {res_lo_lo_hi_78, res_lo_lo_lo_78};
  wire [63:0]   res_lo_hi_lo_78 = {dataGroup_5_78, dataGroup_4_78};
  wire [63:0]   res_lo_hi_hi_78 = {dataGroup_7_78, dataGroup_6_78};
  wire [127:0]  res_lo_hi_78 = {res_lo_hi_hi_78, res_lo_hi_lo_78};
  wire [255:0]  res_lo_78 = {res_lo_hi_78, res_lo_lo_78};
  wire [63:0]   res_hi_lo_lo_78 = {dataGroup_9_78, dataGroup_8_78};
  wire [63:0]   res_hi_lo_hi_78 = {dataGroup_11_78, dataGroup_10_78};
  wire [127:0]  res_hi_lo_78 = {res_hi_lo_hi_78, res_hi_lo_lo_78};
  wire [63:0]   res_hi_hi_lo_78 = {dataGroup_13_78, dataGroup_12_78};
  wire [63:0]   res_hi_hi_hi_78 = {dataGroup_15_78, dataGroup_14_78};
  wire [127:0]  res_hi_hi_78 = {res_hi_hi_hi_78, res_hi_hi_lo_78};
  wire [255:0]  res_hi_78 = {res_hi_hi_78, res_hi_lo_78};
  wire [511:0]  res_152 = {res_hi_78, res_lo_78};
  wire [2047:0] dataGroup_lo_3568 = {dataGroup_lo_hi_3568, dataGroup_lo_lo_3568};
  wire [2047:0] dataGroup_hi_3568 = {dataGroup_hi_hi_3568, dataGroup_hi_lo_3568};
  wire [31:0]   dataGroup_0_79 = dataGroup_lo_3568[63:32];
  wire [2047:0] dataGroup_lo_3569 = {dataGroup_lo_hi_3569, dataGroup_lo_lo_3569};
  wire [2047:0] dataGroup_hi_3569 = {dataGroup_hi_hi_3569, dataGroup_hi_lo_3569};
  wire [31:0]   dataGroup_1_79 = dataGroup_lo_3569[191:160];
  wire [2047:0] dataGroup_lo_3570 = {dataGroup_lo_hi_3570, dataGroup_lo_lo_3570};
  wire [2047:0] dataGroup_hi_3570 = {dataGroup_hi_hi_3570, dataGroup_hi_lo_3570};
  wire [31:0]   dataGroup_2_79 = dataGroup_lo_3570[319:288];
  wire [2047:0] dataGroup_lo_3571 = {dataGroup_lo_hi_3571, dataGroup_lo_lo_3571};
  wire [2047:0] dataGroup_hi_3571 = {dataGroup_hi_hi_3571, dataGroup_hi_lo_3571};
  wire [31:0]   dataGroup_3_79 = dataGroup_lo_3571[447:416];
  wire [2047:0] dataGroup_lo_3572 = {dataGroup_lo_hi_3572, dataGroup_lo_lo_3572};
  wire [2047:0] dataGroup_hi_3572 = {dataGroup_hi_hi_3572, dataGroup_hi_lo_3572};
  wire [31:0]   dataGroup_4_79 = dataGroup_lo_3572[575:544];
  wire [2047:0] dataGroup_lo_3573 = {dataGroup_lo_hi_3573, dataGroup_lo_lo_3573};
  wire [2047:0] dataGroup_hi_3573 = {dataGroup_hi_hi_3573, dataGroup_hi_lo_3573};
  wire [31:0]   dataGroup_5_79 = dataGroup_lo_3573[703:672];
  wire [2047:0] dataGroup_lo_3574 = {dataGroup_lo_hi_3574, dataGroup_lo_lo_3574};
  wire [2047:0] dataGroup_hi_3574 = {dataGroup_hi_hi_3574, dataGroup_hi_lo_3574};
  wire [31:0]   dataGroup_6_79 = dataGroup_lo_3574[831:800];
  wire [2047:0] dataGroup_lo_3575 = {dataGroup_lo_hi_3575, dataGroup_lo_lo_3575};
  wire [2047:0] dataGroup_hi_3575 = {dataGroup_hi_hi_3575, dataGroup_hi_lo_3575};
  wire [31:0]   dataGroup_7_79 = dataGroup_lo_3575[959:928];
  wire [2047:0] dataGroup_lo_3576 = {dataGroup_lo_hi_3576, dataGroup_lo_lo_3576};
  wire [2047:0] dataGroup_hi_3576 = {dataGroup_hi_hi_3576, dataGroup_hi_lo_3576};
  wire [31:0]   dataGroup_8_79 = dataGroup_lo_3576[1087:1056];
  wire [2047:0] dataGroup_lo_3577 = {dataGroup_lo_hi_3577, dataGroup_lo_lo_3577};
  wire [2047:0] dataGroup_hi_3577 = {dataGroup_hi_hi_3577, dataGroup_hi_lo_3577};
  wire [31:0]   dataGroup_9_79 = dataGroup_lo_3577[1215:1184];
  wire [2047:0] dataGroup_lo_3578 = {dataGroup_lo_hi_3578, dataGroup_lo_lo_3578};
  wire [2047:0] dataGroup_hi_3578 = {dataGroup_hi_hi_3578, dataGroup_hi_lo_3578};
  wire [31:0]   dataGroup_10_79 = dataGroup_lo_3578[1343:1312];
  wire [2047:0] dataGroup_lo_3579 = {dataGroup_lo_hi_3579, dataGroup_lo_lo_3579};
  wire [2047:0] dataGroup_hi_3579 = {dataGroup_hi_hi_3579, dataGroup_hi_lo_3579};
  wire [31:0]   dataGroup_11_79 = dataGroup_lo_3579[1471:1440];
  wire [2047:0] dataGroup_lo_3580 = {dataGroup_lo_hi_3580, dataGroup_lo_lo_3580};
  wire [2047:0] dataGroup_hi_3580 = {dataGroup_hi_hi_3580, dataGroup_hi_lo_3580};
  wire [31:0]   dataGroup_12_79 = dataGroup_lo_3580[1599:1568];
  wire [2047:0] dataGroup_lo_3581 = {dataGroup_lo_hi_3581, dataGroup_lo_lo_3581};
  wire [2047:0] dataGroup_hi_3581 = {dataGroup_hi_hi_3581, dataGroup_hi_lo_3581};
  wire [31:0]   dataGroup_13_79 = dataGroup_lo_3581[1727:1696];
  wire [2047:0] dataGroup_lo_3582 = {dataGroup_lo_hi_3582, dataGroup_lo_lo_3582};
  wire [2047:0] dataGroup_hi_3582 = {dataGroup_hi_hi_3582, dataGroup_hi_lo_3582};
  wire [31:0]   dataGroup_14_79 = dataGroup_lo_3582[1855:1824];
  wire [2047:0] dataGroup_lo_3583 = {dataGroup_lo_hi_3583, dataGroup_lo_lo_3583};
  wire [2047:0] dataGroup_hi_3583 = {dataGroup_hi_hi_3583, dataGroup_hi_lo_3583};
  wire [31:0]   dataGroup_15_79 = dataGroup_lo_3583[1983:1952];
  wire [63:0]   res_lo_lo_lo_79 = {dataGroup_1_79, dataGroup_0_79};
  wire [63:0]   res_lo_lo_hi_79 = {dataGroup_3_79, dataGroup_2_79};
  wire [127:0]  res_lo_lo_79 = {res_lo_lo_hi_79, res_lo_lo_lo_79};
  wire [63:0]   res_lo_hi_lo_79 = {dataGroup_5_79, dataGroup_4_79};
  wire [63:0]   res_lo_hi_hi_79 = {dataGroup_7_79, dataGroup_6_79};
  wire [127:0]  res_lo_hi_79 = {res_lo_hi_hi_79, res_lo_hi_lo_79};
  wire [255:0]  res_lo_79 = {res_lo_hi_79, res_lo_lo_79};
  wire [63:0]   res_hi_lo_lo_79 = {dataGroup_9_79, dataGroup_8_79};
  wire [63:0]   res_hi_lo_hi_79 = {dataGroup_11_79, dataGroup_10_79};
  wire [127:0]  res_hi_lo_79 = {res_hi_lo_hi_79, res_hi_lo_lo_79};
  wire [63:0]   res_hi_hi_lo_79 = {dataGroup_13_79, dataGroup_12_79};
  wire [63:0]   res_hi_hi_hi_79 = {dataGroup_15_79, dataGroup_14_79};
  wire [127:0]  res_hi_hi_79 = {res_hi_hi_hi_79, res_hi_hi_lo_79};
  wire [255:0]  res_hi_79 = {res_hi_hi_79, res_hi_lo_79};
  wire [511:0]  res_153 = {res_hi_79, res_lo_79};
  wire [2047:0] dataGroup_lo_3584 = {dataGroup_lo_hi_3584, dataGroup_lo_lo_3584};
  wire [2047:0] dataGroup_hi_3584 = {dataGroup_hi_hi_3584, dataGroup_hi_lo_3584};
  wire [31:0]   dataGroup_0_80 = dataGroup_lo_3584[95:64];
  wire [2047:0] dataGroup_lo_3585 = {dataGroup_lo_hi_3585, dataGroup_lo_lo_3585};
  wire [2047:0] dataGroup_hi_3585 = {dataGroup_hi_hi_3585, dataGroup_hi_lo_3585};
  wire [31:0]   dataGroup_1_80 = dataGroup_lo_3585[223:192];
  wire [2047:0] dataGroup_lo_3586 = {dataGroup_lo_hi_3586, dataGroup_lo_lo_3586};
  wire [2047:0] dataGroup_hi_3586 = {dataGroup_hi_hi_3586, dataGroup_hi_lo_3586};
  wire [31:0]   dataGroup_2_80 = dataGroup_lo_3586[351:320];
  wire [2047:0] dataGroup_lo_3587 = {dataGroup_lo_hi_3587, dataGroup_lo_lo_3587};
  wire [2047:0] dataGroup_hi_3587 = {dataGroup_hi_hi_3587, dataGroup_hi_lo_3587};
  wire [31:0]   dataGroup_3_80 = dataGroup_lo_3587[479:448];
  wire [2047:0] dataGroup_lo_3588 = {dataGroup_lo_hi_3588, dataGroup_lo_lo_3588};
  wire [2047:0] dataGroup_hi_3588 = {dataGroup_hi_hi_3588, dataGroup_hi_lo_3588};
  wire [31:0]   dataGroup_4_80 = dataGroup_lo_3588[607:576];
  wire [2047:0] dataGroup_lo_3589 = {dataGroup_lo_hi_3589, dataGroup_lo_lo_3589};
  wire [2047:0] dataGroup_hi_3589 = {dataGroup_hi_hi_3589, dataGroup_hi_lo_3589};
  wire [31:0]   dataGroup_5_80 = dataGroup_lo_3589[735:704];
  wire [2047:0] dataGroup_lo_3590 = {dataGroup_lo_hi_3590, dataGroup_lo_lo_3590};
  wire [2047:0] dataGroup_hi_3590 = {dataGroup_hi_hi_3590, dataGroup_hi_lo_3590};
  wire [31:0]   dataGroup_6_80 = dataGroup_lo_3590[863:832];
  wire [2047:0] dataGroup_lo_3591 = {dataGroup_lo_hi_3591, dataGroup_lo_lo_3591};
  wire [2047:0] dataGroup_hi_3591 = {dataGroup_hi_hi_3591, dataGroup_hi_lo_3591};
  wire [31:0]   dataGroup_7_80 = dataGroup_lo_3591[991:960];
  wire [2047:0] dataGroup_lo_3592 = {dataGroup_lo_hi_3592, dataGroup_lo_lo_3592};
  wire [2047:0] dataGroup_hi_3592 = {dataGroup_hi_hi_3592, dataGroup_hi_lo_3592};
  wire [31:0]   dataGroup_8_80 = dataGroup_lo_3592[1119:1088];
  wire [2047:0] dataGroup_lo_3593 = {dataGroup_lo_hi_3593, dataGroup_lo_lo_3593};
  wire [2047:0] dataGroup_hi_3593 = {dataGroup_hi_hi_3593, dataGroup_hi_lo_3593};
  wire [31:0]   dataGroup_9_80 = dataGroup_lo_3593[1247:1216];
  wire [2047:0] dataGroup_lo_3594 = {dataGroup_lo_hi_3594, dataGroup_lo_lo_3594};
  wire [2047:0] dataGroup_hi_3594 = {dataGroup_hi_hi_3594, dataGroup_hi_lo_3594};
  wire [31:0]   dataGroup_10_80 = dataGroup_lo_3594[1375:1344];
  wire [2047:0] dataGroup_lo_3595 = {dataGroup_lo_hi_3595, dataGroup_lo_lo_3595};
  wire [2047:0] dataGroup_hi_3595 = {dataGroup_hi_hi_3595, dataGroup_hi_lo_3595};
  wire [31:0]   dataGroup_11_80 = dataGroup_lo_3595[1503:1472];
  wire [2047:0] dataGroup_lo_3596 = {dataGroup_lo_hi_3596, dataGroup_lo_lo_3596};
  wire [2047:0] dataGroup_hi_3596 = {dataGroup_hi_hi_3596, dataGroup_hi_lo_3596};
  wire [31:0]   dataGroup_12_80 = dataGroup_lo_3596[1631:1600];
  wire [2047:0] dataGroup_lo_3597 = {dataGroup_lo_hi_3597, dataGroup_lo_lo_3597};
  wire [2047:0] dataGroup_hi_3597 = {dataGroup_hi_hi_3597, dataGroup_hi_lo_3597};
  wire [31:0]   dataGroup_13_80 = dataGroup_lo_3597[1759:1728];
  wire [2047:0] dataGroup_lo_3598 = {dataGroup_lo_hi_3598, dataGroup_lo_lo_3598};
  wire [2047:0] dataGroup_hi_3598 = {dataGroup_hi_hi_3598, dataGroup_hi_lo_3598};
  wire [31:0]   dataGroup_14_80 = dataGroup_lo_3598[1887:1856];
  wire [2047:0] dataGroup_lo_3599 = {dataGroup_lo_hi_3599, dataGroup_lo_lo_3599};
  wire [2047:0] dataGroup_hi_3599 = {dataGroup_hi_hi_3599, dataGroup_hi_lo_3599};
  wire [31:0]   dataGroup_15_80 = dataGroup_lo_3599[2015:1984];
  wire [63:0]   res_lo_lo_lo_80 = {dataGroup_1_80, dataGroup_0_80};
  wire [63:0]   res_lo_lo_hi_80 = {dataGroup_3_80, dataGroup_2_80};
  wire [127:0]  res_lo_lo_80 = {res_lo_lo_hi_80, res_lo_lo_lo_80};
  wire [63:0]   res_lo_hi_lo_80 = {dataGroup_5_80, dataGroup_4_80};
  wire [63:0]   res_lo_hi_hi_80 = {dataGroup_7_80, dataGroup_6_80};
  wire [127:0]  res_lo_hi_80 = {res_lo_hi_hi_80, res_lo_hi_lo_80};
  wire [255:0]  res_lo_80 = {res_lo_hi_80, res_lo_lo_80};
  wire [63:0]   res_hi_lo_lo_80 = {dataGroup_9_80, dataGroup_8_80};
  wire [63:0]   res_hi_lo_hi_80 = {dataGroup_11_80, dataGroup_10_80};
  wire [127:0]  res_hi_lo_80 = {res_hi_lo_hi_80, res_hi_lo_lo_80};
  wire [63:0]   res_hi_hi_lo_80 = {dataGroup_13_80, dataGroup_12_80};
  wire [63:0]   res_hi_hi_hi_80 = {dataGroup_15_80, dataGroup_14_80};
  wire [127:0]  res_hi_hi_80 = {res_hi_hi_hi_80, res_hi_hi_lo_80};
  wire [255:0]  res_hi_80 = {res_hi_hi_80, res_hi_lo_80};
  wire [511:0]  res_154 = {res_hi_80, res_lo_80};
  wire [2047:0] dataGroup_lo_3600 = {dataGroup_lo_hi_3600, dataGroup_lo_lo_3600};
  wire [2047:0] dataGroup_hi_3600 = {dataGroup_hi_hi_3600, dataGroup_hi_lo_3600};
  wire [31:0]   dataGroup_0_81 = dataGroup_lo_3600[127:96];
  wire [2047:0] dataGroup_lo_3601 = {dataGroup_lo_hi_3601, dataGroup_lo_lo_3601};
  wire [2047:0] dataGroup_hi_3601 = {dataGroup_hi_hi_3601, dataGroup_hi_lo_3601};
  wire [31:0]   dataGroup_1_81 = dataGroup_lo_3601[255:224];
  wire [2047:0] dataGroup_lo_3602 = {dataGroup_lo_hi_3602, dataGroup_lo_lo_3602};
  wire [2047:0] dataGroup_hi_3602 = {dataGroup_hi_hi_3602, dataGroup_hi_lo_3602};
  wire [31:0]   dataGroup_2_81 = dataGroup_lo_3602[383:352];
  wire [2047:0] dataGroup_lo_3603 = {dataGroup_lo_hi_3603, dataGroup_lo_lo_3603};
  wire [2047:0] dataGroup_hi_3603 = {dataGroup_hi_hi_3603, dataGroup_hi_lo_3603};
  wire [31:0]   dataGroup_3_81 = dataGroup_lo_3603[511:480];
  wire [2047:0] dataGroup_lo_3604 = {dataGroup_lo_hi_3604, dataGroup_lo_lo_3604};
  wire [2047:0] dataGroup_hi_3604 = {dataGroup_hi_hi_3604, dataGroup_hi_lo_3604};
  wire [31:0]   dataGroup_4_81 = dataGroup_lo_3604[639:608];
  wire [2047:0] dataGroup_lo_3605 = {dataGroup_lo_hi_3605, dataGroup_lo_lo_3605};
  wire [2047:0] dataGroup_hi_3605 = {dataGroup_hi_hi_3605, dataGroup_hi_lo_3605};
  wire [31:0]   dataGroup_5_81 = dataGroup_lo_3605[767:736];
  wire [2047:0] dataGroup_lo_3606 = {dataGroup_lo_hi_3606, dataGroup_lo_lo_3606};
  wire [2047:0] dataGroup_hi_3606 = {dataGroup_hi_hi_3606, dataGroup_hi_lo_3606};
  wire [31:0]   dataGroup_6_81 = dataGroup_lo_3606[895:864];
  wire [2047:0] dataGroup_lo_3607 = {dataGroup_lo_hi_3607, dataGroup_lo_lo_3607};
  wire [2047:0] dataGroup_hi_3607 = {dataGroup_hi_hi_3607, dataGroup_hi_lo_3607};
  wire [31:0]   dataGroup_7_81 = dataGroup_lo_3607[1023:992];
  wire [2047:0] dataGroup_lo_3608 = {dataGroup_lo_hi_3608, dataGroup_lo_lo_3608};
  wire [2047:0] dataGroup_hi_3608 = {dataGroup_hi_hi_3608, dataGroup_hi_lo_3608};
  wire [31:0]   dataGroup_8_81 = dataGroup_lo_3608[1151:1120];
  wire [2047:0] dataGroup_lo_3609 = {dataGroup_lo_hi_3609, dataGroup_lo_lo_3609};
  wire [2047:0] dataGroup_hi_3609 = {dataGroup_hi_hi_3609, dataGroup_hi_lo_3609};
  wire [31:0]   dataGroup_9_81 = dataGroup_lo_3609[1279:1248];
  wire [2047:0] dataGroup_lo_3610 = {dataGroup_lo_hi_3610, dataGroup_lo_lo_3610};
  wire [2047:0] dataGroup_hi_3610 = {dataGroup_hi_hi_3610, dataGroup_hi_lo_3610};
  wire [31:0]   dataGroup_10_81 = dataGroup_lo_3610[1407:1376];
  wire [2047:0] dataGroup_lo_3611 = {dataGroup_lo_hi_3611, dataGroup_lo_lo_3611};
  wire [2047:0] dataGroup_hi_3611 = {dataGroup_hi_hi_3611, dataGroup_hi_lo_3611};
  wire [31:0]   dataGroup_11_81 = dataGroup_lo_3611[1535:1504];
  wire [2047:0] dataGroup_lo_3612 = {dataGroup_lo_hi_3612, dataGroup_lo_lo_3612};
  wire [2047:0] dataGroup_hi_3612 = {dataGroup_hi_hi_3612, dataGroup_hi_lo_3612};
  wire [31:0]   dataGroup_12_81 = dataGroup_lo_3612[1663:1632];
  wire [2047:0] dataGroup_lo_3613 = {dataGroup_lo_hi_3613, dataGroup_lo_lo_3613};
  wire [2047:0] dataGroup_hi_3613 = {dataGroup_hi_hi_3613, dataGroup_hi_lo_3613};
  wire [31:0]   dataGroup_13_81 = dataGroup_lo_3613[1791:1760];
  wire [2047:0] dataGroup_lo_3614 = {dataGroup_lo_hi_3614, dataGroup_lo_lo_3614};
  wire [2047:0] dataGroup_hi_3614 = {dataGroup_hi_hi_3614, dataGroup_hi_lo_3614};
  wire [31:0]   dataGroup_14_81 = dataGroup_lo_3614[1919:1888];
  wire [2047:0] dataGroup_lo_3615 = {dataGroup_lo_hi_3615, dataGroup_lo_lo_3615};
  wire [2047:0] dataGroup_hi_3615 = {dataGroup_hi_hi_3615, dataGroup_hi_lo_3615};
  wire [31:0]   dataGroup_15_81 = dataGroup_lo_3615[2047:2016];
  wire [63:0]   res_lo_lo_lo_81 = {dataGroup_1_81, dataGroup_0_81};
  wire [63:0]   res_lo_lo_hi_81 = {dataGroup_3_81, dataGroup_2_81};
  wire [127:0]  res_lo_lo_81 = {res_lo_lo_hi_81, res_lo_lo_lo_81};
  wire [63:0]   res_lo_hi_lo_81 = {dataGroup_5_81, dataGroup_4_81};
  wire [63:0]   res_lo_hi_hi_81 = {dataGroup_7_81, dataGroup_6_81};
  wire [127:0]  res_lo_hi_81 = {res_lo_hi_hi_81, res_lo_hi_lo_81};
  wire [255:0]  res_lo_81 = {res_lo_hi_81, res_lo_lo_81};
  wire [63:0]   res_hi_lo_lo_81 = {dataGroup_9_81, dataGroup_8_81};
  wire [63:0]   res_hi_lo_hi_81 = {dataGroup_11_81, dataGroup_10_81};
  wire [127:0]  res_hi_lo_81 = {res_hi_lo_hi_81, res_hi_lo_lo_81};
  wire [63:0]   res_hi_hi_lo_81 = {dataGroup_13_81, dataGroup_12_81};
  wire [63:0]   res_hi_hi_hi_81 = {dataGroup_15_81, dataGroup_14_81};
  wire [127:0]  res_hi_hi_81 = {res_hi_hi_hi_81, res_hi_hi_lo_81};
  wire [255:0]  res_hi_81 = {res_hi_hi_81, res_hi_lo_81};
  wire [511:0]  res_155 = {res_hi_81, res_lo_81};
  wire [1023:0] lo_lo_19 = {res_153, res_152};
  wire [1023:0] lo_hi_19 = {res_155, res_154};
  wire [2047:0] lo_19 = {lo_hi_19, lo_lo_19};
  wire [4095:0] regroupLoadData_2_3 = {2048'h0, lo_19};
  wire [2047:0] dataGroup_lo_3616 = {dataGroup_lo_hi_3616, dataGroup_lo_lo_3616};
  wire [2047:0] dataGroup_hi_3616 = {dataGroup_hi_hi_3616, dataGroup_hi_lo_3616};
  wire [31:0]   dataGroup_0_82 = dataGroup_lo_3616[31:0];
  wire [2047:0] dataGroup_lo_3617 = {dataGroup_lo_hi_3617, dataGroup_lo_lo_3617};
  wire [2047:0] dataGroup_hi_3617 = {dataGroup_hi_hi_3617, dataGroup_hi_lo_3617};
  wire [31:0]   dataGroup_1_82 = dataGroup_lo_3617[191:160];
  wire [2047:0] dataGroup_lo_3618 = {dataGroup_lo_hi_3618, dataGroup_lo_lo_3618};
  wire [2047:0] dataGroup_hi_3618 = {dataGroup_hi_hi_3618, dataGroup_hi_lo_3618};
  wire [31:0]   dataGroup_2_82 = dataGroup_lo_3618[351:320];
  wire [2047:0] dataGroup_lo_3619 = {dataGroup_lo_hi_3619, dataGroup_lo_lo_3619};
  wire [2047:0] dataGroup_hi_3619 = {dataGroup_hi_hi_3619, dataGroup_hi_lo_3619};
  wire [31:0]   dataGroup_3_82 = dataGroup_lo_3619[511:480];
  wire [2047:0] dataGroup_lo_3620 = {dataGroup_lo_hi_3620, dataGroup_lo_lo_3620};
  wire [2047:0] dataGroup_hi_3620 = {dataGroup_hi_hi_3620, dataGroup_hi_lo_3620};
  wire [31:0]   dataGroup_4_82 = dataGroup_lo_3620[671:640];
  wire [2047:0] dataGroup_lo_3621 = {dataGroup_lo_hi_3621, dataGroup_lo_lo_3621};
  wire [2047:0] dataGroup_hi_3621 = {dataGroup_hi_hi_3621, dataGroup_hi_lo_3621};
  wire [31:0]   dataGroup_5_82 = dataGroup_lo_3621[831:800];
  wire [2047:0] dataGroup_lo_3622 = {dataGroup_lo_hi_3622, dataGroup_lo_lo_3622};
  wire [2047:0] dataGroup_hi_3622 = {dataGroup_hi_hi_3622, dataGroup_hi_lo_3622};
  wire [31:0]   dataGroup_6_82 = dataGroup_lo_3622[991:960];
  wire [2047:0] dataGroup_lo_3623 = {dataGroup_lo_hi_3623, dataGroup_lo_lo_3623};
  wire [2047:0] dataGroup_hi_3623 = {dataGroup_hi_hi_3623, dataGroup_hi_lo_3623};
  wire [31:0]   dataGroup_7_82 = dataGroup_lo_3623[1151:1120];
  wire [2047:0] dataGroup_lo_3624 = {dataGroup_lo_hi_3624, dataGroup_lo_lo_3624};
  wire [2047:0] dataGroup_hi_3624 = {dataGroup_hi_hi_3624, dataGroup_hi_lo_3624};
  wire [31:0]   dataGroup_8_82 = dataGroup_lo_3624[1311:1280];
  wire [2047:0] dataGroup_lo_3625 = {dataGroup_lo_hi_3625, dataGroup_lo_lo_3625};
  wire [2047:0] dataGroup_hi_3625 = {dataGroup_hi_hi_3625, dataGroup_hi_lo_3625};
  wire [31:0]   dataGroup_9_82 = dataGroup_lo_3625[1471:1440];
  wire [2047:0] dataGroup_lo_3626 = {dataGroup_lo_hi_3626, dataGroup_lo_lo_3626};
  wire [2047:0] dataGroup_hi_3626 = {dataGroup_hi_hi_3626, dataGroup_hi_lo_3626};
  wire [31:0]   dataGroup_10_82 = dataGroup_lo_3626[1631:1600];
  wire [2047:0] dataGroup_lo_3627 = {dataGroup_lo_hi_3627, dataGroup_lo_lo_3627};
  wire [2047:0] dataGroup_hi_3627 = {dataGroup_hi_hi_3627, dataGroup_hi_lo_3627};
  wire [31:0]   dataGroup_11_82 = dataGroup_lo_3627[1791:1760];
  wire [2047:0] dataGroup_lo_3628 = {dataGroup_lo_hi_3628, dataGroup_lo_lo_3628};
  wire [2047:0] dataGroup_hi_3628 = {dataGroup_hi_hi_3628, dataGroup_hi_lo_3628};
  wire [31:0]   dataGroup_12_82 = dataGroup_lo_3628[1951:1920];
  wire [2047:0] dataGroup_lo_3629 = {dataGroup_lo_hi_3629, dataGroup_lo_lo_3629};
  wire [2047:0] dataGroup_hi_3629 = {dataGroup_hi_hi_3629, dataGroup_hi_lo_3629};
  wire [31:0]   dataGroup_13_82 = dataGroup_hi_3629[63:32];
  wire [2047:0] dataGroup_lo_3630 = {dataGroup_lo_hi_3630, dataGroup_lo_lo_3630};
  wire [2047:0] dataGroup_hi_3630 = {dataGroup_hi_hi_3630, dataGroup_hi_lo_3630};
  wire [31:0]   dataGroup_14_82 = dataGroup_hi_3630[223:192];
  wire [2047:0] dataGroup_lo_3631 = {dataGroup_lo_hi_3631, dataGroup_lo_lo_3631};
  wire [2047:0] dataGroup_hi_3631 = {dataGroup_hi_hi_3631, dataGroup_hi_lo_3631};
  wire [31:0]   dataGroup_15_82 = dataGroup_hi_3631[383:352];
  wire [63:0]   res_lo_lo_lo_82 = {dataGroup_1_82, dataGroup_0_82};
  wire [63:0]   res_lo_lo_hi_82 = {dataGroup_3_82, dataGroup_2_82};
  wire [127:0]  res_lo_lo_82 = {res_lo_lo_hi_82, res_lo_lo_lo_82};
  wire [63:0]   res_lo_hi_lo_82 = {dataGroup_5_82, dataGroup_4_82};
  wire [63:0]   res_lo_hi_hi_82 = {dataGroup_7_82, dataGroup_6_82};
  wire [127:0]  res_lo_hi_82 = {res_lo_hi_hi_82, res_lo_hi_lo_82};
  wire [255:0]  res_lo_82 = {res_lo_hi_82, res_lo_lo_82};
  wire [63:0]   res_hi_lo_lo_82 = {dataGroup_9_82, dataGroup_8_82};
  wire [63:0]   res_hi_lo_hi_82 = {dataGroup_11_82, dataGroup_10_82};
  wire [127:0]  res_hi_lo_82 = {res_hi_lo_hi_82, res_hi_lo_lo_82};
  wire [63:0]   res_hi_hi_lo_82 = {dataGroup_13_82, dataGroup_12_82};
  wire [63:0]   res_hi_hi_hi_82 = {dataGroup_15_82, dataGroup_14_82};
  wire [127:0]  res_hi_hi_82 = {res_hi_hi_hi_82, res_hi_hi_lo_82};
  wire [255:0]  res_hi_82 = {res_hi_hi_82, res_hi_lo_82};
  wire [511:0]  res_160 = {res_hi_82, res_lo_82};
  wire [2047:0] dataGroup_lo_3632 = {dataGroup_lo_hi_3632, dataGroup_lo_lo_3632};
  wire [2047:0] dataGroup_hi_3632 = {dataGroup_hi_hi_3632, dataGroup_hi_lo_3632};
  wire [31:0]   dataGroup_0_83 = dataGroup_lo_3632[63:32];
  wire [2047:0] dataGroup_lo_3633 = {dataGroup_lo_hi_3633, dataGroup_lo_lo_3633};
  wire [2047:0] dataGroup_hi_3633 = {dataGroup_hi_hi_3633, dataGroup_hi_lo_3633};
  wire [31:0]   dataGroup_1_83 = dataGroup_lo_3633[223:192];
  wire [2047:0] dataGroup_lo_3634 = {dataGroup_lo_hi_3634, dataGroup_lo_lo_3634};
  wire [2047:0] dataGroup_hi_3634 = {dataGroup_hi_hi_3634, dataGroup_hi_lo_3634};
  wire [31:0]   dataGroup_2_83 = dataGroup_lo_3634[383:352];
  wire [2047:0] dataGroup_lo_3635 = {dataGroup_lo_hi_3635, dataGroup_lo_lo_3635};
  wire [2047:0] dataGroup_hi_3635 = {dataGroup_hi_hi_3635, dataGroup_hi_lo_3635};
  wire [31:0]   dataGroup_3_83 = dataGroup_lo_3635[543:512];
  wire [2047:0] dataGroup_lo_3636 = {dataGroup_lo_hi_3636, dataGroup_lo_lo_3636};
  wire [2047:0] dataGroup_hi_3636 = {dataGroup_hi_hi_3636, dataGroup_hi_lo_3636};
  wire [31:0]   dataGroup_4_83 = dataGroup_lo_3636[703:672];
  wire [2047:0] dataGroup_lo_3637 = {dataGroup_lo_hi_3637, dataGroup_lo_lo_3637};
  wire [2047:0] dataGroup_hi_3637 = {dataGroup_hi_hi_3637, dataGroup_hi_lo_3637};
  wire [31:0]   dataGroup_5_83 = dataGroup_lo_3637[863:832];
  wire [2047:0] dataGroup_lo_3638 = {dataGroup_lo_hi_3638, dataGroup_lo_lo_3638};
  wire [2047:0] dataGroup_hi_3638 = {dataGroup_hi_hi_3638, dataGroup_hi_lo_3638};
  wire [31:0]   dataGroup_6_83 = dataGroup_lo_3638[1023:992];
  wire [2047:0] dataGroup_lo_3639 = {dataGroup_lo_hi_3639, dataGroup_lo_lo_3639};
  wire [2047:0] dataGroup_hi_3639 = {dataGroup_hi_hi_3639, dataGroup_hi_lo_3639};
  wire [31:0]   dataGroup_7_83 = dataGroup_lo_3639[1183:1152];
  wire [2047:0] dataGroup_lo_3640 = {dataGroup_lo_hi_3640, dataGroup_lo_lo_3640};
  wire [2047:0] dataGroup_hi_3640 = {dataGroup_hi_hi_3640, dataGroup_hi_lo_3640};
  wire [31:0]   dataGroup_8_83 = dataGroup_lo_3640[1343:1312];
  wire [2047:0] dataGroup_lo_3641 = {dataGroup_lo_hi_3641, dataGroup_lo_lo_3641};
  wire [2047:0] dataGroup_hi_3641 = {dataGroup_hi_hi_3641, dataGroup_hi_lo_3641};
  wire [31:0]   dataGroup_9_83 = dataGroup_lo_3641[1503:1472];
  wire [2047:0] dataGroup_lo_3642 = {dataGroup_lo_hi_3642, dataGroup_lo_lo_3642};
  wire [2047:0] dataGroup_hi_3642 = {dataGroup_hi_hi_3642, dataGroup_hi_lo_3642};
  wire [31:0]   dataGroup_10_83 = dataGroup_lo_3642[1663:1632];
  wire [2047:0] dataGroup_lo_3643 = {dataGroup_lo_hi_3643, dataGroup_lo_lo_3643};
  wire [2047:0] dataGroup_hi_3643 = {dataGroup_hi_hi_3643, dataGroup_hi_lo_3643};
  wire [31:0]   dataGroup_11_83 = dataGroup_lo_3643[1823:1792];
  wire [2047:0] dataGroup_lo_3644 = {dataGroup_lo_hi_3644, dataGroup_lo_lo_3644};
  wire [2047:0] dataGroup_hi_3644 = {dataGroup_hi_hi_3644, dataGroup_hi_lo_3644};
  wire [31:0]   dataGroup_12_83 = dataGroup_lo_3644[1983:1952];
  wire [2047:0] dataGroup_lo_3645 = {dataGroup_lo_hi_3645, dataGroup_lo_lo_3645};
  wire [2047:0] dataGroup_hi_3645 = {dataGroup_hi_hi_3645, dataGroup_hi_lo_3645};
  wire [31:0]   dataGroup_13_83 = dataGroup_hi_3645[95:64];
  wire [2047:0] dataGroup_lo_3646 = {dataGroup_lo_hi_3646, dataGroup_lo_lo_3646};
  wire [2047:0] dataGroup_hi_3646 = {dataGroup_hi_hi_3646, dataGroup_hi_lo_3646};
  wire [31:0]   dataGroup_14_83 = dataGroup_hi_3646[255:224];
  wire [2047:0] dataGroup_lo_3647 = {dataGroup_lo_hi_3647, dataGroup_lo_lo_3647};
  wire [2047:0] dataGroup_hi_3647 = {dataGroup_hi_hi_3647, dataGroup_hi_lo_3647};
  wire [31:0]   dataGroup_15_83 = dataGroup_hi_3647[415:384];
  wire [63:0]   res_lo_lo_lo_83 = {dataGroup_1_83, dataGroup_0_83};
  wire [63:0]   res_lo_lo_hi_83 = {dataGroup_3_83, dataGroup_2_83};
  wire [127:0]  res_lo_lo_83 = {res_lo_lo_hi_83, res_lo_lo_lo_83};
  wire [63:0]   res_lo_hi_lo_83 = {dataGroup_5_83, dataGroup_4_83};
  wire [63:0]   res_lo_hi_hi_83 = {dataGroup_7_83, dataGroup_6_83};
  wire [127:0]  res_lo_hi_83 = {res_lo_hi_hi_83, res_lo_hi_lo_83};
  wire [255:0]  res_lo_83 = {res_lo_hi_83, res_lo_lo_83};
  wire [63:0]   res_hi_lo_lo_83 = {dataGroup_9_83, dataGroup_8_83};
  wire [63:0]   res_hi_lo_hi_83 = {dataGroup_11_83, dataGroup_10_83};
  wire [127:0]  res_hi_lo_83 = {res_hi_lo_hi_83, res_hi_lo_lo_83};
  wire [63:0]   res_hi_hi_lo_83 = {dataGroup_13_83, dataGroup_12_83};
  wire [63:0]   res_hi_hi_hi_83 = {dataGroup_15_83, dataGroup_14_83};
  wire [127:0]  res_hi_hi_83 = {res_hi_hi_hi_83, res_hi_hi_lo_83};
  wire [255:0]  res_hi_83 = {res_hi_hi_83, res_hi_lo_83};
  wire [511:0]  res_161 = {res_hi_83, res_lo_83};
  wire [2047:0] dataGroup_lo_3648 = {dataGroup_lo_hi_3648, dataGroup_lo_lo_3648};
  wire [2047:0] dataGroup_hi_3648 = {dataGroup_hi_hi_3648, dataGroup_hi_lo_3648};
  wire [31:0]   dataGroup_0_84 = dataGroup_lo_3648[95:64];
  wire [2047:0] dataGroup_lo_3649 = {dataGroup_lo_hi_3649, dataGroup_lo_lo_3649};
  wire [2047:0] dataGroup_hi_3649 = {dataGroup_hi_hi_3649, dataGroup_hi_lo_3649};
  wire [31:0]   dataGroup_1_84 = dataGroup_lo_3649[255:224];
  wire [2047:0] dataGroup_lo_3650 = {dataGroup_lo_hi_3650, dataGroup_lo_lo_3650};
  wire [2047:0] dataGroup_hi_3650 = {dataGroup_hi_hi_3650, dataGroup_hi_lo_3650};
  wire [31:0]   dataGroup_2_84 = dataGroup_lo_3650[415:384];
  wire [2047:0] dataGroup_lo_3651 = {dataGroup_lo_hi_3651, dataGroup_lo_lo_3651};
  wire [2047:0] dataGroup_hi_3651 = {dataGroup_hi_hi_3651, dataGroup_hi_lo_3651};
  wire [31:0]   dataGroup_3_84 = dataGroup_lo_3651[575:544];
  wire [2047:0] dataGroup_lo_3652 = {dataGroup_lo_hi_3652, dataGroup_lo_lo_3652};
  wire [2047:0] dataGroup_hi_3652 = {dataGroup_hi_hi_3652, dataGroup_hi_lo_3652};
  wire [31:0]   dataGroup_4_84 = dataGroup_lo_3652[735:704];
  wire [2047:0] dataGroup_lo_3653 = {dataGroup_lo_hi_3653, dataGroup_lo_lo_3653};
  wire [2047:0] dataGroup_hi_3653 = {dataGroup_hi_hi_3653, dataGroup_hi_lo_3653};
  wire [31:0]   dataGroup_5_84 = dataGroup_lo_3653[895:864];
  wire [2047:0] dataGroup_lo_3654 = {dataGroup_lo_hi_3654, dataGroup_lo_lo_3654};
  wire [2047:0] dataGroup_hi_3654 = {dataGroup_hi_hi_3654, dataGroup_hi_lo_3654};
  wire [31:0]   dataGroup_6_84 = dataGroup_lo_3654[1055:1024];
  wire [2047:0] dataGroup_lo_3655 = {dataGroup_lo_hi_3655, dataGroup_lo_lo_3655};
  wire [2047:0] dataGroup_hi_3655 = {dataGroup_hi_hi_3655, dataGroup_hi_lo_3655};
  wire [31:0]   dataGroup_7_84 = dataGroup_lo_3655[1215:1184];
  wire [2047:0] dataGroup_lo_3656 = {dataGroup_lo_hi_3656, dataGroup_lo_lo_3656};
  wire [2047:0] dataGroup_hi_3656 = {dataGroup_hi_hi_3656, dataGroup_hi_lo_3656};
  wire [31:0]   dataGroup_8_84 = dataGroup_lo_3656[1375:1344];
  wire [2047:0] dataGroup_lo_3657 = {dataGroup_lo_hi_3657, dataGroup_lo_lo_3657};
  wire [2047:0] dataGroup_hi_3657 = {dataGroup_hi_hi_3657, dataGroup_hi_lo_3657};
  wire [31:0]   dataGroup_9_84 = dataGroup_lo_3657[1535:1504];
  wire [2047:0] dataGroup_lo_3658 = {dataGroup_lo_hi_3658, dataGroup_lo_lo_3658};
  wire [2047:0] dataGroup_hi_3658 = {dataGroup_hi_hi_3658, dataGroup_hi_lo_3658};
  wire [31:0]   dataGroup_10_84 = dataGroup_lo_3658[1695:1664];
  wire [2047:0] dataGroup_lo_3659 = {dataGroup_lo_hi_3659, dataGroup_lo_lo_3659};
  wire [2047:0] dataGroup_hi_3659 = {dataGroup_hi_hi_3659, dataGroup_hi_lo_3659};
  wire [31:0]   dataGroup_11_84 = dataGroup_lo_3659[1855:1824];
  wire [2047:0] dataGroup_lo_3660 = {dataGroup_lo_hi_3660, dataGroup_lo_lo_3660};
  wire [2047:0] dataGroup_hi_3660 = {dataGroup_hi_hi_3660, dataGroup_hi_lo_3660};
  wire [31:0]   dataGroup_12_84 = dataGroup_lo_3660[2015:1984];
  wire [2047:0] dataGroup_lo_3661 = {dataGroup_lo_hi_3661, dataGroup_lo_lo_3661};
  wire [2047:0] dataGroup_hi_3661 = {dataGroup_hi_hi_3661, dataGroup_hi_lo_3661};
  wire [31:0]   dataGroup_13_84 = dataGroup_hi_3661[127:96];
  wire [2047:0] dataGroup_lo_3662 = {dataGroup_lo_hi_3662, dataGroup_lo_lo_3662};
  wire [2047:0] dataGroup_hi_3662 = {dataGroup_hi_hi_3662, dataGroup_hi_lo_3662};
  wire [31:0]   dataGroup_14_84 = dataGroup_hi_3662[287:256];
  wire [2047:0] dataGroup_lo_3663 = {dataGroup_lo_hi_3663, dataGroup_lo_lo_3663};
  wire [2047:0] dataGroup_hi_3663 = {dataGroup_hi_hi_3663, dataGroup_hi_lo_3663};
  wire [31:0]   dataGroup_15_84 = dataGroup_hi_3663[447:416];
  wire [63:0]   res_lo_lo_lo_84 = {dataGroup_1_84, dataGroup_0_84};
  wire [63:0]   res_lo_lo_hi_84 = {dataGroup_3_84, dataGroup_2_84};
  wire [127:0]  res_lo_lo_84 = {res_lo_lo_hi_84, res_lo_lo_lo_84};
  wire [63:0]   res_lo_hi_lo_84 = {dataGroup_5_84, dataGroup_4_84};
  wire [63:0]   res_lo_hi_hi_84 = {dataGroup_7_84, dataGroup_6_84};
  wire [127:0]  res_lo_hi_84 = {res_lo_hi_hi_84, res_lo_hi_lo_84};
  wire [255:0]  res_lo_84 = {res_lo_hi_84, res_lo_lo_84};
  wire [63:0]   res_hi_lo_lo_84 = {dataGroup_9_84, dataGroup_8_84};
  wire [63:0]   res_hi_lo_hi_84 = {dataGroup_11_84, dataGroup_10_84};
  wire [127:0]  res_hi_lo_84 = {res_hi_lo_hi_84, res_hi_lo_lo_84};
  wire [63:0]   res_hi_hi_lo_84 = {dataGroup_13_84, dataGroup_12_84};
  wire [63:0]   res_hi_hi_hi_84 = {dataGroup_15_84, dataGroup_14_84};
  wire [127:0]  res_hi_hi_84 = {res_hi_hi_hi_84, res_hi_hi_lo_84};
  wire [255:0]  res_hi_84 = {res_hi_hi_84, res_hi_lo_84};
  wire [511:0]  res_162 = {res_hi_84, res_lo_84};
  wire [2047:0] dataGroup_lo_3664 = {dataGroup_lo_hi_3664, dataGroup_lo_lo_3664};
  wire [2047:0] dataGroup_hi_3664 = {dataGroup_hi_hi_3664, dataGroup_hi_lo_3664};
  wire [31:0]   dataGroup_0_85 = dataGroup_lo_3664[127:96];
  wire [2047:0] dataGroup_lo_3665 = {dataGroup_lo_hi_3665, dataGroup_lo_lo_3665};
  wire [2047:0] dataGroup_hi_3665 = {dataGroup_hi_hi_3665, dataGroup_hi_lo_3665};
  wire [31:0]   dataGroup_1_85 = dataGroup_lo_3665[287:256];
  wire [2047:0] dataGroup_lo_3666 = {dataGroup_lo_hi_3666, dataGroup_lo_lo_3666};
  wire [2047:0] dataGroup_hi_3666 = {dataGroup_hi_hi_3666, dataGroup_hi_lo_3666};
  wire [31:0]   dataGroup_2_85 = dataGroup_lo_3666[447:416];
  wire [2047:0] dataGroup_lo_3667 = {dataGroup_lo_hi_3667, dataGroup_lo_lo_3667};
  wire [2047:0] dataGroup_hi_3667 = {dataGroup_hi_hi_3667, dataGroup_hi_lo_3667};
  wire [31:0]   dataGroup_3_85 = dataGroup_lo_3667[607:576];
  wire [2047:0] dataGroup_lo_3668 = {dataGroup_lo_hi_3668, dataGroup_lo_lo_3668};
  wire [2047:0] dataGroup_hi_3668 = {dataGroup_hi_hi_3668, dataGroup_hi_lo_3668};
  wire [31:0]   dataGroup_4_85 = dataGroup_lo_3668[767:736];
  wire [2047:0] dataGroup_lo_3669 = {dataGroup_lo_hi_3669, dataGroup_lo_lo_3669};
  wire [2047:0] dataGroup_hi_3669 = {dataGroup_hi_hi_3669, dataGroup_hi_lo_3669};
  wire [31:0]   dataGroup_5_85 = dataGroup_lo_3669[927:896];
  wire [2047:0] dataGroup_lo_3670 = {dataGroup_lo_hi_3670, dataGroup_lo_lo_3670};
  wire [2047:0] dataGroup_hi_3670 = {dataGroup_hi_hi_3670, dataGroup_hi_lo_3670};
  wire [31:0]   dataGroup_6_85 = dataGroup_lo_3670[1087:1056];
  wire [2047:0] dataGroup_lo_3671 = {dataGroup_lo_hi_3671, dataGroup_lo_lo_3671};
  wire [2047:0] dataGroup_hi_3671 = {dataGroup_hi_hi_3671, dataGroup_hi_lo_3671};
  wire [31:0]   dataGroup_7_85 = dataGroup_lo_3671[1247:1216];
  wire [2047:0] dataGroup_lo_3672 = {dataGroup_lo_hi_3672, dataGroup_lo_lo_3672};
  wire [2047:0] dataGroup_hi_3672 = {dataGroup_hi_hi_3672, dataGroup_hi_lo_3672};
  wire [31:0]   dataGroup_8_85 = dataGroup_lo_3672[1407:1376];
  wire [2047:0] dataGroup_lo_3673 = {dataGroup_lo_hi_3673, dataGroup_lo_lo_3673};
  wire [2047:0] dataGroup_hi_3673 = {dataGroup_hi_hi_3673, dataGroup_hi_lo_3673};
  wire [31:0]   dataGroup_9_85 = dataGroup_lo_3673[1567:1536];
  wire [2047:0] dataGroup_lo_3674 = {dataGroup_lo_hi_3674, dataGroup_lo_lo_3674};
  wire [2047:0] dataGroup_hi_3674 = {dataGroup_hi_hi_3674, dataGroup_hi_lo_3674};
  wire [31:0]   dataGroup_10_85 = dataGroup_lo_3674[1727:1696];
  wire [2047:0] dataGroup_lo_3675 = {dataGroup_lo_hi_3675, dataGroup_lo_lo_3675};
  wire [2047:0] dataGroup_hi_3675 = {dataGroup_hi_hi_3675, dataGroup_hi_lo_3675};
  wire [31:0]   dataGroup_11_85 = dataGroup_lo_3675[1887:1856];
  wire [2047:0] dataGroup_lo_3676 = {dataGroup_lo_hi_3676, dataGroup_lo_lo_3676};
  wire [2047:0] dataGroup_hi_3676 = {dataGroup_hi_hi_3676, dataGroup_hi_lo_3676};
  wire [31:0]   dataGroup_12_85 = dataGroup_lo_3676[2047:2016];
  wire [2047:0] dataGroup_lo_3677 = {dataGroup_lo_hi_3677, dataGroup_lo_lo_3677};
  wire [2047:0] dataGroup_hi_3677 = {dataGroup_hi_hi_3677, dataGroup_hi_lo_3677};
  wire [31:0]   dataGroup_13_85 = dataGroup_hi_3677[159:128];
  wire [2047:0] dataGroup_lo_3678 = {dataGroup_lo_hi_3678, dataGroup_lo_lo_3678};
  wire [2047:0] dataGroup_hi_3678 = {dataGroup_hi_hi_3678, dataGroup_hi_lo_3678};
  wire [31:0]   dataGroup_14_85 = dataGroup_hi_3678[319:288];
  wire [2047:0] dataGroup_lo_3679 = {dataGroup_lo_hi_3679, dataGroup_lo_lo_3679};
  wire [2047:0] dataGroup_hi_3679 = {dataGroup_hi_hi_3679, dataGroup_hi_lo_3679};
  wire [31:0]   dataGroup_15_85 = dataGroup_hi_3679[479:448];
  wire [63:0]   res_lo_lo_lo_85 = {dataGroup_1_85, dataGroup_0_85};
  wire [63:0]   res_lo_lo_hi_85 = {dataGroup_3_85, dataGroup_2_85};
  wire [127:0]  res_lo_lo_85 = {res_lo_lo_hi_85, res_lo_lo_lo_85};
  wire [63:0]   res_lo_hi_lo_85 = {dataGroup_5_85, dataGroup_4_85};
  wire [63:0]   res_lo_hi_hi_85 = {dataGroup_7_85, dataGroup_6_85};
  wire [127:0]  res_lo_hi_85 = {res_lo_hi_hi_85, res_lo_hi_lo_85};
  wire [255:0]  res_lo_85 = {res_lo_hi_85, res_lo_lo_85};
  wire [63:0]   res_hi_lo_lo_85 = {dataGroup_9_85, dataGroup_8_85};
  wire [63:0]   res_hi_lo_hi_85 = {dataGroup_11_85, dataGroup_10_85};
  wire [127:0]  res_hi_lo_85 = {res_hi_lo_hi_85, res_hi_lo_lo_85};
  wire [63:0]   res_hi_hi_lo_85 = {dataGroup_13_85, dataGroup_12_85};
  wire [63:0]   res_hi_hi_hi_85 = {dataGroup_15_85, dataGroup_14_85};
  wire [127:0]  res_hi_hi_85 = {res_hi_hi_hi_85, res_hi_hi_lo_85};
  wire [255:0]  res_hi_85 = {res_hi_hi_85, res_hi_lo_85};
  wire [511:0]  res_163 = {res_hi_85, res_lo_85};
  wire [2047:0] dataGroup_lo_3680 = {dataGroup_lo_hi_3680, dataGroup_lo_lo_3680};
  wire [2047:0] dataGroup_hi_3680 = {dataGroup_hi_hi_3680, dataGroup_hi_lo_3680};
  wire [31:0]   dataGroup_0_86 = dataGroup_lo_3680[159:128];
  wire [2047:0] dataGroup_lo_3681 = {dataGroup_lo_hi_3681, dataGroup_lo_lo_3681};
  wire [2047:0] dataGroup_hi_3681 = {dataGroup_hi_hi_3681, dataGroup_hi_lo_3681};
  wire [31:0]   dataGroup_1_86 = dataGroup_lo_3681[319:288];
  wire [2047:0] dataGroup_lo_3682 = {dataGroup_lo_hi_3682, dataGroup_lo_lo_3682};
  wire [2047:0] dataGroup_hi_3682 = {dataGroup_hi_hi_3682, dataGroup_hi_lo_3682};
  wire [31:0]   dataGroup_2_86 = dataGroup_lo_3682[479:448];
  wire [2047:0] dataGroup_lo_3683 = {dataGroup_lo_hi_3683, dataGroup_lo_lo_3683};
  wire [2047:0] dataGroup_hi_3683 = {dataGroup_hi_hi_3683, dataGroup_hi_lo_3683};
  wire [31:0]   dataGroup_3_86 = dataGroup_lo_3683[639:608];
  wire [2047:0] dataGroup_lo_3684 = {dataGroup_lo_hi_3684, dataGroup_lo_lo_3684};
  wire [2047:0] dataGroup_hi_3684 = {dataGroup_hi_hi_3684, dataGroup_hi_lo_3684};
  wire [31:0]   dataGroup_4_86 = dataGroup_lo_3684[799:768];
  wire [2047:0] dataGroup_lo_3685 = {dataGroup_lo_hi_3685, dataGroup_lo_lo_3685};
  wire [2047:0] dataGroup_hi_3685 = {dataGroup_hi_hi_3685, dataGroup_hi_lo_3685};
  wire [31:0]   dataGroup_5_86 = dataGroup_lo_3685[959:928];
  wire [2047:0] dataGroup_lo_3686 = {dataGroup_lo_hi_3686, dataGroup_lo_lo_3686};
  wire [2047:0] dataGroup_hi_3686 = {dataGroup_hi_hi_3686, dataGroup_hi_lo_3686};
  wire [31:0]   dataGroup_6_86 = dataGroup_lo_3686[1119:1088];
  wire [2047:0] dataGroup_lo_3687 = {dataGroup_lo_hi_3687, dataGroup_lo_lo_3687};
  wire [2047:0] dataGroup_hi_3687 = {dataGroup_hi_hi_3687, dataGroup_hi_lo_3687};
  wire [31:0]   dataGroup_7_86 = dataGroup_lo_3687[1279:1248];
  wire [2047:0] dataGroup_lo_3688 = {dataGroup_lo_hi_3688, dataGroup_lo_lo_3688};
  wire [2047:0] dataGroup_hi_3688 = {dataGroup_hi_hi_3688, dataGroup_hi_lo_3688};
  wire [31:0]   dataGroup_8_86 = dataGroup_lo_3688[1439:1408];
  wire [2047:0] dataGroup_lo_3689 = {dataGroup_lo_hi_3689, dataGroup_lo_lo_3689};
  wire [2047:0] dataGroup_hi_3689 = {dataGroup_hi_hi_3689, dataGroup_hi_lo_3689};
  wire [31:0]   dataGroup_9_86 = dataGroup_lo_3689[1599:1568];
  wire [2047:0] dataGroup_lo_3690 = {dataGroup_lo_hi_3690, dataGroup_lo_lo_3690};
  wire [2047:0] dataGroup_hi_3690 = {dataGroup_hi_hi_3690, dataGroup_hi_lo_3690};
  wire [31:0]   dataGroup_10_86 = dataGroup_lo_3690[1759:1728];
  wire [2047:0] dataGroup_lo_3691 = {dataGroup_lo_hi_3691, dataGroup_lo_lo_3691};
  wire [2047:0] dataGroup_hi_3691 = {dataGroup_hi_hi_3691, dataGroup_hi_lo_3691};
  wire [31:0]   dataGroup_11_86 = dataGroup_lo_3691[1919:1888];
  wire [2047:0] dataGroup_lo_3692 = {dataGroup_lo_hi_3692, dataGroup_lo_lo_3692};
  wire [2047:0] dataGroup_hi_3692 = {dataGroup_hi_hi_3692, dataGroup_hi_lo_3692};
  wire [31:0]   dataGroup_12_86 = dataGroup_hi_3692[31:0];
  wire [2047:0] dataGroup_lo_3693 = {dataGroup_lo_hi_3693, dataGroup_lo_lo_3693};
  wire [2047:0] dataGroup_hi_3693 = {dataGroup_hi_hi_3693, dataGroup_hi_lo_3693};
  wire [31:0]   dataGroup_13_86 = dataGroup_hi_3693[191:160];
  wire [2047:0] dataGroup_lo_3694 = {dataGroup_lo_hi_3694, dataGroup_lo_lo_3694};
  wire [2047:0] dataGroup_hi_3694 = {dataGroup_hi_hi_3694, dataGroup_hi_lo_3694};
  wire [31:0]   dataGroup_14_86 = dataGroup_hi_3694[351:320];
  wire [2047:0] dataGroup_lo_3695 = {dataGroup_lo_hi_3695, dataGroup_lo_lo_3695};
  wire [2047:0] dataGroup_hi_3695 = {dataGroup_hi_hi_3695, dataGroup_hi_lo_3695};
  wire [31:0]   dataGroup_15_86 = dataGroup_hi_3695[511:480];
  wire [63:0]   res_lo_lo_lo_86 = {dataGroup_1_86, dataGroup_0_86};
  wire [63:0]   res_lo_lo_hi_86 = {dataGroup_3_86, dataGroup_2_86};
  wire [127:0]  res_lo_lo_86 = {res_lo_lo_hi_86, res_lo_lo_lo_86};
  wire [63:0]   res_lo_hi_lo_86 = {dataGroup_5_86, dataGroup_4_86};
  wire [63:0]   res_lo_hi_hi_86 = {dataGroup_7_86, dataGroup_6_86};
  wire [127:0]  res_lo_hi_86 = {res_lo_hi_hi_86, res_lo_hi_lo_86};
  wire [255:0]  res_lo_86 = {res_lo_hi_86, res_lo_lo_86};
  wire [63:0]   res_hi_lo_lo_86 = {dataGroup_9_86, dataGroup_8_86};
  wire [63:0]   res_hi_lo_hi_86 = {dataGroup_11_86, dataGroup_10_86};
  wire [127:0]  res_hi_lo_86 = {res_hi_lo_hi_86, res_hi_lo_lo_86};
  wire [63:0]   res_hi_hi_lo_86 = {dataGroup_13_86, dataGroup_12_86};
  wire [63:0]   res_hi_hi_hi_86 = {dataGroup_15_86, dataGroup_14_86};
  wire [127:0]  res_hi_hi_86 = {res_hi_hi_hi_86, res_hi_hi_lo_86};
  wire [255:0]  res_hi_86 = {res_hi_hi_86, res_hi_lo_86};
  wire [511:0]  res_164 = {res_hi_86, res_lo_86};
  wire [1023:0] lo_lo_20 = {res_161, res_160};
  wire [1023:0] lo_hi_20 = {res_163, res_162};
  wire [2047:0] lo_20 = {lo_hi_20, lo_lo_20};
  wire [1023:0] hi_lo_20 = {512'h0, res_164};
  wire [2047:0] hi_20 = {1024'h0, hi_lo_20};
  wire [4095:0] regroupLoadData_2_4 = {hi_20, lo_20};
  wire [2047:0] dataGroup_lo_3696 = {dataGroup_lo_hi_3696, dataGroup_lo_lo_3696};
  wire [2047:0] dataGroup_hi_3696 = {dataGroup_hi_hi_3696, dataGroup_hi_lo_3696};
  wire [31:0]   dataGroup_0_87 = dataGroup_lo_3696[31:0];
  wire [2047:0] dataGroup_lo_3697 = {dataGroup_lo_hi_3697, dataGroup_lo_lo_3697};
  wire [2047:0] dataGroup_hi_3697 = {dataGroup_hi_hi_3697, dataGroup_hi_lo_3697};
  wire [31:0]   dataGroup_1_87 = dataGroup_lo_3697[223:192];
  wire [2047:0] dataGroup_lo_3698 = {dataGroup_lo_hi_3698, dataGroup_lo_lo_3698};
  wire [2047:0] dataGroup_hi_3698 = {dataGroup_hi_hi_3698, dataGroup_hi_lo_3698};
  wire [31:0]   dataGroup_2_87 = dataGroup_lo_3698[415:384];
  wire [2047:0] dataGroup_lo_3699 = {dataGroup_lo_hi_3699, dataGroup_lo_lo_3699};
  wire [2047:0] dataGroup_hi_3699 = {dataGroup_hi_hi_3699, dataGroup_hi_lo_3699};
  wire [31:0]   dataGroup_3_87 = dataGroup_lo_3699[607:576];
  wire [2047:0] dataGroup_lo_3700 = {dataGroup_lo_hi_3700, dataGroup_lo_lo_3700};
  wire [2047:0] dataGroup_hi_3700 = {dataGroup_hi_hi_3700, dataGroup_hi_lo_3700};
  wire [31:0]   dataGroup_4_87 = dataGroup_lo_3700[799:768];
  wire [2047:0] dataGroup_lo_3701 = {dataGroup_lo_hi_3701, dataGroup_lo_lo_3701};
  wire [2047:0] dataGroup_hi_3701 = {dataGroup_hi_hi_3701, dataGroup_hi_lo_3701};
  wire [31:0]   dataGroup_5_87 = dataGroup_lo_3701[991:960];
  wire [2047:0] dataGroup_lo_3702 = {dataGroup_lo_hi_3702, dataGroup_lo_lo_3702};
  wire [2047:0] dataGroup_hi_3702 = {dataGroup_hi_hi_3702, dataGroup_hi_lo_3702};
  wire [31:0]   dataGroup_6_87 = dataGroup_lo_3702[1183:1152];
  wire [2047:0] dataGroup_lo_3703 = {dataGroup_lo_hi_3703, dataGroup_lo_lo_3703};
  wire [2047:0] dataGroup_hi_3703 = {dataGroup_hi_hi_3703, dataGroup_hi_lo_3703};
  wire [31:0]   dataGroup_7_87 = dataGroup_lo_3703[1375:1344];
  wire [2047:0] dataGroup_lo_3704 = {dataGroup_lo_hi_3704, dataGroup_lo_lo_3704};
  wire [2047:0] dataGroup_hi_3704 = {dataGroup_hi_hi_3704, dataGroup_hi_lo_3704};
  wire [31:0]   dataGroup_8_87 = dataGroup_lo_3704[1567:1536];
  wire [2047:0] dataGroup_lo_3705 = {dataGroup_lo_hi_3705, dataGroup_lo_lo_3705};
  wire [2047:0] dataGroup_hi_3705 = {dataGroup_hi_hi_3705, dataGroup_hi_lo_3705};
  wire [31:0]   dataGroup_9_87 = dataGroup_lo_3705[1759:1728];
  wire [2047:0] dataGroup_lo_3706 = {dataGroup_lo_hi_3706, dataGroup_lo_lo_3706};
  wire [2047:0] dataGroup_hi_3706 = {dataGroup_hi_hi_3706, dataGroup_hi_lo_3706};
  wire [31:0]   dataGroup_10_87 = dataGroup_lo_3706[1951:1920];
  wire [2047:0] dataGroup_lo_3707 = {dataGroup_lo_hi_3707, dataGroup_lo_lo_3707};
  wire [2047:0] dataGroup_hi_3707 = {dataGroup_hi_hi_3707, dataGroup_hi_lo_3707};
  wire [31:0]   dataGroup_11_87 = dataGroup_hi_3707[95:64];
  wire [2047:0] dataGroup_lo_3708 = {dataGroup_lo_hi_3708, dataGroup_lo_lo_3708};
  wire [2047:0] dataGroup_hi_3708 = {dataGroup_hi_hi_3708, dataGroup_hi_lo_3708};
  wire [31:0]   dataGroup_12_87 = dataGroup_hi_3708[287:256];
  wire [2047:0] dataGroup_lo_3709 = {dataGroup_lo_hi_3709, dataGroup_lo_lo_3709};
  wire [2047:0] dataGroup_hi_3709 = {dataGroup_hi_hi_3709, dataGroup_hi_lo_3709};
  wire [31:0]   dataGroup_13_87 = dataGroup_hi_3709[479:448];
  wire [2047:0] dataGroup_lo_3710 = {dataGroup_lo_hi_3710, dataGroup_lo_lo_3710};
  wire [2047:0] dataGroup_hi_3710 = {dataGroup_hi_hi_3710, dataGroup_hi_lo_3710};
  wire [31:0]   dataGroup_14_87 = dataGroup_hi_3710[671:640];
  wire [2047:0] dataGroup_lo_3711 = {dataGroup_lo_hi_3711, dataGroup_lo_lo_3711};
  wire [2047:0] dataGroup_hi_3711 = {dataGroup_hi_hi_3711, dataGroup_hi_lo_3711};
  wire [31:0]   dataGroup_15_87 = dataGroup_hi_3711[863:832];
  wire [63:0]   res_lo_lo_lo_87 = {dataGroup_1_87, dataGroup_0_87};
  wire [63:0]   res_lo_lo_hi_87 = {dataGroup_3_87, dataGroup_2_87};
  wire [127:0]  res_lo_lo_87 = {res_lo_lo_hi_87, res_lo_lo_lo_87};
  wire [63:0]   res_lo_hi_lo_87 = {dataGroup_5_87, dataGroup_4_87};
  wire [63:0]   res_lo_hi_hi_87 = {dataGroup_7_87, dataGroup_6_87};
  wire [127:0]  res_lo_hi_87 = {res_lo_hi_hi_87, res_lo_hi_lo_87};
  wire [255:0]  res_lo_87 = {res_lo_hi_87, res_lo_lo_87};
  wire [63:0]   res_hi_lo_lo_87 = {dataGroup_9_87, dataGroup_8_87};
  wire [63:0]   res_hi_lo_hi_87 = {dataGroup_11_87, dataGroup_10_87};
  wire [127:0]  res_hi_lo_87 = {res_hi_lo_hi_87, res_hi_lo_lo_87};
  wire [63:0]   res_hi_hi_lo_87 = {dataGroup_13_87, dataGroup_12_87};
  wire [63:0]   res_hi_hi_hi_87 = {dataGroup_15_87, dataGroup_14_87};
  wire [127:0]  res_hi_hi_87 = {res_hi_hi_hi_87, res_hi_hi_lo_87};
  wire [255:0]  res_hi_87 = {res_hi_hi_87, res_hi_lo_87};
  wire [511:0]  res_168 = {res_hi_87, res_lo_87};
  wire [2047:0] dataGroup_lo_3712 = {dataGroup_lo_hi_3712, dataGroup_lo_lo_3712};
  wire [2047:0] dataGroup_hi_3712 = {dataGroup_hi_hi_3712, dataGroup_hi_lo_3712};
  wire [31:0]   dataGroup_0_88 = dataGroup_lo_3712[63:32];
  wire [2047:0] dataGroup_lo_3713 = {dataGroup_lo_hi_3713, dataGroup_lo_lo_3713};
  wire [2047:0] dataGroup_hi_3713 = {dataGroup_hi_hi_3713, dataGroup_hi_lo_3713};
  wire [31:0]   dataGroup_1_88 = dataGroup_lo_3713[255:224];
  wire [2047:0] dataGroup_lo_3714 = {dataGroup_lo_hi_3714, dataGroup_lo_lo_3714};
  wire [2047:0] dataGroup_hi_3714 = {dataGroup_hi_hi_3714, dataGroup_hi_lo_3714};
  wire [31:0]   dataGroup_2_88 = dataGroup_lo_3714[447:416];
  wire [2047:0] dataGroup_lo_3715 = {dataGroup_lo_hi_3715, dataGroup_lo_lo_3715};
  wire [2047:0] dataGroup_hi_3715 = {dataGroup_hi_hi_3715, dataGroup_hi_lo_3715};
  wire [31:0]   dataGroup_3_88 = dataGroup_lo_3715[639:608];
  wire [2047:0] dataGroup_lo_3716 = {dataGroup_lo_hi_3716, dataGroup_lo_lo_3716};
  wire [2047:0] dataGroup_hi_3716 = {dataGroup_hi_hi_3716, dataGroup_hi_lo_3716};
  wire [31:0]   dataGroup_4_88 = dataGroup_lo_3716[831:800];
  wire [2047:0] dataGroup_lo_3717 = {dataGroup_lo_hi_3717, dataGroup_lo_lo_3717};
  wire [2047:0] dataGroup_hi_3717 = {dataGroup_hi_hi_3717, dataGroup_hi_lo_3717};
  wire [31:0]   dataGroup_5_88 = dataGroup_lo_3717[1023:992];
  wire [2047:0] dataGroup_lo_3718 = {dataGroup_lo_hi_3718, dataGroup_lo_lo_3718};
  wire [2047:0] dataGroup_hi_3718 = {dataGroup_hi_hi_3718, dataGroup_hi_lo_3718};
  wire [31:0]   dataGroup_6_88 = dataGroup_lo_3718[1215:1184];
  wire [2047:0] dataGroup_lo_3719 = {dataGroup_lo_hi_3719, dataGroup_lo_lo_3719};
  wire [2047:0] dataGroup_hi_3719 = {dataGroup_hi_hi_3719, dataGroup_hi_lo_3719};
  wire [31:0]   dataGroup_7_88 = dataGroup_lo_3719[1407:1376];
  wire [2047:0] dataGroup_lo_3720 = {dataGroup_lo_hi_3720, dataGroup_lo_lo_3720};
  wire [2047:0] dataGroup_hi_3720 = {dataGroup_hi_hi_3720, dataGroup_hi_lo_3720};
  wire [31:0]   dataGroup_8_88 = dataGroup_lo_3720[1599:1568];
  wire [2047:0] dataGroup_lo_3721 = {dataGroup_lo_hi_3721, dataGroup_lo_lo_3721};
  wire [2047:0] dataGroup_hi_3721 = {dataGroup_hi_hi_3721, dataGroup_hi_lo_3721};
  wire [31:0]   dataGroup_9_88 = dataGroup_lo_3721[1791:1760];
  wire [2047:0] dataGroup_lo_3722 = {dataGroup_lo_hi_3722, dataGroup_lo_lo_3722};
  wire [2047:0] dataGroup_hi_3722 = {dataGroup_hi_hi_3722, dataGroup_hi_lo_3722};
  wire [31:0]   dataGroup_10_88 = dataGroup_lo_3722[1983:1952];
  wire [2047:0] dataGroup_lo_3723 = {dataGroup_lo_hi_3723, dataGroup_lo_lo_3723};
  wire [2047:0] dataGroup_hi_3723 = {dataGroup_hi_hi_3723, dataGroup_hi_lo_3723};
  wire [31:0]   dataGroup_11_88 = dataGroup_hi_3723[127:96];
  wire [2047:0] dataGroup_lo_3724 = {dataGroup_lo_hi_3724, dataGroup_lo_lo_3724};
  wire [2047:0] dataGroup_hi_3724 = {dataGroup_hi_hi_3724, dataGroup_hi_lo_3724};
  wire [31:0]   dataGroup_12_88 = dataGroup_hi_3724[319:288];
  wire [2047:0] dataGroup_lo_3725 = {dataGroup_lo_hi_3725, dataGroup_lo_lo_3725};
  wire [2047:0] dataGroup_hi_3725 = {dataGroup_hi_hi_3725, dataGroup_hi_lo_3725};
  wire [31:0]   dataGroup_13_88 = dataGroup_hi_3725[511:480];
  wire [2047:0] dataGroup_lo_3726 = {dataGroup_lo_hi_3726, dataGroup_lo_lo_3726};
  wire [2047:0] dataGroup_hi_3726 = {dataGroup_hi_hi_3726, dataGroup_hi_lo_3726};
  wire [31:0]   dataGroup_14_88 = dataGroup_hi_3726[703:672];
  wire [2047:0] dataGroup_lo_3727 = {dataGroup_lo_hi_3727, dataGroup_lo_lo_3727};
  wire [2047:0] dataGroup_hi_3727 = {dataGroup_hi_hi_3727, dataGroup_hi_lo_3727};
  wire [31:0]   dataGroup_15_88 = dataGroup_hi_3727[895:864];
  wire [63:0]   res_lo_lo_lo_88 = {dataGroup_1_88, dataGroup_0_88};
  wire [63:0]   res_lo_lo_hi_88 = {dataGroup_3_88, dataGroup_2_88};
  wire [127:0]  res_lo_lo_88 = {res_lo_lo_hi_88, res_lo_lo_lo_88};
  wire [63:0]   res_lo_hi_lo_88 = {dataGroup_5_88, dataGroup_4_88};
  wire [63:0]   res_lo_hi_hi_88 = {dataGroup_7_88, dataGroup_6_88};
  wire [127:0]  res_lo_hi_88 = {res_lo_hi_hi_88, res_lo_hi_lo_88};
  wire [255:0]  res_lo_88 = {res_lo_hi_88, res_lo_lo_88};
  wire [63:0]   res_hi_lo_lo_88 = {dataGroup_9_88, dataGroup_8_88};
  wire [63:0]   res_hi_lo_hi_88 = {dataGroup_11_88, dataGroup_10_88};
  wire [127:0]  res_hi_lo_88 = {res_hi_lo_hi_88, res_hi_lo_lo_88};
  wire [63:0]   res_hi_hi_lo_88 = {dataGroup_13_88, dataGroup_12_88};
  wire [63:0]   res_hi_hi_hi_88 = {dataGroup_15_88, dataGroup_14_88};
  wire [127:0]  res_hi_hi_88 = {res_hi_hi_hi_88, res_hi_hi_lo_88};
  wire [255:0]  res_hi_88 = {res_hi_hi_88, res_hi_lo_88};
  wire [511:0]  res_169 = {res_hi_88, res_lo_88};
  wire [2047:0] dataGroup_lo_3728 = {dataGroup_lo_hi_3728, dataGroup_lo_lo_3728};
  wire [2047:0] dataGroup_hi_3728 = {dataGroup_hi_hi_3728, dataGroup_hi_lo_3728};
  wire [31:0]   dataGroup_0_89 = dataGroup_lo_3728[95:64];
  wire [2047:0] dataGroup_lo_3729 = {dataGroup_lo_hi_3729, dataGroup_lo_lo_3729};
  wire [2047:0] dataGroup_hi_3729 = {dataGroup_hi_hi_3729, dataGroup_hi_lo_3729};
  wire [31:0]   dataGroup_1_89 = dataGroup_lo_3729[287:256];
  wire [2047:0] dataGroup_lo_3730 = {dataGroup_lo_hi_3730, dataGroup_lo_lo_3730};
  wire [2047:0] dataGroup_hi_3730 = {dataGroup_hi_hi_3730, dataGroup_hi_lo_3730};
  wire [31:0]   dataGroup_2_89 = dataGroup_lo_3730[479:448];
  wire [2047:0] dataGroup_lo_3731 = {dataGroup_lo_hi_3731, dataGroup_lo_lo_3731};
  wire [2047:0] dataGroup_hi_3731 = {dataGroup_hi_hi_3731, dataGroup_hi_lo_3731};
  wire [31:0]   dataGroup_3_89 = dataGroup_lo_3731[671:640];
  wire [2047:0] dataGroup_lo_3732 = {dataGroup_lo_hi_3732, dataGroup_lo_lo_3732};
  wire [2047:0] dataGroup_hi_3732 = {dataGroup_hi_hi_3732, dataGroup_hi_lo_3732};
  wire [31:0]   dataGroup_4_89 = dataGroup_lo_3732[863:832];
  wire [2047:0] dataGroup_lo_3733 = {dataGroup_lo_hi_3733, dataGroup_lo_lo_3733};
  wire [2047:0] dataGroup_hi_3733 = {dataGroup_hi_hi_3733, dataGroup_hi_lo_3733};
  wire [31:0]   dataGroup_5_89 = dataGroup_lo_3733[1055:1024];
  wire [2047:0] dataGroup_lo_3734 = {dataGroup_lo_hi_3734, dataGroup_lo_lo_3734};
  wire [2047:0] dataGroup_hi_3734 = {dataGroup_hi_hi_3734, dataGroup_hi_lo_3734};
  wire [31:0]   dataGroup_6_89 = dataGroup_lo_3734[1247:1216];
  wire [2047:0] dataGroup_lo_3735 = {dataGroup_lo_hi_3735, dataGroup_lo_lo_3735};
  wire [2047:0] dataGroup_hi_3735 = {dataGroup_hi_hi_3735, dataGroup_hi_lo_3735};
  wire [31:0]   dataGroup_7_89 = dataGroup_lo_3735[1439:1408];
  wire [2047:0] dataGroup_lo_3736 = {dataGroup_lo_hi_3736, dataGroup_lo_lo_3736};
  wire [2047:0] dataGroup_hi_3736 = {dataGroup_hi_hi_3736, dataGroup_hi_lo_3736};
  wire [31:0]   dataGroup_8_89 = dataGroup_lo_3736[1631:1600];
  wire [2047:0] dataGroup_lo_3737 = {dataGroup_lo_hi_3737, dataGroup_lo_lo_3737};
  wire [2047:0] dataGroup_hi_3737 = {dataGroup_hi_hi_3737, dataGroup_hi_lo_3737};
  wire [31:0]   dataGroup_9_89 = dataGroup_lo_3737[1823:1792];
  wire [2047:0] dataGroup_lo_3738 = {dataGroup_lo_hi_3738, dataGroup_lo_lo_3738};
  wire [2047:0] dataGroup_hi_3738 = {dataGroup_hi_hi_3738, dataGroup_hi_lo_3738};
  wire [31:0]   dataGroup_10_89 = dataGroup_lo_3738[2015:1984];
  wire [2047:0] dataGroup_lo_3739 = {dataGroup_lo_hi_3739, dataGroup_lo_lo_3739};
  wire [2047:0] dataGroup_hi_3739 = {dataGroup_hi_hi_3739, dataGroup_hi_lo_3739};
  wire [31:0]   dataGroup_11_89 = dataGroup_hi_3739[159:128];
  wire [2047:0] dataGroup_lo_3740 = {dataGroup_lo_hi_3740, dataGroup_lo_lo_3740};
  wire [2047:0] dataGroup_hi_3740 = {dataGroup_hi_hi_3740, dataGroup_hi_lo_3740};
  wire [31:0]   dataGroup_12_89 = dataGroup_hi_3740[351:320];
  wire [2047:0] dataGroup_lo_3741 = {dataGroup_lo_hi_3741, dataGroup_lo_lo_3741};
  wire [2047:0] dataGroup_hi_3741 = {dataGroup_hi_hi_3741, dataGroup_hi_lo_3741};
  wire [31:0]   dataGroup_13_89 = dataGroup_hi_3741[543:512];
  wire [2047:0] dataGroup_lo_3742 = {dataGroup_lo_hi_3742, dataGroup_lo_lo_3742};
  wire [2047:0] dataGroup_hi_3742 = {dataGroup_hi_hi_3742, dataGroup_hi_lo_3742};
  wire [31:0]   dataGroup_14_89 = dataGroup_hi_3742[735:704];
  wire [2047:0] dataGroup_lo_3743 = {dataGroup_lo_hi_3743, dataGroup_lo_lo_3743};
  wire [2047:0] dataGroup_hi_3743 = {dataGroup_hi_hi_3743, dataGroup_hi_lo_3743};
  wire [31:0]   dataGroup_15_89 = dataGroup_hi_3743[927:896];
  wire [63:0]   res_lo_lo_lo_89 = {dataGroup_1_89, dataGroup_0_89};
  wire [63:0]   res_lo_lo_hi_89 = {dataGroup_3_89, dataGroup_2_89};
  wire [127:0]  res_lo_lo_89 = {res_lo_lo_hi_89, res_lo_lo_lo_89};
  wire [63:0]   res_lo_hi_lo_89 = {dataGroup_5_89, dataGroup_4_89};
  wire [63:0]   res_lo_hi_hi_89 = {dataGroup_7_89, dataGroup_6_89};
  wire [127:0]  res_lo_hi_89 = {res_lo_hi_hi_89, res_lo_hi_lo_89};
  wire [255:0]  res_lo_89 = {res_lo_hi_89, res_lo_lo_89};
  wire [63:0]   res_hi_lo_lo_89 = {dataGroup_9_89, dataGroup_8_89};
  wire [63:0]   res_hi_lo_hi_89 = {dataGroup_11_89, dataGroup_10_89};
  wire [127:0]  res_hi_lo_89 = {res_hi_lo_hi_89, res_hi_lo_lo_89};
  wire [63:0]   res_hi_hi_lo_89 = {dataGroup_13_89, dataGroup_12_89};
  wire [63:0]   res_hi_hi_hi_89 = {dataGroup_15_89, dataGroup_14_89};
  wire [127:0]  res_hi_hi_89 = {res_hi_hi_hi_89, res_hi_hi_lo_89};
  wire [255:0]  res_hi_89 = {res_hi_hi_89, res_hi_lo_89};
  wire [511:0]  res_170 = {res_hi_89, res_lo_89};
  wire [2047:0] dataGroup_lo_3744 = {dataGroup_lo_hi_3744, dataGroup_lo_lo_3744};
  wire [2047:0] dataGroup_hi_3744 = {dataGroup_hi_hi_3744, dataGroup_hi_lo_3744};
  wire [31:0]   dataGroup_0_90 = dataGroup_lo_3744[127:96];
  wire [2047:0] dataGroup_lo_3745 = {dataGroup_lo_hi_3745, dataGroup_lo_lo_3745};
  wire [2047:0] dataGroup_hi_3745 = {dataGroup_hi_hi_3745, dataGroup_hi_lo_3745};
  wire [31:0]   dataGroup_1_90 = dataGroup_lo_3745[319:288];
  wire [2047:0] dataGroup_lo_3746 = {dataGroup_lo_hi_3746, dataGroup_lo_lo_3746};
  wire [2047:0] dataGroup_hi_3746 = {dataGroup_hi_hi_3746, dataGroup_hi_lo_3746};
  wire [31:0]   dataGroup_2_90 = dataGroup_lo_3746[511:480];
  wire [2047:0] dataGroup_lo_3747 = {dataGroup_lo_hi_3747, dataGroup_lo_lo_3747};
  wire [2047:0] dataGroup_hi_3747 = {dataGroup_hi_hi_3747, dataGroup_hi_lo_3747};
  wire [31:0]   dataGroup_3_90 = dataGroup_lo_3747[703:672];
  wire [2047:0] dataGroup_lo_3748 = {dataGroup_lo_hi_3748, dataGroup_lo_lo_3748};
  wire [2047:0] dataGroup_hi_3748 = {dataGroup_hi_hi_3748, dataGroup_hi_lo_3748};
  wire [31:0]   dataGroup_4_90 = dataGroup_lo_3748[895:864];
  wire [2047:0] dataGroup_lo_3749 = {dataGroup_lo_hi_3749, dataGroup_lo_lo_3749};
  wire [2047:0] dataGroup_hi_3749 = {dataGroup_hi_hi_3749, dataGroup_hi_lo_3749};
  wire [31:0]   dataGroup_5_90 = dataGroup_lo_3749[1087:1056];
  wire [2047:0] dataGroup_lo_3750 = {dataGroup_lo_hi_3750, dataGroup_lo_lo_3750};
  wire [2047:0] dataGroup_hi_3750 = {dataGroup_hi_hi_3750, dataGroup_hi_lo_3750};
  wire [31:0]   dataGroup_6_90 = dataGroup_lo_3750[1279:1248];
  wire [2047:0] dataGroup_lo_3751 = {dataGroup_lo_hi_3751, dataGroup_lo_lo_3751};
  wire [2047:0] dataGroup_hi_3751 = {dataGroup_hi_hi_3751, dataGroup_hi_lo_3751};
  wire [31:0]   dataGroup_7_90 = dataGroup_lo_3751[1471:1440];
  wire [2047:0] dataGroup_lo_3752 = {dataGroup_lo_hi_3752, dataGroup_lo_lo_3752};
  wire [2047:0] dataGroup_hi_3752 = {dataGroup_hi_hi_3752, dataGroup_hi_lo_3752};
  wire [31:0]   dataGroup_8_90 = dataGroup_lo_3752[1663:1632];
  wire [2047:0] dataGroup_lo_3753 = {dataGroup_lo_hi_3753, dataGroup_lo_lo_3753};
  wire [2047:0] dataGroup_hi_3753 = {dataGroup_hi_hi_3753, dataGroup_hi_lo_3753};
  wire [31:0]   dataGroup_9_90 = dataGroup_lo_3753[1855:1824];
  wire [2047:0] dataGroup_lo_3754 = {dataGroup_lo_hi_3754, dataGroup_lo_lo_3754};
  wire [2047:0] dataGroup_hi_3754 = {dataGroup_hi_hi_3754, dataGroup_hi_lo_3754};
  wire [31:0]   dataGroup_10_90 = dataGroup_lo_3754[2047:2016];
  wire [2047:0] dataGroup_lo_3755 = {dataGroup_lo_hi_3755, dataGroup_lo_lo_3755};
  wire [2047:0] dataGroup_hi_3755 = {dataGroup_hi_hi_3755, dataGroup_hi_lo_3755};
  wire [31:0]   dataGroup_11_90 = dataGroup_hi_3755[191:160];
  wire [2047:0] dataGroup_lo_3756 = {dataGroup_lo_hi_3756, dataGroup_lo_lo_3756};
  wire [2047:0] dataGroup_hi_3756 = {dataGroup_hi_hi_3756, dataGroup_hi_lo_3756};
  wire [31:0]   dataGroup_12_90 = dataGroup_hi_3756[383:352];
  wire [2047:0] dataGroup_lo_3757 = {dataGroup_lo_hi_3757, dataGroup_lo_lo_3757};
  wire [2047:0] dataGroup_hi_3757 = {dataGroup_hi_hi_3757, dataGroup_hi_lo_3757};
  wire [31:0]   dataGroup_13_90 = dataGroup_hi_3757[575:544];
  wire [2047:0] dataGroup_lo_3758 = {dataGroup_lo_hi_3758, dataGroup_lo_lo_3758};
  wire [2047:0] dataGroup_hi_3758 = {dataGroup_hi_hi_3758, dataGroup_hi_lo_3758};
  wire [31:0]   dataGroup_14_90 = dataGroup_hi_3758[767:736];
  wire [2047:0] dataGroup_lo_3759 = {dataGroup_lo_hi_3759, dataGroup_lo_lo_3759};
  wire [2047:0] dataGroup_hi_3759 = {dataGroup_hi_hi_3759, dataGroup_hi_lo_3759};
  wire [31:0]   dataGroup_15_90 = dataGroup_hi_3759[959:928];
  wire [63:0]   res_lo_lo_lo_90 = {dataGroup_1_90, dataGroup_0_90};
  wire [63:0]   res_lo_lo_hi_90 = {dataGroup_3_90, dataGroup_2_90};
  wire [127:0]  res_lo_lo_90 = {res_lo_lo_hi_90, res_lo_lo_lo_90};
  wire [63:0]   res_lo_hi_lo_90 = {dataGroup_5_90, dataGroup_4_90};
  wire [63:0]   res_lo_hi_hi_90 = {dataGroup_7_90, dataGroup_6_90};
  wire [127:0]  res_lo_hi_90 = {res_lo_hi_hi_90, res_lo_hi_lo_90};
  wire [255:0]  res_lo_90 = {res_lo_hi_90, res_lo_lo_90};
  wire [63:0]   res_hi_lo_lo_90 = {dataGroup_9_90, dataGroup_8_90};
  wire [63:0]   res_hi_lo_hi_90 = {dataGroup_11_90, dataGroup_10_90};
  wire [127:0]  res_hi_lo_90 = {res_hi_lo_hi_90, res_hi_lo_lo_90};
  wire [63:0]   res_hi_hi_lo_90 = {dataGroup_13_90, dataGroup_12_90};
  wire [63:0]   res_hi_hi_hi_90 = {dataGroup_15_90, dataGroup_14_90};
  wire [127:0]  res_hi_hi_90 = {res_hi_hi_hi_90, res_hi_hi_lo_90};
  wire [255:0]  res_hi_90 = {res_hi_hi_90, res_hi_lo_90};
  wire [511:0]  res_171 = {res_hi_90, res_lo_90};
  wire [2047:0] dataGroup_lo_3760 = {dataGroup_lo_hi_3760, dataGroup_lo_lo_3760};
  wire [2047:0] dataGroup_hi_3760 = {dataGroup_hi_hi_3760, dataGroup_hi_lo_3760};
  wire [31:0]   dataGroup_0_91 = dataGroup_lo_3760[159:128];
  wire [2047:0] dataGroup_lo_3761 = {dataGroup_lo_hi_3761, dataGroup_lo_lo_3761};
  wire [2047:0] dataGroup_hi_3761 = {dataGroup_hi_hi_3761, dataGroup_hi_lo_3761};
  wire [31:0]   dataGroup_1_91 = dataGroup_lo_3761[351:320];
  wire [2047:0] dataGroup_lo_3762 = {dataGroup_lo_hi_3762, dataGroup_lo_lo_3762};
  wire [2047:0] dataGroup_hi_3762 = {dataGroup_hi_hi_3762, dataGroup_hi_lo_3762};
  wire [31:0]   dataGroup_2_91 = dataGroup_lo_3762[543:512];
  wire [2047:0] dataGroup_lo_3763 = {dataGroup_lo_hi_3763, dataGroup_lo_lo_3763};
  wire [2047:0] dataGroup_hi_3763 = {dataGroup_hi_hi_3763, dataGroup_hi_lo_3763};
  wire [31:0]   dataGroup_3_91 = dataGroup_lo_3763[735:704];
  wire [2047:0] dataGroup_lo_3764 = {dataGroup_lo_hi_3764, dataGroup_lo_lo_3764};
  wire [2047:0] dataGroup_hi_3764 = {dataGroup_hi_hi_3764, dataGroup_hi_lo_3764};
  wire [31:0]   dataGroup_4_91 = dataGroup_lo_3764[927:896];
  wire [2047:0] dataGroup_lo_3765 = {dataGroup_lo_hi_3765, dataGroup_lo_lo_3765};
  wire [2047:0] dataGroup_hi_3765 = {dataGroup_hi_hi_3765, dataGroup_hi_lo_3765};
  wire [31:0]   dataGroup_5_91 = dataGroup_lo_3765[1119:1088];
  wire [2047:0] dataGroup_lo_3766 = {dataGroup_lo_hi_3766, dataGroup_lo_lo_3766};
  wire [2047:0] dataGroup_hi_3766 = {dataGroup_hi_hi_3766, dataGroup_hi_lo_3766};
  wire [31:0]   dataGroup_6_91 = dataGroup_lo_3766[1311:1280];
  wire [2047:0] dataGroup_lo_3767 = {dataGroup_lo_hi_3767, dataGroup_lo_lo_3767};
  wire [2047:0] dataGroup_hi_3767 = {dataGroup_hi_hi_3767, dataGroup_hi_lo_3767};
  wire [31:0]   dataGroup_7_91 = dataGroup_lo_3767[1503:1472];
  wire [2047:0] dataGroup_lo_3768 = {dataGroup_lo_hi_3768, dataGroup_lo_lo_3768};
  wire [2047:0] dataGroup_hi_3768 = {dataGroup_hi_hi_3768, dataGroup_hi_lo_3768};
  wire [31:0]   dataGroup_8_91 = dataGroup_lo_3768[1695:1664];
  wire [2047:0] dataGroup_lo_3769 = {dataGroup_lo_hi_3769, dataGroup_lo_lo_3769};
  wire [2047:0] dataGroup_hi_3769 = {dataGroup_hi_hi_3769, dataGroup_hi_lo_3769};
  wire [31:0]   dataGroup_9_91 = dataGroup_lo_3769[1887:1856];
  wire [2047:0] dataGroup_lo_3770 = {dataGroup_lo_hi_3770, dataGroup_lo_lo_3770};
  wire [2047:0] dataGroup_hi_3770 = {dataGroup_hi_hi_3770, dataGroup_hi_lo_3770};
  wire [31:0]   dataGroup_10_91 = dataGroup_hi_3770[31:0];
  wire [2047:0] dataGroup_lo_3771 = {dataGroup_lo_hi_3771, dataGroup_lo_lo_3771};
  wire [2047:0] dataGroup_hi_3771 = {dataGroup_hi_hi_3771, dataGroup_hi_lo_3771};
  wire [31:0]   dataGroup_11_91 = dataGroup_hi_3771[223:192];
  wire [2047:0] dataGroup_lo_3772 = {dataGroup_lo_hi_3772, dataGroup_lo_lo_3772};
  wire [2047:0] dataGroup_hi_3772 = {dataGroup_hi_hi_3772, dataGroup_hi_lo_3772};
  wire [31:0]   dataGroup_12_91 = dataGroup_hi_3772[415:384];
  wire [2047:0] dataGroup_lo_3773 = {dataGroup_lo_hi_3773, dataGroup_lo_lo_3773};
  wire [2047:0] dataGroup_hi_3773 = {dataGroup_hi_hi_3773, dataGroup_hi_lo_3773};
  wire [31:0]   dataGroup_13_91 = dataGroup_hi_3773[607:576];
  wire [2047:0] dataGroup_lo_3774 = {dataGroup_lo_hi_3774, dataGroup_lo_lo_3774};
  wire [2047:0] dataGroup_hi_3774 = {dataGroup_hi_hi_3774, dataGroup_hi_lo_3774};
  wire [31:0]   dataGroup_14_91 = dataGroup_hi_3774[799:768];
  wire [2047:0] dataGroup_lo_3775 = {dataGroup_lo_hi_3775, dataGroup_lo_lo_3775};
  wire [2047:0] dataGroup_hi_3775 = {dataGroup_hi_hi_3775, dataGroup_hi_lo_3775};
  wire [31:0]   dataGroup_15_91 = dataGroup_hi_3775[991:960];
  wire [63:0]   res_lo_lo_lo_91 = {dataGroup_1_91, dataGroup_0_91};
  wire [63:0]   res_lo_lo_hi_91 = {dataGroup_3_91, dataGroup_2_91};
  wire [127:0]  res_lo_lo_91 = {res_lo_lo_hi_91, res_lo_lo_lo_91};
  wire [63:0]   res_lo_hi_lo_91 = {dataGroup_5_91, dataGroup_4_91};
  wire [63:0]   res_lo_hi_hi_91 = {dataGroup_7_91, dataGroup_6_91};
  wire [127:0]  res_lo_hi_91 = {res_lo_hi_hi_91, res_lo_hi_lo_91};
  wire [255:0]  res_lo_91 = {res_lo_hi_91, res_lo_lo_91};
  wire [63:0]   res_hi_lo_lo_91 = {dataGroup_9_91, dataGroup_8_91};
  wire [63:0]   res_hi_lo_hi_91 = {dataGroup_11_91, dataGroup_10_91};
  wire [127:0]  res_hi_lo_91 = {res_hi_lo_hi_91, res_hi_lo_lo_91};
  wire [63:0]   res_hi_hi_lo_91 = {dataGroup_13_91, dataGroup_12_91};
  wire [63:0]   res_hi_hi_hi_91 = {dataGroup_15_91, dataGroup_14_91};
  wire [127:0]  res_hi_hi_91 = {res_hi_hi_hi_91, res_hi_hi_lo_91};
  wire [255:0]  res_hi_91 = {res_hi_hi_91, res_hi_lo_91};
  wire [511:0]  res_172 = {res_hi_91, res_lo_91};
  wire [2047:0] dataGroup_lo_3776 = {dataGroup_lo_hi_3776, dataGroup_lo_lo_3776};
  wire [2047:0] dataGroup_hi_3776 = {dataGroup_hi_hi_3776, dataGroup_hi_lo_3776};
  wire [31:0]   dataGroup_0_92 = dataGroup_lo_3776[191:160];
  wire [2047:0] dataGroup_lo_3777 = {dataGroup_lo_hi_3777, dataGroup_lo_lo_3777};
  wire [2047:0] dataGroup_hi_3777 = {dataGroup_hi_hi_3777, dataGroup_hi_lo_3777};
  wire [31:0]   dataGroup_1_92 = dataGroup_lo_3777[383:352];
  wire [2047:0] dataGroup_lo_3778 = {dataGroup_lo_hi_3778, dataGroup_lo_lo_3778};
  wire [2047:0] dataGroup_hi_3778 = {dataGroup_hi_hi_3778, dataGroup_hi_lo_3778};
  wire [31:0]   dataGroup_2_92 = dataGroup_lo_3778[575:544];
  wire [2047:0] dataGroup_lo_3779 = {dataGroup_lo_hi_3779, dataGroup_lo_lo_3779};
  wire [2047:0] dataGroup_hi_3779 = {dataGroup_hi_hi_3779, dataGroup_hi_lo_3779};
  wire [31:0]   dataGroup_3_92 = dataGroup_lo_3779[767:736];
  wire [2047:0] dataGroup_lo_3780 = {dataGroup_lo_hi_3780, dataGroup_lo_lo_3780};
  wire [2047:0] dataGroup_hi_3780 = {dataGroup_hi_hi_3780, dataGroup_hi_lo_3780};
  wire [31:0]   dataGroup_4_92 = dataGroup_lo_3780[959:928];
  wire [2047:0] dataGroup_lo_3781 = {dataGroup_lo_hi_3781, dataGroup_lo_lo_3781};
  wire [2047:0] dataGroup_hi_3781 = {dataGroup_hi_hi_3781, dataGroup_hi_lo_3781};
  wire [31:0]   dataGroup_5_92 = dataGroup_lo_3781[1151:1120];
  wire [2047:0] dataGroup_lo_3782 = {dataGroup_lo_hi_3782, dataGroup_lo_lo_3782};
  wire [2047:0] dataGroup_hi_3782 = {dataGroup_hi_hi_3782, dataGroup_hi_lo_3782};
  wire [31:0]   dataGroup_6_92 = dataGroup_lo_3782[1343:1312];
  wire [2047:0] dataGroup_lo_3783 = {dataGroup_lo_hi_3783, dataGroup_lo_lo_3783};
  wire [2047:0] dataGroup_hi_3783 = {dataGroup_hi_hi_3783, dataGroup_hi_lo_3783};
  wire [31:0]   dataGroup_7_92 = dataGroup_lo_3783[1535:1504];
  wire [2047:0] dataGroup_lo_3784 = {dataGroup_lo_hi_3784, dataGroup_lo_lo_3784};
  wire [2047:0] dataGroup_hi_3784 = {dataGroup_hi_hi_3784, dataGroup_hi_lo_3784};
  wire [31:0]   dataGroup_8_92 = dataGroup_lo_3784[1727:1696];
  wire [2047:0] dataGroup_lo_3785 = {dataGroup_lo_hi_3785, dataGroup_lo_lo_3785};
  wire [2047:0] dataGroup_hi_3785 = {dataGroup_hi_hi_3785, dataGroup_hi_lo_3785};
  wire [31:0]   dataGroup_9_92 = dataGroup_lo_3785[1919:1888];
  wire [2047:0] dataGroup_lo_3786 = {dataGroup_lo_hi_3786, dataGroup_lo_lo_3786};
  wire [2047:0] dataGroup_hi_3786 = {dataGroup_hi_hi_3786, dataGroup_hi_lo_3786};
  wire [31:0]   dataGroup_10_92 = dataGroup_hi_3786[63:32];
  wire [2047:0] dataGroup_lo_3787 = {dataGroup_lo_hi_3787, dataGroup_lo_lo_3787};
  wire [2047:0] dataGroup_hi_3787 = {dataGroup_hi_hi_3787, dataGroup_hi_lo_3787};
  wire [31:0]   dataGroup_11_92 = dataGroup_hi_3787[255:224];
  wire [2047:0] dataGroup_lo_3788 = {dataGroup_lo_hi_3788, dataGroup_lo_lo_3788};
  wire [2047:0] dataGroup_hi_3788 = {dataGroup_hi_hi_3788, dataGroup_hi_lo_3788};
  wire [31:0]   dataGroup_12_92 = dataGroup_hi_3788[447:416];
  wire [2047:0] dataGroup_lo_3789 = {dataGroup_lo_hi_3789, dataGroup_lo_lo_3789};
  wire [2047:0] dataGroup_hi_3789 = {dataGroup_hi_hi_3789, dataGroup_hi_lo_3789};
  wire [31:0]   dataGroup_13_92 = dataGroup_hi_3789[639:608];
  wire [2047:0] dataGroup_lo_3790 = {dataGroup_lo_hi_3790, dataGroup_lo_lo_3790};
  wire [2047:0] dataGroup_hi_3790 = {dataGroup_hi_hi_3790, dataGroup_hi_lo_3790};
  wire [31:0]   dataGroup_14_92 = dataGroup_hi_3790[831:800];
  wire [2047:0] dataGroup_lo_3791 = {dataGroup_lo_hi_3791, dataGroup_lo_lo_3791};
  wire [2047:0] dataGroup_hi_3791 = {dataGroup_hi_hi_3791, dataGroup_hi_lo_3791};
  wire [31:0]   dataGroup_15_92 = dataGroup_hi_3791[1023:992];
  wire [63:0]   res_lo_lo_lo_92 = {dataGroup_1_92, dataGroup_0_92};
  wire [63:0]   res_lo_lo_hi_92 = {dataGroup_3_92, dataGroup_2_92};
  wire [127:0]  res_lo_lo_92 = {res_lo_lo_hi_92, res_lo_lo_lo_92};
  wire [63:0]   res_lo_hi_lo_92 = {dataGroup_5_92, dataGroup_4_92};
  wire [63:0]   res_lo_hi_hi_92 = {dataGroup_7_92, dataGroup_6_92};
  wire [127:0]  res_lo_hi_92 = {res_lo_hi_hi_92, res_lo_hi_lo_92};
  wire [255:0]  res_lo_92 = {res_lo_hi_92, res_lo_lo_92};
  wire [63:0]   res_hi_lo_lo_92 = {dataGroup_9_92, dataGroup_8_92};
  wire [63:0]   res_hi_lo_hi_92 = {dataGroup_11_92, dataGroup_10_92};
  wire [127:0]  res_hi_lo_92 = {res_hi_lo_hi_92, res_hi_lo_lo_92};
  wire [63:0]   res_hi_hi_lo_92 = {dataGroup_13_92, dataGroup_12_92};
  wire [63:0]   res_hi_hi_hi_92 = {dataGroup_15_92, dataGroup_14_92};
  wire [127:0]  res_hi_hi_92 = {res_hi_hi_hi_92, res_hi_hi_lo_92};
  wire [255:0]  res_hi_92 = {res_hi_hi_92, res_hi_lo_92};
  wire [511:0]  res_173 = {res_hi_92, res_lo_92};
  wire [1023:0] lo_lo_21 = {res_169, res_168};
  wire [1023:0] lo_hi_21 = {res_171, res_170};
  wire [2047:0] lo_21 = {lo_hi_21, lo_lo_21};
  wire [1023:0] hi_lo_21 = {res_173, res_172};
  wire [2047:0] hi_21 = {1024'h0, hi_lo_21};
  wire [4095:0] regroupLoadData_2_5 = {hi_21, lo_21};
  wire [2047:0] dataGroup_lo_3792 = {dataGroup_lo_hi_3792, dataGroup_lo_lo_3792};
  wire [2047:0] dataGroup_hi_3792 = {dataGroup_hi_hi_3792, dataGroup_hi_lo_3792};
  wire [31:0]   dataGroup_0_93 = dataGroup_lo_3792[31:0];
  wire [2047:0] dataGroup_lo_3793 = {dataGroup_lo_hi_3793, dataGroup_lo_lo_3793};
  wire [2047:0] dataGroup_hi_3793 = {dataGroup_hi_hi_3793, dataGroup_hi_lo_3793};
  wire [31:0]   dataGroup_1_93 = dataGroup_lo_3793[255:224];
  wire [2047:0] dataGroup_lo_3794 = {dataGroup_lo_hi_3794, dataGroup_lo_lo_3794};
  wire [2047:0] dataGroup_hi_3794 = {dataGroup_hi_hi_3794, dataGroup_hi_lo_3794};
  wire [31:0]   dataGroup_2_93 = dataGroup_lo_3794[479:448];
  wire [2047:0] dataGroup_lo_3795 = {dataGroup_lo_hi_3795, dataGroup_lo_lo_3795};
  wire [2047:0] dataGroup_hi_3795 = {dataGroup_hi_hi_3795, dataGroup_hi_lo_3795};
  wire [31:0]   dataGroup_3_93 = dataGroup_lo_3795[703:672];
  wire [2047:0] dataGroup_lo_3796 = {dataGroup_lo_hi_3796, dataGroup_lo_lo_3796};
  wire [2047:0] dataGroup_hi_3796 = {dataGroup_hi_hi_3796, dataGroup_hi_lo_3796};
  wire [31:0]   dataGroup_4_93 = dataGroup_lo_3796[927:896];
  wire [2047:0] dataGroup_lo_3797 = {dataGroup_lo_hi_3797, dataGroup_lo_lo_3797};
  wire [2047:0] dataGroup_hi_3797 = {dataGroup_hi_hi_3797, dataGroup_hi_lo_3797};
  wire [31:0]   dataGroup_5_93 = dataGroup_lo_3797[1151:1120];
  wire [2047:0] dataGroup_lo_3798 = {dataGroup_lo_hi_3798, dataGroup_lo_lo_3798};
  wire [2047:0] dataGroup_hi_3798 = {dataGroup_hi_hi_3798, dataGroup_hi_lo_3798};
  wire [31:0]   dataGroup_6_93 = dataGroup_lo_3798[1375:1344];
  wire [2047:0] dataGroup_lo_3799 = {dataGroup_lo_hi_3799, dataGroup_lo_lo_3799};
  wire [2047:0] dataGroup_hi_3799 = {dataGroup_hi_hi_3799, dataGroup_hi_lo_3799};
  wire [31:0]   dataGroup_7_93 = dataGroup_lo_3799[1599:1568];
  wire [2047:0] dataGroup_lo_3800 = {dataGroup_lo_hi_3800, dataGroup_lo_lo_3800};
  wire [2047:0] dataGroup_hi_3800 = {dataGroup_hi_hi_3800, dataGroup_hi_lo_3800};
  wire [31:0]   dataGroup_8_93 = dataGroup_lo_3800[1823:1792];
  wire [2047:0] dataGroup_lo_3801 = {dataGroup_lo_hi_3801, dataGroup_lo_lo_3801};
  wire [2047:0] dataGroup_hi_3801 = {dataGroup_hi_hi_3801, dataGroup_hi_lo_3801};
  wire [31:0]   dataGroup_9_93 = dataGroup_lo_3801[2047:2016];
  wire [2047:0] dataGroup_lo_3802 = {dataGroup_lo_hi_3802, dataGroup_lo_lo_3802};
  wire [2047:0] dataGroup_hi_3802 = {dataGroup_hi_hi_3802, dataGroup_hi_lo_3802};
  wire [31:0]   dataGroup_10_93 = dataGroup_hi_3802[223:192];
  wire [2047:0] dataGroup_lo_3803 = {dataGroup_lo_hi_3803, dataGroup_lo_lo_3803};
  wire [2047:0] dataGroup_hi_3803 = {dataGroup_hi_hi_3803, dataGroup_hi_lo_3803};
  wire [31:0]   dataGroup_11_93 = dataGroup_hi_3803[447:416];
  wire [2047:0] dataGroup_lo_3804 = {dataGroup_lo_hi_3804, dataGroup_lo_lo_3804};
  wire [2047:0] dataGroup_hi_3804 = {dataGroup_hi_hi_3804, dataGroup_hi_lo_3804};
  wire [31:0]   dataGroup_12_93 = dataGroup_hi_3804[671:640];
  wire [2047:0] dataGroup_lo_3805 = {dataGroup_lo_hi_3805, dataGroup_lo_lo_3805};
  wire [2047:0] dataGroup_hi_3805 = {dataGroup_hi_hi_3805, dataGroup_hi_lo_3805};
  wire [31:0]   dataGroup_13_93 = dataGroup_hi_3805[895:864];
  wire [2047:0] dataGroup_lo_3806 = {dataGroup_lo_hi_3806, dataGroup_lo_lo_3806};
  wire [2047:0] dataGroup_hi_3806 = {dataGroup_hi_hi_3806, dataGroup_hi_lo_3806};
  wire [31:0]   dataGroup_14_93 = dataGroup_hi_3806[1119:1088];
  wire [2047:0] dataGroup_lo_3807 = {dataGroup_lo_hi_3807, dataGroup_lo_lo_3807};
  wire [2047:0] dataGroup_hi_3807 = {dataGroup_hi_hi_3807, dataGroup_hi_lo_3807};
  wire [31:0]   dataGroup_15_93 = dataGroup_hi_3807[1343:1312];
  wire [63:0]   res_lo_lo_lo_93 = {dataGroup_1_93, dataGroup_0_93};
  wire [63:0]   res_lo_lo_hi_93 = {dataGroup_3_93, dataGroup_2_93};
  wire [127:0]  res_lo_lo_93 = {res_lo_lo_hi_93, res_lo_lo_lo_93};
  wire [63:0]   res_lo_hi_lo_93 = {dataGroup_5_93, dataGroup_4_93};
  wire [63:0]   res_lo_hi_hi_93 = {dataGroup_7_93, dataGroup_6_93};
  wire [127:0]  res_lo_hi_93 = {res_lo_hi_hi_93, res_lo_hi_lo_93};
  wire [255:0]  res_lo_93 = {res_lo_hi_93, res_lo_lo_93};
  wire [63:0]   res_hi_lo_lo_93 = {dataGroup_9_93, dataGroup_8_93};
  wire [63:0]   res_hi_lo_hi_93 = {dataGroup_11_93, dataGroup_10_93};
  wire [127:0]  res_hi_lo_93 = {res_hi_lo_hi_93, res_hi_lo_lo_93};
  wire [63:0]   res_hi_hi_lo_93 = {dataGroup_13_93, dataGroup_12_93};
  wire [63:0]   res_hi_hi_hi_93 = {dataGroup_15_93, dataGroup_14_93};
  wire [127:0]  res_hi_hi_93 = {res_hi_hi_hi_93, res_hi_hi_lo_93};
  wire [255:0]  res_hi_93 = {res_hi_hi_93, res_hi_lo_93};
  wire [511:0]  res_176 = {res_hi_93, res_lo_93};
  wire [2047:0] dataGroup_lo_3808 = {dataGroup_lo_hi_3808, dataGroup_lo_lo_3808};
  wire [2047:0] dataGroup_hi_3808 = {dataGroup_hi_hi_3808, dataGroup_hi_lo_3808};
  wire [31:0]   dataGroup_0_94 = dataGroup_lo_3808[63:32];
  wire [2047:0] dataGroup_lo_3809 = {dataGroup_lo_hi_3809, dataGroup_lo_lo_3809};
  wire [2047:0] dataGroup_hi_3809 = {dataGroup_hi_hi_3809, dataGroup_hi_lo_3809};
  wire [31:0]   dataGroup_1_94 = dataGroup_lo_3809[287:256];
  wire [2047:0] dataGroup_lo_3810 = {dataGroup_lo_hi_3810, dataGroup_lo_lo_3810};
  wire [2047:0] dataGroup_hi_3810 = {dataGroup_hi_hi_3810, dataGroup_hi_lo_3810};
  wire [31:0]   dataGroup_2_94 = dataGroup_lo_3810[511:480];
  wire [2047:0] dataGroup_lo_3811 = {dataGroup_lo_hi_3811, dataGroup_lo_lo_3811};
  wire [2047:0] dataGroup_hi_3811 = {dataGroup_hi_hi_3811, dataGroup_hi_lo_3811};
  wire [31:0]   dataGroup_3_94 = dataGroup_lo_3811[735:704];
  wire [2047:0] dataGroup_lo_3812 = {dataGroup_lo_hi_3812, dataGroup_lo_lo_3812};
  wire [2047:0] dataGroup_hi_3812 = {dataGroup_hi_hi_3812, dataGroup_hi_lo_3812};
  wire [31:0]   dataGroup_4_94 = dataGroup_lo_3812[959:928];
  wire [2047:0] dataGroup_lo_3813 = {dataGroup_lo_hi_3813, dataGroup_lo_lo_3813};
  wire [2047:0] dataGroup_hi_3813 = {dataGroup_hi_hi_3813, dataGroup_hi_lo_3813};
  wire [31:0]   dataGroup_5_94 = dataGroup_lo_3813[1183:1152];
  wire [2047:0] dataGroup_lo_3814 = {dataGroup_lo_hi_3814, dataGroup_lo_lo_3814};
  wire [2047:0] dataGroup_hi_3814 = {dataGroup_hi_hi_3814, dataGroup_hi_lo_3814};
  wire [31:0]   dataGroup_6_94 = dataGroup_lo_3814[1407:1376];
  wire [2047:0] dataGroup_lo_3815 = {dataGroup_lo_hi_3815, dataGroup_lo_lo_3815};
  wire [2047:0] dataGroup_hi_3815 = {dataGroup_hi_hi_3815, dataGroup_hi_lo_3815};
  wire [31:0]   dataGroup_7_94 = dataGroup_lo_3815[1631:1600];
  wire [2047:0] dataGroup_lo_3816 = {dataGroup_lo_hi_3816, dataGroup_lo_lo_3816};
  wire [2047:0] dataGroup_hi_3816 = {dataGroup_hi_hi_3816, dataGroup_hi_lo_3816};
  wire [31:0]   dataGroup_8_94 = dataGroup_lo_3816[1855:1824];
  wire [2047:0] dataGroup_lo_3817 = {dataGroup_lo_hi_3817, dataGroup_lo_lo_3817};
  wire [2047:0] dataGroup_hi_3817 = {dataGroup_hi_hi_3817, dataGroup_hi_lo_3817};
  wire [31:0]   dataGroup_9_94 = dataGroup_hi_3817[31:0];
  wire [2047:0] dataGroup_lo_3818 = {dataGroup_lo_hi_3818, dataGroup_lo_lo_3818};
  wire [2047:0] dataGroup_hi_3818 = {dataGroup_hi_hi_3818, dataGroup_hi_lo_3818};
  wire [31:0]   dataGroup_10_94 = dataGroup_hi_3818[255:224];
  wire [2047:0] dataGroup_lo_3819 = {dataGroup_lo_hi_3819, dataGroup_lo_lo_3819};
  wire [2047:0] dataGroup_hi_3819 = {dataGroup_hi_hi_3819, dataGroup_hi_lo_3819};
  wire [31:0]   dataGroup_11_94 = dataGroup_hi_3819[479:448];
  wire [2047:0] dataGroup_lo_3820 = {dataGroup_lo_hi_3820, dataGroup_lo_lo_3820};
  wire [2047:0] dataGroup_hi_3820 = {dataGroup_hi_hi_3820, dataGroup_hi_lo_3820};
  wire [31:0]   dataGroup_12_94 = dataGroup_hi_3820[703:672];
  wire [2047:0] dataGroup_lo_3821 = {dataGroup_lo_hi_3821, dataGroup_lo_lo_3821};
  wire [2047:0] dataGroup_hi_3821 = {dataGroup_hi_hi_3821, dataGroup_hi_lo_3821};
  wire [31:0]   dataGroup_13_94 = dataGroup_hi_3821[927:896];
  wire [2047:0] dataGroup_lo_3822 = {dataGroup_lo_hi_3822, dataGroup_lo_lo_3822};
  wire [2047:0] dataGroup_hi_3822 = {dataGroup_hi_hi_3822, dataGroup_hi_lo_3822};
  wire [31:0]   dataGroup_14_94 = dataGroup_hi_3822[1151:1120];
  wire [2047:0] dataGroup_lo_3823 = {dataGroup_lo_hi_3823, dataGroup_lo_lo_3823};
  wire [2047:0] dataGroup_hi_3823 = {dataGroup_hi_hi_3823, dataGroup_hi_lo_3823};
  wire [31:0]   dataGroup_15_94 = dataGroup_hi_3823[1375:1344];
  wire [63:0]   res_lo_lo_lo_94 = {dataGroup_1_94, dataGroup_0_94};
  wire [63:0]   res_lo_lo_hi_94 = {dataGroup_3_94, dataGroup_2_94};
  wire [127:0]  res_lo_lo_94 = {res_lo_lo_hi_94, res_lo_lo_lo_94};
  wire [63:0]   res_lo_hi_lo_94 = {dataGroup_5_94, dataGroup_4_94};
  wire [63:0]   res_lo_hi_hi_94 = {dataGroup_7_94, dataGroup_6_94};
  wire [127:0]  res_lo_hi_94 = {res_lo_hi_hi_94, res_lo_hi_lo_94};
  wire [255:0]  res_lo_94 = {res_lo_hi_94, res_lo_lo_94};
  wire [63:0]   res_hi_lo_lo_94 = {dataGroup_9_94, dataGroup_8_94};
  wire [63:0]   res_hi_lo_hi_94 = {dataGroup_11_94, dataGroup_10_94};
  wire [127:0]  res_hi_lo_94 = {res_hi_lo_hi_94, res_hi_lo_lo_94};
  wire [63:0]   res_hi_hi_lo_94 = {dataGroup_13_94, dataGroup_12_94};
  wire [63:0]   res_hi_hi_hi_94 = {dataGroup_15_94, dataGroup_14_94};
  wire [127:0]  res_hi_hi_94 = {res_hi_hi_hi_94, res_hi_hi_lo_94};
  wire [255:0]  res_hi_94 = {res_hi_hi_94, res_hi_lo_94};
  wire [511:0]  res_177 = {res_hi_94, res_lo_94};
  wire [2047:0] dataGroup_lo_3824 = {dataGroup_lo_hi_3824, dataGroup_lo_lo_3824};
  wire [2047:0] dataGroup_hi_3824 = {dataGroup_hi_hi_3824, dataGroup_hi_lo_3824};
  wire [31:0]   dataGroup_0_95 = dataGroup_lo_3824[95:64];
  wire [2047:0] dataGroup_lo_3825 = {dataGroup_lo_hi_3825, dataGroup_lo_lo_3825};
  wire [2047:0] dataGroup_hi_3825 = {dataGroup_hi_hi_3825, dataGroup_hi_lo_3825};
  wire [31:0]   dataGroup_1_95 = dataGroup_lo_3825[319:288];
  wire [2047:0] dataGroup_lo_3826 = {dataGroup_lo_hi_3826, dataGroup_lo_lo_3826};
  wire [2047:0] dataGroup_hi_3826 = {dataGroup_hi_hi_3826, dataGroup_hi_lo_3826};
  wire [31:0]   dataGroup_2_95 = dataGroup_lo_3826[543:512];
  wire [2047:0] dataGroup_lo_3827 = {dataGroup_lo_hi_3827, dataGroup_lo_lo_3827};
  wire [2047:0] dataGroup_hi_3827 = {dataGroup_hi_hi_3827, dataGroup_hi_lo_3827};
  wire [31:0]   dataGroup_3_95 = dataGroup_lo_3827[767:736];
  wire [2047:0] dataGroup_lo_3828 = {dataGroup_lo_hi_3828, dataGroup_lo_lo_3828};
  wire [2047:0] dataGroup_hi_3828 = {dataGroup_hi_hi_3828, dataGroup_hi_lo_3828};
  wire [31:0]   dataGroup_4_95 = dataGroup_lo_3828[991:960];
  wire [2047:0] dataGroup_lo_3829 = {dataGroup_lo_hi_3829, dataGroup_lo_lo_3829};
  wire [2047:0] dataGroup_hi_3829 = {dataGroup_hi_hi_3829, dataGroup_hi_lo_3829};
  wire [31:0]   dataGroup_5_95 = dataGroup_lo_3829[1215:1184];
  wire [2047:0] dataGroup_lo_3830 = {dataGroup_lo_hi_3830, dataGroup_lo_lo_3830};
  wire [2047:0] dataGroup_hi_3830 = {dataGroup_hi_hi_3830, dataGroup_hi_lo_3830};
  wire [31:0]   dataGroup_6_95 = dataGroup_lo_3830[1439:1408];
  wire [2047:0] dataGroup_lo_3831 = {dataGroup_lo_hi_3831, dataGroup_lo_lo_3831};
  wire [2047:0] dataGroup_hi_3831 = {dataGroup_hi_hi_3831, dataGroup_hi_lo_3831};
  wire [31:0]   dataGroup_7_95 = dataGroup_lo_3831[1663:1632];
  wire [2047:0] dataGroup_lo_3832 = {dataGroup_lo_hi_3832, dataGroup_lo_lo_3832};
  wire [2047:0] dataGroup_hi_3832 = {dataGroup_hi_hi_3832, dataGroup_hi_lo_3832};
  wire [31:0]   dataGroup_8_95 = dataGroup_lo_3832[1887:1856];
  wire [2047:0] dataGroup_lo_3833 = {dataGroup_lo_hi_3833, dataGroup_lo_lo_3833};
  wire [2047:0] dataGroup_hi_3833 = {dataGroup_hi_hi_3833, dataGroup_hi_lo_3833};
  wire [31:0]   dataGroup_9_95 = dataGroup_hi_3833[63:32];
  wire [2047:0] dataGroup_lo_3834 = {dataGroup_lo_hi_3834, dataGroup_lo_lo_3834};
  wire [2047:0] dataGroup_hi_3834 = {dataGroup_hi_hi_3834, dataGroup_hi_lo_3834};
  wire [31:0]   dataGroup_10_95 = dataGroup_hi_3834[287:256];
  wire [2047:0] dataGroup_lo_3835 = {dataGroup_lo_hi_3835, dataGroup_lo_lo_3835};
  wire [2047:0] dataGroup_hi_3835 = {dataGroup_hi_hi_3835, dataGroup_hi_lo_3835};
  wire [31:0]   dataGroup_11_95 = dataGroup_hi_3835[511:480];
  wire [2047:0] dataGroup_lo_3836 = {dataGroup_lo_hi_3836, dataGroup_lo_lo_3836};
  wire [2047:0] dataGroup_hi_3836 = {dataGroup_hi_hi_3836, dataGroup_hi_lo_3836};
  wire [31:0]   dataGroup_12_95 = dataGroup_hi_3836[735:704];
  wire [2047:0] dataGroup_lo_3837 = {dataGroup_lo_hi_3837, dataGroup_lo_lo_3837};
  wire [2047:0] dataGroup_hi_3837 = {dataGroup_hi_hi_3837, dataGroup_hi_lo_3837};
  wire [31:0]   dataGroup_13_95 = dataGroup_hi_3837[959:928];
  wire [2047:0] dataGroup_lo_3838 = {dataGroup_lo_hi_3838, dataGroup_lo_lo_3838};
  wire [2047:0] dataGroup_hi_3838 = {dataGroup_hi_hi_3838, dataGroup_hi_lo_3838};
  wire [31:0]   dataGroup_14_95 = dataGroup_hi_3838[1183:1152];
  wire [2047:0] dataGroup_lo_3839 = {dataGroup_lo_hi_3839, dataGroup_lo_lo_3839};
  wire [2047:0] dataGroup_hi_3839 = {dataGroup_hi_hi_3839, dataGroup_hi_lo_3839};
  wire [31:0]   dataGroup_15_95 = dataGroup_hi_3839[1407:1376];
  wire [63:0]   res_lo_lo_lo_95 = {dataGroup_1_95, dataGroup_0_95};
  wire [63:0]   res_lo_lo_hi_95 = {dataGroup_3_95, dataGroup_2_95};
  wire [127:0]  res_lo_lo_95 = {res_lo_lo_hi_95, res_lo_lo_lo_95};
  wire [63:0]   res_lo_hi_lo_95 = {dataGroup_5_95, dataGroup_4_95};
  wire [63:0]   res_lo_hi_hi_95 = {dataGroup_7_95, dataGroup_6_95};
  wire [127:0]  res_lo_hi_95 = {res_lo_hi_hi_95, res_lo_hi_lo_95};
  wire [255:0]  res_lo_95 = {res_lo_hi_95, res_lo_lo_95};
  wire [63:0]   res_hi_lo_lo_95 = {dataGroup_9_95, dataGroup_8_95};
  wire [63:0]   res_hi_lo_hi_95 = {dataGroup_11_95, dataGroup_10_95};
  wire [127:0]  res_hi_lo_95 = {res_hi_lo_hi_95, res_hi_lo_lo_95};
  wire [63:0]   res_hi_hi_lo_95 = {dataGroup_13_95, dataGroup_12_95};
  wire [63:0]   res_hi_hi_hi_95 = {dataGroup_15_95, dataGroup_14_95};
  wire [127:0]  res_hi_hi_95 = {res_hi_hi_hi_95, res_hi_hi_lo_95};
  wire [255:0]  res_hi_95 = {res_hi_hi_95, res_hi_lo_95};
  wire [511:0]  res_178 = {res_hi_95, res_lo_95};
  wire [2047:0] dataGroup_lo_3840 = {dataGroup_lo_hi_3840, dataGroup_lo_lo_3840};
  wire [2047:0] dataGroup_hi_3840 = {dataGroup_hi_hi_3840, dataGroup_hi_lo_3840};
  wire [31:0]   dataGroup_0_96 = dataGroup_lo_3840[127:96];
  wire [2047:0] dataGroup_lo_3841 = {dataGroup_lo_hi_3841, dataGroup_lo_lo_3841};
  wire [2047:0] dataGroup_hi_3841 = {dataGroup_hi_hi_3841, dataGroup_hi_lo_3841};
  wire [31:0]   dataGroup_1_96 = dataGroup_lo_3841[351:320];
  wire [2047:0] dataGroup_lo_3842 = {dataGroup_lo_hi_3842, dataGroup_lo_lo_3842};
  wire [2047:0] dataGroup_hi_3842 = {dataGroup_hi_hi_3842, dataGroup_hi_lo_3842};
  wire [31:0]   dataGroup_2_96 = dataGroup_lo_3842[575:544];
  wire [2047:0] dataGroup_lo_3843 = {dataGroup_lo_hi_3843, dataGroup_lo_lo_3843};
  wire [2047:0] dataGroup_hi_3843 = {dataGroup_hi_hi_3843, dataGroup_hi_lo_3843};
  wire [31:0]   dataGroup_3_96 = dataGroup_lo_3843[799:768];
  wire [2047:0] dataGroup_lo_3844 = {dataGroup_lo_hi_3844, dataGroup_lo_lo_3844};
  wire [2047:0] dataGroup_hi_3844 = {dataGroup_hi_hi_3844, dataGroup_hi_lo_3844};
  wire [31:0]   dataGroup_4_96 = dataGroup_lo_3844[1023:992];
  wire [2047:0] dataGroup_lo_3845 = {dataGroup_lo_hi_3845, dataGroup_lo_lo_3845};
  wire [2047:0] dataGroup_hi_3845 = {dataGroup_hi_hi_3845, dataGroup_hi_lo_3845};
  wire [31:0]   dataGroup_5_96 = dataGroup_lo_3845[1247:1216];
  wire [2047:0] dataGroup_lo_3846 = {dataGroup_lo_hi_3846, dataGroup_lo_lo_3846};
  wire [2047:0] dataGroup_hi_3846 = {dataGroup_hi_hi_3846, dataGroup_hi_lo_3846};
  wire [31:0]   dataGroup_6_96 = dataGroup_lo_3846[1471:1440];
  wire [2047:0] dataGroup_lo_3847 = {dataGroup_lo_hi_3847, dataGroup_lo_lo_3847};
  wire [2047:0] dataGroup_hi_3847 = {dataGroup_hi_hi_3847, dataGroup_hi_lo_3847};
  wire [31:0]   dataGroup_7_96 = dataGroup_lo_3847[1695:1664];
  wire [2047:0] dataGroup_lo_3848 = {dataGroup_lo_hi_3848, dataGroup_lo_lo_3848};
  wire [2047:0] dataGroup_hi_3848 = {dataGroup_hi_hi_3848, dataGroup_hi_lo_3848};
  wire [31:0]   dataGroup_8_96 = dataGroup_lo_3848[1919:1888];
  wire [2047:0] dataGroup_lo_3849 = {dataGroup_lo_hi_3849, dataGroup_lo_lo_3849};
  wire [2047:0] dataGroup_hi_3849 = {dataGroup_hi_hi_3849, dataGroup_hi_lo_3849};
  wire [31:0]   dataGroup_9_96 = dataGroup_hi_3849[95:64];
  wire [2047:0] dataGroup_lo_3850 = {dataGroup_lo_hi_3850, dataGroup_lo_lo_3850};
  wire [2047:0] dataGroup_hi_3850 = {dataGroup_hi_hi_3850, dataGroup_hi_lo_3850};
  wire [31:0]   dataGroup_10_96 = dataGroup_hi_3850[319:288];
  wire [2047:0] dataGroup_lo_3851 = {dataGroup_lo_hi_3851, dataGroup_lo_lo_3851};
  wire [2047:0] dataGroup_hi_3851 = {dataGroup_hi_hi_3851, dataGroup_hi_lo_3851};
  wire [31:0]   dataGroup_11_96 = dataGroup_hi_3851[543:512];
  wire [2047:0] dataGroup_lo_3852 = {dataGroup_lo_hi_3852, dataGroup_lo_lo_3852};
  wire [2047:0] dataGroup_hi_3852 = {dataGroup_hi_hi_3852, dataGroup_hi_lo_3852};
  wire [31:0]   dataGroup_12_96 = dataGroup_hi_3852[767:736];
  wire [2047:0] dataGroup_lo_3853 = {dataGroup_lo_hi_3853, dataGroup_lo_lo_3853};
  wire [2047:0] dataGroup_hi_3853 = {dataGroup_hi_hi_3853, dataGroup_hi_lo_3853};
  wire [31:0]   dataGroup_13_96 = dataGroup_hi_3853[991:960];
  wire [2047:0] dataGroup_lo_3854 = {dataGroup_lo_hi_3854, dataGroup_lo_lo_3854};
  wire [2047:0] dataGroup_hi_3854 = {dataGroup_hi_hi_3854, dataGroup_hi_lo_3854};
  wire [31:0]   dataGroup_14_96 = dataGroup_hi_3854[1215:1184];
  wire [2047:0] dataGroup_lo_3855 = {dataGroup_lo_hi_3855, dataGroup_lo_lo_3855};
  wire [2047:0] dataGroup_hi_3855 = {dataGroup_hi_hi_3855, dataGroup_hi_lo_3855};
  wire [31:0]   dataGroup_15_96 = dataGroup_hi_3855[1439:1408];
  wire [63:0]   res_lo_lo_lo_96 = {dataGroup_1_96, dataGroup_0_96};
  wire [63:0]   res_lo_lo_hi_96 = {dataGroup_3_96, dataGroup_2_96};
  wire [127:0]  res_lo_lo_96 = {res_lo_lo_hi_96, res_lo_lo_lo_96};
  wire [63:0]   res_lo_hi_lo_96 = {dataGroup_5_96, dataGroup_4_96};
  wire [63:0]   res_lo_hi_hi_96 = {dataGroup_7_96, dataGroup_6_96};
  wire [127:0]  res_lo_hi_96 = {res_lo_hi_hi_96, res_lo_hi_lo_96};
  wire [255:0]  res_lo_96 = {res_lo_hi_96, res_lo_lo_96};
  wire [63:0]   res_hi_lo_lo_96 = {dataGroup_9_96, dataGroup_8_96};
  wire [63:0]   res_hi_lo_hi_96 = {dataGroup_11_96, dataGroup_10_96};
  wire [127:0]  res_hi_lo_96 = {res_hi_lo_hi_96, res_hi_lo_lo_96};
  wire [63:0]   res_hi_hi_lo_96 = {dataGroup_13_96, dataGroup_12_96};
  wire [63:0]   res_hi_hi_hi_96 = {dataGroup_15_96, dataGroup_14_96};
  wire [127:0]  res_hi_hi_96 = {res_hi_hi_hi_96, res_hi_hi_lo_96};
  wire [255:0]  res_hi_96 = {res_hi_hi_96, res_hi_lo_96};
  wire [511:0]  res_179 = {res_hi_96, res_lo_96};
  wire [2047:0] dataGroup_lo_3856 = {dataGroup_lo_hi_3856, dataGroup_lo_lo_3856};
  wire [2047:0] dataGroup_hi_3856 = {dataGroup_hi_hi_3856, dataGroup_hi_lo_3856};
  wire [31:0]   dataGroup_0_97 = dataGroup_lo_3856[159:128];
  wire [2047:0] dataGroup_lo_3857 = {dataGroup_lo_hi_3857, dataGroup_lo_lo_3857};
  wire [2047:0] dataGroup_hi_3857 = {dataGroup_hi_hi_3857, dataGroup_hi_lo_3857};
  wire [31:0]   dataGroup_1_97 = dataGroup_lo_3857[383:352];
  wire [2047:0] dataGroup_lo_3858 = {dataGroup_lo_hi_3858, dataGroup_lo_lo_3858};
  wire [2047:0] dataGroup_hi_3858 = {dataGroup_hi_hi_3858, dataGroup_hi_lo_3858};
  wire [31:0]   dataGroup_2_97 = dataGroup_lo_3858[607:576];
  wire [2047:0] dataGroup_lo_3859 = {dataGroup_lo_hi_3859, dataGroup_lo_lo_3859};
  wire [2047:0] dataGroup_hi_3859 = {dataGroup_hi_hi_3859, dataGroup_hi_lo_3859};
  wire [31:0]   dataGroup_3_97 = dataGroup_lo_3859[831:800];
  wire [2047:0] dataGroup_lo_3860 = {dataGroup_lo_hi_3860, dataGroup_lo_lo_3860};
  wire [2047:0] dataGroup_hi_3860 = {dataGroup_hi_hi_3860, dataGroup_hi_lo_3860};
  wire [31:0]   dataGroup_4_97 = dataGroup_lo_3860[1055:1024];
  wire [2047:0] dataGroup_lo_3861 = {dataGroup_lo_hi_3861, dataGroup_lo_lo_3861};
  wire [2047:0] dataGroup_hi_3861 = {dataGroup_hi_hi_3861, dataGroup_hi_lo_3861};
  wire [31:0]   dataGroup_5_97 = dataGroup_lo_3861[1279:1248];
  wire [2047:0] dataGroup_lo_3862 = {dataGroup_lo_hi_3862, dataGroup_lo_lo_3862};
  wire [2047:0] dataGroup_hi_3862 = {dataGroup_hi_hi_3862, dataGroup_hi_lo_3862};
  wire [31:0]   dataGroup_6_97 = dataGroup_lo_3862[1503:1472];
  wire [2047:0] dataGroup_lo_3863 = {dataGroup_lo_hi_3863, dataGroup_lo_lo_3863};
  wire [2047:0] dataGroup_hi_3863 = {dataGroup_hi_hi_3863, dataGroup_hi_lo_3863};
  wire [31:0]   dataGroup_7_97 = dataGroup_lo_3863[1727:1696];
  wire [2047:0] dataGroup_lo_3864 = {dataGroup_lo_hi_3864, dataGroup_lo_lo_3864};
  wire [2047:0] dataGroup_hi_3864 = {dataGroup_hi_hi_3864, dataGroup_hi_lo_3864};
  wire [31:0]   dataGroup_8_97 = dataGroup_lo_3864[1951:1920];
  wire [2047:0] dataGroup_lo_3865 = {dataGroup_lo_hi_3865, dataGroup_lo_lo_3865};
  wire [2047:0] dataGroup_hi_3865 = {dataGroup_hi_hi_3865, dataGroup_hi_lo_3865};
  wire [31:0]   dataGroup_9_97 = dataGroup_hi_3865[127:96];
  wire [2047:0] dataGroup_lo_3866 = {dataGroup_lo_hi_3866, dataGroup_lo_lo_3866};
  wire [2047:0] dataGroup_hi_3866 = {dataGroup_hi_hi_3866, dataGroup_hi_lo_3866};
  wire [31:0]   dataGroup_10_97 = dataGroup_hi_3866[351:320];
  wire [2047:0] dataGroup_lo_3867 = {dataGroup_lo_hi_3867, dataGroup_lo_lo_3867};
  wire [2047:0] dataGroup_hi_3867 = {dataGroup_hi_hi_3867, dataGroup_hi_lo_3867};
  wire [31:0]   dataGroup_11_97 = dataGroup_hi_3867[575:544];
  wire [2047:0] dataGroup_lo_3868 = {dataGroup_lo_hi_3868, dataGroup_lo_lo_3868};
  wire [2047:0] dataGroup_hi_3868 = {dataGroup_hi_hi_3868, dataGroup_hi_lo_3868};
  wire [31:0]   dataGroup_12_97 = dataGroup_hi_3868[799:768];
  wire [2047:0] dataGroup_lo_3869 = {dataGroup_lo_hi_3869, dataGroup_lo_lo_3869};
  wire [2047:0] dataGroup_hi_3869 = {dataGroup_hi_hi_3869, dataGroup_hi_lo_3869};
  wire [31:0]   dataGroup_13_97 = dataGroup_hi_3869[1023:992];
  wire [2047:0] dataGroup_lo_3870 = {dataGroup_lo_hi_3870, dataGroup_lo_lo_3870};
  wire [2047:0] dataGroup_hi_3870 = {dataGroup_hi_hi_3870, dataGroup_hi_lo_3870};
  wire [31:0]   dataGroup_14_97 = dataGroup_hi_3870[1247:1216];
  wire [2047:0] dataGroup_lo_3871 = {dataGroup_lo_hi_3871, dataGroup_lo_lo_3871};
  wire [2047:0] dataGroup_hi_3871 = {dataGroup_hi_hi_3871, dataGroup_hi_lo_3871};
  wire [31:0]   dataGroup_15_97 = dataGroup_hi_3871[1471:1440];
  wire [63:0]   res_lo_lo_lo_97 = {dataGroup_1_97, dataGroup_0_97};
  wire [63:0]   res_lo_lo_hi_97 = {dataGroup_3_97, dataGroup_2_97};
  wire [127:0]  res_lo_lo_97 = {res_lo_lo_hi_97, res_lo_lo_lo_97};
  wire [63:0]   res_lo_hi_lo_97 = {dataGroup_5_97, dataGroup_4_97};
  wire [63:0]   res_lo_hi_hi_97 = {dataGroup_7_97, dataGroup_6_97};
  wire [127:0]  res_lo_hi_97 = {res_lo_hi_hi_97, res_lo_hi_lo_97};
  wire [255:0]  res_lo_97 = {res_lo_hi_97, res_lo_lo_97};
  wire [63:0]   res_hi_lo_lo_97 = {dataGroup_9_97, dataGroup_8_97};
  wire [63:0]   res_hi_lo_hi_97 = {dataGroup_11_97, dataGroup_10_97};
  wire [127:0]  res_hi_lo_97 = {res_hi_lo_hi_97, res_hi_lo_lo_97};
  wire [63:0]   res_hi_hi_lo_97 = {dataGroup_13_97, dataGroup_12_97};
  wire [63:0]   res_hi_hi_hi_97 = {dataGroup_15_97, dataGroup_14_97};
  wire [127:0]  res_hi_hi_97 = {res_hi_hi_hi_97, res_hi_hi_lo_97};
  wire [255:0]  res_hi_97 = {res_hi_hi_97, res_hi_lo_97};
  wire [511:0]  res_180 = {res_hi_97, res_lo_97};
  wire [2047:0] dataGroup_lo_3872 = {dataGroup_lo_hi_3872, dataGroup_lo_lo_3872};
  wire [2047:0] dataGroup_hi_3872 = {dataGroup_hi_hi_3872, dataGroup_hi_lo_3872};
  wire [31:0]   dataGroup_0_98 = dataGroup_lo_3872[191:160];
  wire [2047:0] dataGroup_lo_3873 = {dataGroup_lo_hi_3873, dataGroup_lo_lo_3873};
  wire [2047:0] dataGroup_hi_3873 = {dataGroup_hi_hi_3873, dataGroup_hi_lo_3873};
  wire [31:0]   dataGroup_1_98 = dataGroup_lo_3873[415:384];
  wire [2047:0] dataGroup_lo_3874 = {dataGroup_lo_hi_3874, dataGroup_lo_lo_3874};
  wire [2047:0] dataGroup_hi_3874 = {dataGroup_hi_hi_3874, dataGroup_hi_lo_3874};
  wire [31:0]   dataGroup_2_98 = dataGroup_lo_3874[639:608];
  wire [2047:0] dataGroup_lo_3875 = {dataGroup_lo_hi_3875, dataGroup_lo_lo_3875};
  wire [2047:0] dataGroup_hi_3875 = {dataGroup_hi_hi_3875, dataGroup_hi_lo_3875};
  wire [31:0]   dataGroup_3_98 = dataGroup_lo_3875[863:832];
  wire [2047:0] dataGroup_lo_3876 = {dataGroup_lo_hi_3876, dataGroup_lo_lo_3876};
  wire [2047:0] dataGroup_hi_3876 = {dataGroup_hi_hi_3876, dataGroup_hi_lo_3876};
  wire [31:0]   dataGroup_4_98 = dataGroup_lo_3876[1087:1056];
  wire [2047:0] dataGroup_lo_3877 = {dataGroup_lo_hi_3877, dataGroup_lo_lo_3877};
  wire [2047:0] dataGroup_hi_3877 = {dataGroup_hi_hi_3877, dataGroup_hi_lo_3877};
  wire [31:0]   dataGroup_5_98 = dataGroup_lo_3877[1311:1280];
  wire [2047:0] dataGroup_lo_3878 = {dataGroup_lo_hi_3878, dataGroup_lo_lo_3878};
  wire [2047:0] dataGroup_hi_3878 = {dataGroup_hi_hi_3878, dataGroup_hi_lo_3878};
  wire [31:0]   dataGroup_6_98 = dataGroup_lo_3878[1535:1504];
  wire [2047:0] dataGroup_lo_3879 = {dataGroup_lo_hi_3879, dataGroup_lo_lo_3879};
  wire [2047:0] dataGroup_hi_3879 = {dataGroup_hi_hi_3879, dataGroup_hi_lo_3879};
  wire [31:0]   dataGroup_7_98 = dataGroup_lo_3879[1759:1728];
  wire [2047:0] dataGroup_lo_3880 = {dataGroup_lo_hi_3880, dataGroup_lo_lo_3880};
  wire [2047:0] dataGroup_hi_3880 = {dataGroup_hi_hi_3880, dataGroup_hi_lo_3880};
  wire [31:0]   dataGroup_8_98 = dataGroup_lo_3880[1983:1952];
  wire [2047:0] dataGroup_lo_3881 = {dataGroup_lo_hi_3881, dataGroup_lo_lo_3881};
  wire [2047:0] dataGroup_hi_3881 = {dataGroup_hi_hi_3881, dataGroup_hi_lo_3881};
  wire [31:0]   dataGroup_9_98 = dataGroup_hi_3881[159:128];
  wire [2047:0] dataGroup_lo_3882 = {dataGroup_lo_hi_3882, dataGroup_lo_lo_3882};
  wire [2047:0] dataGroup_hi_3882 = {dataGroup_hi_hi_3882, dataGroup_hi_lo_3882};
  wire [31:0]   dataGroup_10_98 = dataGroup_hi_3882[383:352];
  wire [2047:0] dataGroup_lo_3883 = {dataGroup_lo_hi_3883, dataGroup_lo_lo_3883};
  wire [2047:0] dataGroup_hi_3883 = {dataGroup_hi_hi_3883, dataGroup_hi_lo_3883};
  wire [31:0]   dataGroup_11_98 = dataGroup_hi_3883[607:576];
  wire [2047:0] dataGroup_lo_3884 = {dataGroup_lo_hi_3884, dataGroup_lo_lo_3884};
  wire [2047:0] dataGroup_hi_3884 = {dataGroup_hi_hi_3884, dataGroup_hi_lo_3884};
  wire [31:0]   dataGroup_12_98 = dataGroup_hi_3884[831:800];
  wire [2047:0] dataGroup_lo_3885 = {dataGroup_lo_hi_3885, dataGroup_lo_lo_3885};
  wire [2047:0] dataGroup_hi_3885 = {dataGroup_hi_hi_3885, dataGroup_hi_lo_3885};
  wire [31:0]   dataGroup_13_98 = dataGroup_hi_3885[1055:1024];
  wire [2047:0] dataGroup_lo_3886 = {dataGroup_lo_hi_3886, dataGroup_lo_lo_3886};
  wire [2047:0] dataGroup_hi_3886 = {dataGroup_hi_hi_3886, dataGroup_hi_lo_3886};
  wire [31:0]   dataGroup_14_98 = dataGroup_hi_3886[1279:1248];
  wire [2047:0] dataGroup_lo_3887 = {dataGroup_lo_hi_3887, dataGroup_lo_lo_3887};
  wire [2047:0] dataGroup_hi_3887 = {dataGroup_hi_hi_3887, dataGroup_hi_lo_3887};
  wire [31:0]   dataGroup_15_98 = dataGroup_hi_3887[1503:1472];
  wire [63:0]   res_lo_lo_lo_98 = {dataGroup_1_98, dataGroup_0_98};
  wire [63:0]   res_lo_lo_hi_98 = {dataGroup_3_98, dataGroup_2_98};
  wire [127:0]  res_lo_lo_98 = {res_lo_lo_hi_98, res_lo_lo_lo_98};
  wire [63:0]   res_lo_hi_lo_98 = {dataGroup_5_98, dataGroup_4_98};
  wire [63:0]   res_lo_hi_hi_98 = {dataGroup_7_98, dataGroup_6_98};
  wire [127:0]  res_lo_hi_98 = {res_lo_hi_hi_98, res_lo_hi_lo_98};
  wire [255:0]  res_lo_98 = {res_lo_hi_98, res_lo_lo_98};
  wire [63:0]   res_hi_lo_lo_98 = {dataGroup_9_98, dataGroup_8_98};
  wire [63:0]   res_hi_lo_hi_98 = {dataGroup_11_98, dataGroup_10_98};
  wire [127:0]  res_hi_lo_98 = {res_hi_lo_hi_98, res_hi_lo_lo_98};
  wire [63:0]   res_hi_hi_lo_98 = {dataGroup_13_98, dataGroup_12_98};
  wire [63:0]   res_hi_hi_hi_98 = {dataGroup_15_98, dataGroup_14_98};
  wire [127:0]  res_hi_hi_98 = {res_hi_hi_hi_98, res_hi_hi_lo_98};
  wire [255:0]  res_hi_98 = {res_hi_hi_98, res_hi_lo_98};
  wire [511:0]  res_181 = {res_hi_98, res_lo_98};
  wire [2047:0] dataGroup_lo_3888 = {dataGroup_lo_hi_3888, dataGroup_lo_lo_3888};
  wire [2047:0] dataGroup_hi_3888 = {dataGroup_hi_hi_3888, dataGroup_hi_lo_3888};
  wire [31:0]   dataGroup_0_99 = dataGroup_lo_3888[223:192];
  wire [2047:0] dataGroup_lo_3889 = {dataGroup_lo_hi_3889, dataGroup_lo_lo_3889};
  wire [2047:0] dataGroup_hi_3889 = {dataGroup_hi_hi_3889, dataGroup_hi_lo_3889};
  wire [31:0]   dataGroup_1_99 = dataGroup_lo_3889[447:416];
  wire [2047:0] dataGroup_lo_3890 = {dataGroup_lo_hi_3890, dataGroup_lo_lo_3890};
  wire [2047:0] dataGroup_hi_3890 = {dataGroup_hi_hi_3890, dataGroup_hi_lo_3890};
  wire [31:0]   dataGroup_2_99 = dataGroup_lo_3890[671:640];
  wire [2047:0] dataGroup_lo_3891 = {dataGroup_lo_hi_3891, dataGroup_lo_lo_3891};
  wire [2047:0] dataGroup_hi_3891 = {dataGroup_hi_hi_3891, dataGroup_hi_lo_3891};
  wire [31:0]   dataGroup_3_99 = dataGroup_lo_3891[895:864];
  wire [2047:0] dataGroup_lo_3892 = {dataGroup_lo_hi_3892, dataGroup_lo_lo_3892};
  wire [2047:0] dataGroup_hi_3892 = {dataGroup_hi_hi_3892, dataGroup_hi_lo_3892};
  wire [31:0]   dataGroup_4_99 = dataGroup_lo_3892[1119:1088];
  wire [2047:0] dataGroup_lo_3893 = {dataGroup_lo_hi_3893, dataGroup_lo_lo_3893};
  wire [2047:0] dataGroup_hi_3893 = {dataGroup_hi_hi_3893, dataGroup_hi_lo_3893};
  wire [31:0]   dataGroup_5_99 = dataGroup_lo_3893[1343:1312];
  wire [2047:0] dataGroup_lo_3894 = {dataGroup_lo_hi_3894, dataGroup_lo_lo_3894};
  wire [2047:0] dataGroup_hi_3894 = {dataGroup_hi_hi_3894, dataGroup_hi_lo_3894};
  wire [31:0]   dataGroup_6_99 = dataGroup_lo_3894[1567:1536];
  wire [2047:0] dataGroup_lo_3895 = {dataGroup_lo_hi_3895, dataGroup_lo_lo_3895};
  wire [2047:0] dataGroup_hi_3895 = {dataGroup_hi_hi_3895, dataGroup_hi_lo_3895};
  wire [31:0]   dataGroup_7_99 = dataGroup_lo_3895[1791:1760];
  wire [2047:0] dataGroup_lo_3896 = {dataGroup_lo_hi_3896, dataGroup_lo_lo_3896};
  wire [2047:0] dataGroup_hi_3896 = {dataGroup_hi_hi_3896, dataGroup_hi_lo_3896};
  wire [31:0]   dataGroup_8_99 = dataGroup_lo_3896[2015:1984];
  wire [2047:0] dataGroup_lo_3897 = {dataGroup_lo_hi_3897, dataGroup_lo_lo_3897};
  wire [2047:0] dataGroup_hi_3897 = {dataGroup_hi_hi_3897, dataGroup_hi_lo_3897};
  wire [31:0]   dataGroup_9_99 = dataGroup_hi_3897[191:160];
  wire [2047:0] dataGroup_lo_3898 = {dataGroup_lo_hi_3898, dataGroup_lo_lo_3898};
  wire [2047:0] dataGroup_hi_3898 = {dataGroup_hi_hi_3898, dataGroup_hi_lo_3898};
  wire [31:0]   dataGroup_10_99 = dataGroup_hi_3898[415:384];
  wire [2047:0] dataGroup_lo_3899 = {dataGroup_lo_hi_3899, dataGroup_lo_lo_3899};
  wire [2047:0] dataGroup_hi_3899 = {dataGroup_hi_hi_3899, dataGroup_hi_lo_3899};
  wire [31:0]   dataGroup_11_99 = dataGroup_hi_3899[639:608];
  wire [2047:0] dataGroup_lo_3900 = {dataGroup_lo_hi_3900, dataGroup_lo_lo_3900};
  wire [2047:0] dataGroup_hi_3900 = {dataGroup_hi_hi_3900, dataGroup_hi_lo_3900};
  wire [31:0]   dataGroup_12_99 = dataGroup_hi_3900[863:832];
  wire [2047:0] dataGroup_lo_3901 = {dataGroup_lo_hi_3901, dataGroup_lo_lo_3901};
  wire [2047:0] dataGroup_hi_3901 = {dataGroup_hi_hi_3901, dataGroup_hi_lo_3901};
  wire [31:0]   dataGroup_13_99 = dataGroup_hi_3901[1087:1056];
  wire [2047:0] dataGroup_lo_3902 = {dataGroup_lo_hi_3902, dataGroup_lo_lo_3902};
  wire [2047:0] dataGroup_hi_3902 = {dataGroup_hi_hi_3902, dataGroup_hi_lo_3902};
  wire [31:0]   dataGroup_14_99 = dataGroup_hi_3902[1311:1280];
  wire [2047:0] dataGroup_lo_3903 = {dataGroup_lo_hi_3903, dataGroup_lo_lo_3903};
  wire [2047:0] dataGroup_hi_3903 = {dataGroup_hi_hi_3903, dataGroup_hi_lo_3903};
  wire [31:0]   dataGroup_15_99 = dataGroup_hi_3903[1535:1504];
  wire [63:0]   res_lo_lo_lo_99 = {dataGroup_1_99, dataGroup_0_99};
  wire [63:0]   res_lo_lo_hi_99 = {dataGroup_3_99, dataGroup_2_99};
  wire [127:0]  res_lo_lo_99 = {res_lo_lo_hi_99, res_lo_lo_lo_99};
  wire [63:0]   res_lo_hi_lo_99 = {dataGroup_5_99, dataGroup_4_99};
  wire [63:0]   res_lo_hi_hi_99 = {dataGroup_7_99, dataGroup_6_99};
  wire [127:0]  res_lo_hi_99 = {res_lo_hi_hi_99, res_lo_hi_lo_99};
  wire [255:0]  res_lo_99 = {res_lo_hi_99, res_lo_lo_99};
  wire [63:0]   res_hi_lo_lo_99 = {dataGroup_9_99, dataGroup_8_99};
  wire [63:0]   res_hi_lo_hi_99 = {dataGroup_11_99, dataGroup_10_99};
  wire [127:0]  res_hi_lo_99 = {res_hi_lo_hi_99, res_hi_lo_lo_99};
  wire [63:0]   res_hi_hi_lo_99 = {dataGroup_13_99, dataGroup_12_99};
  wire [63:0]   res_hi_hi_hi_99 = {dataGroup_15_99, dataGroup_14_99};
  wire [127:0]  res_hi_hi_99 = {res_hi_hi_hi_99, res_hi_hi_lo_99};
  wire [255:0]  res_hi_99 = {res_hi_hi_99, res_hi_lo_99};
  wire [511:0]  res_182 = {res_hi_99, res_lo_99};
  wire [1023:0] lo_lo_22 = {res_177, res_176};
  wire [1023:0] lo_hi_22 = {res_179, res_178};
  wire [2047:0] lo_22 = {lo_hi_22, lo_lo_22};
  wire [1023:0] hi_lo_22 = {res_181, res_180};
  wire [1023:0] hi_hi_22 = {512'h0, res_182};
  wire [2047:0] hi_22 = {hi_hi_22, hi_lo_22};
  wire [4095:0] regroupLoadData_2_6 = {hi_22, lo_22};
  wire [2047:0] dataGroup_lo_3904 = {dataGroup_lo_hi_3904, dataGroup_lo_lo_3904};
  wire [2047:0] dataGroup_hi_3904 = {dataGroup_hi_hi_3904, dataGroup_hi_lo_3904};
  wire [31:0]   dataGroup_0_100 = dataGroup_lo_3904[31:0];
  wire [2047:0] dataGroup_lo_3905 = {dataGroup_lo_hi_3905, dataGroup_lo_lo_3905};
  wire [2047:0] dataGroup_hi_3905 = {dataGroup_hi_hi_3905, dataGroup_hi_lo_3905};
  wire [31:0]   dataGroup_1_100 = dataGroup_lo_3905[287:256];
  wire [2047:0] dataGroup_lo_3906 = {dataGroup_lo_hi_3906, dataGroup_lo_lo_3906};
  wire [2047:0] dataGroup_hi_3906 = {dataGroup_hi_hi_3906, dataGroup_hi_lo_3906};
  wire [31:0]   dataGroup_2_100 = dataGroup_lo_3906[543:512];
  wire [2047:0] dataGroup_lo_3907 = {dataGroup_lo_hi_3907, dataGroup_lo_lo_3907};
  wire [2047:0] dataGroup_hi_3907 = {dataGroup_hi_hi_3907, dataGroup_hi_lo_3907};
  wire [31:0]   dataGroup_3_100 = dataGroup_lo_3907[799:768];
  wire [2047:0] dataGroup_lo_3908 = {dataGroup_lo_hi_3908, dataGroup_lo_lo_3908};
  wire [2047:0] dataGroup_hi_3908 = {dataGroup_hi_hi_3908, dataGroup_hi_lo_3908};
  wire [31:0]   dataGroup_4_100 = dataGroup_lo_3908[1055:1024];
  wire [2047:0] dataGroup_lo_3909 = {dataGroup_lo_hi_3909, dataGroup_lo_lo_3909};
  wire [2047:0] dataGroup_hi_3909 = {dataGroup_hi_hi_3909, dataGroup_hi_lo_3909};
  wire [31:0]   dataGroup_5_100 = dataGroup_lo_3909[1311:1280];
  wire [2047:0] dataGroup_lo_3910 = {dataGroup_lo_hi_3910, dataGroup_lo_lo_3910};
  wire [2047:0] dataGroup_hi_3910 = {dataGroup_hi_hi_3910, dataGroup_hi_lo_3910};
  wire [31:0]   dataGroup_6_100 = dataGroup_lo_3910[1567:1536];
  wire [2047:0] dataGroup_lo_3911 = {dataGroup_lo_hi_3911, dataGroup_lo_lo_3911};
  wire [2047:0] dataGroup_hi_3911 = {dataGroup_hi_hi_3911, dataGroup_hi_lo_3911};
  wire [31:0]   dataGroup_7_100 = dataGroup_lo_3911[1823:1792];
  wire [2047:0] dataGroup_lo_3912 = {dataGroup_lo_hi_3912, dataGroup_lo_lo_3912};
  wire [2047:0] dataGroup_hi_3912 = {dataGroup_hi_hi_3912, dataGroup_hi_lo_3912};
  wire [31:0]   dataGroup_8_100 = dataGroup_hi_3912[31:0];
  wire [2047:0] dataGroup_lo_3913 = {dataGroup_lo_hi_3913, dataGroup_lo_lo_3913};
  wire [2047:0] dataGroup_hi_3913 = {dataGroup_hi_hi_3913, dataGroup_hi_lo_3913};
  wire [31:0]   dataGroup_9_100 = dataGroup_hi_3913[287:256];
  wire [2047:0] dataGroup_lo_3914 = {dataGroup_lo_hi_3914, dataGroup_lo_lo_3914};
  wire [2047:0] dataGroup_hi_3914 = {dataGroup_hi_hi_3914, dataGroup_hi_lo_3914};
  wire [31:0]   dataGroup_10_100 = dataGroup_hi_3914[543:512];
  wire [2047:0] dataGroup_lo_3915 = {dataGroup_lo_hi_3915, dataGroup_lo_lo_3915};
  wire [2047:0] dataGroup_hi_3915 = {dataGroup_hi_hi_3915, dataGroup_hi_lo_3915};
  wire [31:0]   dataGroup_11_100 = dataGroup_hi_3915[799:768];
  wire [2047:0] dataGroup_lo_3916 = {dataGroup_lo_hi_3916, dataGroup_lo_lo_3916};
  wire [2047:0] dataGroup_hi_3916 = {dataGroup_hi_hi_3916, dataGroup_hi_lo_3916};
  wire [31:0]   dataGroup_12_100 = dataGroup_hi_3916[1055:1024];
  wire [2047:0] dataGroup_lo_3917 = {dataGroup_lo_hi_3917, dataGroup_lo_lo_3917};
  wire [2047:0] dataGroup_hi_3917 = {dataGroup_hi_hi_3917, dataGroup_hi_lo_3917};
  wire [31:0]   dataGroup_13_100 = dataGroup_hi_3917[1311:1280];
  wire [2047:0] dataGroup_lo_3918 = {dataGroup_lo_hi_3918, dataGroup_lo_lo_3918};
  wire [2047:0] dataGroup_hi_3918 = {dataGroup_hi_hi_3918, dataGroup_hi_lo_3918};
  wire [31:0]   dataGroup_14_100 = dataGroup_hi_3918[1567:1536];
  wire [2047:0] dataGroup_lo_3919 = {dataGroup_lo_hi_3919, dataGroup_lo_lo_3919};
  wire [2047:0] dataGroup_hi_3919 = {dataGroup_hi_hi_3919, dataGroup_hi_lo_3919};
  wire [31:0]   dataGroup_15_100 = dataGroup_hi_3919[1823:1792];
  wire [63:0]   res_lo_lo_lo_100 = {dataGroup_1_100, dataGroup_0_100};
  wire [63:0]   res_lo_lo_hi_100 = {dataGroup_3_100, dataGroup_2_100};
  wire [127:0]  res_lo_lo_100 = {res_lo_lo_hi_100, res_lo_lo_lo_100};
  wire [63:0]   res_lo_hi_lo_100 = {dataGroup_5_100, dataGroup_4_100};
  wire [63:0]   res_lo_hi_hi_100 = {dataGroup_7_100, dataGroup_6_100};
  wire [127:0]  res_lo_hi_100 = {res_lo_hi_hi_100, res_lo_hi_lo_100};
  wire [255:0]  res_lo_100 = {res_lo_hi_100, res_lo_lo_100};
  wire [63:0]   res_hi_lo_lo_100 = {dataGroup_9_100, dataGroup_8_100};
  wire [63:0]   res_hi_lo_hi_100 = {dataGroup_11_100, dataGroup_10_100};
  wire [127:0]  res_hi_lo_100 = {res_hi_lo_hi_100, res_hi_lo_lo_100};
  wire [63:0]   res_hi_hi_lo_100 = {dataGroup_13_100, dataGroup_12_100};
  wire [63:0]   res_hi_hi_hi_100 = {dataGroup_15_100, dataGroup_14_100};
  wire [127:0]  res_hi_hi_100 = {res_hi_hi_hi_100, res_hi_hi_lo_100};
  wire [255:0]  res_hi_100 = {res_hi_hi_100, res_hi_lo_100};
  wire [511:0]  res_184 = {res_hi_100, res_lo_100};
  wire [2047:0] dataGroup_lo_3920 = {dataGroup_lo_hi_3920, dataGroup_lo_lo_3920};
  wire [2047:0] dataGroup_hi_3920 = {dataGroup_hi_hi_3920, dataGroup_hi_lo_3920};
  wire [31:0]   dataGroup_0_101 = dataGroup_lo_3920[63:32];
  wire [2047:0] dataGroup_lo_3921 = {dataGroup_lo_hi_3921, dataGroup_lo_lo_3921};
  wire [2047:0] dataGroup_hi_3921 = {dataGroup_hi_hi_3921, dataGroup_hi_lo_3921};
  wire [31:0]   dataGroup_1_101 = dataGroup_lo_3921[319:288];
  wire [2047:0] dataGroup_lo_3922 = {dataGroup_lo_hi_3922, dataGroup_lo_lo_3922};
  wire [2047:0] dataGroup_hi_3922 = {dataGroup_hi_hi_3922, dataGroup_hi_lo_3922};
  wire [31:0]   dataGroup_2_101 = dataGroup_lo_3922[575:544];
  wire [2047:0] dataGroup_lo_3923 = {dataGroup_lo_hi_3923, dataGroup_lo_lo_3923};
  wire [2047:0] dataGroup_hi_3923 = {dataGroup_hi_hi_3923, dataGroup_hi_lo_3923};
  wire [31:0]   dataGroup_3_101 = dataGroup_lo_3923[831:800];
  wire [2047:0] dataGroup_lo_3924 = {dataGroup_lo_hi_3924, dataGroup_lo_lo_3924};
  wire [2047:0] dataGroup_hi_3924 = {dataGroup_hi_hi_3924, dataGroup_hi_lo_3924};
  wire [31:0]   dataGroup_4_101 = dataGroup_lo_3924[1087:1056];
  wire [2047:0] dataGroup_lo_3925 = {dataGroup_lo_hi_3925, dataGroup_lo_lo_3925};
  wire [2047:0] dataGroup_hi_3925 = {dataGroup_hi_hi_3925, dataGroup_hi_lo_3925};
  wire [31:0]   dataGroup_5_101 = dataGroup_lo_3925[1343:1312];
  wire [2047:0] dataGroup_lo_3926 = {dataGroup_lo_hi_3926, dataGroup_lo_lo_3926};
  wire [2047:0] dataGroup_hi_3926 = {dataGroup_hi_hi_3926, dataGroup_hi_lo_3926};
  wire [31:0]   dataGroup_6_101 = dataGroup_lo_3926[1599:1568];
  wire [2047:0] dataGroup_lo_3927 = {dataGroup_lo_hi_3927, dataGroup_lo_lo_3927};
  wire [2047:0] dataGroup_hi_3927 = {dataGroup_hi_hi_3927, dataGroup_hi_lo_3927};
  wire [31:0]   dataGroup_7_101 = dataGroup_lo_3927[1855:1824];
  wire [2047:0] dataGroup_lo_3928 = {dataGroup_lo_hi_3928, dataGroup_lo_lo_3928};
  wire [2047:0] dataGroup_hi_3928 = {dataGroup_hi_hi_3928, dataGroup_hi_lo_3928};
  wire [31:0]   dataGroup_8_101 = dataGroup_hi_3928[63:32];
  wire [2047:0] dataGroup_lo_3929 = {dataGroup_lo_hi_3929, dataGroup_lo_lo_3929};
  wire [2047:0] dataGroup_hi_3929 = {dataGroup_hi_hi_3929, dataGroup_hi_lo_3929};
  wire [31:0]   dataGroup_9_101 = dataGroup_hi_3929[319:288];
  wire [2047:0] dataGroup_lo_3930 = {dataGroup_lo_hi_3930, dataGroup_lo_lo_3930};
  wire [2047:0] dataGroup_hi_3930 = {dataGroup_hi_hi_3930, dataGroup_hi_lo_3930};
  wire [31:0]   dataGroup_10_101 = dataGroup_hi_3930[575:544];
  wire [2047:0] dataGroup_lo_3931 = {dataGroup_lo_hi_3931, dataGroup_lo_lo_3931};
  wire [2047:0] dataGroup_hi_3931 = {dataGroup_hi_hi_3931, dataGroup_hi_lo_3931};
  wire [31:0]   dataGroup_11_101 = dataGroup_hi_3931[831:800];
  wire [2047:0] dataGroup_lo_3932 = {dataGroup_lo_hi_3932, dataGroup_lo_lo_3932};
  wire [2047:0] dataGroup_hi_3932 = {dataGroup_hi_hi_3932, dataGroup_hi_lo_3932};
  wire [31:0]   dataGroup_12_101 = dataGroup_hi_3932[1087:1056];
  wire [2047:0] dataGroup_lo_3933 = {dataGroup_lo_hi_3933, dataGroup_lo_lo_3933};
  wire [2047:0] dataGroup_hi_3933 = {dataGroup_hi_hi_3933, dataGroup_hi_lo_3933};
  wire [31:0]   dataGroup_13_101 = dataGroup_hi_3933[1343:1312];
  wire [2047:0] dataGroup_lo_3934 = {dataGroup_lo_hi_3934, dataGroup_lo_lo_3934};
  wire [2047:0] dataGroup_hi_3934 = {dataGroup_hi_hi_3934, dataGroup_hi_lo_3934};
  wire [31:0]   dataGroup_14_101 = dataGroup_hi_3934[1599:1568];
  wire [2047:0] dataGroup_lo_3935 = {dataGroup_lo_hi_3935, dataGroup_lo_lo_3935};
  wire [2047:0] dataGroup_hi_3935 = {dataGroup_hi_hi_3935, dataGroup_hi_lo_3935};
  wire [31:0]   dataGroup_15_101 = dataGroup_hi_3935[1855:1824];
  wire [63:0]   res_lo_lo_lo_101 = {dataGroup_1_101, dataGroup_0_101};
  wire [63:0]   res_lo_lo_hi_101 = {dataGroup_3_101, dataGroup_2_101};
  wire [127:0]  res_lo_lo_101 = {res_lo_lo_hi_101, res_lo_lo_lo_101};
  wire [63:0]   res_lo_hi_lo_101 = {dataGroup_5_101, dataGroup_4_101};
  wire [63:0]   res_lo_hi_hi_101 = {dataGroup_7_101, dataGroup_6_101};
  wire [127:0]  res_lo_hi_101 = {res_lo_hi_hi_101, res_lo_hi_lo_101};
  wire [255:0]  res_lo_101 = {res_lo_hi_101, res_lo_lo_101};
  wire [63:0]   res_hi_lo_lo_101 = {dataGroup_9_101, dataGroup_8_101};
  wire [63:0]   res_hi_lo_hi_101 = {dataGroup_11_101, dataGroup_10_101};
  wire [127:0]  res_hi_lo_101 = {res_hi_lo_hi_101, res_hi_lo_lo_101};
  wire [63:0]   res_hi_hi_lo_101 = {dataGroup_13_101, dataGroup_12_101};
  wire [63:0]   res_hi_hi_hi_101 = {dataGroup_15_101, dataGroup_14_101};
  wire [127:0]  res_hi_hi_101 = {res_hi_hi_hi_101, res_hi_hi_lo_101};
  wire [255:0]  res_hi_101 = {res_hi_hi_101, res_hi_lo_101};
  wire [511:0]  res_185 = {res_hi_101, res_lo_101};
  wire [2047:0] dataGroup_lo_3936 = {dataGroup_lo_hi_3936, dataGroup_lo_lo_3936};
  wire [2047:0] dataGroup_hi_3936 = {dataGroup_hi_hi_3936, dataGroup_hi_lo_3936};
  wire [31:0]   dataGroup_0_102 = dataGroup_lo_3936[95:64];
  wire [2047:0] dataGroup_lo_3937 = {dataGroup_lo_hi_3937, dataGroup_lo_lo_3937};
  wire [2047:0] dataGroup_hi_3937 = {dataGroup_hi_hi_3937, dataGroup_hi_lo_3937};
  wire [31:0]   dataGroup_1_102 = dataGroup_lo_3937[351:320];
  wire [2047:0] dataGroup_lo_3938 = {dataGroup_lo_hi_3938, dataGroup_lo_lo_3938};
  wire [2047:0] dataGroup_hi_3938 = {dataGroup_hi_hi_3938, dataGroup_hi_lo_3938};
  wire [31:0]   dataGroup_2_102 = dataGroup_lo_3938[607:576];
  wire [2047:0] dataGroup_lo_3939 = {dataGroup_lo_hi_3939, dataGroup_lo_lo_3939};
  wire [2047:0] dataGroup_hi_3939 = {dataGroup_hi_hi_3939, dataGroup_hi_lo_3939};
  wire [31:0]   dataGroup_3_102 = dataGroup_lo_3939[863:832];
  wire [2047:0] dataGroup_lo_3940 = {dataGroup_lo_hi_3940, dataGroup_lo_lo_3940};
  wire [2047:0] dataGroup_hi_3940 = {dataGroup_hi_hi_3940, dataGroup_hi_lo_3940};
  wire [31:0]   dataGroup_4_102 = dataGroup_lo_3940[1119:1088];
  wire [2047:0] dataGroup_lo_3941 = {dataGroup_lo_hi_3941, dataGroup_lo_lo_3941};
  wire [2047:0] dataGroup_hi_3941 = {dataGroup_hi_hi_3941, dataGroup_hi_lo_3941};
  wire [31:0]   dataGroup_5_102 = dataGroup_lo_3941[1375:1344];
  wire [2047:0] dataGroup_lo_3942 = {dataGroup_lo_hi_3942, dataGroup_lo_lo_3942};
  wire [2047:0] dataGroup_hi_3942 = {dataGroup_hi_hi_3942, dataGroup_hi_lo_3942};
  wire [31:0]   dataGroup_6_102 = dataGroup_lo_3942[1631:1600];
  wire [2047:0] dataGroup_lo_3943 = {dataGroup_lo_hi_3943, dataGroup_lo_lo_3943};
  wire [2047:0] dataGroup_hi_3943 = {dataGroup_hi_hi_3943, dataGroup_hi_lo_3943};
  wire [31:0]   dataGroup_7_102 = dataGroup_lo_3943[1887:1856];
  wire [2047:0] dataGroup_lo_3944 = {dataGroup_lo_hi_3944, dataGroup_lo_lo_3944};
  wire [2047:0] dataGroup_hi_3944 = {dataGroup_hi_hi_3944, dataGroup_hi_lo_3944};
  wire [31:0]   dataGroup_8_102 = dataGroup_hi_3944[95:64];
  wire [2047:0] dataGroup_lo_3945 = {dataGroup_lo_hi_3945, dataGroup_lo_lo_3945};
  wire [2047:0] dataGroup_hi_3945 = {dataGroup_hi_hi_3945, dataGroup_hi_lo_3945};
  wire [31:0]   dataGroup_9_102 = dataGroup_hi_3945[351:320];
  wire [2047:0] dataGroup_lo_3946 = {dataGroup_lo_hi_3946, dataGroup_lo_lo_3946};
  wire [2047:0] dataGroup_hi_3946 = {dataGroup_hi_hi_3946, dataGroup_hi_lo_3946};
  wire [31:0]   dataGroup_10_102 = dataGroup_hi_3946[607:576];
  wire [2047:0] dataGroup_lo_3947 = {dataGroup_lo_hi_3947, dataGroup_lo_lo_3947};
  wire [2047:0] dataGroup_hi_3947 = {dataGroup_hi_hi_3947, dataGroup_hi_lo_3947};
  wire [31:0]   dataGroup_11_102 = dataGroup_hi_3947[863:832];
  wire [2047:0] dataGroup_lo_3948 = {dataGroup_lo_hi_3948, dataGroup_lo_lo_3948};
  wire [2047:0] dataGroup_hi_3948 = {dataGroup_hi_hi_3948, dataGroup_hi_lo_3948};
  wire [31:0]   dataGroup_12_102 = dataGroup_hi_3948[1119:1088];
  wire [2047:0] dataGroup_lo_3949 = {dataGroup_lo_hi_3949, dataGroup_lo_lo_3949};
  wire [2047:0] dataGroup_hi_3949 = {dataGroup_hi_hi_3949, dataGroup_hi_lo_3949};
  wire [31:0]   dataGroup_13_102 = dataGroup_hi_3949[1375:1344];
  wire [2047:0] dataGroup_lo_3950 = {dataGroup_lo_hi_3950, dataGroup_lo_lo_3950};
  wire [2047:0] dataGroup_hi_3950 = {dataGroup_hi_hi_3950, dataGroup_hi_lo_3950};
  wire [31:0]   dataGroup_14_102 = dataGroup_hi_3950[1631:1600];
  wire [2047:0] dataGroup_lo_3951 = {dataGroup_lo_hi_3951, dataGroup_lo_lo_3951};
  wire [2047:0] dataGroup_hi_3951 = {dataGroup_hi_hi_3951, dataGroup_hi_lo_3951};
  wire [31:0]   dataGroup_15_102 = dataGroup_hi_3951[1887:1856];
  wire [63:0]   res_lo_lo_lo_102 = {dataGroup_1_102, dataGroup_0_102};
  wire [63:0]   res_lo_lo_hi_102 = {dataGroup_3_102, dataGroup_2_102};
  wire [127:0]  res_lo_lo_102 = {res_lo_lo_hi_102, res_lo_lo_lo_102};
  wire [63:0]   res_lo_hi_lo_102 = {dataGroup_5_102, dataGroup_4_102};
  wire [63:0]   res_lo_hi_hi_102 = {dataGroup_7_102, dataGroup_6_102};
  wire [127:0]  res_lo_hi_102 = {res_lo_hi_hi_102, res_lo_hi_lo_102};
  wire [255:0]  res_lo_102 = {res_lo_hi_102, res_lo_lo_102};
  wire [63:0]   res_hi_lo_lo_102 = {dataGroup_9_102, dataGroup_8_102};
  wire [63:0]   res_hi_lo_hi_102 = {dataGroup_11_102, dataGroup_10_102};
  wire [127:0]  res_hi_lo_102 = {res_hi_lo_hi_102, res_hi_lo_lo_102};
  wire [63:0]   res_hi_hi_lo_102 = {dataGroup_13_102, dataGroup_12_102};
  wire [63:0]   res_hi_hi_hi_102 = {dataGroup_15_102, dataGroup_14_102};
  wire [127:0]  res_hi_hi_102 = {res_hi_hi_hi_102, res_hi_hi_lo_102};
  wire [255:0]  res_hi_102 = {res_hi_hi_102, res_hi_lo_102};
  wire [511:0]  res_186 = {res_hi_102, res_lo_102};
  wire [2047:0] dataGroup_lo_3952 = {dataGroup_lo_hi_3952, dataGroup_lo_lo_3952};
  wire [2047:0] dataGroup_hi_3952 = {dataGroup_hi_hi_3952, dataGroup_hi_lo_3952};
  wire [31:0]   dataGroup_0_103 = dataGroup_lo_3952[127:96];
  wire [2047:0] dataGroup_lo_3953 = {dataGroup_lo_hi_3953, dataGroup_lo_lo_3953};
  wire [2047:0] dataGroup_hi_3953 = {dataGroup_hi_hi_3953, dataGroup_hi_lo_3953};
  wire [31:0]   dataGroup_1_103 = dataGroup_lo_3953[383:352];
  wire [2047:0] dataGroup_lo_3954 = {dataGroup_lo_hi_3954, dataGroup_lo_lo_3954};
  wire [2047:0] dataGroup_hi_3954 = {dataGroup_hi_hi_3954, dataGroup_hi_lo_3954};
  wire [31:0]   dataGroup_2_103 = dataGroup_lo_3954[639:608];
  wire [2047:0] dataGroup_lo_3955 = {dataGroup_lo_hi_3955, dataGroup_lo_lo_3955};
  wire [2047:0] dataGroup_hi_3955 = {dataGroup_hi_hi_3955, dataGroup_hi_lo_3955};
  wire [31:0]   dataGroup_3_103 = dataGroup_lo_3955[895:864];
  wire [2047:0] dataGroup_lo_3956 = {dataGroup_lo_hi_3956, dataGroup_lo_lo_3956};
  wire [2047:0] dataGroup_hi_3956 = {dataGroup_hi_hi_3956, dataGroup_hi_lo_3956};
  wire [31:0]   dataGroup_4_103 = dataGroup_lo_3956[1151:1120];
  wire [2047:0] dataGroup_lo_3957 = {dataGroup_lo_hi_3957, dataGroup_lo_lo_3957};
  wire [2047:0] dataGroup_hi_3957 = {dataGroup_hi_hi_3957, dataGroup_hi_lo_3957};
  wire [31:0]   dataGroup_5_103 = dataGroup_lo_3957[1407:1376];
  wire [2047:0] dataGroup_lo_3958 = {dataGroup_lo_hi_3958, dataGroup_lo_lo_3958};
  wire [2047:0] dataGroup_hi_3958 = {dataGroup_hi_hi_3958, dataGroup_hi_lo_3958};
  wire [31:0]   dataGroup_6_103 = dataGroup_lo_3958[1663:1632];
  wire [2047:0] dataGroup_lo_3959 = {dataGroup_lo_hi_3959, dataGroup_lo_lo_3959};
  wire [2047:0] dataGroup_hi_3959 = {dataGroup_hi_hi_3959, dataGroup_hi_lo_3959};
  wire [31:0]   dataGroup_7_103 = dataGroup_lo_3959[1919:1888];
  wire [2047:0] dataGroup_lo_3960 = {dataGroup_lo_hi_3960, dataGroup_lo_lo_3960};
  wire [2047:0] dataGroup_hi_3960 = {dataGroup_hi_hi_3960, dataGroup_hi_lo_3960};
  wire [31:0]   dataGroup_8_103 = dataGroup_hi_3960[127:96];
  wire [2047:0] dataGroup_lo_3961 = {dataGroup_lo_hi_3961, dataGroup_lo_lo_3961};
  wire [2047:0] dataGroup_hi_3961 = {dataGroup_hi_hi_3961, dataGroup_hi_lo_3961};
  wire [31:0]   dataGroup_9_103 = dataGroup_hi_3961[383:352];
  wire [2047:0] dataGroup_lo_3962 = {dataGroup_lo_hi_3962, dataGroup_lo_lo_3962};
  wire [2047:0] dataGroup_hi_3962 = {dataGroup_hi_hi_3962, dataGroup_hi_lo_3962};
  wire [31:0]   dataGroup_10_103 = dataGroup_hi_3962[639:608];
  wire [2047:0] dataGroup_lo_3963 = {dataGroup_lo_hi_3963, dataGroup_lo_lo_3963};
  wire [2047:0] dataGroup_hi_3963 = {dataGroup_hi_hi_3963, dataGroup_hi_lo_3963};
  wire [31:0]   dataGroup_11_103 = dataGroup_hi_3963[895:864];
  wire [2047:0] dataGroup_lo_3964 = {dataGroup_lo_hi_3964, dataGroup_lo_lo_3964};
  wire [2047:0] dataGroup_hi_3964 = {dataGroup_hi_hi_3964, dataGroup_hi_lo_3964};
  wire [31:0]   dataGroup_12_103 = dataGroup_hi_3964[1151:1120];
  wire [2047:0] dataGroup_lo_3965 = {dataGroup_lo_hi_3965, dataGroup_lo_lo_3965};
  wire [2047:0] dataGroup_hi_3965 = {dataGroup_hi_hi_3965, dataGroup_hi_lo_3965};
  wire [31:0]   dataGroup_13_103 = dataGroup_hi_3965[1407:1376];
  wire [2047:0] dataGroup_lo_3966 = {dataGroup_lo_hi_3966, dataGroup_lo_lo_3966};
  wire [2047:0] dataGroup_hi_3966 = {dataGroup_hi_hi_3966, dataGroup_hi_lo_3966};
  wire [31:0]   dataGroup_14_103 = dataGroup_hi_3966[1663:1632];
  wire [2047:0] dataGroup_lo_3967 = {dataGroup_lo_hi_3967, dataGroup_lo_lo_3967};
  wire [2047:0] dataGroup_hi_3967 = {dataGroup_hi_hi_3967, dataGroup_hi_lo_3967};
  wire [31:0]   dataGroup_15_103 = dataGroup_hi_3967[1919:1888];
  wire [63:0]   res_lo_lo_lo_103 = {dataGroup_1_103, dataGroup_0_103};
  wire [63:0]   res_lo_lo_hi_103 = {dataGroup_3_103, dataGroup_2_103};
  wire [127:0]  res_lo_lo_103 = {res_lo_lo_hi_103, res_lo_lo_lo_103};
  wire [63:0]   res_lo_hi_lo_103 = {dataGroup_5_103, dataGroup_4_103};
  wire [63:0]   res_lo_hi_hi_103 = {dataGroup_7_103, dataGroup_6_103};
  wire [127:0]  res_lo_hi_103 = {res_lo_hi_hi_103, res_lo_hi_lo_103};
  wire [255:0]  res_lo_103 = {res_lo_hi_103, res_lo_lo_103};
  wire [63:0]   res_hi_lo_lo_103 = {dataGroup_9_103, dataGroup_8_103};
  wire [63:0]   res_hi_lo_hi_103 = {dataGroup_11_103, dataGroup_10_103};
  wire [127:0]  res_hi_lo_103 = {res_hi_lo_hi_103, res_hi_lo_lo_103};
  wire [63:0]   res_hi_hi_lo_103 = {dataGroup_13_103, dataGroup_12_103};
  wire [63:0]   res_hi_hi_hi_103 = {dataGroup_15_103, dataGroup_14_103};
  wire [127:0]  res_hi_hi_103 = {res_hi_hi_hi_103, res_hi_hi_lo_103};
  wire [255:0]  res_hi_103 = {res_hi_hi_103, res_hi_lo_103};
  wire [511:0]  res_187 = {res_hi_103, res_lo_103};
  wire [2047:0] dataGroup_lo_3968 = {dataGroup_lo_hi_3968, dataGroup_lo_lo_3968};
  wire [2047:0] dataGroup_hi_3968 = {dataGroup_hi_hi_3968, dataGroup_hi_lo_3968};
  wire [31:0]   dataGroup_0_104 = dataGroup_lo_3968[159:128];
  wire [2047:0] dataGroup_lo_3969 = {dataGroup_lo_hi_3969, dataGroup_lo_lo_3969};
  wire [2047:0] dataGroup_hi_3969 = {dataGroup_hi_hi_3969, dataGroup_hi_lo_3969};
  wire [31:0]   dataGroup_1_104 = dataGroup_lo_3969[415:384];
  wire [2047:0] dataGroup_lo_3970 = {dataGroup_lo_hi_3970, dataGroup_lo_lo_3970};
  wire [2047:0] dataGroup_hi_3970 = {dataGroup_hi_hi_3970, dataGroup_hi_lo_3970};
  wire [31:0]   dataGroup_2_104 = dataGroup_lo_3970[671:640];
  wire [2047:0] dataGroup_lo_3971 = {dataGroup_lo_hi_3971, dataGroup_lo_lo_3971};
  wire [2047:0] dataGroup_hi_3971 = {dataGroup_hi_hi_3971, dataGroup_hi_lo_3971};
  wire [31:0]   dataGroup_3_104 = dataGroup_lo_3971[927:896];
  wire [2047:0] dataGroup_lo_3972 = {dataGroup_lo_hi_3972, dataGroup_lo_lo_3972};
  wire [2047:0] dataGroup_hi_3972 = {dataGroup_hi_hi_3972, dataGroup_hi_lo_3972};
  wire [31:0]   dataGroup_4_104 = dataGroup_lo_3972[1183:1152];
  wire [2047:0] dataGroup_lo_3973 = {dataGroup_lo_hi_3973, dataGroup_lo_lo_3973};
  wire [2047:0] dataGroup_hi_3973 = {dataGroup_hi_hi_3973, dataGroup_hi_lo_3973};
  wire [31:0]   dataGroup_5_104 = dataGroup_lo_3973[1439:1408];
  wire [2047:0] dataGroup_lo_3974 = {dataGroup_lo_hi_3974, dataGroup_lo_lo_3974};
  wire [2047:0] dataGroup_hi_3974 = {dataGroup_hi_hi_3974, dataGroup_hi_lo_3974};
  wire [31:0]   dataGroup_6_104 = dataGroup_lo_3974[1695:1664];
  wire [2047:0] dataGroup_lo_3975 = {dataGroup_lo_hi_3975, dataGroup_lo_lo_3975};
  wire [2047:0] dataGroup_hi_3975 = {dataGroup_hi_hi_3975, dataGroup_hi_lo_3975};
  wire [31:0]   dataGroup_7_104 = dataGroup_lo_3975[1951:1920];
  wire [2047:0] dataGroup_lo_3976 = {dataGroup_lo_hi_3976, dataGroup_lo_lo_3976};
  wire [2047:0] dataGroup_hi_3976 = {dataGroup_hi_hi_3976, dataGroup_hi_lo_3976};
  wire [31:0]   dataGroup_8_104 = dataGroup_hi_3976[159:128];
  wire [2047:0] dataGroup_lo_3977 = {dataGroup_lo_hi_3977, dataGroup_lo_lo_3977};
  wire [2047:0] dataGroup_hi_3977 = {dataGroup_hi_hi_3977, dataGroup_hi_lo_3977};
  wire [31:0]   dataGroup_9_104 = dataGroup_hi_3977[415:384];
  wire [2047:0] dataGroup_lo_3978 = {dataGroup_lo_hi_3978, dataGroup_lo_lo_3978};
  wire [2047:0] dataGroup_hi_3978 = {dataGroup_hi_hi_3978, dataGroup_hi_lo_3978};
  wire [31:0]   dataGroup_10_104 = dataGroup_hi_3978[671:640];
  wire [2047:0] dataGroup_lo_3979 = {dataGroup_lo_hi_3979, dataGroup_lo_lo_3979};
  wire [2047:0] dataGroup_hi_3979 = {dataGroup_hi_hi_3979, dataGroup_hi_lo_3979};
  wire [31:0]   dataGroup_11_104 = dataGroup_hi_3979[927:896];
  wire [2047:0] dataGroup_lo_3980 = {dataGroup_lo_hi_3980, dataGroup_lo_lo_3980};
  wire [2047:0] dataGroup_hi_3980 = {dataGroup_hi_hi_3980, dataGroup_hi_lo_3980};
  wire [31:0]   dataGroup_12_104 = dataGroup_hi_3980[1183:1152];
  wire [2047:0] dataGroup_lo_3981 = {dataGroup_lo_hi_3981, dataGroup_lo_lo_3981};
  wire [2047:0] dataGroup_hi_3981 = {dataGroup_hi_hi_3981, dataGroup_hi_lo_3981};
  wire [31:0]   dataGroup_13_104 = dataGroup_hi_3981[1439:1408];
  wire [2047:0] dataGroup_lo_3982 = {dataGroup_lo_hi_3982, dataGroup_lo_lo_3982};
  wire [2047:0] dataGroup_hi_3982 = {dataGroup_hi_hi_3982, dataGroup_hi_lo_3982};
  wire [31:0]   dataGroup_14_104 = dataGroup_hi_3982[1695:1664];
  wire [2047:0] dataGroup_lo_3983 = {dataGroup_lo_hi_3983, dataGroup_lo_lo_3983};
  wire [2047:0] dataGroup_hi_3983 = {dataGroup_hi_hi_3983, dataGroup_hi_lo_3983};
  wire [31:0]   dataGroup_15_104 = dataGroup_hi_3983[1951:1920];
  wire [63:0]   res_lo_lo_lo_104 = {dataGroup_1_104, dataGroup_0_104};
  wire [63:0]   res_lo_lo_hi_104 = {dataGroup_3_104, dataGroup_2_104};
  wire [127:0]  res_lo_lo_104 = {res_lo_lo_hi_104, res_lo_lo_lo_104};
  wire [63:0]   res_lo_hi_lo_104 = {dataGroup_5_104, dataGroup_4_104};
  wire [63:0]   res_lo_hi_hi_104 = {dataGroup_7_104, dataGroup_6_104};
  wire [127:0]  res_lo_hi_104 = {res_lo_hi_hi_104, res_lo_hi_lo_104};
  wire [255:0]  res_lo_104 = {res_lo_hi_104, res_lo_lo_104};
  wire [63:0]   res_hi_lo_lo_104 = {dataGroup_9_104, dataGroup_8_104};
  wire [63:0]   res_hi_lo_hi_104 = {dataGroup_11_104, dataGroup_10_104};
  wire [127:0]  res_hi_lo_104 = {res_hi_lo_hi_104, res_hi_lo_lo_104};
  wire [63:0]   res_hi_hi_lo_104 = {dataGroup_13_104, dataGroup_12_104};
  wire [63:0]   res_hi_hi_hi_104 = {dataGroup_15_104, dataGroup_14_104};
  wire [127:0]  res_hi_hi_104 = {res_hi_hi_hi_104, res_hi_hi_lo_104};
  wire [255:0]  res_hi_104 = {res_hi_hi_104, res_hi_lo_104};
  wire [511:0]  res_188 = {res_hi_104, res_lo_104};
  wire [2047:0] dataGroup_lo_3984 = {dataGroup_lo_hi_3984, dataGroup_lo_lo_3984};
  wire [2047:0] dataGroup_hi_3984 = {dataGroup_hi_hi_3984, dataGroup_hi_lo_3984};
  wire [31:0]   dataGroup_0_105 = dataGroup_lo_3984[191:160];
  wire [2047:0] dataGroup_lo_3985 = {dataGroup_lo_hi_3985, dataGroup_lo_lo_3985};
  wire [2047:0] dataGroup_hi_3985 = {dataGroup_hi_hi_3985, dataGroup_hi_lo_3985};
  wire [31:0]   dataGroup_1_105 = dataGroup_lo_3985[447:416];
  wire [2047:0] dataGroup_lo_3986 = {dataGroup_lo_hi_3986, dataGroup_lo_lo_3986};
  wire [2047:0] dataGroup_hi_3986 = {dataGroup_hi_hi_3986, dataGroup_hi_lo_3986};
  wire [31:0]   dataGroup_2_105 = dataGroup_lo_3986[703:672];
  wire [2047:0] dataGroup_lo_3987 = {dataGroup_lo_hi_3987, dataGroup_lo_lo_3987};
  wire [2047:0] dataGroup_hi_3987 = {dataGroup_hi_hi_3987, dataGroup_hi_lo_3987};
  wire [31:0]   dataGroup_3_105 = dataGroup_lo_3987[959:928];
  wire [2047:0] dataGroup_lo_3988 = {dataGroup_lo_hi_3988, dataGroup_lo_lo_3988};
  wire [2047:0] dataGroup_hi_3988 = {dataGroup_hi_hi_3988, dataGroup_hi_lo_3988};
  wire [31:0]   dataGroup_4_105 = dataGroup_lo_3988[1215:1184];
  wire [2047:0] dataGroup_lo_3989 = {dataGroup_lo_hi_3989, dataGroup_lo_lo_3989};
  wire [2047:0] dataGroup_hi_3989 = {dataGroup_hi_hi_3989, dataGroup_hi_lo_3989};
  wire [31:0]   dataGroup_5_105 = dataGroup_lo_3989[1471:1440];
  wire [2047:0] dataGroup_lo_3990 = {dataGroup_lo_hi_3990, dataGroup_lo_lo_3990};
  wire [2047:0] dataGroup_hi_3990 = {dataGroup_hi_hi_3990, dataGroup_hi_lo_3990};
  wire [31:0]   dataGroup_6_105 = dataGroup_lo_3990[1727:1696];
  wire [2047:0] dataGroup_lo_3991 = {dataGroup_lo_hi_3991, dataGroup_lo_lo_3991};
  wire [2047:0] dataGroup_hi_3991 = {dataGroup_hi_hi_3991, dataGroup_hi_lo_3991};
  wire [31:0]   dataGroup_7_105 = dataGroup_lo_3991[1983:1952];
  wire [2047:0] dataGroup_lo_3992 = {dataGroup_lo_hi_3992, dataGroup_lo_lo_3992};
  wire [2047:0] dataGroup_hi_3992 = {dataGroup_hi_hi_3992, dataGroup_hi_lo_3992};
  wire [31:0]   dataGroup_8_105 = dataGroup_hi_3992[191:160];
  wire [2047:0] dataGroup_lo_3993 = {dataGroup_lo_hi_3993, dataGroup_lo_lo_3993};
  wire [2047:0] dataGroup_hi_3993 = {dataGroup_hi_hi_3993, dataGroup_hi_lo_3993};
  wire [31:0]   dataGroup_9_105 = dataGroup_hi_3993[447:416];
  wire [2047:0] dataGroup_lo_3994 = {dataGroup_lo_hi_3994, dataGroup_lo_lo_3994};
  wire [2047:0] dataGroup_hi_3994 = {dataGroup_hi_hi_3994, dataGroup_hi_lo_3994};
  wire [31:0]   dataGroup_10_105 = dataGroup_hi_3994[703:672];
  wire [2047:0] dataGroup_lo_3995 = {dataGroup_lo_hi_3995, dataGroup_lo_lo_3995};
  wire [2047:0] dataGroup_hi_3995 = {dataGroup_hi_hi_3995, dataGroup_hi_lo_3995};
  wire [31:0]   dataGroup_11_105 = dataGroup_hi_3995[959:928];
  wire [2047:0] dataGroup_lo_3996 = {dataGroup_lo_hi_3996, dataGroup_lo_lo_3996};
  wire [2047:0] dataGroup_hi_3996 = {dataGroup_hi_hi_3996, dataGroup_hi_lo_3996};
  wire [31:0]   dataGroup_12_105 = dataGroup_hi_3996[1215:1184];
  wire [2047:0] dataGroup_lo_3997 = {dataGroup_lo_hi_3997, dataGroup_lo_lo_3997};
  wire [2047:0] dataGroup_hi_3997 = {dataGroup_hi_hi_3997, dataGroup_hi_lo_3997};
  wire [31:0]   dataGroup_13_105 = dataGroup_hi_3997[1471:1440];
  wire [2047:0] dataGroup_lo_3998 = {dataGroup_lo_hi_3998, dataGroup_lo_lo_3998};
  wire [2047:0] dataGroup_hi_3998 = {dataGroup_hi_hi_3998, dataGroup_hi_lo_3998};
  wire [31:0]   dataGroup_14_105 = dataGroup_hi_3998[1727:1696];
  wire [2047:0] dataGroup_lo_3999 = {dataGroup_lo_hi_3999, dataGroup_lo_lo_3999};
  wire [2047:0] dataGroup_hi_3999 = {dataGroup_hi_hi_3999, dataGroup_hi_lo_3999};
  wire [31:0]   dataGroup_15_105 = dataGroup_hi_3999[1983:1952];
  wire [63:0]   res_lo_lo_lo_105 = {dataGroup_1_105, dataGroup_0_105};
  wire [63:0]   res_lo_lo_hi_105 = {dataGroup_3_105, dataGroup_2_105};
  wire [127:0]  res_lo_lo_105 = {res_lo_lo_hi_105, res_lo_lo_lo_105};
  wire [63:0]   res_lo_hi_lo_105 = {dataGroup_5_105, dataGroup_4_105};
  wire [63:0]   res_lo_hi_hi_105 = {dataGroup_7_105, dataGroup_6_105};
  wire [127:0]  res_lo_hi_105 = {res_lo_hi_hi_105, res_lo_hi_lo_105};
  wire [255:0]  res_lo_105 = {res_lo_hi_105, res_lo_lo_105};
  wire [63:0]   res_hi_lo_lo_105 = {dataGroup_9_105, dataGroup_8_105};
  wire [63:0]   res_hi_lo_hi_105 = {dataGroup_11_105, dataGroup_10_105};
  wire [127:0]  res_hi_lo_105 = {res_hi_lo_hi_105, res_hi_lo_lo_105};
  wire [63:0]   res_hi_hi_lo_105 = {dataGroup_13_105, dataGroup_12_105};
  wire [63:0]   res_hi_hi_hi_105 = {dataGroup_15_105, dataGroup_14_105};
  wire [127:0]  res_hi_hi_105 = {res_hi_hi_hi_105, res_hi_hi_lo_105};
  wire [255:0]  res_hi_105 = {res_hi_hi_105, res_hi_lo_105};
  wire [511:0]  res_189 = {res_hi_105, res_lo_105};
  wire [2047:0] dataGroup_lo_4000 = {dataGroup_lo_hi_4000, dataGroup_lo_lo_4000};
  wire [2047:0] dataGroup_hi_4000 = {dataGroup_hi_hi_4000, dataGroup_hi_lo_4000};
  wire [31:0]   dataGroup_0_106 = dataGroup_lo_4000[223:192];
  wire [2047:0] dataGroup_lo_4001 = {dataGroup_lo_hi_4001, dataGroup_lo_lo_4001};
  wire [2047:0] dataGroup_hi_4001 = {dataGroup_hi_hi_4001, dataGroup_hi_lo_4001};
  wire [31:0]   dataGroup_1_106 = dataGroup_lo_4001[479:448];
  wire [2047:0] dataGroup_lo_4002 = {dataGroup_lo_hi_4002, dataGroup_lo_lo_4002};
  wire [2047:0] dataGroup_hi_4002 = {dataGroup_hi_hi_4002, dataGroup_hi_lo_4002};
  wire [31:0]   dataGroup_2_106 = dataGroup_lo_4002[735:704];
  wire [2047:0] dataGroup_lo_4003 = {dataGroup_lo_hi_4003, dataGroup_lo_lo_4003};
  wire [2047:0] dataGroup_hi_4003 = {dataGroup_hi_hi_4003, dataGroup_hi_lo_4003};
  wire [31:0]   dataGroup_3_106 = dataGroup_lo_4003[991:960];
  wire [2047:0] dataGroup_lo_4004 = {dataGroup_lo_hi_4004, dataGroup_lo_lo_4004};
  wire [2047:0] dataGroup_hi_4004 = {dataGroup_hi_hi_4004, dataGroup_hi_lo_4004};
  wire [31:0]   dataGroup_4_106 = dataGroup_lo_4004[1247:1216];
  wire [2047:0] dataGroup_lo_4005 = {dataGroup_lo_hi_4005, dataGroup_lo_lo_4005};
  wire [2047:0] dataGroup_hi_4005 = {dataGroup_hi_hi_4005, dataGroup_hi_lo_4005};
  wire [31:0]   dataGroup_5_106 = dataGroup_lo_4005[1503:1472];
  wire [2047:0] dataGroup_lo_4006 = {dataGroup_lo_hi_4006, dataGroup_lo_lo_4006};
  wire [2047:0] dataGroup_hi_4006 = {dataGroup_hi_hi_4006, dataGroup_hi_lo_4006};
  wire [31:0]   dataGroup_6_106 = dataGroup_lo_4006[1759:1728];
  wire [2047:0] dataGroup_lo_4007 = {dataGroup_lo_hi_4007, dataGroup_lo_lo_4007};
  wire [2047:0] dataGroup_hi_4007 = {dataGroup_hi_hi_4007, dataGroup_hi_lo_4007};
  wire [31:0]   dataGroup_7_106 = dataGroup_lo_4007[2015:1984];
  wire [2047:0] dataGroup_lo_4008 = {dataGroup_lo_hi_4008, dataGroup_lo_lo_4008};
  wire [2047:0] dataGroup_hi_4008 = {dataGroup_hi_hi_4008, dataGroup_hi_lo_4008};
  wire [31:0]   dataGroup_8_106 = dataGroup_hi_4008[223:192];
  wire [2047:0] dataGroup_lo_4009 = {dataGroup_lo_hi_4009, dataGroup_lo_lo_4009};
  wire [2047:0] dataGroup_hi_4009 = {dataGroup_hi_hi_4009, dataGroup_hi_lo_4009};
  wire [31:0]   dataGroup_9_106 = dataGroup_hi_4009[479:448];
  wire [2047:0] dataGroup_lo_4010 = {dataGroup_lo_hi_4010, dataGroup_lo_lo_4010};
  wire [2047:0] dataGroup_hi_4010 = {dataGroup_hi_hi_4010, dataGroup_hi_lo_4010};
  wire [31:0]   dataGroup_10_106 = dataGroup_hi_4010[735:704];
  wire [2047:0] dataGroup_lo_4011 = {dataGroup_lo_hi_4011, dataGroup_lo_lo_4011};
  wire [2047:0] dataGroup_hi_4011 = {dataGroup_hi_hi_4011, dataGroup_hi_lo_4011};
  wire [31:0]   dataGroup_11_106 = dataGroup_hi_4011[991:960];
  wire [2047:0] dataGroup_lo_4012 = {dataGroup_lo_hi_4012, dataGroup_lo_lo_4012};
  wire [2047:0] dataGroup_hi_4012 = {dataGroup_hi_hi_4012, dataGroup_hi_lo_4012};
  wire [31:0]   dataGroup_12_106 = dataGroup_hi_4012[1247:1216];
  wire [2047:0] dataGroup_lo_4013 = {dataGroup_lo_hi_4013, dataGroup_lo_lo_4013};
  wire [2047:0] dataGroup_hi_4013 = {dataGroup_hi_hi_4013, dataGroup_hi_lo_4013};
  wire [31:0]   dataGroup_13_106 = dataGroup_hi_4013[1503:1472];
  wire [2047:0] dataGroup_lo_4014 = {dataGroup_lo_hi_4014, dataGroup_lo_lo_4014};
  wire [2047:0] dataGroup_hi_4014 = {dataGroup_hi_hi_4014, dataGroup_hi_lo_4014};
  wire [31:0]   dataGroup_14_106 = dataGroup_hi_4014[1759:1728];
  wire [2047:0] dataGroup_lo_4015 = {dataGroup_lo_hi_4015, dataGroup_lo_lo_4015};
  wire [2047:0] dataGroup_hi_4015 = {dataGroup_hi_hi_4015, dataGroup_hi_lo_4015};
  wire [31:0]   dataGroup_15_106 = dataGroup_hi_4015[2015:1984];
  wire [63:0]   res_lo_lo_lo_106 = {dataGroup_1_106, dataGroup_0_106};
  wire [63:0]   res_lo_lo_hi_106 = {dataGroup_3_106, dataGroup_2_106};
  wire [127:0]  res_lo_lo_106 = {res_lo_lo_hi_106, res_lo_lo_lo_106};
  wire [63:0]   res_lo_hi_lo_106 = {dataGroup_5_106, dataGroup_4_106};
  wire [63:0]   res_lo_hi_hi_106 = {dataGroup_7_106, dataGroup_6_106};
  wire [127:0]  res_lo_hi_106 = {res_lo_hi_hi_106, res_lo_hi_lo_106};
  wire [255:0]  res_lo_106 = {res_lo_hi_106, res_lo_lo_106};
  wire [63:0]   res_hi_lo_lo_106 = {dataGroup_9_106, dataGroup_8_106};
  wire [63:0]   res_hi_lo_hi_106 = {dataGroup_11_106, dataGroup_10_106};
  wire [127:0]  res_hi_lo_106 = {res_hi_lo_hi_106, res_hi_lo_lo_106};
  wire [63:0]   res_hi_hi_lo_106 = {dataGroup_13_106, dataGroup_12_106};
  wire [63:0]   res_hi_hi_hi_106 = {dataGroup_15_106, dataGroup_14_106};
  wire [127:0]  res_hi_hi_106 = {res_hi_hi_hi_106, res_hi_hi_lo_106};
  wire [255:0]  res_hi_106 = {res_hi_hi_106, res_hi_lo_106};
  wire [511:0]  res_190 = {res_hi_106, res_lo_106};
  wire [2047:0] dataGroup_lo_4016 = {dataGroup_lo_hi_4016, dataGroup_lo_lo_4016};
  wire [2047:0] dataGroup_hi_4016 = {dataGroup_hi_hi_4016, dataGroup_hi_lo_4016};
  wire [31:0]   dataGroup_0_107 = dataGroup_lo_4016[255:224];
  wire [2047:0] dataGroup_lo_4017 = {dataGroup_lo_hi_4017, dataGroup_lo_lo_4017};
  wire [2047:0] dataGroup_hi_4017 = {dataGroup_hi_hi_4017, dataGroup_hi_lo_4017};
  wire [31:0]   dataGroup_1_107 = dataGroup_lo_4017[511:480];
  wire [2047:0] dataGroup_lo_4018 = {dataGroup_lo_hi_4018, dataGroup_lo_lo_4018};
  wire [2047:0] dataGroup_hi_4018 = {dataGroup_hi_hi_4018, dataGroup_hi_lo_4018};
  wire [31:0]   dataGroup_2_107 = dataGroup_lo_4018[767:736];
  wire [2047:0] dataGroup_lo_4019 = {dataGroup_lo_hi_4019, dataGroup_lo_lo_4019};
  wire [2047:0] dataGroup_hi_4019 = {dataGroup_hi_hi_4019, dataGroup_hi_lo_4019};
  wire [31:0]   dataGroup_3_107 = dataGroup_lo_4019[1023:992];
  wire [2047:0] dataGroup_lo_4020 = {dataGroup_lo_hi_4020, dataGroup_lo_lo_4020};
  wire [2047:0] dataGroup_hi_4020 = {dataGroup_hi_hi_4020, dataGroup_hi_lo_4020};
  wire [31:0]   dataGroup_4_107 = dataGroup_lo_4020[1279:1248];
  wire [2047:0] dataGroup_lo_4021 = {dataGroup_lo_hi_4021, dataGroup_lo_lo_4021};
  wire [2047:0] dataGroup_hi_4021 = {dataGroup_hi_hi_4021, dataGroup_hi_lo_4021};
  wire [31:0]   dataGroup_5_107 = dataGroup_lo_4021[1535:1504];
  wire [2047:0] dataGroup_lo_4022 = {dataGroup_lo_hi_4022, dataGroup_lo_lo_4022};
  wire [2047:0] dataGroup_hi_4022 = {dataGroup_hi_hi_4022, dataGroup_hi_lo_4022};
  wire [31:0]   dataGroup_6_107 = dataGroup_lo_4022[1791:1760];
  wire [2047:0] dataGroup_lo_4023 = {dataGroup_lo_hi_4023, dataGroup_lo_lo_4023};
  wire [2047:0] dataGroup_hi_4023 = {dataGroup_hi_hi_4023, dataGroup_hi_lo_4023};
  wire [31:0]   dataGroup_7_107 = dataGroup_lo_4023[2047:2016];
  wire [2047:0] dataGroup_lo_4024 = {dataGroup_lo_hi_4024, dataGroup_lo_lo_4024};
  wire [2047:0] dataGroup_hi_4024 = {dataGroup_hi_hi_4024, dataGroup_hi_lo_4024};
  wire [31:0]   dataGroup_8_107 = dataGroup_hi_4024[255:224];
  wire [2047:0] dataGroup_lo_4025 = {dataGroup_lo_hi_4025, dataGroup_lo_lo_4025};
  wire [2047:0] dataGroup_hi_4025 = {dataGroup_hi_hi_4025, dataGroup_hi_lo_4025};
  wire [31:0]   dataGroup_9_107 = dataGroup_hi_4025[511:480];
  wire [2047:0] dataGroup_lo_4026 = {dataGroup_lo_hi_4026, dataGroup_lo_lo_4026};
  wire [2047:0] dataGroup_hi_4026 = {dataGroup_hi_hi_4026, dataGroup_hi_lo_4026};
  wire [31:0]   dataGroup_10_107 = dataGroup_hi_4026[767:736];
  wire [2047:0] dataGroup_lo_4027 = {dataGroup_lo_hi_4027, dataGroup_lo_lo_4027};
  wire [2047:0] dataGroup_hi_4027 = {dataGroup_hi_hi_4027, dataGroup_hi_lo_4027};
  wire [31:0]   dataGroup_11_107 = dataGroup_hi_4027[1023:992];
  wire [2047:0] dataGroup_lo_4028 = {dataGroup_lo_hi_4028, dataGroup_lo_lo_4028};
  wire [2047:0] dataGroup_hi_4028 = {dataGroup_hi_hi_4028, dataGroup_hi_lo_4028};
  wire [31:0]   dataGroup_12_107 = dataGroup_hi_4028[1279:1248];
  wire [2047:0] dataGroup_lo_4029 = {dataGroup_lo_hi_4029, dataGroup_lo_lo_4029};
  wire [2047:0] dataGroup_hi_4029 = {dataGroup_hi_hi_4029, dataGroup_hi_lo_4029};
  wire [31:0]   dataGroup_13_107 = dataGroup_hi_4029[1535:1504];
  wire [2047:0] dataGroup_lo_4030 = {dataGroup_lo_hi_4030, dataGroup_lo_lo_4030};
  wire [2047:0] dataGroup_hi_4030 = {dataGroup_hi_hi_4030, dataGroup_hi_lo_4030};
  wire [31:0]   dataGroup_14_107 = dataGroup_hi_4030[1791:1760];
  wire [2047:0] dataGroup_lo_4031 = {dataGroup_lo_hi_4031, dataGroup_lo_lo_4031};
  wire [2047:0] dataGroup_hi_4031 = {dataGroup_hi_hi_4031, dataGroup_hi_lo_4031};
  wire [31:0]   dataGroup_15_107 = dataGroup_hi_4031[2047:2016];
  wire [63:0]   res_lo_lo_lo_107 = {dataGroup_1_107, dataGroup_0_107};
  wire [63:0]   res_lo_lo_hi_107 = {dataGroup_3_107, dataGroup_2_107};
  wire [127:0]  res_lo_lo_107 = {res_lo_lo_hi_107, res_lo_lo_lo_107};
  wire [63:0]   res_lo_hi_lo_107 = {dataGroup_5_107, dataGroup_4_107};
  wire [63:0]   res_lo_hi_hi_107 = {dataGroup_7_107, dataGroup_6_107};
  wire [127:0]  res_lo_hi_107 = {res_lo_hi_hi_107, res_lo_hi_lo_107};
  wire [255:0]  res_lo_107 = {res_lo_hi_107, res_lo_lo_107};
  wire [63:0]   res_hi_lo_lo_107 = {dataGroup_9_107, dataGroup_8_107};
  wire [63:0]   res_hi_lo_hi_107 = {dataGroup_11_107, dataGroup_10_107};
  wire [127:0]  res_hi_lo_107 = {res_hi_lo_hi_107, res_hi_lo_lo_107};
  wire [63:0]   res_hi_hi_lo_107 = {dataGroup_13_107, dataGroup_12_107};
  wire [63:0]   res_hi_hi_hi_107 = {dataGroup_15_107, dataGroup_14_107};
  wire [127:0]  res_hi_hi_107 = {res_hi_hi_hi_107, res_hi_hi_lo_107};
  wire [255:0]  res_hi_107 = {res_hi_hi_107, res_hi_lo_107};
  wire [511:0]  res_191 = {res_hi_107, res_lo_107};
  wire [1023:0] lo_lo_23 = {res_185, res_184};
  wire [1023:0] lo_hi_23 = {res_187, res_186};
  wire [2047:0] lo_23 = {lo_hi_23, lo_lo_23};
  wire [1023:0] hi_lo_23 = {res_189, res_188};
  wire [1023:0] hi_hi_23 = {res_191, res_190};
  wire [2047:0] hi_23 = {hi_hi_23, hi_lo_23};
  wire [4095:0] regroupLoadData_2_7 = {hi_23, lo_23};
  wire          vrfWritePort_0_valid_0 = accessState_0 & writeReadyReg;
  wire [3:0]    vrfWritePort_0_bits_mask_0 = maskForGroup[3:0];
  wire [3:0]    vrfWritePort_1_bits_mask_0 = maskForGroup[7:4];
  wire [3:0]    vrfWritePort_2_bits_mask_0 = maskForGroup[11:8];
  wire [3:0]    vrfWritePort_3_bits_mask_0 = maskForGroup[15:12];
  wire [3:0]    vrfWritePort_4_bits_mask_0 = maskForGroup[19:16];
  wire [3:0]    vrfWritePort_5_bits_mask_0 = maskForGroup[23:20];
  wire [3:0]    vrfWritePort_6_bits_mask_0 = maskForGroup[27:24];
  wire [3:0]    vrfWritePort_7_bits_mask_0 = maskForGroup[31:28];
  wire [3:0]    vrfWritePort_8_bits_mask_0 = maskForGroup[35:32];
  wire [3:0]    vrfWritePort_9_bits_mask_0 = maskForGroup[39:36];
  wire [3:0]    vrfWritePort_10_bits_mask_0 = maskForGroup[43:40];
  wire [3:0]    vrfWritePort_11_bits_mask_0 = maskForGroup[47:44];
  wire [3:0]    vrfWritePort_12_bits_mask_0 = maskForGroup[51:48];
  wire [3:0]    vrfWritePort_13_bits_mask_0 = maskForGroup[55:52];
  wire [3:0]    vrfWritePort_14_bits_mask_0 = maskForGroup[59:56];
  wire [3:0]    vrfWritePort_15_bits_mask_0 = maskForGroup[63:60];
  wire [7:0]    _vrfWritePort_15_bits_data_T = 8'h1 << accessPtr;
  wire [31:0]   vrfWritePort_0_bits_data_0 =
    (_vrfWritePort_15_bits_data_T[0] ? accessData_0[31:0] : 32'h0) | (_vrfWritePort_15_bits_data_T[1] ? accessData_1[31:0] : 32'h0) | (_vrfWritePort_15_bits_data_T[2] ? accessData_2[31:0] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[3] ? accessData_3[31:0] : 32'h0) | (_vrfWritePort_15_bits_data_T[4] ? accessData_4[31:0] : 32'h0) | (_vrfWritePort_15_bits_data_T[5] ? accessData_5[31:0] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[6] ? accessData_6[31:0] : 32'h0) | (_vrfWritePort_15_bits_data_T[7] ? accessData_7[31:0] : 32'h0);
  wire          vrfWritePort_0_bits_offset_0 = dataGroup[0];
  wire          vrfWritePort_1_bits_offset_0 = dataGroup[0];
  wire          vrfWritePort_2_bits_offset_0 = dataGroup[0];
  wire          vrfWritePort_3_bits_offset_0 = dataGroup[0];
  wire          vrfWritePort_4_bits_offset_0 = dataGroup[0];
  wire          vrfWritePort_5_bits_offset_0 = dataGroup[0];
  wire          vrfWritePort_6_bits_offset_0 = dataGroup[0];
  wire          vrfWritePort_7_bits_offset_0 = dataGroup[0];
  wire          vrfWritePort_8_bits_offset_0 = dataGroup[0];
  wire          vrfWritePort_9_bits_offset_0 = dataGroup[0];
  wire          vrfWritePort_10_bits_offset_0 = dataGroup[0];
  wire          vrfWritePort_11_bits_offset_0 = dataGroup[0];
  wire          vrfWritePort_12_bits_offset_0 = dataGroup[0];
  wire          vrfWritePort_13_bits_offset_0 = dataGroup[0];
  wire          vrfWritePort_14_bits_offset_0 = dataGroup[0];
  wire          vrfWritePort_15_bits_offset_0 = dataGroup[0];
  wire [4:0]    _GEN_9 = {2'h0, accessPtr} * {1'h0, segmentInstructionIndexInterval} + {2'h0, dataGroup[3:1]};
  wire [4:0]    vrfWritePort_0_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_9;
  assign accessStateUpdate_0 = ~(vrfWritePort_0_ready_0 & vrfWritePort_0_valid_0) & accessState_0;
  wire          vrfWritePort_1_valid_0 = accessState_1 & writeReadyReg;
  wire [31:0]   vrfWritePort_1_bits_data_0 =
    (_vrfWritePort_15_bits_data_T[0] ? accessData_0[63:32] : 32'h0) | (_vrfWritePort_15_bits_data_T[1] ? accessData_1[63:32] : 32'h0) | (_vrfWritePort_15_bits_data_T[2] ? accessData_2[63:32] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[3] ? accessData_3[63:32] : 32'h0) | (_vrfWritePort_15_bits_data_T[4] ? accessData_4[63:32] : 32'h0) | (_vrfWritePort_15_bits_data_T[5] ? accessData_5[63:32] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[6] ? accessData_6[63:32] : 32'h0) | (_vrfWritePort_15_bits_data_T[7] ? accessData_7[63:32] : 32'h0);
  wire [4:0]    vrfWritePort_1_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_9;
  assign accessStateUpdate_1 = ~(vrfWritePort_1_ready_0 & vrfWritePort_1_valid_0) & accessState_1;
  wire          vrfWritePort_2_valid_0 = accessState_2 & writeReadyReg;
  wire [31:0]   vrfWritePort_2_bits_data_0 =
    (_vrfWritePort_15_bits_data_T[0] ? accessData_0[95:64] : 32'h0) | (_vrfWritePort_15_bits_data_T[1] ? accessData_1[95:64] : 32'h0) | (_vrfWritePort_15_bits_data_T[2] ? accessData_2[95:64] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[3] ? accessData_3[95:64] : 32'h0) | (_vrfWritePort_15_bits_data_T[4] ? accessData_4[95:64] : 32'h0) | (_vrfWritePort_15_bits_data_T[5] ? accessData_5[95:64] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[6] ? accessData_6[95:64] : 32'h0) | (_vrfWritePort_15_bits_data_T[7] ? accessData_7[95:64] : 32'h0);
  wire [4:0]    vrfWritePort_2_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_9;
  assign accessStateUpdate_2 = ~(vrfWritePort_2_ready_0 & vrfWritePort_2_valid_0) & accessState_2;
  wire          vrfWritePort_3_valid_0 = accessState_3 & writeReadyReg;
  wire [31:0]   vrfWritePort_3_bits_data_0 =
    (_vrfWritePort_15_bits_data_T[0] ? accessData_0[127:96] : 32'h0) | (_vrfWritePort_15_bits_data_T[1] ? accessData_1[127:96] : 32'h0) | (_vrfWritePort_15_bits_data_T[2] ? accessData_2[127:96] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[3] ? accessData_3[127:96] : 32'h0) | (_vrfWritePort_15_bits_data_T[4] ? accessData_4[127:96] : 32'h0) | (_vrfWritePort_15_bits_data_T[5] ? accessData_5[127:96] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[6] ? accessData_6[127:96] : 32'h0) | (_vrfWritePort_15_bits_data_T[7] ? accessData_7[127:96] : 32'h0);
  wire [4:0]    vrfWritePort_3_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_9;
  assign accessStateUpdate_3 = ~(vrfWritePort_3_ready_0 & vrfWritePort_3_valid_0) & accessState_3;
  wire          vrfWritePort_4_valid_0 = accessState_4 & writeReadyReg;
  wire [31:0]   vrfWritePort_4_bits_data_0 =
    (_vrfWritePort_15_bits_data_T[0] ? accessData_0[159:128] : 32'h0) | (_vrfWritePort_15_bits_data_T[1] ? accessData_1[159:128] : 32'h0) | (_vrfWritePort_15_bits_data_T[2] ? accessData_2[159:128] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[3] ? accessData_3[159:128] : 32'h0) | (_vrfWritePort_15_bits_data_T[4] ? accessData_4[159:128] : 32'h0) | (_vrfWritePort_15_bits_data_T[5] ? accessData_5[159:128] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[6] ? accessData_6[159:128] : 32'h0) | (_vrfWritePort_15_bits_data_T[7] ? accessData_7[159:128] : 32'h0);
  wire [4:0]    vrfWritePort_4_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_9;
  assign accessStateUpdate_4 = ~(vrfWritePort_4_ready_0 & vrfWritePort_4_valid_0) & accessState_4;
  wire          vrfWritePort_5_valid_0 = accessState_5 & writeReadyReg;
  wire [31:0]   vrfWritePort_5_bits_data_0 =
    (_vrfWritePort_15_bits_data_T[0] ? accessData_0[191:160] : 32'h0) | (_vrfWritePort_15_bits_data_T[1] ? accessData_1[191:160] : 32'h0) | (_vrfWritePort_15_bits_data_T[2] ? accessData_2[191:160] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[3] ? accessData_3[191:160] : 32'h0) | (_vrfWritePort_15_bits_data_T[4] ? accessData_4[191:160] : 32'h0) | (_vrfWritePort_15_bits_data_T[5] ? accessData_5[191:160] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[6] ? accessData_6[191:160] : 32'h0) | (_vrfWritePort_15_bits_data_T[7] ? accessData_7[191:160] : 32'h0);
  wire [4:0]    vrfWritePort_5_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_9;
  assign accessStateUpdate_5 = ~(vrfWritePort_5_ready_0 & vrfWritePort_5_valid_0) & accessState_5;
  wire          vrfWritePort_6_valid_0 = accessState_6 & writeReadyReg;
  wire [31:0]   vrfWritePort_6_bits_data_0 =
    (_vrfWritePort_15_bits_data_T[0] ? accessData_0[223:192] : 32'h0) | (_vrfWritePort_15_bits_data_T[1] ? accessData_1[223:192] : 32'h0) | (_vrfWritePort_15_bits_data_T[2] ? accessData_2[223:192] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[3] ? accessData_3[223:192] : 32'h0) | (_vrfWritePort_15_bits_data_T[4] ? accessData_4[223:192] : 32'h0) | (_vrfWritePort_15_bits_data_T[5] ? accessData_5[223:192] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[6] ? accessData_6[223:192] : 32'h0) | (_vrfWritePort_15_bits_data_T[7] ? accessData_7[223:192] : 32'h0);
  wire [4:0]    vrfWritePort_6_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_9;
  assign accessStateUpdate_6 = ~(vrfWritePort_6_ready_0 & vrfWritePort_6_valid_0) & accessState_6;
  wire          vrfWritePort_7_valid_0 = accessState_7 & writeReadyReg;
  wire [31:0]   vrfWritePort_7_bits_data_0 =
    (_vrfWritePort_15_bits_data_T[0] ? accessData_0[255:224] : 32'h0) | (_vrfWritePort_15_bits_data_T[1] ? accessData_1[255:224] : 32'h0) | (_vrfWritePort_15_bits_data_T[2] ? accessData_2[255:224] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[3] ? accessData_3[255:224] : 32'h0) | (_vrfWritePort_15_bits_data_T[4] ? accessData_4[255:224] : 32'h0) | (_vrfWritePort_15_bits_data_T[5] ? accessData_5[255:224] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[6] ? accessData_6[255:224] : 32'h0) | (_vrfWritePort_15_bits_data_T[7] ? accessData_7[255:224] : 32'h0);
  wire [4:0]    vrfWritePort_7_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_9;
  assign accessStateUpdate_7 = ~(vrfWritePort_7_ready_0 & vrfWritePort_7_valid_0) & accessState_7;
  wire          vrfWritePort_8_valid_0 = accessState_8 & writeReadyReg;
  wire [31:0]   vrfWritePort_8_bits_data_0 =
    (_vrfWritePort_15_bits_data_T[0] ? accessData_0[287:256] : 32'h0) | (_vrfWritePort_15_bits_data_T[1] ? accessData_1[287:256] : 32'h0) | (_vrfWritePort_15_bits_data_T[2] ? accessData_2[287:256] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[3] ? accessData_3[287:256] : 32'h0) | (_vrfWritePort_15_bits_data_T[4] ? accessData_4[287:256] : 32'h0) | (_vrfWritePort_15_bits_data_T[5] ? accessData_5[287:256] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[6] ? accessData_6[287:256] : 32'h0) | (_vrfWritePort_15_bits_data_T[7] ? accessData_7[287:256] : 32'h0);
  wire [4:0]    vrfWritePort_8_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_9;
  assign accessStateUpdate_8 = ~(vrfWritePort_8_ready_0 & vrfWritePort_8_valid_0) & accessState_8;
  wire          vrfWritePort_9_valid_0 = accessState_9 & writeReadyReg;
  wire [31:0]   vrfWritePort_9_bits_data_0 =
    (_vrfWritePort_15_bits_data_T[0] ? accessData_0[319:288] : 32'h0) | (_vrfWritePort_15_bits_data_T[1] ? accessData_1[319:288] : 32'h0) | (_vrfWritePort_15_bits_data_T[2] ? accessData_2[319:288] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[3] ? accessData_3[319:288] : 32'h0) | (_vrfWritePort_15_bits_data_T[4] ? accessData_4[319:288] : 32'h0) | (_vrfWritePort_15_bits_data_T[5] ? accessData_5[319:288] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[6] ? accessData_6[319:288] : 32'h0) | (_vrfWritePort_15_bits_data_T[7] ? accessData_7[319:288] : 32'h0);
  wire [4:0]    vrfWritePort_9_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_9;
  assign accessStateUpdate_9 = ~(vrfWritePort_9_ready_0 & vrfWritePort_9_valid_0) & accessState_9;
  wire          vrfWritePort_10_valid_0 = accessState_10 & writeReadyReg;
  wire [31:0]   vrfWritePort_10_bits_data_0 =
    (_vrfWritePort_15_bits_data_T[0] ? accessData_0[351:320] : 32'h0) | (_vrfWritePort_15_bits_data_T[1] ? accessData_1[351:320] : 32'h0) | (_vrfWritePort_15_bits_data_T[2] ? accessData_2[351:320] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[3] ? accessData_3[351:320] : 32'h0) | (_vrfWritePort_15_bits_data_T[4] ? accessData_4[351:320] : 32'h0) | (_vrfWritePort_15_bits_data_T[5] ? accessData_5[351:320] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[6] ? accessData_6[351:320] : 32'h0) | (_vrfWritePort_15_bits_data_T[7] ? accessData_7[351:320] : 32'h0);
  wire [4:0]    vrfWritePort_10_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_9;
  assign accessStateUpdate_10 = ~(vrfWritePort_10_ready_0 & vrfWritePort_10_valid_0) & accessState_10;
  wire          vrfWritePort_11_valid_0 = accessState_11 & writeReadyReg;
  wire [31:0]   vrfWritePort_11_bits_data_0 =
    (_vrfWritePort_15_bits_data_T[0] ? accessData_0[383:352] : 32'h0) | (_vrfWritePort_15_bits_data_T[1] ? accessData_1[383:352] : 32'h0) | (_vrfWritePort_15_bits_data_T[2] ? accessData_2[383:352] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[3] ? accessData_3[383:352] : 32'h0) | (_vrfWritePort_15_bits_data_T[4] ? accessData_4[383:352] : 32'h0) | (_vrfWritePort_15_bits_data_T[5] ? accessData_5[383:352] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[6] ? accessData_6[383:352] : 32'h0) | (_vrfWritePort_15_bits_data_T[7] ? accessData_7[383:352] : 32'h0);
  wire [4:0]    vrfWritePort_11_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_9;
  assign accessStateUpdate_11 = ~(vrfWritePort_11_ready_0 & vrfWritePort_11_valid_0) & accessState_11;
  wire          vrfWritePort_12_valid_0 = accessState_12 & writeReadyReg;
  wire [31:0]   vrfWritePort_12_bits_data_0 =
    (_vrfWritePort_15_bits_data_T[0] ? accessData_0[415:384] : 32'h0) | (_vrfWritePort_15_bits_data_T[1] ? accessData_1[415:384] : 32'h0) | (_vrfWritePort_15_bits_data_T[2] ? accessData_2[415:384] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[3] ? accessData_3[415:384] : 32'h0) | (_vrfWritePort_15_bits_data_T[4] ? accessData_4[415:384] : 32'h0) | (_vrfWritePort_15_bits_data_T[5] ? accessData_5[415:384] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[6] ? accessData_6[415:384] : 32'h0) | (_vrfWritePort_15_bits_data_T[7] ? accessData_7[415:384] : 32'h0);
  wire [4:0]    vrfWritePort_12_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_9;
  assign accessStateUpdate_12 = ~(vrfWritePort_12_ready_0 & vrfWritePort_12_valid_0) & accessState_12;
  wire          vrfWritePort_13_valid_0 = accessState_13 & writeReadyReg;
  wire [31:0]   vrfWritePort_13_bits_data_0 =
    (_vrfWritePort_15_bits_data_T[0] ? accessData_0[447:416] : 32'h0) | (_vrfWritePort_15_bits_data_T[1] ? accessData_1[447:416] : 32'h0) | (_vrfWritePort_15_bits_data_T[2] ? accessData_2[447:416] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[3] ? accessData_3[447:416] : 32'h0) | (_vrfWritePort_15_bits_data_T[4] ? accessData_4[447:416] : 32'h0) | (_vrfWritePort_15_bits_data_T[5] ? accessData_5[447:416] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[6] ? accessData_6[447:416] : 32'h0) | (_vrfWritePort_15_bits_data_T[7] ? accessData_7[447:416] : 32'h0);
  wire [4:0]    vrfWritePort_13_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_9;
  assign accessStateUpdate_13 = ~(vrfWritePort_13_ready_0 & vrfWritePort_13_valid_0) & accessState_13;
  wire          vrfWritePort_14_valid_0 = accessState_14 & writeReadyReg;
  wire [31:0]   vrfWritePort_14_bits_data_0 =
    (_vrfWritePort_15_bits_data_T[0] ? accessData_0[479:448] : 32'h0) | (_vrfWritePort_15_bits_data_T[1] ? accessData_1[479:448] : 32'h0) | (_vrfWritePort_15_bits_data_T[2] ? accessData_2[479:448] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[3] ? accessData_3[479:448] : 32'h0) | (_vrfWritePort_15_bits_data_T[4] ? accessData_4[479:448] : 32'h0) | (_vrfWritePort_15_bits_data_T[5] ? accessData_5[479:448] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[6] ? accessData_6[479:448] : 32'h0) | (_vrfWritePort_15_bits_data_T[7] ? accessData_7[479:448] : 32'h0);
  wire [4:0]    vrfWritePort_14_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_9;
  assign accessStateUpdate_14 = ~(vrfWritePort_14_ready_0 & vrfWritePort_14_valid_0) & accessState_14;
  wire          vrfWritePort_15_valid_0 = accessState_15 & writeReadyReg;
  wire [31:0]   vrfWritePort_15_bits_data_0 =
    (_vrfWritePort_15_bits_data_T[0] ? accessData_0[511:480] : 32'h0) | (_vrfWritePort_15_bits_data_T[1] ? accessData_1[511:480] : 32'h0) | (_vrfWritePort_15_bits_data_T[2] ? accessData_2[511:480] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[3] ? accessData_3[511:480] : 32'h0) | (_vrfWritePort_15_bits_data_T[4] ? accessData_4[511:480] : 32'h0) | (_vrfWritePort_15_bits_data_T[5] ? accessData_5[511:480] : 32'h0)
    | (_vrfWritePort_15_bits_data_T[6] ? accessData_6[511:480] : 32'h0) | (_vrfWritePort_15_bits_data_T[7] ? accessData_7[511:480] : 32'h0);
  wire [4:0]    vrfWritePort_15_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_9;
  assign accessStateUpdate_15 = ~(vrfWritePort_15_ready_0 & vrfWritePort_15_valid_0) & accessState_15;
  reg           sendStateReg_0;
  reg           sendStateReg_1;
  reg           sendStateReg_2;
  reg           sendStateReg_3;
  reg           sendStateReg_4;
  reg           sendStateReg_5;
  reg           sendStateReg_6;
  reg           sendStateReg_7;
  reg           sendStateReg_8;
  reg           sendStateReg_9;
  reg           sendStateReg_10;
  reg           sendStateReg_11;
  reg           sendStateReg_12;
  reg           sendStateReg_13;
  reg           sendStateReg_14;
  reg           sendStateReg_15;
  wire          lastCacheRequest = lastRequest & _lastCacheRequest_T;
  reg           lastCacheRequestReg;
  reg           lastCacheLineAckReg;
  wire          bufferClear = ~(memResponse_valid_0 | alignedDequeue_valid | bufferFull | ~writeStageReady);
  wire          _status_idle_output = lastCacheRequestReg & lastCacheLineAckReg & bufferClear & ~sendRequest;
  reg           idleNext;
  always @(posedge clock) begin
    if (reset) begin
      lsuRequestReg_instructionInformation_nf <= 3'h0;
      lsuRequestReg_instructionInformation_mew <= 1'h0;
      lsuRequestReg_instructionInformation_mop <= 2'h0;
      lsuRequestReg_instructionInformation_lumop <= 5'h0;
      lsuRequestReg_instructionInformation_eew <= 2'h0;
      lsuRequestReg_instructionInformation_vs3 <= 5'h0;
      lsuRequestReg_instructionInformation_isStore <= 1'h0;
      lsuRequestReg_instructionInformation_maskedLoadStore <= 1'h0;
      lsuRequestReg_rs1Data <= 32'h0;
      lsuRequestReg_rs2Data <= 32'h0;
      lsuRequestReg_instructionIndex <= 3'h0;
      csrInterfaceReg_vl <= 11'h0;
      csrInterfaceReg_vStart <= 11'h0;
      csrInterfaceReg_vlmul <= 3'h0;
      csrInterfaceReg_vSew <= 2'h0;
      csrInterfaceReg_vxrm <= 2'h0;
      csrInterfaceReg_vta <= 1'h0;
      csrInterfaceReg_vma <= 1'h0;
      requestFireNext <= 1'h0;
      dataEEW <= 2'h0;
      maskReg <= 64'h0;
      needAmend <= 1'h0;
      lastMaskAmendReg <= 63'h0;
      maskGroupCounter <= 4'h0;
      maskCounterInGroup <= 2'h0;
      maskForGroup <= 64'h0;
      isLastMaskGroup <= 1'h0;
      accessData_0 <= 512'h0;
      accessData_1 <= 512'h0;
      accessData_2 <= 512'h0;
      accessData_3 <= 512'h0;
      accessData_4 <= 512'h0;
      accessData_5 <= 512'h0;
      accessData_6 <= 512'h0;
      accessData_7 <= 512'h0;
      accessPtr <= 3'h0;
      accessState_0 <= 1'h0;
      accessState_1 <= 1'h0;
      accessState_2 <= 1'h0;
      accessState_3 <= 1'h0;
      accessState_4 <= 1'h0;
      accessState_5 <= 1'h0;
      accessState_6 <= 1'h0;
      accessState_7 <= 1'h0;
      accessState_8 <= 1'h0;
      accessState_9 <= 1'h0;
      accessState_10 <= 1'h0;
      accessState_11 <= 1'h0;
      accessState_12 <= 1'h0;
      accessState_13 <= 1'h0;
      accessState_14 <= 1'h0;
      accessState_15 <= 1'h0;
      dataGroup <= 4'h0;
      dataBuffer_0 <= 512'h0;
      dataBuffer_1 <= 512'h0;
      dataBuffer_2 <= 512'h0;
      dataBuffer_3 <= 512'h0;
      dataBuffer_4 <= 512'h0;
      dataBuffer_5 <= 512'h0;
      dataBuffer_6 <= 512'h0;
      dataBuffer_7 <= 512'h0;
      bufferBaseCacheLineIndex <= 5'h0;
      cacheLineIndexInBuffer <= 3'h0;
      segmentInstructionIndexInterval <= 4'h0;
      lastWriteVrfIndexReg <= 12'h0;
      lastCacheNeedPush <= 1'h0;
      cacheLineNumberReg <= 12'h0;
      sendRequest <= 1'h0;
      writeReadyReg <= 1'h0;
      unalignedCacheLine_valid <= 1'h0;
      unalignedCacheLine_bits_data <= 512'h0;
      unalignedCacheLine_bits_index <= 5'h0;
      bufferFull <= 1'h0;
      waitForFirstDataGroup <= 1'h0;
      sendStateReg_0 <= 1'h0;
      sendStateReg_1 <= 1'h0;
      sendStateReg_2 <= 1'h0;
      sendStateReg_3 <= 1'h0;
      sendStateReg_4 <= 1'h0;
      sendStateReg_5 <= 1'h0;
      sendStateReg_6 <= 1'h0;
      sendStateReg_7 <= 1'h0;
      sendStateReg_8 <= 1'h0;
      sendStateReg_9 <= 1'h0;
      sendStateReg_10 <= 1'h0;
      sendStateReg_11 <= 1'h0;
      sendStateReg_12 <= 1'h0;
      sendStateReg_13 <= 1'h0;
      sendStateReg_14 <= 1'h0;
      sendStateReg_15 <= 1'h0;
      lastCacheRequestReg <= 1'h1;
      lastCacheLineAckReg <= 1'h1;
      idleNext <= 1'h1;
    end
    else begin
      automatic logic _GEN_10 = bufferDequeueFire | accessStateCheck & ~lastPtr;
      if (lsuRequest_valid) begin
        lsuRequestReg_instructionInformation_nf <= nfCorrection;
        lsuRequestReg_instructionInformation_mew <= ~invalidInstruction & lsuRequest_bits_instructionInformation_mew;
        lsuRequestReg_instructionInformation_mop <= invalidInstruction ? 2'h0 : lsuRequest_bits_instructionInformation_mop;
        lsuRequestReg_instructionInformation_lumop <= invalidInstruction ? 5'h0 : lsuRequest_bits_instructionInformation_lumop;
        lsuRequestReg_instructionInformation_eew <= invalidInstruction ? 2'h0 : lsuRequest_bits_instructionInformation_eew;
        lsuRequestReg_instructionInformation_vs3 <= invalidInstruction ? 5'h0 : lsuRequest_bits_instructionInformation_vs3;
        lsuRequestReg_instructionInformation_isStore <= ~invalidInstruction & lsuRequest_bits_instructionInformation_isStore;
        lsuRequestReg_instructionInformation_maskedLoadStore <= ~invalidInstruction & lsuRequest_bits_instructionInformation_maskedLoadStore;
        lsuRequestReg_rs1Data <= invalidInstruction ? 32'h0 : lsuRequest_bits_rs1Data;
        lsuRequestReg_rs2Data <= invalidInstruction ? 32'h0 : lsuRequest_bits_rs2Data;
        lsuRequestReg_instructionIndex <= lsuRequest_bits_instructionIndex;
        csrInterfaceReg_vl <= csrInterface_vl;
        csrInterfaceReg_vStart <= csrInterface_vStart;
        csrInterfaceReg_vlmul <= csrInterface_vlmul;
        csrInterfaceReg_vSew <= csrInterface_vSew;
        csrInterfaceReg_vxrm <= csrInterface_vxrm;
        csrInterfaceReg_vta <= csrInterface_vta;
        csrInterfaceReg_vma <= csrInterface_vma;
        dataEEW <= lsuRequest_bits_instructionInformation_eew;
        needAmend <= |(csrInterface_vl[5:0]);
        lastMaskAmendReg <= lastMaskAmend;
        segmentInstructionIndexInterval <= csrInterface_vlmul[2] ? 4'h1 : 4'h1 << csrInterface_vlmul[1:0];
        lastWriteVrfIndexReg <= lastWriteVrfIndex;
        lastCacheNeedPush <= lastCacheLineIndex == lastWriteVrfIndex;
        cacheLineNumberReg <= lastCacheLineIndex;
      end
      requestFireNext <= lsuRequest_valid;
      if (_maskSelect_valid_output | lsuRequest_valid) begin
        maskReg <= maskAmend;
        isLastMaskGroup <= lsuRequest_valid ? csrInterface_vl[10:6] == 5'h0 : {1'h0, _maskSelect_bits_output} == csrInterfaceReg_vl[10:6];
      end
      if (bufferDequeueFire & isLastDataGroup)
        maskGroupCounter <= nextMaskGroup;
      else if (lsuRequest_valid)
        maskGroupCounter <= 4'h0;
      if (lsuRequest_valid | bufferDequeueFire) begin
        maskCounterInGroup <= isLastDataGroup | lsuRequest_valid ? 2'h0 : nextMaskCount;
        waitForFirstDataGroup <= lsuRequest_valid;
      end
      if (bufferDequeueFire) begin
        automatic logic [7:0]    _GEN_11;
        automatic logic [4095:0] _GEN_12;
        _GEN_11 = 8'h1 << lsuRequestReg_instructionInformation_nf;
        _GEN_12 =
          (dataEEWOH[0]
             ? (_GEN_11[0] ? regroupLoadData_0_0 : 4096'h0) | (_GEN_11[1] ? regroupLoadData_0_1 : 4096'h0) | (_GEN_11[2] ? regroupLoadData_0_2 : 4096'h0) | (_GEN_11[3] ? regroupLoadData_0_3 : 4096'h0)
               | (_GEN_11[4] ? regroupLoadData_0_4 : 4096'h0) | (_GEN_11[5] ? regroupLoadData_0_5 : 4096'h0) | (_GEN_11[6] ? regroupLoadData_0_6 : 4096'h0) | (_GEN_11[7] ? regroupLoadData_0_7 : 4096'h0)
             : 4096'h0)
          | (dataEEWOH[1]
               ? (_GEN_11[0] ? regroupLoadData_1_0 : 4096'h0) | (_GEN_11[1] ? regroupLoadData_1_1 : 4096'h0) | (_GEN_11[2] ? regroupLoadData_1_2 : 4096'h0) | (_GEN_11[3] ? regroupLoadData_1_3 : 4096'h0)
                 | (_GEN_11[4] ? regroupLoadData_1_4 : 4096'h0) | (_GEN_11[5] ? regroupLoadData_1_5 : 4096'h0) | (_GEN_11[6] ? regroupLoadData_1_6 : 4096'h0) | (_GEN_11[7] ? regroupLoadData_1_7 : 4096'h0)
               : 4096'h0)
          | (dataEEWOH[2]
               ? (_GEN_11[0] ? regroupLoadData_2_0 : 4096'h0) | (_GEN_11[1] ? regroupLoadData_2_1 : 4096'h0) | (_GEN_11[2] ? regroupLoadData_2_2 : 4096'h0) | (_GEN_11[3] ? regroupLoadData_2_3 : 4096'h0)
                 | (_GEN_11[4] ? regroupLoadData_2_4 : 4096'h0) | (_GEN_11[5] ? regroupLoadData_2_5 : 4096'h0) | (_GEN_11[6] ? regroupLoadData_2_6 : 4096'h0) | (_GEN_11[7] ? regroupLoadData_2_7 : 4096'h0)
               : 4096'h0);
        maskForGroup <= maskForGroupWire;
        accessData_0 <= _GEN_12[511:0];
        accessData_1 <= _GEN_12[1023:512];
        accessData_2 <= _GEN_12[1535:1024];
        accessData_3 <= _GEN_12[2047:1536];
        accessData_4 <= _GEN_12[2559:2048];
        accessData_5 <= _GEN_12[3071:2560];
        accessData_6 <= _GEN_12[3583:3072];
        accessData_7 <= _GEN_12[4095:3584];
        dataGroup <= waitForFirstDataGroup ? 4'h0 : dataGroup + 4'h1;
        sendStateReg_0 <= initSendState_0;
        sendStateReg_1 <= initSendState_1;
        sendStateReg_2 <= initSendState_2;
        sendStateReg_3 <= initSendState_3;
        sendStateReg_4 <= initSendState_4;
        sendStateReg_5 <= initSendState_5;
        sendStateReg_6 <= initSendState_6;
        sendStateReg_7 <= initSendState_7;
        sendStateReg_8 <= initSendState_8;
        sendStateReg_9 <= initSendState_9;
        sendStateReg_10 <= initSendState_10;
        sendStateReg_11 <= initSendState_11;
        sendStateReg_12 <= initSendState_12;
        sendStateReg_13 <= initSendState_13;
        sendStateReg_14 <= initSendState_14;
        sendStateReg_15 <= initSendState_15;
      end
      if (_GEN_10)
        accessPtr <= bufferDequeueFire ? lsuRequestReg_instructionInformation_nf : accessPtr - 3'h1;
      accessState_0 <= _GEN_10 ? (bufferDequeueFire ? initSendState_0 : sendStateReg_0) : accessStateUpdate_0;
      accessState_1 <= _GEN_10 ? (bufferDequeueFire ? initSendState_1 : sendStateReg_1) : accessStateUpdate_1;
      accessState_2 <= _GEN_10 ? (bufferDequeueFire ? initSendState_2 : sendStateReg_2) : accessStateUpdate_2;
      accessState_3 <= _GEN_10 ? (bufferDequeueFire ? initSendState_3 : sendStateReg_3) : accessStateUpdate_3;
      accessState_4 <= _GEN_10 ? (bufferDequeueFire ? initSendState_4 : sendStateReg_4) : accessStateUpdate_4;
      accessState_5 <= _GEN_10 ? (bufferDequeueFire ? initSendState_5 : sendStateReg_5) : accessStateUpdate_5;
      accessState_6 <= _GEN_10 ? (bufferDequeueFire ? initSendState_6 : sendStateReg_6) : accessStateUpdate_6;
      accessState_7 <= _GEN_10 ? (bufferDequeueFire ? initSendState_7 : sendStateReg_7) : accessStateUpdate_7;
      accessState_8 <= _GEN_10 ? (bufferDequeueFire ? initSendState_8 : sendStateReg_8) : accessStateUpdate_8;
      accessState_9 <= _GEN_10 ? (bufferDequeueFire ? initSendState_9 : sendStateReg_9) : accessStateUpdate_9;
      accessState_10 <= _GEN_10 ? (bufferDequeueFire ? initSendState_10 : sendStateReg_10) : accessStateUpdate_10;
      accessState_11 <= _GEN_10 ? (bufferDequeueFire ? initSendState_11 : sendStateReg_11) : accessStateUpdate_11;
      accessState_12 <= _GEN_10 ? (bufferDequeueFire ? initSendState_12 : sendStateReg_12) : accessStateUpdate_12;
      accessState_13 <= _GEN_10 ? (bufferDequeueFire ? initSendState_13 : sendStateReg_13) : accessStateUpdate_13;
      accessState_14 <= _GEN_10 ? (bufferDequeueFire ? initSendState_14 : sendStateReg_14) : accessStateUpdate_14;
      accessState_15 <= _GEN_10 ? (bufferDequeueFire ? initSendState_15 : sendStateReg_15) : accessStateUpdate_15;
      if (bufferEnqueueSelect[0])
        dataBuffer_0 <= alignedDequeue_bits_data;
      if (bufferEnqueueSelect[1])
        dataBuffer_1 <= alignedDequeue_bits_data;
      if (bufferEnqueueSelect[2])
        dataBuffer_2 <= alignedDequeue_bits_data;
      if (bufferEnqueueSelect[3])
        dataBuffer_3 <= alignedDequeue_bits_data;
      if (bufferEnqueueSelect[4])
        dataBuffer_4 <= alignedDequeue_bits_data;
      if (bufferEnqueueSelect[5])
        dataBuffer_5 <= alignedDequeue_bits_data;
      if (bufferEnqueueSelect[6])
        dataBuffer_6 <= alignedDequeue_bits_data;
      if (bufferEnqueueSelect[7])
        dataBuffer_7 <= alignedDequeue_bits_data;
      if (_bufferTailFire_T & cacheLineIndexInBuffer == 3'h0)
        bufferBaseCacheLineIndex <= alignedDequeue_bits_index;
      if (_bufferTailFire_T | bufferDequeueFire)
        cacheLineIndexInBuffer <= bufferDequeueFire ? 3'h0 : cacheLineIndexInBuffer + 3'h1;
      if (validInstruction | _lastCacheRequest_T & lastRequest)
        sendRequest <= lsuRequest_valid & (|csrInterface_vl);
      writeReadyReg <= ~lsuRequest_valid;
      if (unalignedEnqueueFire ^ _bufferTailFire_T | lsuRequest_valid)
        unalignedCacheLine_valid <= unalignedEnqueueFire;
      if (unalignedEnqueueFire) begin
        unalignedCacheLine_bits_data <= memResponse_bits_data_0;
        unalignedCacheLine_bits_index <= nextIndex;
      end
      if (bufferTailFire | bufferDequeueFire)
        bufferFull <= ~bufferDequeueFire;
      if (lastCacheRequest | validInstruction)
        lastCacheRequestReg <= lastCacheRequest;
      if (anyLastCacheLineAck | validInstruction)
        lastCacheLineAckReg <= anyLastCacheLineAck;
      idleNext <= _status_idle_output;
    end
    invalidInstructionNext <= invalidInstruction & lsuRequest_valid;
    if (_lastCacheRequest_T | lsuRequest_valid)
      cacheLineIndex <= lsuRequest_valid ? 5'h0 : nextCacheLineIndex;
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:284];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [8:0] i = 9'h0; i < 9'h11D; i += 9'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        lsuRequestReg_instructionInformation_nf = _RANDOM[9'h0][2:0];
        lsuRequestReg_instructionInformation_mew = _RANDOM[9'h0][3];
        lsuRequestReg_instructionInformation_mop = _RANDOM[9'h0][5:4];
        lsuRequestReg_instructionInformation_lumop = _RANDOM[9'h0][10:6];
        lsuRequestReg_instructionInformation_eew = _RANDOM[9'h0][12:11];
        lsuRequestReg_instructionInformation_vs3 = _RANDOM[9'h0][17:13];
        lsuRequestReg_instructionInformation_isStore = _RANDOM[9'h0][18];
        lsuRequestReg_instructionInformation_maskedLoadStore = _RANDOM[9'h0][19];
        lsuRequestReg_rs1Data = {_RANDOM[9'h0][31:20], _RANDOM[9'h1][19:0]};
        lsuRequestReg_rs2Data = {_RANDOM[9'h1][31:20], _RANDOM[9'h2][19:0]};
        lsuRequestReg_instructionIndex = _RANDOM[9'h2][22:20];
        csrInterfaceReg_vl = {_RANDOM[9'h2][31:23], _RANDOM[9'h3][1:0]};
        csrInterfaceReg_vStart = _RANDOM[9'h3][12:2];
        csrInterfaceReg_vlmul = _RANDOM[9'h3][15:13];
        csrInterfaceReg_vSew = _RANDOM[9'h3][17:16];
        csrInterfaceReg_vxrm = _RANDOM[9'h3][19:18];
        csrInterfaceReg_vta = _RANDOM[9'h3][20];
        csrInterfaceReg_vma = _RANDOM[9'h3][21];
        requestFireNext = _RANDOM[9'h3][22];
        dataEEW = _RANDOM[9'h3][24:23];
        maskReg = {_RANDOM[9'h3][31:25], _RANDOM[9'h4], _RANDOM[9'h5][24:0]};
        needAmend = _RANDOM[9'h5][25];
        lastMaskAmendReg = {_RANDOM[9'h5][31:26], _RANDOM[9'h6], _RANDOM[9'h7][24:0]};
        maskGroupCounter = _RANDOM[9'h7][28:25];
        maskCounterInGroup = _RANDOM[9'h7][30:29];
        maskForGroup = {_RANDOM[9'h7][31], _RANDOM[9'h8], _RANDOM[9'h9][30:0]};
        isLastMaskGroup = _RANDOM[9'h9][31];
        accessData_0 =
          {_RANDOM[9'hA],
           _RANDOM[9'hB],
           _RANDOM[9'hC],
           _RANDOM[9'hD],
           _RANDOM[9'hE],
           _RANDOM[9'hF],
           _RANDOM[9'h10],
           _RANDOM[9'h11],
           _RANDOM[9'h12],
           _RANDOM[9'h13],
           _RANDOM[9'h14],
           _RANDOM[9'h15],
           _RANDOM[9'h16],
           _RANDOM[9'h17],
           _RANDOM[9'h18],
           _RANDOM[9'h19]};
        accessData_1 =
          {_RANDOM[9'h1A],
           _RANDOM[9'h1B],
           _RANDOM[9'h1C],
           _RANDOM[9'h1D],
           _RANDOM[9'h1E],
           _RANDOM[9'h1F],
           _RANDOM[9'h20],
           _RANDOM[9'h21],
           _RANDOM[9'h22],
           _RANDOM[9'h23],
           _RANDOM[9'h24],
           _RANDOM[9'h25],
           _RANDOM[9'h26],
           _RANDOM[9'h27],
           _RANDOM[9'h28],
           _RANDOM[9'h29]};
        accessData_2 =
          {_RANDOM[9'h2A],
           _RANDOM[9'h2B],
           _RANDOM[9'h2C],
           _RANDOM[9'h2D],
           _RANDOM[9'h2E],
           _RANDOM[9'h2F],
           _RANDOM[9'h30],
           _RANDOM[9'h31],
           _RANDOM[9'h32],
           _RANDOM[9'h33],
           _RANDOM[9'h34],
           _RANDOM[9'h35],
           _RANDOM[9'h36],
           _RANDOM[9'h37],
           _RANDOM[9'h38],
           _RANDOM[9'h39]};
        accessData_3 =
          {_RANDOM[9'h3A],
           _RANDOM[9'h3B],
           _RANDOM[9'h3C],
           _RANDOM[9'h3D],
           _RANDOM[9'h3E],
           _RANDOM[9'h3F],
           _RANDOM[9'h40],
           _RANDOM[9'h41],
           _RANDOM[9'h42],
           _RANDOM[9'h43],
           _RANDOM[9'h44],
           _RANDOM[9'h45],
           _RANDOM[9'h46],
           _RANDOM[9'h47],
           _RANDOM[9'h48],
           _RANDOM[9'h49]};
        accessData_4 =
          {_RANDOM[9'h4A],
           _RANDOM[9'h4B],
           _RANDOM[9'h4C],
           _RANDOM[9'h4D],
           _RANDOM[9'h4E],
           _RANDOM[9'h4F],
           _RANDOM[9'h50],
           _RANDOM[9'h51],
           _RANDOM[9'h52],
           _RANDOM[9'h53],
           _RANDOM[9'h54],
           _RANDOM[9'h55],
           _RANDOM[9'h56],
           _RANDOM[9'h57],
           _RANDOM[9'h58],
           _RANDOM[9'h59]};
        accessData_5 =
          {_RANDOM[9'h5A],
           _RANDOM[9'h5B],
           _RANDOM[9'h5C],
           _RANDOM[9'h5D],
           _RANDOM[9'h5E],
           _RANDOM[9'h5F],
           _RANDOM[9'h60],
           _RANDOM[9'h61],
           _RANDOM[9'h62],
           _RANDOM[9'h63],
           _RANDOM[9'h64],
           _RANDOM[9'h65],
           _RANDOM[9'h66],
           _RANDOM[9'h67],
           _RANDOM[9'h68],
           _RANDOM[9'h69]};
        accessData_6 =
          {_RANDOM[9'h6A],
           _RANDOM[9'h6B],
           _RANDOM[9'h6C],
           _RANDOM[9'h6D],
           _RANDOM[9'h6E],
           _RANDOM[9'h6F],
           _RANDOM[9'h70],
           _RANDOM[9'h71],
           _RANDOM[9'h72],
           _RANDOM[9'h73],
           _RANDOM[9'h74],
           _RANDOM[9'h75],
           _RANDOM[9'h76],
           _RANDOM[9'h77],
           _RANDOM[9'h78],
           _RANDOM[9'h79]};
        accessData_7 =
          {_RANDOM[9'h7A],
           _RANDOM[9'h7B],
           _RANDOM[9'h7C],
           _RANDOM[9'h7D],
           _RANDOM[9'h7E],
           _RANDOM[9'h7F],
           _RANDOM[9'h80],
           _RANDOM[9'h81],
           _RANDOM[9'h82],
           _RANDOM[9'h83],
           _RANDOM[9'h84],
           _RANDOM[9'h85],
           _RANDOM[9'h86],
           _RANDOM[9'h87],
           _RANDOM[9'h88],
           _RANDOM[9'h89]};
        accessPtr = _RANDOM[9'h8A][2:0];
        accessState_0 = _RANDOM[9'h8A][3];
        accessState_1 = _RANDOM[9'h8A][4];
        accessState_2 = _RANDOM[9'h8A][5];
        accessState_3 = _RANDOM[9'h8A][6];
        accessState_4 = _RANDOM[9'h8A][7];
        accessState_5 = _RANDOM[9'h8A][8];
        accessState_6 = _RANDOM[9'h8A][9];
        accessState_7 = _RANDOM[9'h8A][10];
        accessState_8 = _RANDOM[9'h8A][11];
        accessState_9 = _RANDOM[9'h8A][12];
        accessState_10 = _RANDOM[9'h8A][13];
        accessState_11 = _RANDOM[9'h8A][14];
        accessState_12 = _RANDOM[9'h8A][15];
        accessState_13 = _RANDOM[9'h8A][16];
        accessState_14 = _RANDOM[9'h8A][17];
        accessState_15 = _RANDOM[9'h8A][18];
        dataGroup = _RANDOM[9'h8A][22:19];
        dataBuffer_0 =
          {_RANDOM[9'h8A][31:23],
           _RANDOM[9'h8B],
           _RANDOM[9'h8C],
           _RANDOM[9'h8D],
           _RANDOM[9'h8E],
           _RANDOM[9'h8F],
           _RANDOM[9'h90],
           _RANDOM[9'h91],
           _RANDOM[9'h92],
           _RANDOM[9'h93],
           _RANDOM[9'h94],
           _RANDOM[9'h95],
           _RANDOM[9'h96],
           _RANDOM[9'h97],
           _RANDOM[9'h98],
           _RANDOM[9'h99],
           _RANDOM[9'h9A][22:0]};
        dataBuffer_1 =
          {_RANDOM[9'h9A][31:23],
           _RANDOM[9'h9B],
           _RANDOM[9'h9C],
           _RANDOM[9'h9D],
           _RANDOM[9'h9E],
           _RANDOM[9'h9F],
           _RANDOM[9'hA0],
           _RANDOM[9'hA1],
           _RANDOM[9'hA2],
           _RANDOM[9'hA3],
           _RANDOM[9'hA4],
           _RANDOM[9'hA5],
           _RANDOM[9'hA6],
           _RANDOM[9'hA7],
           _RANDOM[9'hA8],
           _RANDOM[9'hA9],
           _RANDOM[9'hAA][22:0]};
        dataBuffer_2 =
          {_RANDOM[9'hAA][31:23],
           _RANDOM[9'hAB],
           _RANDOM[9'hAC],
           _RANDOM[9'hAD],
           _RANDOM[9'hAE],
           _RANDOM[9'hAF],
           _RANDOM[9'hB0],
           _RANDOM[9'hB1],
           _RANDOM[9'hB2],
           _RANDOM[9'hB3],
           _RANDOM[9'hB4],
           _RANDOM[9'hB5],
           _RANDOM[9'hB6],
           _RANDOM[9'hB7],
           _RANDOM[9'hB8],
           _RANDOM[9'hB9],
           _RANDOM[9'hBA][22:0]};
        dataBuffer_3 =
          {_RANDOM[9'hBA][31:23],
           _RANDOM[9'hBB],
           _RANDOM[9'hBC],
           _RANDOM[9'hBD],
           _RANDOM[9'hBE],
           _RANDOM[9'hBF],
           _RANDOM[9'hC0],
           _RANDOM[9'hC1],
           _RANDOM[9'hC2],
           _RANDOM[9'hC3],
           _RANDOM[9'hC4],
           _RANDOM[9'hC5],
           _RANDOM[9'hC6],
           _RANDOM[9'hC7],
           _RANDOM[9'hC8],
           _RANDOM[9'hC9],
           _RANDOM[9'hCA][22:0]};
        dataBuffer_4 =
          {_RANDOM[9'hCA][31:23],
           _RANDOM[9'hCB],
           _RANDOM[9'hCC],
           _RANDOM[9'hCD],
           _RANDOM[9'hCE],
           _RANDOM[9'hCF],
           _RANDOM[9'hD0],
           _RANDOM[9'hD1],
           _RANDOM[9'hD2],
           _RANDOM[9'hD3],
           _RANDOM[9'hD4],
           _RANDOM[9'hD5],
           _RANDOM[9'hD6],
           _RANDOM[9'hD7],
           _RANDOM[9'hD8],
           _RANDOM[9'hD9],
           _RANDOM[9'hDA][22:0]};
        dataBuffer_5 =
          {_RANDOM[9'hDA][31:23],
           _RANDOM[9'hDB],
           _RANDOM[9'hDC],
           _RANDOM[9'hDD],
           _RANDOM[9'hDE],
           _RANDOM[9'hDF],
           _RANDOM[9'hE0],
           _RANDOM[9'hE1],
           _RANDOM[9'hE2],
           _RANDOM[9'hE3],
           _RANDOM[9'hE4],
           _RANDOM[9'hE5],
           _RANDOM[9'hE6],
           _RANDOM[9'hE7],
           _RANDOM[9'hE8],
           _RANDOM[9'hE9],
           _RANDOM[9'hEA][22:0]};
        dataBuffer_6 =
          {_RANDOM[9'hEA][31:23],
           _RANDOM[9'hEB],
           _RANDOM[9'hEC],
           _RANDOM[9'hED],
           _RANDOM[9'hEE],
           _RANDOM[9'hEF],
           _RANDOM[9'hF0],
           _RANDOM[9'hF1],
           _RANDOM[9'hF2],
           _RANDOM[9'hF3],
           _RANDOM[9'hF4],
           _RANDOM[9'hF5],
           _RANDOM[9'hF6],
           _RANDOM[9'hF7],
           _RANDOM[9'hF8],
           _RANDOM[9'hF9],
           _RANDOM[9'hFA][22:0]};
        dataBuffer_7 =
          {_RANDOM[9'hFA][31:23],
           _RANDOM[9'hFB],
           _RANDOM[9'hFC],
           _RANDOM[9'hFD],
           _RANDOM[9'hFE],
           _RANDOM[9'hFF],
           _RANDOM[9'h100],
           _RANDOM[9'h101],
           _RANDOM[9'h102],
           _RANDOM[9'h103],
           _RANDOM[9'h104],
           _RANDOM[9'h105],
           _RANDOM[9'h106],
           _RANDOM[9'h107],
           _RANDOM[9'h108],
           _RANDOM[9'h109],
           _RANDOM[9'h10A][22:0]};
        bufferBaseCacheLineIndex = _RANDOM[9'h10A][27:23];
        cacheLineIndexInBuffer = _RANDOM[9'h10A][30:28];
        invalidInstructionNext = _RANDOM[9'h10A][31];
        segmentInstructionIndexInterval = _RANDOM[9'h10B][3:0];
        lastWriteVrfIndexReg = _RANDOM[9'h10B][15:4];
        lastCacheNeedPush = _RANDOM[9'h10B][16];
        cacheLineNumberReg = _RANDOM[9'h10B][28:17];
        cacheLineIndex = {_RANDOM[9'h10B][31:29], _RANDOM[9'h10C][1:0]};
        sendRequest = _RANDOM[9'h10C][2];
        writeReadyReg = _RANDOM[9'h10C][3];
        unalignedCacheLine_valid = _RANDOM[9'h10C][4];
        unalignedCacheLine_bits_data =
          {_RANDOM[9'h10C][31:5],
           _RANDOM[9'h10D],
           _RANDOM[9'h10E],
           _RANDOM[9'h10F],
           _RANDOM[9'h110],
           _RANDOM[9'h111],
           _RANDOM[9'h112],
           _RANDOM[9'h113],
           _RANDOM[9'h114],
           _RANDOM[9'h115],
           _RANDOM[9'h116],
           _RANDOM[9'h117],
           _RANDOM[9'h118],
           _RANDOM[9'h119],
           _RANDOM[9'h11A],
           _RANDOM[9'h11B],
           _RANDOM[9'h11C][4:0]};
        unalignedCacheLine_bits_index = _RANDOM[9'h11C][9:5];
        bufferFull = _RANDOM[9'h11C][10];
        waitForFirstDataGroup = _RANDOM[9'h11C][11];
        sendStateReg_0 = _RANDOM[9'h11C][12];
        sendStateReg_1 = _RANDOM[9'h11C][13];
        sendStateReg_2 = _RANDOM[9'h11C][14];
        sendStateReg_3 = _RANDOM[9'h11C][15];
        sendStateReg_4 = _RANDOM[9'h11C][16];
        sendStateReg_5 = _RANDOM[9'h11C][17];
        sendStateReg_6 = _RANDOM[9'h11C][18];
        sendStateReg_7 = _RANDOM[9'h11C][19];
        sendStateReg_8 = _RANDOM[9'h11C][20];
        sendStateReg_9 = _RANDOM[9'h11C][21];
        sendStateReg_10 = _RANDOM[9'h11C][22];
        sendStateReg_11 = _RANDOM[9'h11C][23];
        sendStateReg_12 = _RANDOM[9'h11C][24];
        sendStateReg_13 = _RANDOM[9'h11C][25];
        sendStateReg_14 = _RANDOM[9'h11C][26];
        sendStateReg_15 = _RANDOM[9'h11C][27];
        lastCacheRequestReg = _RANDOM[9'h11C][28];
        lastCacheLineAckReg = _RANDOM[9'h11C][29];
        idleNext = _RANDOM[9'h11C][30];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  assign maskSelect_valid = _maskSelect_valid_output;
  assign maskSelect_bits = _maskSelect_bits_output;
  assign memRequest_valid = memRequest_valid_0;
  assign memRequest_bits_src = memRequest_bits_src_0;
  assign memRequest_bits_address = memRequest_bits_address_0;
  assign memResponse_ready = memResponse_ready_0;
  assign status_idle = _status_idle_output;
  assign status_last = ~idleNext & _status_idle_output | invalidInstructionNext;
  assign status_instructionIndex = lsuRequestReg_instructionIndex;
  assign status_changeMaskGroup = _maskSelect_valid_output & ~lsuRequest_valid;
  assign status_startAddress = requestAddress;
  assign status_endAddress = {lsuRequestReg_rs1Data[31:6] + {14'h0, cacheLineNumberReg}, 6'h0};
  assign vrfWritePort_0_valid = vrfWritePort_0_valid_0;
  assign vrfWritePort_0_bits_vd = vrfWritePort_0_bits_vd_0;
  assign vrfWritePort_0_bits_offset = vrfWritePort_0_bits_offset_0;
  assign vrfWritePort_0_bits_mask = vrfWritePort_0_bits_mask_0;
  assign vrfWritePort_0_bits_data = vrfWritePort_0_bits_data_0;
  assign vrfWritePort_0_bits_instructionIndex = vrfWritePort_0_bits_instructionIndex_0;
  assign vrfWritePort_1_valid = vrfWritePort_1_valid_0;
  assign vrfWritePort_1_bits_vd = vrfWritePort_1_bits_vd_0;
  assign vrfWritePort_1_bits_offset = vrfWritePort_1_bits_offset_0;
  assign vrfWritePort_1_bits_mask = vrfWritePort_1_bits_mask_0;
  assign vrfWritePort_1_bits_data = vrfWritePort_1_bits_data_0;
  assign vrfWritePort_1_bits_instructionIndex = vrfWritePort_1_bits_instructionIndex_0;
  assign vrfWritePort_2_valid = vrfWritePort_2_valid_0;
  assign vrfWritePort_2_bits_vd = vrfWritePort_2_bits_vd_0;
  assign vrfWritePort_2_bits_offset = vrfWritePort_2_bits_offset_0;
  assign vrfWritePort_2_bits_mask = vrfWritePort_2_bits_mask_0;
  assign vrfWritePort_2_bits_data = vrfWritePort_2_bits_data_0;
  assign vrfWritePort_2_bits_instructionIndex = vrfWritePort_2_bits_instructionIndex_0;
  assign vrfWritePort_3_valid = vrfWritePort_3_valid_0;
  assign vrfWritePort_3_bits_vd = vrfWritePort_3_bits_vd_0;
  assign vrfWritePort_3_bits_offset = vrfWritePort_3_bits_offset_0;
  assign vrfWritePort_3_bits_mask = vrfWritePort_3_bits_mask_0;
  assign vrfWritePort_3_bits_data = vrfWritePort_3_bits_data_0;
  assign vrfWritePort_3_bits_instructionIndex = vrfWritePort_3_bits_instructionIndex_0;
  assign vrfWritePort_4_valid = vrfWritePort_4_valid_0;
  assign vrfWritePort_4_bits_vd = vrfWritePort_4_bits_vd_0;
  assign vrfWritePort_4_bits_offset = vrfWritePort_4_bits_offset_0;
  assign vrfWritePort_4_bits_mask = vrfWritePort_4_bits_mask_0;
  assign vrfWritePort_4_bits_data = vrfWritePort_4_bits_data_0;
  assign vrfWritePort_4_bits_instructionIndex = vrfWritePort_4_bits_instructionIndex_0;
  assign vrfWritePort_5_valid = vrfWritePort_5_valid_0;
  assign vrfWritePort_5_bits_vd = vrfWritePort_5_bits_vd_0;
  assign vrfWritePort_5_bits_offset = vrfWritePort_5_bits_offset_0;
  assign vrfWritePort_5_bits_mask = vrfWritePort_5_bits_mask_0;
  assign vrfWritePort_5_bits_data = vrfWritePort_5_bits_data_0;
  assign vrfWritePort_5_bits_instructionIndex = vrfWritePort_5_bits_instructionIndex_0;
  assign vrfWritePort_6_valid = vrfWritePort_6_valid_0;
  assign vrfWritePort_6_bits_vd = vrfWritePort_6_bits_vd_0;
  assign vrfWritePort_6_bits_offset = vrfWritePort_6_bits_offset_0;
  assign vrfWritePort_6_bits_mask = vrfWritePort_6_bits_mask_0;
  assign vrfWritePort_6_bits_data = vrfWritePort_6_bits_data_0;
  assign vrfWritePort_6_bits_instructionIndex = vrfWritePort_6_bits_instructionIndex_0;
  assign vrfWritePort_7_valid = vrfWritePort_7_valid_0;
  assign vrfWritePort_7_bits_vd = vrfWritePort_7_bits_vd_0;
  assign vrfWritePort_7_bits_offset = vrfWritePort_7_bits_offset_0;
  assign vrfWritePort_7_bits_mask = vrfWritePort_7_bits_mask_0;
  assign vrfWritePort_7_bits_data = vrfWritePort_7_bits_data_0;
  assign vrfWritePort_7_bits_instructionIndex = vrfWritePort_7_bits_instructionIndex_0;
  assign vrfWritePort_8_valid = vrfWritePort_8_valid_0;
  assign vrfWritePort_8_bits_vd = vrfWritePort_8_bits_vd_0;
  assign vrfWritePort_8_bits_offset = vrfWritePort_8_bits_offset_0;
  assign vrfWritePort_8_bits_mask = vrfWritePort_8_bits_mask_0;
  assign vrfWritePort_8_bits_data = vrfWritePort_8_bits_data_0;
  assign vrfWritePort_8_bits_instructionIndex = vrfWritePort_8_bits_instructionIndex_0;
  assign vrfWritePort_9_valid = vrfWritePort_9_valid_0;
  assign vrfWritePort_9_bits_vd = vrfWritePort_9_bits_vd_0;
  assign vrfWritePort_9_bits_offset = vrfWritePort_9_bits_offset_0;
  assign vrfWritePort_9_bits_mask = vrfWritePort_9_bits_mask_0;
  assign vrfWritePort_9_bits_data = vrfWritePort_9_bits_data_0;
  assign vrfWritePort_9_bits_instructionIndex = vrfWritePort_9_bits_instructionIndex_0;
  assign vrfWritePort_10_valid = vrfWritePort_10_valid_0;
  assign vrfWritePort_10_bits_vd = vrfWritePort_10_bits_vd_0;
  assign vrfWritePort_10_bits_offset = vrfWritePort_10_bits_offset_0;
  assign vrfWritePort_10_bits_mask = vrfWritePort_10_bits_mask_0;
  assign vrfWritePort_10_bits_data = vrfWritePort_10_bits_data_0;
  assign vrfWritePort_10_bits_instructionIndex = vrfWritePort_10_bits_instructionIndex_0;
  assign vrfWritePort_11_valid = vrfWritePort_11_valid_0;
  assign vrfWritePort_11_bits_vd = vrfWritePort_11_bits_vd_0;
  assign vrfWritePort_11_bits_offset = vrfWritePort_11_bits_offset_0;
  assign vrfWritePort_11_bits_mask = vrfWritePort_11_bits_mask_0;
  assign vrfWritePort_11_bits_data = vrfWritePort_11_bits_data_0;
  assign vrfWritePort_11_bits_instructionIndex = vrfWritePort_11_bits_instructionIndex_0;
  assign vrfWritePort_12_valid = vrfWritePort_12_valid_0;
  assign vrfWritePort_12_bits_vd = vrfWritePort_12_bits_vd_0;
  assign vrfWritePort_12_bits_offset = vrfWritePort_12_bits_offset_0;
  assign vrfWritePort_12_bits_mask = vrfWritePort_12_bits_mask_0;
  assign vrfWritePort_12_bits_data = vrfWritePort_12_bits_data_0;
  assign vrfWritePort_12_bits_instructionIndex = vrfWritePort_12_bits_instructionIndex_0;
  assign vrfWritePort_13_valid = vrfWritePort_13_valid_0;
  assign vrfWritePort_13_bits_vd = vrfWritePort_13_bits_vd_0;
  assign vrfWritePort_13_bits_offset = vrfWritePort_13_bits_offset_0;
  assign vrfWritePort_13_bits_mask = vrfWritePort_13_bits_mask_0;
  assign vrfWritePort_13_bits_data = vrfWritePort_13_bits_data_0;
  assign vrfWritePort_13_bits_instructionIndex = vrfWritePort_13_bits_instructionIndex_0;
  assign vrfWritePort_14_valid = vrfWritePort_14_valid_0;
  assign vrfWritePort_14_bits_vd = vrfWritePort_14_bits_vd_0;
  assign vrfWritePort_14_bits_offset = vrfWritePort_14_bits_offset_0;
  assign vrfWritePort_14_bits_mask = vrfWritePort_14_bits_mask_0;
  assign vrfWritePort_14_bits_data = vrfWritePort_14_bits_data_0;
  assign vrfWritePort_14_bits_instructionIndex = vrfWritePort_14_bits_instructionIndex_0;
  assign vrfWritePort_15_valid = vrfWritePort_15_valid_0;
  assign vrfWritePort_15_bits_vd = vrfWritePort_15_bits_vd_0;
  assign vrfWritePort_15_bits_offset = vrfWritePort_15_bits_offset_0;
  assign vrfWritePort_15_bits_mask = vrfWritePort_15_bits_mask_0;
  assign vrfWritePort_15_bits_data = vrfWritePort_15_bits_data_0;
  assign vrfWritePort_15_bits_instructionIndex = vrfWritePort_15_bits_instructionIndex_0;
endmodule

