
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module StoreUnit(
  input          clock,
                 reset,
                 lsuRequest_valid,
  input  [2:0]   lsuRequest_bits_instructionInformation_nf,
  input          lsuRequest_bits_instructionInformation_mew,
  input  [1:0]   lsuRequest_bits_instructionInformation_mop,
  input  [4:0]   lsuRequest_bits_instructionInformation_lumop,
  input  [1:0]   lsuRequest_bits_instructionInformation_eew,
  input  [4:0]   lsuRequest_bits_instructionInformation_vs3,
  input          lsuRequest_bits_instructionInformation_isStore,
                 lsuRequest_bits_instructionInformation_maskedLoadStore,
  input  [31:0]  lsuRequest_bits_rs1Data,
                 lsuRequest_bits_rs2Data,
  input  [2:0]   lsuRequest_bits_instructionIndex,
  input  [12:0]  csrInterface_vl,
                 csrInterface_vStart,
  input  [2:0]   csrInterface_vlmul,
  input  [1:0]   csrInterface_vSew,
                 csrInterface_vxrm,
  input          csrInterface_vta,
                 csrInterface_vma,
  input  [15:0]  maskInput,
  output         maskSelect_valid,
  output [7:0]   maskSelect_bits,
  input          memRequest_ready,
  output         memRequest_valid,
  output [127:0] memRequest_bits_data,
  output [15:0]  memRequest_bits_mask,
  output [8:0]   memRequest_bits_index,
  output [31:0]  memRequest_bits_address,
  output         status_idle,
                 status_last,
  output [2:0]   status_instructionIndex,
  output         status_changeMaskGroup,
  output [31:0]  status_startAddress,
                 status_endAddress,
  input          vrfReadDataPorts_0_ready,
  output         vrfReadDataPorts_0_valid,
  output [4:0]   vrfReadDataPorts_0_bits_vs,
                 vrfReadDataPorts_0_bits_offset,
  output [2:0]   vrfReadDataPorts_0_bits_instructionIndex,
  input          vrfReadDataPorts_1_ready,
  output         vrfReadDataPorts_1_valid,
  output [4:0]   vrfReadDataPorts_1_bits_vs,
                 vrfReadDataPorts_1_bits_offset,
  output [2:0]   vrfReadDataPorts_1_bits_instructionIndex,
  input          vrfReadDataPorts_2_ready,
  output         vrfReadDataPorts_2_valid,
  output [4:0]   vrfReadDataPorts_2_bits_vs,
                 vrfReadDataPorts_2_bits_offset,
  output [2:0]   vrfReadDataPorts_2_bits_instructionIndex,
  input          vrfReadDataPorts_3_ready,
  output         vrfReadDataPorts_3_valid,
  output [4:0]   vrfReadDataPorts_3_bits_vs,
                 vrfReadDataPorts_3_bits_offset,
  output [2:0]   vrfReadDataPorts_3_bits_instructionIndex,
  input          vrfReadResults_0_valid,
  input  [31:0]  vrfReadResults_0_bits,
  input          vrfReadResults_1_valid,
  input  [31:0]  vrfReadResults_1_bits,
  input          vrfReadResults_2_valid,
  input  [31:0]  vrfReadResults_2_bits,
  input          vrfReadResults_3_valid,
  input  [31:0]  vrfReadResults_3_bits,
  input          storeResponse
);

  wire             _addressQueue_fifo_empty;
  wire             _addressQueue_fifo_full;
  wire             _addressQueue_fifo_error;
  wire             _vrfReadQueueVec_fifo_3_empty;
  wire             _vrfReadQueueVec_fifo_3_full;
  wire             _vrfReadQueueVec_fifo_3_error;
  wire [31:0]      _vrfReadQueueVec_fifo_3_data_out;
  wire             _vrfReadQueueVec_fifo_2_empty;
  wire             _vrfReadQueueVec_fifo_2_full;
  wire             _vrfReadQueueVec_fifo_2_error;
  wire [31:0]      _vrfReadQueueVec_fifo_2_data_out;
  wire             _vrfReadQueueVec_fifo_1_empty;
  wire             _vrfReadQueueVec_fifo_1_full;
  wire             _vrfReadQueueVec_fifo_1_error;
  wire [31:0]      _vrfReadQueueVec_fifo_1_data_out;
  wire             _vrfReadQueueVec_fifo_empty;
  wire             _vrfReadQueueVec_fifo_full;
  wire             _vrfReadQueueVec_fifo_error;
  wire [31:0]      _vrfReadQueueVec_fifo_data_out;
  wire             addressQueue_almostFull;
  wire             addressQueue_almostEmpty;
  wire             vrfReadQueueVec_3_almostFull;
  wire             vrfReadQueueVec_3_almostEmpty;
  wire             vrfReadQueueVec_2_almostFull;
  wire             vrfReadQueueVec_2_almostEmpty;
  wire             vrfReadQueueVec_1_almostFull;
  wire             vrfReadQueueVec_1_almostEmpty;
  wire             vrfReadQueueVec_0_almostFull;
  wire             vrfReadQueueVec_0_almostEmpty;
  wire             memRequest_ready_0 = memRequest_ready;
  wire             vrfReadDataPorts_0_ready_0 = vrfReadDataPorts_0_ready;
  wire             vrfReadDataPorts_1_ready_0 = vrfReadDataPorts_1_ready;
  wire             vrfReadDataPorts_2_ready_0 = vrfReadDataPorts_2_ready;
  wire             vrfReadDataPorts_3_ready_0 = vrfReadDataPorts_3_ready;
  wire             vrfReadQueueVec_0_enq_valid = vrfReadResults_0_valid;
  wire [31:0]      vrfReadQueueVec_0_enq_bits = vrfReadResults_0_bits;
  wire             vrfReadQueueVec_1_enq_valid = vrfReadResults_1_valid;
  wire [31:0]      vrfReadQueueVec_1_enq_bits = vrfReadResults_1_bits;
  wire             vrfReadQueueVec_2_enq_valid = vrfReadResults_2_valid;
  wire [31:0]      vrfReadQueueVec_2_enq_bits = vrfReadResults_2_bits;
  wire             vrfReadQueueVec_3_enq_valid = vrfReadResults_3_valid;
  wire [31:0]      vrfReadQueueVec_3_enq_bits = vrfReadResults_3_bits;
  wire             addressQueue_deq_ready = storeResponse;
  wire [1:0]       accessStateCheck_lo = 2'h0;
  wire [1:0]       accessStateCheck_hi = 2'h0;
  wire             accessStateCheck = 1'h1;
  wire             accessStateUpdate_0 = 1'h0;
  wire             accessStateUpdate_1 = 1'h0;
  wire             accessStateUpdate_2 = 1'h0;
  wire             accessStateUpdate_3 = 1'h0;
  wire [511:0]     hi = 512'h0;
  wire [511:0]     hi_1 = 512'h0;
  wire [511:0]     hi_2 = 512'h0;
  wire [511:0]     hi_3 = 512'h0;
  wire [511:0]     hi_8 = 512'h0;
  wire [511:0]     hi_9 = 512'h0;
  wire [511:0]     hi_10 = 512'h0;
  wire [511:0]     hi_11 = 512'h0;
  wire [511:0]     hi_16 = 512'h0;
  wire [511:0]     hi_17 = 512'h0;
  wire [511:0]     hi_18 = 512'h0;
  wire [511:0]     hi_19 = 512'h0;
  wire [255:0]     lo_hi = 256'h0;
  wire [255:0]     hi_lo = 256'h0;
  wire [255:0]     hi_hi = 256'h0;
  wire [255:0]     lo_hi_1 = 256'h0;
  wire [255:0]     hi_lo_1 = 256'h0;
  wire [255:0]     hi_hi_1 = 256'h0;
  wire [255:0]     hi_lo_2 = 256'h0;
  wire [255:0]     hi_hi_2 = 256'h0;
  wire [255:0]     hi_lo_3 = 256'h0;
  wire [255:0]     hi_hi_3 = 256'h0;
  wire [255:0]     hi_hi_4 = 256'h0;
  wire [255:0]     hi_hi_5 = 256'h0;
  wire [255:0]     lo_hi_8 = 256'h0;
  wire [255:0]     hi_lo_8 = 256'h0;
  wire [255:0]     hi_hi_8 = 256'h0;
  wire [255:0]     lo_hi_9 = 256'h0;
  wire [255:0]     hi_lo_9 = 256'h0;
  wire [255:0]     hi_hi_9 = 256'h0;
  wire [255:0]     hi_lo_10 = 256'h0;
  wire [255:0]     hi_hi_10 = 256'h0;
  wire [255:0]     hi_lo_11 = 256'h0;
  wire [255:0]     hi_hi_11 = 256'h0;
  wire [255:0]     hi_hi_12 = 256'h0;
  wire [255:0]     hi_hi_13 = 256'h0;
  wire [255:0]     lo_hi_16 = 256'h0;
  wire [255:0]     hi_lo_16 = 256'h0;
  wire [255:0]     hi_hi_16 = 256'h0;
  wire [255:0]     lo_hi_17 = 256'h0;
  wire [255:0]     hi_lo_17 = 256'h0;
  wire [255:0]     hi_hi_17 = 256'h0;
  wire [255:0]     hi_lo_18 = 256'h0;
  wire [255:0]     hi_hi_18 = 256'h0;
  wire [255:0]     hi_lo_19 = 256'h0;
  wire [255:0]     hi_hi_19 = 256'h0;
  wire [255:0]     hi_hi_20 = 256'h0;
  wire [255:0]     hi_hi_21 = 256'h0;
  wire [127:0]     res_1 = 128'h0;
  wire [127:0]     res_2 = 128'h0;
  wire [127:0]     res_3 = 128'h0;
  wire [127:0]     res_4 = 128'h0;
  wire [127:0]     res_5 = 128'h0;
  wire [127:0]     res_6 = 128'h0;
  wire [127:0]     res_7 = 128'h0;
  wire [127:0]     res_10 = 128'h0;
  wire [127:0]     res_11 = 128'h0;
  wire [127:0]     res_12 = 128'h0;
  wire [127:0]     res_13 = 128'h0;
  wire [127:0]     res_14 = 128'h0;
  wire [127:0]     res_15 = 128'h0;
  wire [127:0]     res_19 = 128'h0;
  wire [127:0]     res_20 = 128'h0;
  wire [127:0]     res_21 = 128'h0;
  wire [127:0]     res_22 = 128'h0;
  wire [127:0]     res_23 = 128'h0;
  wire [127:0]     res_28 = 128'h0;
  wire [127:0]     res_29 = 128'h0;
  wire [127:0]     res_30 = 128'h0;
  wire [127:0]     res_31 = 128'h0;
  wire [127:0]     res_37 = 128'h0;
  wire [127:0]     res_38 = 128'h0;
  wire [127:0]     res_39 = 128'h0;
  wire [127:0]     res_46 = 128'h0;
  wire [127:0]     res_47 = 128'h0;
  wire [127:0]     res_55 = 128'h0;
  wire [127:0]     res_65 = 128'h0;
  wire [127:0]     res_66 = 128'h0;
  wire [127:0]     res_67 = 128'h0;
  wire [127:0]     res_68 = 128'h0;
  wire [127:0]     res_69 = 128'h0;
  wire [127:0]     res_70 = 128'h0;
  wire [127:0]     res_71 = 128'h0;
  wire [127:0]     res_74 = 128'h0;
  wire [127:0]     res_75 = 128'h0;
  wire [127:0]     res_76 = 128'h0;
  wire [127:0]     res_77 = 128'h0;
  wire [127:0]     res_78 = 128'h0;
  wire [127:0]     res_79 = 128'h0;
  wire [127:0]     res_83 = 128'h0;
  wire [127:0]     res_84 = 128'h0;
  wire [127:0]     res_85 = 128'h0;
  wire [127:0]     res_86 = 128'h0;
  wire [127:0]     res_87 = 128'h0;
  wire [127:0]     res_92 = 128'h0;
  wire [127:0]     res_93 = 128'h0;
  wire [127:0]     res_94 = 128'h0;
  wire [127:0]     res_95 = 128'h0;
  wire [127:0]     res_101 = 128'h0;
  wire [127:0]     res_102 = 128'h0;
  wire [127:0]     res_103 = 128'h0;
  wire [127:0]     res_110 = 128'h0;
  wire [127:0]     res_111 = 128'h0;
  wire [127:0]     res_119 = 128'h0;
  wire [127:0]     res_129 = 128'h0;
  wire [127:0]     res_130 = 128'h0;
  wire [127:0]     res_131 = 128'h0;
  wire [127:0]     res_132 = 128'h0;
  wire [127:0]     res_133 = 128'h0;
  wire [127:0]     res_134 = 128'h0;
  wire [127:0]     res_135 = 128'h0;
  wire [127:0]     res_138 = 128'h0;
  wire [127:0]     res_139 = 128'h0;
  wire [127:0]     res_140 = 128'h0;
  wire [127:0]     res_141 = 128'h0;
  wire [127:0]     res_142 = 128'h0;
  wire [127:0]     res_143 = 128'h0;
  wire [127:0]     res_147 = 128'h0;
  wire [127:0]     res_148 = 128'h0;
  wire [127:0]     res_149 = 128'h0;
  wire [127:0]     res_150 = 128'h0;
  wire [127:0]     res_151 = 128'h0;
  wire [127:0]     res_156 = 128'h0;
  wire [127:0]     res_157 = 128'h0;
  wire [127:0]     res_158 = 128'h0;
  wire [127:0]     res_159 = 128'h0;
  wire [127:0]     res_165 = 128'h0;
  wire [127:0]     res_166 = 128'h0;
  wire [127:0]     res_167 = 128'h0;
  wire [127:0]     res_174 = 128'h0;
  wire [127:0]     res_175 = 128'h0;
  wire [127:0]     res_183 = 128'h0;
  wire [1:0]       vrfReadDataPorts_0_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_1_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_2_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_3_bits_readSource = 2'h2;
  wire [31:0]      alignedDequeueAddress;
  reg  [2:0]       lsuRequestReg_instructionInformation_nf;
  reg              lsuRequestReg_instructionInformation_mew;
  reg  [1:0]       lsuRequestReg_instructionInformation_mop;
  reg  [4:0]       lsuRequestReg_instructionInformation_lumop;
  reg  [1:0]       lsuRequestReg_instructionInformation_eew;
  reg  [4:0]       lsuRequestReg_instructionInformation_vs3;
  reg              lsuRequestReg_instructionInformation_isStore;
  reg              lsuRequestReg_instructionInformation_maskedLoadStore;
  reg  [31:0]      lsuRequestReg_rs1Data;
  reg  [31:0]      lsuRequestReg_rs2Data;
  reg  [2:0]       lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_0_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_1_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_2_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_3_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  reg  [12:0]      csrInterfaceReg_vl;
  reg  [12:0]      csrInterfaceReg_vStart;
  reg  [2:0]       csrInterfaceReg_vlmul;
  reg  [1:0]       csrInterfaceReg_vSew;
  reg  [1:0]       csrInterfaceReg_vxrm;
  reg              csrInterfaceReg_vta;
  reg              csrInterfaceReg_vma;
  reg              requestFireNext;
  reg  [1:0]       dataEEW;
  wire [3:0]       _dataEEWOH_T = 4'h1 << dataEEW;
  wire [2:0]       dataEEWOH = _dataEEWOH_T[2:0];
  wire             isMaskType = lsuRequest_valid ? lsuRequest_bits_instructionInformation_maskedLoadStore : lsuRequestReg_instructionInformation_maskedLoadStore;
  wire [15:0]      maskAmend = isMaskType ? maskInput : 16'hFFFF;
  reg  [15:0]      maskReg;
  wire [15:0]      _lastMaskAmend_T_1 = 16'h1 << csrInterface_vl[3:0];
  wire [13:0]      _GEN = _lastMaskAmend_T_1[14:1] | _lastMaskAmend_T_1[15:2];
  wire [12:0]      _GEN_0 = _GEN[12:0] | {_lastMaskAmend_T_1[15], _GEN[13:2]};
  wire [10:0]      _GEN_1 = _GEN_0[10:0] | {_lastMaskAmend_T_1[15], _GEN[13], _GEN_0[12:4]};
  wire [14:0]      lastMaskAmend = {_lastMaskAmend_T_1[15], _GEN[13], _GEN_0[12:11], _GEN_1[10:7], _GEN_1[6:0] | {_lastMaskAmend_T_1[15], _GEN[13], _GEN_0[12:11], _GEN_1[10:8]}};
  reg              needAmend;
  reg  [14:0]      lastMaskAmendReg;
  wire [1:0]       countEndForGroup = {1'h0, dataEEWOH[1]} | {2{dataEEWOH[2]}};
  reg  [7:0]       maskGroupCounter;
  wire [7:0]       nextMaskGroup = maskGroupCounter + 8'h1;
  reg  [1:0]       maskCounterInGroup;
  wire [1:0]       nextMaskCount = maskCounterInGroup + 2'h1;
  wire             isLastDataGroup = maskCounterInGroup == countEndForGroup;
  wire [7:0]       _maskSelect_bits_output = lsuRequest_valid ? 8'h0 : nextMaskGroup;
  reg              isLastMaskGroup;
  wire [15:0]      maskWire = maskReg & (needAmend & isLastMaskGroup ? {1'h0, lastMaskAmendReg} : 16'hFFFF);
  wire [3:0]       maskForGroupWire_lo_lo_lo = {{2{maskWire[1]}}, {2{maskWire[0]}}};
  wire [3:0]       maskForGroupWire_lo_lo_hi = {{2{maskWire[3]}}, {2{maskWire[2]}}};
  wire [7:0]       maskForGroupWire_lo_lo = {maskForGroupWire_lo_lo_hi, maskForGroupWire_lo_lo_lo};
  wire [3:0]       maskForGroupWire_lo_hi_lo = {{2{maskWire[5]}}, {2{maskWire[4]}}};
  wire [3:0]       maskForGroupWire_lo_hi_hi = {{2{maskWire[7]}}, {2{maskWire[6]}}};
  wire [7:0]       maskForGroupWire_lo_hi = {maskForGroupWire_lo_hi_hi, maskForGroupWire_lo_hi_lo};
  wire [15:0]      maskForGroupWire_lo = {maskForGroupWire_lo_hi, maskForGroupWire_lo_lo};
  wire [3:0]       maskForGroupWire_hi_lo_lo = {{2{maskWire[9]}}, {2{maskWire[8]}}};
  wire [3:0]       maskForGroupWire_hi_lo_hi = {{2{maskWire[11]}}, {2{maskWire[10]}}};
  wire [7:0]       maskForGroupWire_hi_lo = {maskForGroupWire_hi_lo_hi, maskForGroupWire_hi_lo_lo};
  wire [3:0]       maskForGroupWire_hi_hi_lo = {{2{maskWire[13]}}, {2{maskWire[12]}}};
  wire [3:0]       maskForGroupWire_hi_hi_hi = {{2{maskWire[15]}}, {2{maskWire[14]}}};
  wire [7:0]       maskForGroupWire_hi_hi = {maskForGroupWire_hi_hi_hi, maskForGroupWire_hi_hi_lo};
  wire [15:0]      maskForGroupWire_hi = {maskForGroupWire_hi_hi, maskForGroupWire_hi_lo};
  wire [3:0]       maskForGroupWire_lo_lo_lo_1 = {{2{maskWire[1]}}, {2{maskWire[0]}}};
  wire [3:0]       maskForGroupWire_lo_lo_hi_1 = {{2{maskWire[3]}}, {2{maskWire[2]}}};
  wire [7:0]       maskForGroupWire_lo_lo_1 = {maskForGroupWire_lo_lo_hi_1, maskForGroupWire_lo_lo_lo_1};
  wire [3:0]       maskForGroupWire_lo_hi_lo_1 = {{2{maskWire[5]}}, {2{maskWire[4]}}};
  wire [3:0]       maskForGroupWire_lo_hi_hi_1 = {{2{maskWire[7]}}, {2{maskWire[6]}}};
  wire [7:0]       maskForGroupWire_lo_hi_1 = {maskForGroupWire_lo_hi_hi_1, maskForGroupWire_lo_hi_lo_1};
  wire [15:0]      maskForGroupWire_lo_1 = {maskForGroupWire_lo_hi_1, maskForGroupWire_lo_lo_1};
  wire [3:0]       maskForGroupWire_hi_lo_lo_1 = {{2{maskWire[9]}}, {2{maskWire[8]}}};
  wire [3:0]       maskForGroupWire_hi_lo_hi_1 = {{2{maskWire[11]}}, {2{maskWire[10]}}};
  wire [7:0]       maskForGroupWire_hi_lo_1 = {maskForGroupWire_hi_lo_hi_1, maskForGroupWire_hi_lo_lo_1};
  wire [3:0]       maskForGroupWire_hi_hi_lo_1 = {{2{maskWire[13]}}, {2{maskWire[12]}}};
  wire [3:0]       maskForGroupWire_hi_hi_hi_1 = {{2{maskWire[15]}}, {2{maskWire[14]}}};
  wire [7:0]       maskForGroupWire_hi_hi_1 = {maskForGroupWire_hi_hi_hi_1, maskForGroupWire_hi_hi_lo_1};
  wire [15:0]      maskForGroupWire_hi_1 = {maskForGroupWire_hi_hi_1, maskForGroupWire_hi_lo_1};
  wire [3:0]       _maskForGroupWire_T_69 = 4'h1 << maskCounterInGroup;
  wire [7:0]       maskForGroupWire_lo_lo_lo_2 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]       maskForGroupWire_lo_lo_hi_2 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]      maskForGroupWire_lo_lo_2 = {maskForGroupWire_lo_lo_hi_2, maskForGroupWire_lo_lo_lo_2};
  wire [7:0]       maskForGroupWire_lo_hi_lo_2 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]       maskForGroupWire_lo_hi_hi_2 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]      maskForGroupWire_lo_hi_2 = {maskForGroupWire_lo_hi_hi_2, maskForGroupWire_lo_hi_lo_2};
  wire [31:0]      maskForGroupWire_lo_2 = {maskForGroupWire_lo_hi_2, maskForGroupWire_lo_lo_2};
  wire [7:0]       maskForGroupWire_hi_lo_lo_2 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]       maskForGroupWire_hi_lo_hi_2 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]      maskForGroupWire_hi_lo_2 = {maskForGroupWire_hi_lo_hi_2, maskForGroupWire_hi_lo_lo_2};
  wire [7:0]       maskForGroupWire_hi_hi_lo_2 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]       maskForGroupWire_hi_hi_hi_2 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]      maskForGroupWire_hi_hi_2 = {maskForGroupWire_hi_hi_hi_2, maskForGroupWire_hi_hi_lo_2};
  wire [31:0]      maskForGroupWire_hi_2 = {maskForGroupWire_hi_hi_2, maskForGroupWire_hi_lo_2};
  wire [7:0]       maskForGroupWire_lo_lo_lo_3 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]       maskForGroupWire_lo_lo_hi_3 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]      maskForGroupWire_lo_lo_3 = {maskForGroupWire_lo_lo_hi_3, maskForGroupWire_lo_lo_lo_3};
  wire [7:0]       maskForGroupWire_lo_hi_lo_3 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]       maskForGroupWire_lo_hi_hi_3 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]      maskForGroupWire_lo_hi_3 = {maskForGroupWire_lo_hi_hi_3, maskForGroupWire_lo_hi_lo_3};
  wire [31:0]      maskForGroupWire_lo_3 = {maskForGroupWire_lo_hi_3, maskForGroupWire_lo_lo_3};
  wire [7:0]       maskForGroupWire_hi_lo_lo_3 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]       maskForGroupWire_hi_lo_hi_3 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]      maskForGroupWire_hi_lo_3 = {maskForGroupWire_hi_lo_hi_3, maskForGroupWire_hi_lo_lo_3};
  wire [7:0]       maskForGroupWire_hi_hi_lo_3 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]       maskForGroupWire_hi_hi_hi_3 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]      maskForGroupWire_hi_hi_3 = {maskForGroupWire_hi_hi_hi_3, maskForGroupWire_hi_hi_lo_3};
  wire [31:0]      maskForGroupWire_hi_3 = {maskForGroupWire_hi_hi_3, maskForGroupWire_hi_lo_3};
  wire [7:0]       maskForGroupWire_lo_lo_lo_4 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]       maskForGroupWire_lo_lo_hi_4 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]      maskForGroupWire_lo_lo_4 = {maskForGroupWire_lo_lo_hi_4, maskForGroupWire_lo_lo_lo_4};
  wire [7:0]       maskForGroupWire_lo_hi_lo_4 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]       maskForGroupWire_lo_hi_hi_4 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]      maskForGroupWire_lo_hi_4 = {maskForGroupWire_lo_hi_hi_4, maskForGroupWire_lo_hi_lo_4};
  wire [31:0]      maskForGroupWire_lo_4 = {maskForGroupWire_lo_hi_4, maskForGroupWire_lo_lo_4};
  wire [7:0]       maskForGroupWire_hi_lo_lo_4 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]       maskForGroupWire_hi_lo_hi_4 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]      maskForGroupWire_hi_lo_4 = {maskForGroupWire_hi_lo_hi_4, maskForGroupWire_hi_lo_lo_4};
  wire [7:0]       maskForGroupWire_hi_hi_lo_4 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]       maskForGroupWire_hi_hi_hi_4 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]      maskForGroupWire_hi_hi_4 = {maskForGroupWire_hi_hi_hi_4, maskForGroupWire_hi_hi_lo_4};
  wire [31:0]      maskForGroupWire_hi_4 = {maskForGroupWire_hi_hi_4, maskForGroupWire_hi_lo_4};
  wire [7:0]       maskForGroupWire_lo_lo_lo_5 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]       maskForGroupWire_lo_lo_hi_5 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]      maskForGroupWire_lo_lo_5 = {maskForGroupWire_lo_lo_hi_5, maskForGroupWire_lo_lo_lo_5};
  wire [7:0]       maskForGroupWire_lo_hi_lo_5 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]       maskForGroupWire_lo_hi_hi_5 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]      maskForGroupWire_lo_hi_5 = {maskForGroupWire_lo_hi_hi_5, maskForGroupWire_lo_hi_lo_5};
  wire [31:0]      maskForGroupWire_lo_5 = {maskForGroupWire_lo_hi_5, maskForGroupWire_lo_lo_5};
  wire [7:0]       maskForGroupWire_hi_lo_lo_5 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]       maskForGroupWire_hi_lo_hi_5 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]      maskForGroupWire_hi_lo_5 = {maskForGroupWire_hi_lo_hi_5, maskForGroupWire_hi_lo_lo_5};
  wire [7:0]       maskForGroupWire_hi_hi_lo_5 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]       maskForGroupWire_hi_hi_hi_5 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]      maskForGroupWire_hi_hi_5 = {maskForGroupWire_hi_hi_hi_5, maskForGroupWire_hi_hi_lo_5};
  wire [31:0]      maskForGroupWire_hi_5 = {maskForGroupWire_hi_hi_5, maskForGroupWire_hi_lo_5};
  wire [15:0]      maskForGroupWire =
    (dataEEWOH[0] ? maskWire : 16'h0) | (dataEEWOH[1] ? (maskCounterInGroup[0] ? maskForGroupWire_hi : maskForGroupWire_lo_1) : 16'h0)
    | (dataEEWOH[2]
         ? (_maskForGroupWire_T_69[0] ? maskForGroupWire_lo_2[15:0] : 16'h0) | (_maskForGroupWire_T_69[1] ? maskForGroupWire_lo_3[31:16] : 16'h0) | (_maskForGroupWire_T_69[2] ? maskForGroupWire_hi_4[15:0] : 16'h0)
           | (_maskForGroupWire_T_69[3] ? maskForGroupWire_hi_5[31:16] : 16'h0)
         : 16'h0);
  wire [1:0]       initSendState_lo = maskForGroupWire[1:0];
  wire [1:0]       fillBySeg_lo_lo_lo = maskForGroupWire[1:0];
  wire [1:0]       initSendState_hi = maskForGroupWire[3:2];
  wire [1:0]       fillBySeg_lo_lo_hi = maskForGroupWire[3:2];
  wire             initSendState_0 = |{initSendState_hi, initSendState_lo};
  wire [1:0]       initSendState_lo_1 = maskForGroupWire[5:4];
  wire [1:0]       fillBySeg_lo_hi_lo = maskForGroupWire[5:4];
  wire [1:0]       initSendState_hi_1 = maskForGroupWire[7:6];
  wire [1:0]       fillBySeg_lo_hi_hi = maskForGroupWire[7:6];
  wire             initSendState_1 = |{initSendState_hi_1, initSendState_lo_1};
  wire [1:0]       initSendState_lo_2 = maskForGroupWire[9:8];
  wire [1:0]       fillBySeg_hi_lo_lo = maskForGroupWire[9:8];
  wire [1:0]       initSendState_hi_2 = maskForGroupWire[11:10];
  wire [1:0]       fillBySeg_hi_lo_hi = maskForGroupWire[11:10];
  wire             initSendState_2 = |{initSendState_hi_2, initSendState_lo_2};
  wire [1:0]       initSendState_lo_3 = maskForGroupWire[13:12];
  wire [1:0]       fillBySeg_hi_hi_lo = maskForGroupWire[13:12];
  wire [1:0]       initSendState_hi_3 = maskForGroupWire[15:14];
  wire [1:0]       fillBySeg_hi_hi_hi = maskForGroupWire[15:14];
  wire             initSendState_3 = |{initSendState_hi_3, initSendState_lo_3};
  reg  [127:0]     accessData_0;
  wire [127:0]     accessDataUpdate_1 = accessData_0;
  reg  [127:0]     accessData_1;
  wire [127:0]     accessDataUpdate_2 = accessData_1;
  reg  [127:0]     accessData_2;
  wire [127:0]     accessDataUpdate_3 = accessData_2;
  reg  [127:0]     accessData_3;
  wire [127:0]     accessDataUpdate_4 = accessData_3;
  reg  [127:0]     accessData_4;
  wire [127:0]     accessDataUpdate_5 = accessData_4;
  reg  [127:0]     accessData_5;
  wire [127:0]     accessDataUpdate_6 = accessData_5;
  reg  [127:0]     accessData_6;
  wire [127:0]     accessDataUpdate_7 = accessData_6;
  reg  [127:0]     accessData_7;
  reg  [2:0]       accessPtr;
  reg  [7:0]       dataGroup;
  reg  [127:0]     dataBuffer_0;
  reg  [127:0]     dataBuffer_1;
  reg  [127:0]     dataBuffer_2;
  reg  [127:0]     dataBuffer_3;
  reg  [127:0]     dataBuffer_4;
  reg  [127:0]     dataBuffer_5;
  reg  [127:0]     dataBuffer_6;
  reg  [127:0]     dataBuffer_7;
  reg  [8:0]       bufferBaseCacheLineIndex;
  wire [8:0]       memRequest_bits_index_0 = bufferBaseCacheLineIndex;
  reg  [2:0]       cacheLineIndexInBuffer;
  wire [3:0]       initOffset = lsuRequestReg_rs1Data[3:0];
  wire             invalidInstruction = csrInterface_vl == 13'h0;
  reg              invalidInstructionNext;
  wire             wholeType = lsuRequest_bits_instructionInformation_lumop[3];
  wire [2:0]       nfCorrection = wholeType ? 3'h0 : lsuRequest_bits_instructionInformation_nf;
  reg  [3:0]       segmentInstructionIndexInterval;
  wire [19:0]      bytePerInstruction = {3'h0, {13'h0, {1'h0, nfCorrection} + 4'h1} * {4'h0, csrInterface_vl}} << lsuRequest_bits_instructionInformation_eew;
  wire [19:0]      accessMemSize = bytePerInstruction + {16'h0, lsuRequest_bits_rs1Data[3:0]};
  wire [15:0]      lastCacheLineIndex = accessMemSize[19:4] - {15'h0, accessMemSize[3:0] == 4'h0};
  wire [15:0]      lastWriteVrfIndex = bytePerInstruction[19:4] - {15'h0, bytePerInstruction[3:0] == 4'h0};
  reg  [15:0]      lastWriteVrfIndexReg;
  reg              lastCacheNeedPush;
  reg  [15:0]      cacheLineNumberReg;
  wire [15:0]      dataByteSize = {3'h0, csrInterface_vl} << lsuRequest_bits_instructionInformation_eew;
  wire [11:0]      lastDataGroupForInstruction = dataByteSize[15:4] - {11'h0, dataByteSize[3:0] == 4'h0};
  reg  [11:0]      lastDataGroupReg;
  wire [7:0]       nextDataGroup = lsuRequest_valid ? 8'h0 : dataGroup + 8'h1;
  wire             isLastRead = {4'h0, dataGroup} == lastDataGroupReg;
  reg              hazardCheck;
  wire             accessBufferEnqueueFire;
  wire             vrfReadQueueVec_0_deq_ready;
  wire             vrfReadQueueVec_0_enq_ready = ~_vrfReadQueueVec_fifo_full | vrfReadQueueVec_0_deq_ready;
  wire             vrfReadQueueVec_0_deq_valid = ~_vrfReadQueueVec_fifo_empty | vrfReadQueueVec_0_enq_valid;
  wire [31:0]      vrfReadQueueVec_0_deq_bits = _vrfReadQueueVec_fifo_empty ? vrfReadQueueVec_0_enq_bits : _vrfReadQueueVec_fifo_data_out;
  wire             vrfReadQueueVec_1_deq_ready;
  wire             vrfReadQueueVec_1_enq_ready = ~_vrfReadQueueVec_fifo_1_full | vrfReadQueueVec_1_deq_ready;
  wire             vrfReadQueueVec_1_deq_valid = ~_vrfReadQueueVec_fifo_1_empty | vrfReadQueueVec_1_enq_valid;
  wire [31:0]      vrfReadQueueVec_1_deq_bits = _vrfReadQueueVec_fifo_1_empty ? vrfReadQueueVec_1_enq_bits : _vrfReadQueueVec_fifo_1_data_out;
  wire             vrfReadQueueVec_2_deq_ready;
  wire             vrfReadQueueVec_2_enq_ready = ~_vrfReadQueueVec_fifo_2_full | vrfReadQueueVec_2_deq_ready;
  wire             vrfReadQueueVec_2_deq_valid = ~_vrfReadQueueVec_fifo_2_empty | vrfReadQueueVec_2_enq_valid;
  wire [31:0]      vrfReadQueueVec_2_deq_bits = _vrfReadQueueVec_fifo_2_empty ? vrfReadQueueVec_2_enq_bits : _vrfReadQueueVec_fifo_2_data_out;
  wire             vrfReadQueueVec_3_deq_ready;
  wire             vrfReadQueueVec_3_enq_ready = ~_vrfReadQueueVec_fifo_3_full | vrfReadQueueVec_3_deq_ready;
  wire             vrfReadQueueVec_3_deq_valid = ~_vrfReadQueueVec_fifo_3_empty | vrfReadQueueVec_3_enq_valid;
  wire [31:0]      vrfReadQueueVec_3_deq_bits = _vrfReadQueueVec_fifo_3_empty ? vrfReadQueueVec_3_enq_bits : _vrfReadQueueVec_fifo_3_data_out;
  reg  [2:0]       readStageValid_segPtr;
  reg  [7:0]       readStageValid_readCount;
  reg              readStageValid_stageValid;
  wire             readStageValid_lastReadPtr = readStageValid_segPtr == 3'h0;
  wire [7:0]       readStageValid_nextReadCount = lsuRequest_valid ? 8'h0 : readStageValid_readCount + 8'h1;
  wire             readStageValid_lastReadGroup = {4'h0, readStageValid_readCount} == lastDataGroupReg;
  wire             vrfReadDataPorts_0_valid_0;
  wire             _readStageValid_T_11 = vrfReadDataPorts_0_ready_0 & vrfReadDataPorts_0_valid_0;
  reg  [3:0]       readStageValid_readCounter;
  wire [3:0]       readStageValid_counterChange = _readStageValid_T_11 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_0_valid_0 = readStageValid_stageValid & ~(readStageValid_readCounter[3]);
  wire [4:0]       _GEN_2 = {1'h0, segmentInstructionIndexInterval};
  wire [4:0]       vrfReadDataPorts_0_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr} * _GEN_2 + {2'h0, readStageValid_readCount[7:5]};
  wire [4:0]       vrfReadDataPorts_0_bits_offset_0 = readStageValid_readCount[4:0];
  reg  [2:0]       readStageValid_segPtr_1;
  reg  [7:0]       readStageValid_readCount_1;
  reg              readStageValid_stageValid_1;
  wire             readStageValid_lastReadPtr_1 = readStageValid_segPtr_1 == 3'h0;
  wire [7:0]       readStageValid_nextReadCount_1 = lsuRequest_valid ? 8'h0 : readStageValid_readCount_1 + 8'h1;
  wire             readStageValid_lastReadGroup_1 = {4'h0, readStageValid_readCount_1} == lastDataGroupReg;
  wire             vrfReadDataPorts_1_valid_0;
  wire             _readStageValid_T_30 = vrfReadDataPorts_1_ready_0 & vrfReadDataPorts_1_valid_0;
  reg  [3:0]       readStageValid_readCounter_1;
  wire [3:0]       readStageValid_counterChange_1 = _readStageValid_T_30 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_1_valid_0 = readStageValid_stageValid_1 & ~(readStageValid_readCounter_1[3]);
  wire [4:0]       vrfReadDataPorts_1_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_1} * _GEN_2 + {2'h0, readStageValid_readCount_1[7:5]};
  wire [4:0]       vrfReadDataPorts_1_bits_offset_0 = readStageValid_readCount_1[4:0];
  reg  [2:0]       readStageValid_segPtr_2;
  reg  [7:0]       readStageValid_readCount_2;
  reg              readStageValid_stageValid_2;
  wire             readStageValid_lastReadPtr_2 = readStageValid_segPtr_2 == 3'h0;
  wire [7:0]       readStageValid_nextReadCount_2 = lsuRequest_valid ? 8'h0 : readStageValid_readCount_2 + 8'h1;
  wire             readStageValid_lastReadGroup_2 = {4'h0, readStageValid_readCount_2} == lastDataGroupReg;
  wire             vrfReadDataPorts_2_valid_0;
  wire             _readStageValid_T_49 = vrfReadDataPorts_2_ready_0 & vrfReadDataPorts_2_valid_0;
  reg  [3:0]       readStageValid_readCounter_2;
  wire [3:0]       readStageValid_counterChange_2 = _readStageValid_T_49 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_2_valid_0 = readStageValid_stageValid_2 & ~(readStageValid_readCounter_2[3]);
  wire [4:0]       vrfReadDataPorts_2_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_2} * _GEN_2 + {2'h0, readStageValid_readCount_2[7:5]};
  wire [4:0]       vrfReadDataPorts_2_bits_offset_0 = readStageValid_readCount_2[4:0];
  reg  [2:0]       readStageValid_segPtr_3;
  reg  [7:0]       readStageValid_readCount_3;
  reg              readStageValid_stageValid_3;
  wire             readStageValid_lastReadPtr_3 = readStageValid_segPtr_3 == 3'h0;
  wire [7:0]       readStageValid_nextReadCount_3 = lsuRequest_valid ? 8'h0 : readStageValid_readCount_3 + 8'h1;
  wire             readStageValid_lastReadGroup_3 = {4'h0, readStageValid_readCount_3} == lastDataGroupReg;
  wire             vrfReadDataPorts_3_valid_0;
  wire             _readStageValid_T_68 = vrfReadDataPorts_3_ready_0 & vrfReadDataPorts_3_valid_0;
  reg  [3:0]       readStageValid_readCounter_3;
  wire [3:0]       readStageValid_counterChange_3 = _readStageValid_T_68 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_3_valid_0 = readStageValid_stageValid_3 & ~(readStageValid_readCounter_3[3]);
  wire [4:0]       vrfReadDataPorts_3_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_3} * _GEN_2 + {2'h0, readStageValid_readCount_3[7:5]};
  wire [4:0]       vrfReadDataPorts_3_bits_offset_0 = readStageValid_readCount_3[4:0];
  wire             readStageValid =
    |{readStageValid_stageValid, readStageValid_readCounter, readStageValid_stageValid_1, readStageValid_readCounter_1, readStageValid_stageValid_2, readStageValid_readCounter_2, readStageValid_stageValid_3, readStageValid_readCounter_3};
  reg              bufferFull;
  wire             accessBufferDequeueReady;
  wire             accessBufferEnqueueReady = ~bufferFull | accessBufferDequeueReady;
  wire             accessBufferEnqueueValid = vrfReadQueueVec_0_deq_valid & vrfReadQueueVec_1_deq_valid & vrfReadQueueVec_2_deq_valid & vrfReadQueueVec_3_deq_valid;
  wire             readQueueClear = ~(vrfReadQueueVec_0_deq_valid | vrfReadQueueVec_1_deq_valid | vrfReadQueueVec_2_deq_valid | vrfReadQueueVec_3_deq_valid);
  assign accessBufferEnqueueFire = accessBufferEnqueueValid & accessBufferEnqueueReady;
  assign vrfReadQueueVec_0_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_1_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_2_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_3_deq_ready = accessBufferEnqueueFire;
  wire             lastPtr = accessPtr == 3'h0;
  wire             lastPtrEnq = lastPtr & accessBufferEnqueueFire;
  wire             accessBufferDequeueValid = bufferFull | lastPtrEnq;
  wire             accessBufferDequeueFire = accessBufferDequeueValid & accessBufferDequeueReady;
  wire [63:0]      accessDataUpdate_lo = {vrfReadQueueVec_1_deq_bits, vrfReadQueueVec_0_deq_bits};
  wire [63:0]      accessDataUpdate_hi = {vrfReadQueueVec_3_deq_bits, vrfReadQueueVec_2_deq_bits};
  wire [127:0]     accessDataUpdate_0 = {accessDataUpdate_hi, accessDataUpdate_lo};
  reg              bufferValid;
  reg  [15:0]      maskForBufferData_0;
  reg  [15:0]      maskForBufferData_1;
  reg  [15:0]      maskForBufferData_2;
  reg  [15:0]      maskForBufferData_3;
  reg  [15:0]      maskForBufferData_4;
  reg  [15:0]      maskForBufferData_5;
  reg  [15:0]      maskForBufferData_6;
  reg  [15:0]      maskForBufferData_7;
  reg              lastDataGroupInDataBuffer;
  wire             memRequest_valid_0;
  wire             _addressQueue_enq_valid_T = memRequest_ready_0 & memRequest_valid_0;
  wire             alignedDequeueFire;
  assign alignedDequeueFire = _addressQueue_enq_valid_T;
  wire             addressQueue_enq_valid;
  assign addressQueue_enq_valid = _addressQueue_enq_valid_T;
  reg  [127:0]     cacheLineTemp;
  reg  [15:0]      maskTemp;
  reg              canSendTail;
  wire             isLastCacheLineInBuffer = cacheLineIndexInBuffer == lsuRequestReg_instructionInformation_nf;
  wire             bufferWillClear = alignedDequeueFire & isLastCacheLineInBuffer;
  wire             addressQueue_enq_ready;
  wire             addressQueueFree;
  assign accessBufferDequeueReady = ~bufferValid | memRequest_ready_0 & isLastCacheLineInBuffer & addressQueueFree;
  wire [127:0]     bufferStageEnqueueData_0 = bufferFull ? accessData_0 : accessDataUpdate_0;
  wire [127:0]     bufferStageEnqueueData_1 = bufferFull ? accessData_1 : accessDataUpdate_1;
  wire [127:0]     bufferStageEnqueueData_2 = bufferFull ? accessData_2 : accessDataUpdate_2;
  wire [127:0]     bufferStageEnqueueData_3 = bufferFull ? accessData_3 : accessDataUpdate_3;
  wire [127:0]     bufferStageEnqueueData_4 = bufferFull ? accessData_4 : accessDataUpdate_4;
  wire [127:0]     bufferStageEnqueueData_5 = bufferFull ? accessData_5 : accessDataUpdate_5;
  wire [127:0]     bufferStageEnqueueData_6 = bufferFull ? accessData_6 : accessDataUpdate_6;
  wire [127:0]     bufferStageEnqueueData_7 = bufferFull ? accessData_7 : accessDataUpdate_7;
  wire [7:0]       _fillBySeg_T = 8'h1 << lsuRequestReg_instructionInformation_nf;
  wire [3:0]       fillBySeg_lo_lo = {fillBySeg_lo_lo_hi, fillBySeg_lo_lo_lo};
  wire [3:0]       fillBySeg_lo_hi = {fillBySeg_lo_hi_hi, fillBySeg_lo_hi_lo};
  wire [7:0]       fillBySeg_lo = {fillBySeg_lo_hi, fillBySeg_lo_lo};
  wire [3:0]       fillBySeg_hi_lo = {fillBySeg_hi_lo_hi, fillBySeg_hi_lo_lo};
  wire [3:0]       fillBySeg_hi_hi = {fillBySeg_hi_hi_hi, fillBySeg_hi_hi_lo};
  wire [7:0]       fillBySeg_hi = {fillBySeg_hi_hi, fillBySeg_hi_lo};
  wire [3:0]       fillBySeg_lo_lo_lo_1 = {{2{maskForGroupWire[1]}}, {2{maskForGroupWire[0]}}};
  wire [3:0]       fillBySeg_lo_lo_hi_1 = {{2{maskForGroupWire[3]}}, {2{maskForGroupWire[2]}}};
  wire [7:0]       fillBySeg_lo_lo_1 = {fillBySeg_lo_lo_hi_1, fillBySeg_lo_lo_lo_1};
  wire [3:0]       fillBySeg_lo_hi_lo_1 = {{2{maskForGroupWire[5]}}, {2{maskForGroupWire[4]}}};
  wire [3:0]       fillBySeg_lo_hi_hi_1 = {{2{maskForGroupWire[7]}}, {2{maskForGroupWire[6]}}};
  wire [7:0]       fillBySeg_lo_hi_1 = {fillBySeg_lo_hi_hi_1, fillBySeg_lo_hi_lo_1};
  wire [15:0]      fillBySeg_lo_1 = {fillBySeg_lo_hi_1, fillBySeg_lo_lo_1};
  wire [3:0]       fillBySeg_hi_lo_lo_1 = {{2{maskForGroupWire[9]}}, {2{maskForGroupWire[8]}}};
  wire [3:0]       fillBySeg_hi_lo_hi_1 = {{2{maskForGroupWire[11]}}, {2{maskForGroupWire[10]}}};
  wire [7:0]       fillBySeg_hi_lo_1 = {fillBySeg_hi_lo_hi_1, fillBySeg_hi_lo_lo_1};
  wire [3:0]       fillBySeg_hi_hi_lo_1 = {{2{maskForGroupWire[13]}}, {2{maskForGroupWire[12]}}};
  wire [3:0]       fillBySeg_hi_hi_hi_1 = {{2{maskForGroupWire[15]}}, {2{maskForGroupWire[14]}}};
  wire [7:0]       fillBySeg_hi_hi_1 = {fillBySeg_hi_hi_hi_1, fillBySeg_hi_hi_lo_1};
  wire [15:0]      fillBySeg_hi_1 = {fillBySeg_hi_hi_1, fillBySeg_hi_lo_1};
  wire [5:0]       fillBySeg_lo_lo_lo_2 = {{3{maskForGroupWire[1]}}, {3{maskForGroupWire[0]}}};
  wire [5:0]       fillBySeg_lo_lo_hi_2 = {{3{maskForGroupWire[3]}}, {3{maskForGroupWire[2]}}};
  wire [11:0]      fillBySeg_lo_lo_2 = {fillBySeg_lo_lo_hi_2, fillBySeg_lo_lo_lo_2};
  wire [5:0]       fillBySeg_lo_hi_lo_2 = {{3{maskForGroupWire[5]}}, {3{maskForGroupWire[4]}}};
  wire [5:0]       fillBySeg_lo_hi_hi_2 = {{3{maskForGroupWire[7]}}, {3{maskForGroupWire[6]}}};
  wire [11:0]      fillBySeg_lo_hi_2 = {fillBySeg_lo_hi_hi_2, fillBySeg_lo_hi_lo_2};
  wire [23:0]      fillBySeg_lo_2 = {fillBySeg_lo_hi_2, fillBySeg_lo_lo_2};
  wire [5:0]       fillBySeg_hi_lo_lo_2 = {{3{maskForGroupWire[9]}}, {3{maskForGroupWire[8]}}};
  wire [5:0]       fillBySeg_hi_lo_hi_2 = {{3{maskForGroupWire[11]}}, {3{maskForGroupWire[10]}}};
  wire [11:0]      fillBySeg_hi_lo_2 = {fillBySeg_hi_lo_hi_2, fillBySeg_hi_lo_lo_2};
  wire [5:0]       fillBySeg_hi_hi_lo_2 = {{3{maskForGroupWire[13]}}, {3{maskForGroupWire[12]}}};
  wire [5:0]       fillBySeg_hi_hi_hi_2 = {{3{maskForGroupWire[15]}}, {3{maskForGroupWire[14]}}};
  wire [11:0]      fillBySeg_hi_hi_2 = {fillBySeg_hi_hi_hi_2, fillBySeg_hi_hi_lo_2};
  wire [23:0]      fillBySeg_hi_2 = {fillBySeg_hi_hi_2, fillBySeg_hi_lo_2};
  wire [7:0]       fillBySeg_lo_lo_lo_3 = {{4{maskForGroupWire[1]}}, {4{maskForGroupWire[0]}}};
  wire [7:0]       fillBySeg_lo_lo_hi_3 = {{4{maskForGroupWire[3]}}, {4{maskForGroupWire[2]}}};
  wire [15:0]      fillBySeg_lo_lo_3 = {fillBySeg_lo_lo_hi_3, fillBySeg_lo_lo_lo_3};
  wire [7:0]       fillBySeg_lo_hi_lo_3 = {{4{maskForGroupWire[5]}}, {4{maskForGroupWire[4]}}};
  wire [7:0]       fillBySeg_lo_hi_hi_3 = {{4{maskForGroupWire[7]}}, {4{maskForGroupWire[6]}}};
  wire [15:0]      fillBySeg_lo_hi_3 = {fillBySeg_lo_hi_hi_3, fillBySeg_lo_hi_lo_3};
  wire [31:0]      fillBySeg_lo_3 = {fillBySeg_lo_hi_3, fillBySeg_lo_lo_3};
  wire [7:0]       fillBySeg_hi_lo_lo_3 = {{4{maskForGroupWire[9]}}, {4{maskForGroupWire[8]}}};
  wire [7:0]       fillBySeg_hi_lo_hi_3 = {{4{maskForGroupWire[11]}}, {4{maskForGroupWire[10]}}};
  wire [15:0]      fillBySeg_hi_lo_3 = {fillBySeg_hi_lo_hi_3, fillBySeg_hi_lo_lo_3};
  wire [7:0]       fillBySeg_hi_hi_lo_3 = {{4{maskForGroupWire[13]}}, {4{maskForGroupWire[12]}}};
  wire [7:0]       fillBySeg_hi_hi_hi_3 = {{4{maskForGroupWire[15]}}, {4{maskForGroupWire[14]}}};
  wire [15:0]      fillBySeg_hi_hi_3 = {fillBySeg_hi_hi_hi_3, fillBySeg_hi_hi_lo_3};
  wire [31:0]      fillBySeg_hi_3 = {fillBySeg_hi_hi_3, fillBySeg_hi_lo_3};
  wire [9:0]       fillBySeg_lo_lo_lo_4 = {{5{maskForGroupWire[1]}}, {5{maskForGroupWire[0]}}};
  wire [9:0]       fillBySeg_lo_lo_hi_4 = {{5{maskForGroupWire[3]}}, {5{maskForGroupWire[2]}}};
  wire [19:0]      fillBySeg_lo_lo_4 = {fillBySeg_lo_lo_hi_4, fillBySeg_lo_lo_lo_4};
  wire [9:0]       fillBySeg_lo_hi_lo_4 = {{5{maskForGroupWire[5]}}, {5{maskForGroupWire[4]}}};
  wire [9:0]       fillBySeg_lo_hi_hi_4 = {{5{maskForGroupWire[7]}}, {5{maskForGroupWire[6]}}};
  wire [19:0]      fillBySeg_lo_hi_4 = {fillBySeg_lo_hi_hi_4, fillBySeg_lo_hi_lo_4};
  wire [39:0]      fillBySeg_lo_4 = {fillBySeg_lo_hi_4, fillBySeg_lo_lo_4};
  wire [9:0]       fillBySeg_hi_lo_lo_4 = {{5{maskForGroupWire[9]}}, {5{maskForGroupWire[8]}}};
  wire [9:0]       fillBySeg_hi_lo_hi_4 = {{5{maskForGroupWire[11]}}, {5{maskForGroupWire[10]}}};
  wire [19:0]      fillBySeg_hi_lo_4 = {fillBySeg_hi_lo_hi_4, fillBySeg_hi_lo_lo_4};
  wire [9:0]       fillBySeg_hi_hi_lo_4 = {{5{maskForGroupWire[13]}}, {5{maskForGroupWire[12]}}};
  wire [9:0]       fillBySeg_hi_hi_hi_4 = {{5{maskForGroupWire[15]}}, {5{maskForGroupWire[14]}}};
  wire [19:0]      fillBySeg_hi_hi_4 = {fillBySeg_hi_hi_hi_4, fillBySeg_hi_hi_lo_4};
  wire [39:0]      fillBySeg_hi_4 = {fillBySeg_hi_hi_4, fillBySeg_hi_lo_4};
  wire [11:0]      fillBySeg_lo_lo_lo_5 = {{6{maskForGroupWire[1]}}, {6{maskForGroupWire[0]}}};
  wire [11:0]      fillBySeg_lo_lo_hi_5 = {{6{maskForGroupWire[3]}}, {6{maskForGroupWire[2]}}};
  wire [23:0]      fillBySeg_lo_lo_5 = {fillBySeg_lo_lo_hi_5, fillBySeg_lo_lo_lo_5};
  wire [11:0]      fillBySeg_lo_hi_lo_5 = {{6{maskForGroupWire[5]}}, {6{maskForGroupWire[4]}}};
  wire [11:0]      fillBySeg_lo_hi_hi_5 = {{6{maskForGroupWire[7]}}, {6{maskForGroupWire[6]}}};
  wire [23:0]      fillBySeg_lo_hi_5 = {fillBySeg_lo_hi_hi_5, fillBySeg_lo_hi_lo_5};
  wire [47:0]      fillBySeg_lo_5 = {fillBySeg_lo_hi_5, fillBySeg_lo_lo_5};
  wire [11:0]      fillBySeg_hi_lo_lo_5 = {{6{maskForGroupWire[9]}}, {6{maskForGroupWire[8]}}};
  wire [11:0]      fillBySeg_hi_lo_hi_5 = {{6{maskForGroupWire[11]}}, {6{maskForGroupWire[10]}}};
  wire [23:0]      fillBySeg_hi_lo_5 = {fillBySeg_hi_lo_hi_5, fillBySeg_hi_lo_lo_5};
  wire [11:0]      fillBySeg_hi_hi_lo_5 = {{6{maskForGroupWire[13]}}, {6{maskForGroupWire[12]}}};
  wire [11:0]      fillBySeg_hi_hi_hi_5 = {{6{maskForGroupWire[15]}}, {6{maskForGroupWire[14]}}};
  wire [23:0]      fillBySeg_hi_hi_5 = {fillBySeg_hi_hi_hi_5, fillBySeg_hi_hi_lo_5};
  wire [47:0]      fillBySeg_hi_5 = {fillBySeg_hi_hi_5, fillBySeg_hi_lo_5};
  wire [13:0]      fillBySeg_lo_lo_lo_6 = {{7{maskForGroupWire[1]}}, {7{maskForGroupWire[0]}}};
  wire [13:0]      fillBySeg_lo_lo_hi_6 = {{7{maskForGroupWire[3]}}, {7{maskForGroupWire[2]}}};
  wire [27:0]      fillBySeg_lo_lo_6 = {fillBySeg_lo_lo_hi_6, fillBySeg_lo_lo_lo_6};
  wire [13:0]      fillBySeg_lo_hi_lo_6 = {{7{maskForGroupWire[5]}}, {7{maskForGroupWire[4]}}};
  wire [13:0]      fillBySeg_lo_hi_hi_6 = {{7{maskForGroupWire[7]}}, {7{maskForGroupWire[6]}}};
  wire [27:0]      fillBySeg_lo_hi_6 = {fillBySeg_lo_hi_hi_6, fillBySeg_lo_hi_lo_6};
  wire [55:0]      fillBySeg_lo_6 = {fillBySeg_lo_hi_6, fillBySeg_lo_lo_6};
  wire [13:0]      fillBySeg_hi_lo_lo_6 = {{7{maskForGroupWire[9]}}, {7{maskForGroupWire[8]}}};
  wire [13:0]      fillBySeg_hi_lo_hi_6 = {{7{maskForGroupWire[11]}}, {7{maskForGroupWire[10]}}};
  wire [27:0]      fillBySeg_hi_lo_6 = {fillBySeg_hi_lo_hi_6, fillBySeg_hi_lo_lo_6};
  wire [13:0]      fillBySeg_hi_hi_lo_6 = {{7{maskForGroupWire[13]}}, {7{maskForGroupWire[12]}}};
  wire [13:0]      fillBySeg_hi_hi_hi_6 = {{7{maskForGroupWire[15]}}, {7{maskForGroupWire[14]}}};
  wire [27:0]      fillBySeg_hi_hi_6 = {fillBySeg_hi_hi_hi_6, fillBySeg_hi_hi_lo_6};
  wire [55:0]      fillBySeg_hi_6 = {fillBySeg_hi_hi_6, fillBySeg_hi_lo_6};
  wire [15:0]      fillBySeg_lo_lo_lo_7 = {{8{maskForGroupWire[1]}}, {8{maskForGroupWire[0]}}};
  wire [15:0]      fillBySeg_lo_lo_hi_7 = {{8{maskForGroupWire[3]}}, {8{maskForGroupWire[2]}}};
  wire [31:0]      fillBySeg_lo_lo_7 = {fillBySeg_lo_lo_hi_7, fillBySeg_lo_lo_lo_7};
  wire [15:0]      fillBySeg_lo_hi_lo_7 = {{8{maskForGroupWire[5]}}, {8{maskForGroupWire[4]}}};
  wire [15:0]      fillBySeg_lo_hi_hi_7 = {{8{maskForGroupWire[7]}}, {8{maskForGroupWire[6]}}};
  wire [31:0]      fillBySeg_lo_hi_7 = {fillBySeg_lo_hi_hi_7, fillBySeg_lo_hi_lo_7};
  wire [63:0]      fillBySeg_lo_7 = {fillBySeg_lo_hi_7, fillBySeg_lo_lo_7};
  wire [15:0]      fillBySeg_hi_lo_lo_7 = {{8{maskForGroupWire[9]}}, {8{maskForGroupWire[8]}}};
  wire [15:0]      fillBySeg_hi_lo_hi_7 = {{8{maskForGroupWire[11]}}, {8{maskForGroupWire[10]}}};
  wire [31:0]      fillBySeg_hi_lo_7 = {fillBySeg_hi_lo_hi_7, fillBySeg_hi_lo_lo_7};
  wire [15:0]      fillBySeg_hi_hi_lo_7 = {{8{maskForGroupWire[13]}}, {8{maskForGroupWire[12]}}};
  wire [15:0]      fillBySeg_hi_hi_hi_7 = {{8{maskForGroupWire[15]}}, {8{maskForGroupWire[14]}}};
  wire [31:0]      fillBySeg_hi_hi_7 = {fillBySeg_hi_hi_hi_7, fillBySeg_hi_hi_lo_7};
  wire [63:0]      fillBySeg_hi_7 = {fillBySeg_hi_hi_7, fillBySeg_hi_lo_7};
  wire [127:0]     fillBySeg =
    {16'h0,
     {16'h0,
      {16'h0,
       {16'h0,
        {16'h0, {16'h0, {16'h0, _fillBySeg_T[0] ? {fillBySeg_hi, fillBySeg_lo} : 16'h0} | (_fillBySeg_T[1] ? {fillBySeg_hi_1, fillBySeg_lo_1} : 32'h0)} | (_fillBySeg_T[2] ? {fillBySeg_hi_2, fillBySeg_lo_2} : 48'h0)}
          | (_fillBySeg_T[3] ? {fillBySeg_hi_3, fillBySeg_lo_3} : 64'h0)} | (_fillBySeg_T[4] ? {fillBySeg_hi_4, fillBySeg_lo_4} : 80'h0)} | (_fillBySeg_T[5] ? {fillBySeg_hi_5, fillBySeg_lo_5} : 96'h0)}
       | (_fillBySeg_T[6] ? {fillBySeg_hi_6, fillBySeg_lo_6} : 112'h0)} | (_fillBySeg_T[7] ? {fillBySeg_hi_7, fillBySeg_lo_7} : 128'h0);
  wire [7:0]       dataRegroupBySew_0_0 = bufferStageEnqueueData_0[7:0];
  wire [7:0]       dataRegroupBySew_0_1 = bufferStageEnqueueData_0[15:8];
  wire [7:0]       dataRegroupBySew_0_2 = bufferStageEnqueueData_0[23:16];
  wire [7:0]       dataRegroupBySew_0_3 = bufferStageEnqueueData_0[31:24];
  wire [7:0]       dataRegroupBySew_0_4 = bufferStageEnqueueData_0[39:32];
  wire [7:0]       dataRegroupBySew_0_5 = bufferStageEnqueueData_0[47:40];
  wire [7:0]       dataRegroupBySew_0_6 = bufferStageEnqueueData_0[55:48];
  wire [7:0]       dataRegroupBySew_0_7 = bufferStageEnqueueData_0[63:56];
  wire [7:0]       dataRegroupBySew_0_8 = bufferStageEnqueueData_0[71:64];
  wire [7:0]       dataRegroupBySew_0_9 = bufferStageEnqueueData_0[79:72];
  wire [7:0]       dataRegroupBySew_0_10 = bufferStageEnqueueData_0[87:80];
  wire [7:0]       dataRegroupBySew_0_11 = bufferStageEnqueueData_0[95:88];
  wire [7:0]       dataRegroupBySew_0_12 = bufferStageEnqueueData_0[103:96];
  wire [7:0]       dataRegroupBySew_0_13 = bufferStageEnqueueData_0[111:104];
  wire [7:0]       dataRegroupBySew_0_14 = bufferStageEnqueueData_0[119:112];
  wire [7:0]       dataRegroupBySew_0_15 = bufferStageEnqueueData_0[127:120];
  wire [7:0]       dataRegroupBySew_1_0 = bufferStageEnqueueData_1[7:0];
  wire [7:0]       dataRegroupBySew_1_1 = bufferStageEnqueueData_1[15:8];
  wire [7:0]       dataRegroupBySew_1_2 = bufferStageEnqueueData_1[23:16];
  wire [7:0]       dataRegroupBySew_1_3 = bufferStageEnqueueData_1[31:24];
  wire [7:0]       dataRegroupBySew_1_4 = bufferStageEnqueueData_1[39:32];
  wire [7:0]       dataRegroupBySew_1_5 = bufferStageEnqueueData_1[47:40];
  wire [7:0]       dataRegroupBySew_1_6 = bufferStageEnqueueData_1[55:48];
  wire [7:0]       dataRegroupBySew_1_7 = bufferStageEnqueueData_1[63:56];
  wire [7:0]       dataRegroupBySew_1_8 = bufferStageEnqueueData_1[71:64];
  wire [7:0]       dataRegroupBySew_1_9 = bufferStageEnqueueData_1[79:72];
  wire [7:0]       dataRegroupBySew_1_10 = bufferStageEnqueueData_1[87:80];
  wire [7:0]       dataRegroupBySew_1_11 = bufferStageEnqueueData_1[95:88];
  wire [7:0]       dataRegroupBySew_1_12 = bufferStageEnqueueData_1[103:96];
  wire [7:0]       dataRegroupBySew_1_13 = bufferStageEnqueueData_1[111:104];
  wire [7:0]       dataRegroupBySew_1_14 = bufferStageEnqueueData_1[119:112];
  wire [7:0]       dataRegroupBySew_1_15 = bufferStageEnqueueData_1[127:120];
  wire [7:0]       dataRegroupBySew_2_0 = bufferStageEnqueueData_2[7:0];
  wire [7:0]       dataRegroupBySew_2_1 = bufferStageEnqueueData_2[15:8];
  wire [7:0]       dataRegroupBySew_2_2 = bufferStageEnqueueData_2[23:16];
  wire [7:0]       dataRegroupBySew_2_3 = bufferStageEnqueueData_2[31:24];
  wire [7:0]       dataRegroupBySew_2_4 = bufferStageEnqueueData_2[39:32];
  wire [7:0]       dataRegroupBySew_2_5 = bufferStageEnqueueData_2[47:40];
  wire [7:0]       dataRegroupBySew_2_6 = bufferStageEnqueueData_2[55:48];
  wire [7:0]       dataRegroupBySew_2_7 = bufferStageEnqueueData_2[63:56];
  wire [7:0]       dataRegroupBySew_2_8 = bufferStageEnqueueData_2[71:64];
  wire [7:0]       dataRegroupBySew_2_9 = bufferStageEnqueueData_2[79:72];
  wire [7:0]       dataRegroupBySew_2_10 = bufferStageEnqueueData_2[87:80];
  wire [7:0]       dataRegroupBySew_2_11 = bufferStageEnqueueData_2[95:88];
  wire [7:0]       dataRegroupBySew_2_12 = bufferStageEnqueueData_2[103:96];
  wire [7:0]       dataRegroupBySew_2_13 = bufferStageEnqueueData_2[111:104];
  wire [7:0]       dataRegroupBySew_2_14 = bufferStageEnqueueData_2[119:112];
  wire [7:0]       dataRegroupBySew_2_15 = bufferStageEnqueueData_2[127:120];
  wire [7:0]       dataRegroupBySew_3_0 = bufferStageEnqueueData_3[7:0];
  wire [7:0]       dataRegroupBySew_3_1 = bufferStageEnqueueData_3[15:8];
  wire [7:0]       dataRegroupBySew_3_2 = bufferStageEnqueueData_3[23:16];
  wire [7:0]       dataRegroupBySew_3_3 = bufferStageEnqueueData_3[31:24];
  wire [7:0]       dataRegroupBySew_3_4 = bufferStageEnqueueData_3[39:32];
  wire [7:0]       dataRegroupBySew_3_5 = bufferStageEnqueueData_3[47:40];
  wire [7:0]       dataRegroupBySew_3_6 = bufferStageEnqueueData_3[55:48];
  wire [7:0]       dataRegroupBySew_3_7 = bufferStageEnqueueData_3[63:56];
  wire [7:0]       dataRegroupBySew_3_8 = bufferStageEnqueueData_3[71:64];
  wire [7:0]       dataRegroupBySew_3_9 = bufferStageEnqueueData_3[79:72];
  wire [7:0]       dataRegroupBySew_3_10 = bufferStageEnqueueData_3[87:80];
  wire [7:0]       dataRegroupBySew_3_11 = bufferStageEnqueueData_3[95:88];
  wire [7:0]       dataRegroupBySew_3_12 = bufferStageEnqueueData_3[103:96];
  wire [7:0]       dataRegroupBySew_3_13 = bufferStageEnqueueData_3[111:104];
  wire [7:0]       dataRegroupBySew_3_14 = bufferStageEnqueueData_3[119:112];
  wire [7:0]       dataRegroupBySew_3_15 = bufferStageEnqueueData_3[127:120];
  wire [7:0]       dataRegroupBySew_4_0 = bufferStageEnqueueData_4[7:0];
  wire [7:0]       dataRegroupBySew_4_1 = bufferStageEnqueueData_4[15:8];
  wire [7:0]       dataRegroupBySew_4_2 = bufferStageEnqueueData_4[23:16];
  wire [7:0]       dataRegroupBySew_4_3 = bufferStageEnqueueData_4[31:24];
  wire [7:0]       dataRegroupBySew_4_4 = bufferStageEnqueueData_4[39:32];
  wire [7:0]       dataRegroupBySew_4_5 = bufferStageEnqueueData_4[47:40];
  wire [7:0]       dataRegroupBySew_4_6 = bufferStageEnqueueData_4[55:48];
  wire [7:0]       dataRegroupBySew_4_7 = bufferStageEnqueueData_4[63:56];
  wire [7:0]       dataRegroupBySew_4_8 = bufferStageEnqueueData_4[71:64];
  wire [7:0]       dataRegroupBySew_4_9 = bufferStageEnqueueData_4[79:72];
  wire [7:0]       dataRegroupBySew_4_10 = bufferStageEnqueueData_4[87:80];
  wire [7:0]       dataRegroupBySew_4_11 = bufferStageEnqueueData_4[95:88];
  wire [7:0]       dataRegroupBySew_4_12 = bufferStageEnqueueData_4[103:96];
  wire [7:0]       dataRegroupBySew_4_13 = bufferStageEnqueueData_4[111:104];
  wire [7:0]       dataRegroupBySew_4_14 = bufferStageEnqueueData_4[119:112];
  wire [7:0]       dataRegroupBySew_4_15 = bufferStageEnqueueData_4[127:120];
  wire [7:0]       dataRegroupBySew_5_0 = bufferStageEnqueueData_5[7:0];
  wire [7:0]       dataRegroupBySew_5_1 = bufferStageEnqueueData_5[15:8];
  wire [7:0]       dataRegroupBySew_5_2 = bufferStageEnqueueData_5[23:16];
  wire [7:0]       dataRegroupBySew_5_3 = bufferStageEnqueueData_5[31:24];
  wire [7:0]       dataRegroupBySew_5_4 = bufferStageEnqueueData_5[39:32];
  wire [7:0]       dataRegroupBySew_5_5 = bufferStageEnqueueData_5[47:40];
  wire [7:0]       dataRegroupBySew_5_6 = bufferStageEnqueueData_5[55:48];
  wire [7:0]       dataRegroupBySew_5_7 = bufferStageEnqueueData_5[63:56];
  wire [7:0]       dataRegroupBySew_5_8 = bufferStageEnqueueData_5[71:64];
  wire [7:0]       dataRegroupBySew_5_9 = bufferStageEnqueueData_5[79:72];
  wire [7:0]       dataRegroupBySew_5_10 = bufferStageEnqueueData_5[87:80];
  wire [7:0]       dataRegroupBySew_5_11 = bufferStageEnqueueData_5[95:88];
  wire [7:0]       dataRegroupBySew_5_12 = bufferStageEnqueueData_5[103:96];
  wire [7:0]       dataRegroupBySew_5_13 = bufferStageEnqueueData_5[111:104];
  wire [7:0]       dataRegroupBySew_5_14 = bufferStageEnqueueData_5[119:112];
  wire [7:0]       dataRegroupBySew_5_15 = bufferStageEnqueueData_5[127:120];
  wire [7:0]       dataRegroupBySew_6_0 = bufferStageEnqueueData_6[7:0];
  wire [7:0]       dataRegroupBySew_6_1 = bufferStageEnqueueData_6[15:8];
  wire [7:0]       dataRegroupBySew_6_2 = bufferStageEnqueueData_6[23:16];
  wire [7:0]       dataRegroupBySew_6_3 = bufferStageEnqueueData_6[31:24];
  wire [7:0]       dataRegroupBySew_6_4 = bufferStageEnqueueData_6[39:32];
  wire [7:0]       dataRegroupBySew_6_5 = bufferStageEnqueueData_6[47:40];
  wire [7:0]       dataRegroupBySew_6_6 = bufferStageEnqueueData_6[55:48];
  wire [7:0]       dataRegroupBySew_6_7 = bufferStageEnqueueData_6[63:56];
  wire [7:0]       dataRegroupBySew_6_8 = bufferStageEnqueueData_6[71:64];
  wire [7:0]       dataRegroupBySew_6_9 = bufferStageEnqueueData_6[79:72];
  wire [7:0]       dataRegroupBySew_6_10 = bufferStageEnqueueData_6[87:80];
  wire [7:0]       dataRegroupBySew_6_11 = bufferStageEnqueueData_6[95:88];
  wire [7:0]       dataRegroupBySew_6_12 = bufferStageEnqueueData_6[103:96];
  wire [7:0]       dataRegroupBySew_6_13 = bufferStageEnqueueData_6[111:104];
  wire [7:0]       dataRegroupBySew_6_14 = bufferStageEnqueueData_6[119:112];
  wire [7:0]       dataRegroupBySew_6_15 = bufferStageEnqueueData_6[127:120];
  wire [7:0]       dataRegroupBySew_7_0 = bufferStageEnqueueData_7[7:0];
  wire [7:0]       dataRegroupBySew_7_1 = bufferStageEnqueueData_7[15:8];
  wire [7:0]       dataRegroupBySew_7_2 = bufferStageEnqueueData_7[23:16];
  wire [7:0]       dataRegroupBySew_7_3 = bufferStageEnqueueData_7[31:24];
  wire [7:0]       dataRegroupBySew_7_4 = bufferStageEnqueueData_7[39:32];
  wire [7:0]       dataRegroupBySew_7_5 = bufferStageEnqueueData_7[47:40];
  wire [7:0]       dataRegroupBySew_7_6 = bufferStageEnqueueData_7[55:48];
  wire [7:0]       dataRegroupBySew_7_7 = bufferStageEnqueueData_7[63:56];
  wire [7:0]       dataRegroupBySew_7_8 = bufferStageEnqueueData_7[71:64];
  wire [7:0]       dataRegroupBySew_7_9 = bufferStageEnqueueData_7[79:72];
  wire [7:0]       dataRegroupBySew_7_10 = bufferStageEnqueueData_7[87:80];
  wire [7:0]       dataRegroupBySew_7_11 = bufferStageEnqueueData_7[95:88];
  wire [7:0]       dataRegroupBySew_7_12 = bufferStageEnqueueData_7[103:96];
  wire [7:0]       dataRegroupBySew_7_13 = bufferStageEnqueueData_7[111:104];
  wire [7:0]       dataRegroupBySew_7_14 = bufferStageEnqueueData_7[119:112];
  wire [7:0]       dataRegroupBySew_7_15 = bufferStageEnqueueData_7[127:120];
  wire [15:0]      dataInMem_lo_lo_lo = {dataRegroupBySew_0_1, dataRegroupBySew_0_0};
  wire [15:0]      dataInMem_lo_lo_hi = {dataRegroupBySew_0_3, dataRegroupBySew_0_2};
  wire [31:0]      dataInMem_lo_lo = {dataInMem_lo_lo_hi, dataInMem_lo_lo_lo};
  wire [15:0]      dataInMem_lo_hi_lo = {dataRegroupBySew_0_5, dataRegroupBySew_0_4};
  wire [15:0]      dataInMem_lo_hi_hi = {dataRegroupBySew_0_7, dataRegroupBySew_0_6};
  wire [31:0]      dataInMem_lo_hi = {dataInMem_lo_hi_hi, dataInMem_lo_hi_lo};
  wire [63:0]      dataInMem_lo = {dataInMem_lo_hi, dataInMem_lo_lo};
  wire [15:0]      dataInMem_hi_lo_lo = {dataRegroupBySew_0_9, dataRegroupBySew_0_8};
  wire [15:0]      dataInMem_hi_lo_hi = {dataRegroupBySew_0_11, dataRegroupBySew_0_10};
  wire [31:0]      dataInMem_hi_lo = {dataInMem_hi_lo_hi, dataInMem_hi_lo_lo};
  wire [15:0]      dataInMem_hi_hi_lo = {dataRegroupBySew_0_13, dataRegroupBySew_0_12};
  wire [15:0]      dataInMem_hi_hi_hi = {dataRegroupBySew_0_15, dataRegroupBySew_0_14};
  wire [31:0]      dataInMem_hi_hi = {dataInMem_hi_hi_hi, dataInMem_hi_hi_lo};
  wire [63:0]      dataInMem_hi = {dataInMem_hi_hi, dataInMem_hi_lo};
  wire [127:0]     dataInMem = {dataInMem_hi, dataInMem_lo};
  wire [127:0]     regroupCacheLine_0 = dataInMem;
  wire [127:0]     res = regroupCacheLine_0;
  wire [255:0]     lo_lo = {128'h0, res};
  wire [511:0]     lo = {256'h0, lo_lo};
  wire [1023:0]    regroupLoadData_0_0 = {512'h0, lo};
  wire [31:0]      dataInMem_lo_lo_lo_1 = {dataRegroupBySew_1_1, dataRegroupBySew_0_1, dataRegroupBySew_1_0, dataRegroupBySew_0_0};
  wire [31:0]      dataInMem_lo_lo_hi_1 = {dataRegroupBySew_1_3, dataRegroupBySew_0_3, dataRegroupBySew_1_2, dataRegroupBySew_0_2};
  wire [63:0]      dataInMem_lo_lo_1 = {dataInMem_lo_lo_hi_1, dataInMem_lo_lo_lo_1};
  wire [31:0]      dataInMem_lo_hi_lo_1 = {dataRegroupBySew_1_5, dataRegroupBySew_0_5, dataRegroupBySew_1_4, dataRegroupBySew_0_4};
  wire [31:0]      dataInMem_lo_hi_hi_1 = {dataRegroupBySew_1_7, dataRegroupBySew_0_7, dataRegroupBySew_1_6, dataRegroupBySew_0_6};
  wire [63:0]      dataInMem_lo_hi_1 = {dataInMem_lo_hi_hi_1, dataInMem_lo_hi_lo_1};
  wire [127:0]     dataInMem_lo_1 = {dataInMem_lo_hi_1, dataInMem_lo_lo_1};
  wire [31:0]      dataInMem_hi_lo_lo_1 = {dataRegroupBySew_1_9, dataRegroupBySew_0_9, dataRegroupBySew_1_8, dataRegroupBySew_0_8};
  wire [31:0]      dataInMem_hi_lo_hi_1 = {dataRegroupBySew_1_11, dataRegroupBySew_0_11, dataRegroupBySew_1_10, dataRegroupBySew_0_10};
  wire [63:0]      dataInMem_hi_lo_1 = {dataInMem_hi_lo_hi_1, dataInMem_hi_lo_lo_1};
  wire [31:0]      dataInMem_hi_hi_lo_1 = {dataRegroupBySew_1_13, dataRegroupBySew_0_13, dataRegroupBySew_1_12, dataRegroupBySew_0_12};
  wire [31:0]      dataInMem_hi_hi_hi_1 = {dataRegroupBySew_1_15, dataRegroupBySew_0_15, dataRegroupBySew_1_14, dataRegroupBySew_0_14};
  wire [63:0]      dataInMem_hi_hi_1 = {dataInMem_hi_hi_hi_1, dataInMem_hi_hi_lo_1};
  wire [127:0]     dataInMem_hi_1 = {dataInMem_hi_hi_1, dataInMem_hi_lo_1};
  wire [255:0]     dataInMem_1 = {dataInMem_hi_1, dataInMem_lo_1};
  wire [127:0]     regroupCacheLine_1_0 = dataInMem_1[127:0];
  wire [127:0]     regroupCacheLine_1_1 = dataInMem_1[255:128];
  wire [127:0]     res_8 = regroupCacheLine_1_0;
  wire [127:0]     res_9 = regroupCacheLine_1_1;
  wire [255:0]     lo_lo_1 = {res_9, res_8};
  wire [511:0]     lo_1 = {256'h0, lo_lo_1};
  wire [1023:0]    regroupLoadData_0_1 = {512'h0, lo_1};
  wire [15:0]      _GEN_3 = {dataRegroupBySew_2_0, dataRegroupBySew_1_0};
  wire [15:0]      dataInMem_hi_2;
  assign dataInMem_hi_2 = _GEN_3;
  wire [15:0]      dataInMem_lo_hi_5;
  assign dataInMem_lo_hi_5 = _GEN_3;
  wire [15:0]      dataInMem_lo_hi_22;
  assign dataInMem_lo_hi_22 = _GEN_3;
  wire [15:0]      _GEN_4 = {dataRegroupBySew_2_1, dataRegroupBySew_1_1};
  wire [15:0]      dataInMem_hi_3;
  assign dataInMem_hi_3 = _GEN_4;
  wire [15:0]      dataInMem_lo_hi_6;
  assign dataInMem_lo_hi_6 = _GEN_4;
  wire [15:0]      dataInMem_lo_hi_23;
  assign dataInMem_lo_hi_23 = _GEN_4;
  wire [15:0]      _GEN_5 = {dataRegroupBySew_2_2, dataRegroupBySew_1_2};
  wire [15:0]      dataInMem_hi_4;
  assign dataInMem_hi_4 = _GEN_5;
  wire [15:0]      dataInMem_lo_hi_7;
  assign dataInMem_lo_hi_7 = _GEN_5;
  wire [15:0]      dataInMem_lo_hi_24;
  assign dataInMem_lo_hi_24 = _GEN_5;
  wire [15:0]      _GEN_6 = {dataRegroupBySew_2_3, dataRegroupBySew_1_3};
  wire [15:0]      dataInMem_hi_5;
  assign dataInMem_hi_5 = _GEN_6;
  wire [15:0]      dataInMem_lo_hi_8;
  assign dataInMem_lo_hi_8 = _GEN_6;
  wire [15:0]      dataInMem_lo_hi_25;
  assign dataInMem_lo_hi_25 = _GEN_6;
  wire [15:0]      _GEN_7 = {dataRegroupBySew_2_4, dataRegroupBySew_1_4};
  wire [15:0]      dataInMem_hi_6;
  assign dataInMem_hi_6 = _GEN_7;
  wire [15:0]      dataInMem_lo_hi_9;
  assign dataInMem_lo_hi_9 = _GEN_7;
  wire [15:0]      dataInMem_lo_hi_26;
  assign dataInMem_lo_hi_26 = _GEN_7;
  wire [15:0]      _GEN_8 = {dataRegroupBySew_2_5, dataRegroupBySew_1_5};
  wire [15:0]      dataInMem_hi_7;
  assign dataInMem_hi_7 = _GEN_8;
  wire [15:0]      dataInMem_lo_hi_10;
  assign dataInMem_lo_hi_10 = _GEN_8;
  wire [15:0]      dataInMem_lo_hi_27;
  assign dataInMem_lo_hi_27 = _GEN_8;
  wire [15:0]      _GEN_9 = {dataRegroupBySew_2_6, dataRegroupBySew_1_6};
  wire [15:0]      dataInMem_hi_8;
  assign dataInMem_hi_8 = _GEN_9;
  wire [15:0]      dataInMem_lo_hi_11;
  assign dataInMem_lo_hi_11 = _GEN_9;
  wire [15:0]      dataInMem_lo_hi_28;
  assign dataInMem_lo_hi_28 = _GEN_9;
  wire [15:0]      _GEN_10 = {dataRegroupBySew_2_7, dataRegroupBySew_1_7};
  wire [15:0]      dataInMem_hi_9;
  assign dataInMem_hi_9 = _GEN_10;
  wire [15:0]      dataInMem_lo_hi_12;
  assign dataInMem_lo_hi_12 = _GEN_10;
  wire [15:0]      dataInMem_lo_hi_29;
  assign dataInMem_lo_hi_29 = _GEN_10;
  wire [15:0]      _GEN_11 = {dataRegroupBySew_2_8, dataRegroupBySew_1_8};
  wire [15:0]      dataInMem_hi_10;
  assign dataInMem_hi_10 = _GEN_11;
  wire [15:0]      dataInMem_lo_hi_13;
  assign dataInMem_lo_hi_13 = _GEN_11;
  wire [15:0]      dataInMem_lo_hi_30;
  assign dataInMem_lo_hi_30 = _GEN_11;
  wire [15:0]      _GEN_12 = {dataRegroupBySew_2_9, dataRegroupBySew_1_9};
  wire [15:0]      dataInMem_hi_11;
  assign dataInMem_hi_11 = _GEN_12;
  wire [15:0]      dataInMem_lo_hi_14;
  assign dataInMem_lo_hi_14 = _GEN_12;
  wire [15:0]      dataInMem_lo_hi_31;
  assign dataInMem_lo_hi_31 = _GEN_12;
  wire [15:0]      _GEN_13 = {dataRegroupBySew_2_10, dataRegroupBySew_1_10};
  wire [15:0]      dataInMem_hi_12;
  assign dataInMem_hi_12 = _GEN_13;
  wire [15:0]      dataInMem_lo_hi_15;
  assign dataInMem_lo_hi_15 = _GEN_13;
  wire [15:0]      dataInMem_lo_hi_32;
  assign dataInMem_lo_hi_32 = _GEN_13;
  wire [15:0]      _GEN_14 = {dataRegroupBySew_2_11, dataRegroupBySew_1_11};
  wire [15:0]      dataInMem_hi_13;
  assign dataInMem_hi_13 = _GEN_14;
  wire [15:0]      dataInMem_lo_hi_16;
  assign dataInMem_lo_hi_16 = _GEN_14;
  wire [15:0]      dataInMem_lo_hi_33;
  assign dataInMem_lo_hi_33 = _GEN_14;
  wire [15:0]      _GEN_15 = {dataRegroupBySew_2_12, dataRegroupBySew_1_12};
  wire [15:0]      dataInMem_hi_14;
  assign dataInMem_hi_14 = _GEN_15;
  wire [15:0]      dataInMem_lo_hi_17;
  assign dataInMem_lo_hi_17 = _GEN_15;
  wire [15:0]      dataInMem_lo_hi_34;
  assign dataInMem_lo_hi_34 = _GEN_15;
  wire [15:0]      _GEN_16 = {dataRegroupBySew_2_13, dataRegroupBySew_1_13};
  wire [15:0]      dataInMem_hi_15;
  assign dataInMem_hi_15 = _GEN_16;
  wire [15:0]      dataInMem_lo_hi_18;
  assign dataInMem_lo_hi_18 = _GEN_16;
  wire [15:0]      dataInMem_lo_hi_35;
  assign dataInMem_lo_hi_35 = _GEN_16;
  wire [15:0]      _GEN_17 = {dataRegroupBySew_2_14, dataRegroupBySew_1_14};
  wire [15:0]      dataInMem_hi_16;
  assign dataInMem_hi_16 = _GEN_17;
  wire [15:0]      dataInMem_lo_hi_19;
  assign dataInMem_lo_hi_19 = _GEN_17;
  wire [15:0]      dataInMem_lo_hi_36;
  assign dataInMem_lo_hi_36 = _GEN_17;
  wire [15:0]      _GEN_18 = {dataRegroupBySew_2_15, dataRegroupBySew_1_15};
  wire [15:0]      dataInMem_hi_17;
  assign dataInMem_hi_17 = _GEN_18;
  wire [15:0]      dataInMem_lo_hi_20;
  assign dataInMem_lo_hi_20 = _GEN_18;
  wire [15:0]      dataInMem_lo_hi_37;
  assign dataInMem_lo_hi_37 = _GEN_18;
  wire [47:0]      dataInMem_lo_lo_lo_2 = {dataInMem_hi_3, dataRegroupBySew_0_1, dataInMem_hi_2, dataRegroupBySew_0_0};
  wire [47:0]      dataInMem_lo_lo_hi_2 = {dataInMem_hi_5, dataRegroupBySew_0_3, dataInMem_hi_4, dataRegroupBySew_0_2};
  wire [95:0]      dataInMem_lo_lo_2 = {dataInMem_lo_lo_hi_2, dataInMem_lo_lo_lo_2};
  wire [47:0]      dataInMem_lo_hi_lo_2 = {dataInMem_hi_7, dataRegroupBySew_0_5, dataInMem_hi_6, dataRegroupBySew_0_4};
  wire [47:0]      dataInMem_lo_hi_hi_2 = {dataInMem_hi_9, dataRegroupBySew_0_7, dataInMem_hi_8, dataRegroupBySew_0_6};
  wire [95:0]      dataInMem_lo_hi_2 = {dataInMem_lo_hi_hi_2, dataInMem_lo_hi_lo_2};
  wire [191:0]     dataInMem_lo_2 = {dataInMem_lo_hi_2, dataInMem_lo_lo_2};
  wire [47:0]      dataInMem_hi_lo_lo_2 = {dataInMem_hi_11, dataRegroupBySew_0_9, dataInMem_hi_10, dataRegroupBySew_0_8};
  wire [47:0]      dataInMem_hi_lo_hi_2 = {dataInMem_hi_13, dataRegroupBySew_0_11, dataInMem_hi_12, dataRegroupBySew_0_10};
  wire [95:0]      dataInMem_hi_lo_2 = {dataInMem_hi_lo_hi_2, dataInMem_hi_lo_lo_2};
  wire [47:0]      dataInMem_hi_hi_lo_2 = {dataInMem_hi_15, dataRegroupBySew_0_13, dataInMem_hi_14, dataRegroupBySew_0_12};
  wire [47:0]      dataInMem_hi_hi_hi_2 = {dataInMem_hi_17, dataRegroupBySew_0_15, dataInMem_hi_16, dataRegroupBySew_0_14};
  wire [95:0]      dataInMem_hi_hi_2 = {dataInMem_hi_hi_hi_2, dataInMem_hi_hi_lo_2};
  wire [191:0]     dataInMem_hi_18 = {dataInMem_hi_hi_2, dataInMem_hi_lo_2};
  wire [383:0]     dataInMem_2 = {dataInMem_hi_18, dataInMem_lo_2};
  wire [127:0]     regroupCacheLine_2_0 = dataInMem_2[127:0];
  wire [127:0]     regroupCacheLine_2_1 = dataInMem_2[255:128];
  wire [127:0]     regroupCacheLine_2_2 = dataInMem_2[383:256];
  wire [127:0]     res_16 = regroupCacheLine_2_0;
  wire [127:0]     res_17 = regroupCacheLine_2_1;
  wire [127:0]     res_18 = regroupCacheLine_2_2;
  wire [255:0]     lo_lo_2 = {res_17, res_16};
  wire [255:0]     lo_hi_2 = {128'h0, res_18};
  wire [511:0]     lo_2 = {lo_hi_2, lo_lo_2};
  wire [1023:0]    regroupLoadData_0_2 = {512'h0, lo_2};
  wire [15:0]      _GEN_19 = {dataRegroupBySew_1_0, dataRegroupBySew_0_0};
  wire [15:0]      dataInMem_lo_3;
  assign dataInMem_lo_3 = _GEN_19;
  wire [15:0]      dataInMem_lo_20;
  assign dataInMem_lo_20 = _GEN_19;
  wire [15:0]      dataInMem_lo_lo_7;
  assign dataInMem_lo_lo_7 = _GEN_19;
  wire [15:0]      _GEN_20 = {dataRegroupBySew_3_0, dataRegroupBySew_2_0};
  wire [15:0]      dataInMem_hi_19;
  assign dataInMem_hi_19 = _GEN_20;
  wire [15:0]      dataInMem_lo_hi_39;
  assign dataInMem_lo_hi_39 = _GEN_20;
  wire [15:0]      _GEN_21 = {dataRegroupBySew_1_1, dataRegroupBySew_0_1};
  wire [15:0]      dataInMem_lo_4;
  assign dataInMem_lo_4 = _GEN_21;
  wire [15:0]      dataInMem_lo_21;
  assign dataInMem_lo_21 = _GEN_21;
  wire [15:0]      dataInMem_lo_lo_8;
  assign dataInMem_lo_lo_8 = _GEN_21;
  wire [15:0]      _GEN_22 = {dataRegroupBySew_3_1, dataRegroupBySew_2_1};
  wire [15:0]      dataInMem_hi_20;
  assign dataInMem_hi_20 = _GEN_22;
  wire [15:0]      dataInMem_lo_hi_40;
  assign dataInMem_lo_hi_40 = _GEN_22;
  wire [15:0]      _GEN_23 = {dataRegroupBySew_1_2, dataRegroupBySew_0_2};
  wire [15:0]      dataInMem_lo_5;
  assign dataInMem_lo_5 = _GEN_23;
  wire [15:0]      dataInMem_lo_22;
  assign dataInMem_lo_22 = _GEN_23;
  wire [15:0]      dataInMem_lo_lo_9;
  assign dataInMem_lo_lo_9 = _GEN_23;
  wire [15:0]      _GEN_24 = {dataRegroupBySew_3_2, dataRegroupBySew_2_2};
  wire [15:0]      dataInMem_hi_21;
  assign dataInMem_hi_21 = _GEN_24;
  wire [15:0]      dataInMem_lo_hi_41;
  assign dataInMem_lo_hi_41 = _GEN_24;
  wire [15:0]      _GEN_25 = {dataRegroupBySew_1_3, dataRegroupBySew_0_3};
  wire [15:0]      dataInMem_lo_6;
  assign dataInMem_lo_6 = _GEN_25;
  wire [15:0]      dataInMem_lo_23;
  assign dataInMem_lo_23 = _GEN_25;
  wire [15:0]      dataInMem_lo_lo_10;
  assign dataInMem_lo_lo_10 = _GEN_25;
  wire [15:0]      _GEN_26 = {dataRegroupBySew_3_3, dataRegroupBySew_2_3};
  wire [15:0]      dataInMem_hi_22;
  assign dataInMem_hi_22 = _GEN_26;
  wire [15:0]      dataInMem_lo_hi_42;
  assign dataInMem_lo_hi_42 = _GEN_26;
  wire [15:0]      _GEN_27 = {dataRegroupBySew_1_4, dataRegroupBySew_0_4};
  wire [15:0]      dataInMem_lo_7;
  assign dataInMem_lo_7 = _GEN_27;
  wire [15:0]      dataInMem_lo_24;
  assign dataInMem_lo_24 = _GEN_27;
  wire [15:0]      dataInMem_lo_lo_11;
  assign dataInMem_lo_lo_11 = _GEN_27;
  wire [15:0]      _GEN_28 = {dataRegroupBySew_3_4, dataRegroupBySew_2_4};
  wire [15:0]      dataInMem_hi_23;
  assign dataInMem_hi_23 = _GEN_28;
  wire [15:0]      dataInMem_lo_hi_43;
  assign dataInMem_lo_hi_43 = _GEN_28;
  wire [15:0]      _GEN_29 = {dataRegroupBySew_1_5, dataRegroupBySew_0_5};
  wire [15:0]      dataInMem_lo_8;
  assign dataInMem_lo_8 = _GEN_29;
  wire [15:0]      dataInMem_lo_25;
  assign dataInMem_lo_25 = _GEN_29;
  wire [15:0]      dataInMem_lo_lo_12;
  assign dataInMem_lo_lo_12 = _GEN_29;
  wire [15:0]      _GEN_30 = {dataRegroupBySew_3_5, dataRegroupBySew_2_5};
  wire [15:0]      dataInMem_hi_24;
  assign dataInMem_hi_24 = _GEN_30;
  wire [15:0]      dataInMem_lo_hi_44;
  assign dataInMem_lo_hi_44 = _GEN_30;
  wire [15:0]      _GEN_31 = {dataRegroupBySew_1_6, dataRegroupBySew_0_6};
  wire [15:0]      dataInMem_lo_9;
  assign dataInMem_lo_9 = _GEN_31;
  wire [15:0]      dataInMem_lo_26;
  assign dataInMem_lo_26 = _GEN_31;
  wire [15:0]      dataInMem_lo_lo_13;
  assign dataInMem_lo_lo_13 = _GEN_31;
  wire [15:0]      _GEN_32 = {dataRegroupBySew_3_6, dataRegroupBySew_2_6};
  wire [15:0]      dataInMem_hi_25;
  assign dataInMem_hi_25 = _GEN_32;
  wire [15:0]      dataInMem_lo_hi_45;
  assign dataInMem_lo_hi_45 = _GEN_32;
  wire [15:0]      _GEN_33 = {dataRegroupBySew_1_7, dataRegroupBySew_0_7};
  wire [15:0]      dataInMem_lo_10;
  assign dataInMem_lo_10 = _GEN_33;
  wire [15:0]      dataInMem_lo_27;
  assign dataInMem_lo_27 = _GEN_33;
  wire [15:0]      dataInMem_lo_lo_14;
  assign dataInMem_lo_lo_14 = _GEN_33;
  wire [15:0]      _GEN_34 = {dataRegroupBySew_3_7, dataRegroupBySew_2_7};
  wire [15:0]      dataInMem_hi_26;
  assign dataInMem_hi_26 = _GEN_34;
  wire [15:0]      dataInMem_lo_hi_46;
  assign dataInMem_lo_hi_46 = _GEN_34;
  wire [15:0]      _GEN_35 = {dataRegroupBySew_1_8, dataRegroupBySew_0_8};
  wire [15:0]      dataInMem_lo_11;
  assign dataInMem_lo_11 = _GEN_35;
  wire [15:0]      dataInMem_lo_28;
  assign dataInMem_lo_28 = _GEN_35;
  wire [15:0]      dataInMem_lo_lo_15;
  assign dataInMem_lo_lo_15 = _GEN_35;
  wire [15:0]      _GEN_36 = {dataRegroupBySew_3_8, dataRegroupBySew_2_8};
  wire [15:0]      dataInMem_hi_27;
  assign dataInMem_hi_27 = _GEN_36;
  wire [15:0]      dataInMem_lo_hi_47;
  assign dataInMem_lo_hi_47 = _GEN_36;
  wire [15:0]      _GEN_37 = {dataRegroupBySew_1_9, dataRegroupBySew_0_9};
  wire [15:0]      dataInMem_lo_12;
  assign dataInMem_lo_12 = _GEN_37;
  wire [15:0]      dataInMem_lo_29;
  assign dataInMem_lo_29 = _GEN_37;
  wire [15:0]      dataInMem_lo_lo_16;
  assign dataInMem_lo_lo_16 = _GEN_37;
  wire [15:0]      _GEN_38 = {dataRegroupBySew_3_9, dataRegroupBySew_2_9};
  wire [15:0]      dataInMem_hi_28;
  assign dataInMem_hi_28 = _GEN_38;
  wire [15:0]      dataInMem_lo_hi_48;
  assign dataInMem_lo_hi_48 = _GEN_38;
  wire [15:0]      _GEN_39 = {dataRegroupBySew_1_10, dataRegroupBySew_0_10};
  wire [15:0]      dataInMem_lo_13;
  assign dataInMem_lo_13 = _GEN_39;
  wire [15:0]      dataInMem_lo_30;
  assign dataInMem_lo_30 = _GEN_39;
  wire [15:0]      dataInMem_lo_lo_17;
  assign dataInMem_lo_lo_17 = _GEN_39;
  wire [15:0]      _GEN_40 = {dataRegroupBySew_3_10, dataRegroupBySew_2_10};
  wire [15:0]      dataInMem_hi_29;
  assign dataInMem_hi_29 = _GEN_40;
  wire [15:0]      dataInMem_lo_hi_49;
  assign dataInMem_lo_hi_49 = _GEN_40;
  wire [15:0]      _GEN_41 = {dataRegroupBySew_1_11, dataRegroupBySew_0_11};
  wire [15:0]      dataInMem_lo_14;
  assign dataInMem_lo_14 = _GEN_41;
  wire [15:0]      dataInMem_lo_31;
  assign dataInMem_lo_31 = _GEN_41;
  wire [15:0]      dataInMem_lo_lo_18;
  assign dataInMem_lo_lo_18 = _GEN_41;
  wire [15:0]      _GEN_42 = {dataRegroupBySew_3_11, dataRegroupBySew_2_11};
  wire [15:0]      dataInMem_hi_30;
  assign dataInMem_hi_30 = _GEN_42;
  wire [15:0]      dataInMem_lo_hi_50;
  assign dataInMem_lo_hi_50 = _GEN_42;
  wire [15:0]      _GEN_43 = {dataRegroupBySew_1_12, dataRegroupBySew_0_12};
  wire [15:0]      dataInMem_lo_15;
  assign dataInMem_lo_15 = _GEN_43;
  wire [15:0]      dataInMem_lo_32;
  assign dataInMem_lo_32 = _GEN_43;
  wire [15:0]      dataInMem_lo_lo_19;
  assign dataInMem_lo_lo_19 = _GEN_43;
  wire [15:0]      _GEN_44 = {dataRegroupBySew_3_12, dataRegroupBySew_2_12};
  wire [15:0]      dataInMem_hi_31;
  assign dataInMem_hi_31 = _GEN_44;
  wire [15:0]      dataInMem_lo_hi_51;
  assign dataInMem_lo_hi_51 = _GEN_44;
  wire [15:0]      _GEN_45 = {dataRegroupBySew_1_13, dataRegroupBySew_0_13};
  wire [15:0]      dataInMem_lo_16;
  assign dataInMem_lo_16 = _GEN_45;
  wire [15:0]      dataInMem_lo_33;
  assign dataInMem_lo_33 = _GEN_45;
  wire [15:0]      dataInMem_lo_lo_20;
  assign dataInMem_lo_lo_20 = _GEN_45;
  wire [15:0]      _GEN_46 = {dataRegroupBySew_3_13, dataRegroupBySew_2_13};
  wire [15:0]      dataInMem_hi_32;
  assign dataInMem_hi_32 = _GEN_46;
  wire [15:0]      dataInMem_lo_hi_52;
  assign dataInMem_lo_hi_52 = _GEN_46;
  wire [15:0]      _GEN_47 = {dataRegroupBySew_1_14, dataRegroupBySew_0_14};
  wire [15:0]      dataInMem_lo_17;
  assign dataInMem_lo_17 = _GEN_47;
  wire [15:0]      dataInMem_lo_34;
  assign dataInMem_lo_34 = _GEN_47;
  wire [15:0]      dataInMem_lo_lo_21;
  assign dataInMem_lo_lo_21 = _GEN_47;
  wire [15:0]      _GEN_48 = {dataRegroupBySew_3_14, dataRegroupBySew_2_14};
  wire [15:0]      dataInMem_hi_33;
  assign dataInMem_hi_33 = _GEN_48;
  wire [15:0]      dataInMem_lo_hi_53;
  assign dataInMem_lo_hi_53 = _GEN_48;
  wire [15:0]      _GEN_49 = {dataRegroupBySew_1_15, dataRegroupBySew_0_15};
  wire [15:0]      dataInMem_lo_18;
  assign dataInMem_lo_18 = _GEN_49;
  wire [15:0]      dataInMem_lo_35;
  assign dataInMem_lo_35 = _GEN_49;
  wire [15:0]      dataInMem_lo_lo_22;
  assign dataInMem_lo_lo_22 = _GEN_49;
  wire [15:0]      _GEN_50 = {dataRegroupBySew_3_15, dataRegroupBySew_2_15};
  wire [15:0]      dataInMem_hi_34;
  assign dataInMem_hi_34 = _GEN_50;
  wire [15:0]      dataInMem_lo_hi_54;
  assign dataInMem_lo_hi_54 = _GEN_50;
  wire [63:0]      dataInMem_lo_lo_lo_3 = {dataInMem_hi_20, dataInMem_lo_4, dataInMem_hi_19, dataInMem_lo_3};
  wire [63:0]      dataInMem_lo_lo_hi_3 = {dataInMem_hi_22, dataInMem_lo_6, dataInMem_hi_21, dataInMem_lo_5};
  wire [127:0]     dataInMem_lo_lo_3 = {dataInMem_lo_lo_hi_3, dataInMem_lo_lo_lo_3};
  wire [63:0]      dataInMem_lo_hi_lo_3 = {dataInMem_hi_24, dataInMem_lo_8, dataInMem_hi_23, dataInMem_lo_7};
  wire [63:0]      dataInMem_lo_hi_hi_3 = {dataInMem_hi_26, dataInMem_lo_10, dataInMem_hi_25, dataInMem_lo_9};
  wire [127:0]     dataInMem_lo_hi_3 = {dataInMem_lo_hi_hi_3, dataInMem_lo_hi_lo_3};
  wire [255:0]     dataInMem_lo_19 = {dataInMem_lo_hi_3, dataInMem_lo_lo_3};
  wire [63:0]      dataInMem_hi_lo_lo_3 = {dataInMem_hi_28, dataInMem_lo_12, dataInMem_hi_27, dataInMem_lo_11};
  wire [63:0]      dataInMem_hi_lo_hi_3 = {dataInMem_hi_30, dataInMem_lo_14, dataInMem_hi_29, dataInMem_lo_13};
  wire [127:0]     dataInMem_hi_lo_3 = {dataInMem_hi_lo_hi_3, dataInMem_hi_lo_lo_3};
  wire [63:0]      dataInMem_hi_hi_lo_3 = {dataInMem_hi_32, dataInMem_lo_16, dataInMem_hi_31, dataInMem_lo_15};
  wire [63:0]      dataInMem_hi_hi_hi_3 = {dataInMem_hi_34, dataInMem_lo_18, dataInMem_hi_33, dataInMem_lo_17};
  wire [127:0]     dataInMem_hi_hi_3 = {dataInMem_hi_hi_hi_3, dataInMem_hi_hi_lo_3};
  wire [255:0]     dataInMem_hi_35 = {dataInMem_hi_hi_3, dataInMem_hi_lo_3};
  wire [511:0]     dataInMem_3 = {dataInMem_hi_35, dataInMem_lo_19};
  wire [127:0]     regroupCacheLine_3_0 = dataInMem_3[127:0];
  wire [127:0]     regroupCacheLine_3_1 = dataInMem_3[255:128];
  wire [127:0]     regroupCacheLine_3_2 = dataInMem_3[383:256];
  wire [127:0]     regroupCacheLine_3_3 = dataInMem_3[511:384];
  wire [127:0]     res_24 = regroupCacheLine_3_0;
  wire [127:0]     res_25 = regroupCacheLine_3_1;
  wire [127:0]     res_26 = regroupCacheLine_3_2;
  wire [127:0]     res_27 = regroupCacheLine_3_3;
  wire [255:0]     lo_lo_3 = {res_25, res_24};
  wire [255:0]     lo_hi_3 = {res_27, res_26};
  wire [511:0]     lo_3 = {lo_hi_3, lo_lo_3};
  wire [1023:0]    regroupLoadData_0_3 = {512'h0, lo_3};
  wire [15:0]      _GEN_51 = {dataRegroupBySew_4_0, dataRegroupBySew_3_0};
  wire [15:0]      dataInMem_hi_hi_4;
  assign dataInMem_hi_hi_4 = _GEN_51;
  wire [15:0]      dataInMem_hi_lo_6;
  assign dataInMem_hi_lo_6 = _GEN_51;
  wire [23:0]      dataInMem_hi_36 = {dataInMem_hi_hi_4, dataRegroupBySew_2_0};
  wire [15:0]      _GEN_52 = {dataRegroupBySew_4_1, dataRegroupBySew_3_1};
  wire [15:0]      dataInMem_hi_hi_5;
  assign dataInMem_hi_hi_5 = _GEN_52;
  wire [15:0]      dataInMem_hi_lo_7;
  assign dataInMem_hi_lo_7 = _GEN_52;
  wire [23:0]      dataInMem_hi_37 = {dataInMem_hi_hi_5, dataRegroupBySew_2_1};
  wire [15:0]      _GEN_53 = {dataRegroupBySew_4_2, dataRegroupBySew_3_2};
  wire [15:0]      dataInMem_hi_hi_6;
  assign dataInMem_hi_hi_6 = _GEN_53;
  wire [15:0]      dataInMem_hi_lo_8;
  assign dataInMem_hi_lo_8 = _GEN_53;
  wire [23:0]      dataInMem_hi_38 = {dataInMem_hi_hi_6, dataRegroupBySew_2_2};
  wire [15:0]      _GEN_54 = {dataRegroupBySew_4_3, dataRegroupBySew_3_3};
  wire [15:0]      dataInMem_hi_hi_7;
  assign dataInMem_hi_hi_7 = _GEN_54;
  wire [15:0]      dataInMem_hi_lo_9;
  assign dataInMem_hi_lo_9 = _GEN_54;
  wire [23:0]      dataInMem_hi_39 = {dataInMem_hi_hi_7, dataRegroupBySew_2_3};
  wire [15:0]      _GEN_55 = {dataRegroupBySew_4_4, dataRegroupBySew_3_4};
  wire [15:0]      dataInMem_hi_hi_8;
  assign dataInMem_hi_hi_8 = _GEN_55;
  wire [15:0]      dataInMem_hi_lo_10;
  assign dataInMem_hi_lo_10 = _GEN_55;
  wire [23:0]      dataInMem_hi_40 = {dataInMem_hi_hi_8, dataRegroupBySew_2_4};
  wire [15:0]      _GEN_56 = {dataRegroupBySew_4_5, dataRegroupBySew_3_5};
  wire [15:0]      dataInMem_hi_hi_9;
  assign dataInMem_hi_hi_9 = _GEN_56;
  wire [15:0]      dataInMem_hi_lo_11;
  assign dataInMem_hi_lo_11 = _GEN_56;
  wire [23:0]      dataInMem_hi_41 = {dataInMem_hi_hi_9, dataRegroupBySew_2_5};
  wire [15:0]      _GEN_57 = {dataRegroupBySew_4_6, dataRegroupBySew_3_6};
  wire [15:0]      dataInMem_hi_hi_10;
  assign dataInMem_hi_hi_10 = _GEN_57;
  wire [15:0]      dataInMem_hi_lo_12;
  assign dataInMem_hi_lo_12 = _GEN_57;
  wire [23:0]      dataInMem_hi_42 = {dataInMem_hi_hi_10, dataRegroupBySew_2_6};
  wire [15:0]      _GEN_58 = {dataRegroupBySew_4_7, dataRegroupBySew_3_7};
  wire [15:0]      dataInMem_hi_hi_11;
  assign dataInMem_hi_hi_11 = _GEN_58;
  wire [15:0]      dataInMem_hi_lo_13;
  assign dataInMem_hi_lo_13 = _GEN_58;
  wire [23:0]      dataInMem_hi_43 = {dataInMem_hi_hi_11, dataRegroupBySew_2_7};
  wire [15:0]      _GEN_59 = {dataRegroupBySew_4_8, dataRegroupBySew_3_8};
  wire [15:0]      dataInMem_hi_hi_12;
  assign dataInMem_hi_hi_12 = _GEN_59;
  wire [15:0]      dataInMem_hi_lo_14;
  assign dataInMem_hi_lo_14 = _GEN_59;
  wire [23:0]      dataInMem_hi_44 = {dataInMem_hi_hi_12, dataRegroupBySew_2_8};
  wire [15:0]      _GEN_60 = {dataRegroupBySew_4_9, dataRegroupBySew_3_9};
  wire [15:0]      dataInMem_hi_hi_13;
  assign dataInMem_hi_hi_13 = _GEN_60;
  wire [15:0]      dataInMem_hi_lo_15;
  assign dataInMem_hi_lo_15 = _GEN_60;
  wire [23:0]      dataInMem_hi_45 = {dataInMem_hi_hi_13, dataRegroupBySew_2_9};
  wire [15:0]      _GEN_61 = {dataRegroupBySew_4_10, dataRegroupBySew_3_10};
  wire [15:0]      dataInMem_hi_hi_14;
  assign dataInMem_hi_hi_14 = _GEN_61;
  wire [15:0]      dataInMem_hi_lo_16;
  assign dataInMem_hi_lo_16 = _GEN_61;
  wire [23:0]      dataInMem_hi_46 = {dataInMem_hi_hi_14, dataRegroupBySew_2_10};
  wire [15:0]      _GEN_62 = {dataRegroupBySew_4_11, dataRegroupBySew_3_11};
  wire [15:0]      dataInMem_hi_hi_15;
  assign dataInMem_hi_hi_15 = _GEN_62;
  wire [15:0]      dataInMem_hi_lo_17;
  assign dataInMem_hi_lo_17 = _GEN_62;
  wire [23:0]      dataInMem_hi_47 = {dataInMem_hi_hi_15, dataRegroupBySew_2_11};
  wire [15:0]      _GEN_63 = {dataRegroupBySew_4_12, dataRegroupBySew_3_12};
  wire [15:0]      dataInMem_hi_hi_16;
  assign dataInMem_hi_hi_16 = _GEN_63;
  wire [15:0]      dataInMem_hi_lo_18;
  assign dataInMem_hi_lo_18 = _GEN_63;
  wire [23:0]      dataInMem_hi_48 = {dataInMem_hi_hi_16, dataRegroupBySew_2_12};
  wire [15:0]      _GEN_64 = {dataRegroupBySew_4_13, dataRegroupBySew_3_13};
  wire [15:0]      dataInMem_hi_hi_17;
  assign dataInMem_hi_hi_17 = _GEN_64;
  wire [15:0]      dataInMem_hi_lo_19;
  assign dataInMem_hi_lo_19 = _GEN_64;
  wire [23:0]      dataInMem_hi_49 = {dataInMem_hi_hi_17, dataRegroupBySew_2_13};
  wire [15:0]      _GEN_65 = {dataRegroupBySew_4_14, dataRegroupBySew_3_14};
  wire [15:0]      dataInMem_hi_hi_18;
  assign dataInMem_hi_hi_18 = _GEN_65;
  wire [15:0]      dataInMem_hi_lo_20;
  assign dataInMem_hi_lo_20 = _GEN_65;
  wire [23:0]      dataInMem_hi_50 = {dataInMem_hi_hi_18, dataRegroupBySew_2_14};
  wire [15:0]      _GEN_66 = {dataRegroupBySew_4_15, dataRegroupBySew_3_15};
  wire [15:0]      dataInMem_hi_hi_19;
  assign dataInMem_hi_hi_19 = _GEN_66;
  wire [15:0]      dataInMem_hi_lo_21;
  assign dataInMem_hi_lo_21 = _GEN_66;
  wire [23:0]      dataInMem_hi_51 = {dataInMem_hi_hi_19, dataRegroupBySew_2_15};
  wire [79:0]      dataInMem_lo_lo_lo_4 = {dataInMem_hi_37, dataInMem_lo_21, dataInMem_hi_36, dataInMem_lo_20};
  wire [79:0]      dataInMem_lo_lo_hi_4 = {dataInMem_hi_39, dataInMem_lo_23, dataInMem_hi_38, dataInMem_lo_22};
  wire [159:0]     dataInMem_lo_lo_4 = {dataInMem_lo_lo_hi_4, dataInMem_lo_lo_lo_4};
  wire [79:0]      dataInMem_lo_hi_lo_4 = {dataInMem_hi_41, dataInMem_lo_25, dataInMem_hi_40, dataInMem_lo_24};
  wire [79:0]      dataInMem_lo_hi_hi_4 = {dataInMem_hi_43, dataInMem_lo_27, dataInMem_hi_42, dataInMem_lo_26};
  wire [159:0]     dataInMem_lo_hi_4 = {dataInMem_lo_hi_hi_4, dataInMem_lo_hi_lo_4};
  wire [319:0]     dataInMem_lo_36 = {dataInMem_lo_hi_4, dataInMem_lo_lo_4};
  wire [79:0]      dataInMem_hi_lo_lo_4 = {dataInMem_hi_45, dataInMem_lo_29, dataInMem_hi_44, dataInMem_lo_28};
  wire [79:0]      dataInMem_hi_lo_hi_4 = {dataInMem_hi_47, dataInMem_lo_31, dataInMem_hi_46, dataInMem_lo_30};
  wire [159:0]     dataInMem_hi_lo_4 = {dataInMem_hi_lo_hi_4, dataInMem_hi_lo_lo_4};
  wire [79:0]      dataInMem_hi_hi_lo_4 = {dataInMem_hi_49, dataInMem_lo_33, dataInMem_hi_48, dataInMem_lo_32};
  wire [79:0]      dataInMem_hi_hi_hi_4 = {dataInMem_hi_51, dataInMem_lo_35, dataInMem_hi_50, dataInMem_lo_34};
  wire [159:0]     dataInMem_hi_hi_20 = {dataInMem_hi_hi_hi_4, dataInMem_hi_hi_lo_4};
  wire [319:0]     dataInMem_hi_52 = {dataInMem_hi_hi_20, dataInMem_hi_lo_4};
  wire [639:0]     dataInMem_4 = {dataInMem_hi_52, dataInMem_lo_36};
  wire [127:0]     regroupCacheLine_4_0 = dataInMem_4[127:0];
  wire [127:0]     regroupCacheLine_4_1 = dataInMem_4[255:128];
  wire [127:0]     regroupCacheLine_4_2 = dataInMem_4[383:256];
  wire [127:0]     regroupCacheLine_4_3 = dataInMem_4[511:384];
  wire [127:0]     regroupCacheLine_4_4 = dataInMem_4[639:512];
  wire [127:0]     res_32 = regroupCacheLine_4_0;
  wire [127:0]     res_33 = regroupCacheLine_4_1;
  wire [127:0]     res_34 = regroupCacheLine_4_2;
  wire [127:0]     res_35 = regroupCacheLine_4_3;
  wire [127:0]     res_36 = regroupCacheLine_4_4;
  wire [255:0]     lo_lo_4 = {res_33, res_32};
  wire [255:0]     lo_hi_4 = {res_35, res_34};
  wire [511:0]     lo_4 = {lo_hi_4, lo_lo_4};
  wire [255:0]     hi_lo_4 = {128'h0, res_36};
  wire [511:0]     hi_4 = {256'h0, hi_lo_4};
  wire [1023:0]    regroupLoadData_0_4 = {hi_4, lo_4};
  wire [23:0]      dataInMem_lo_37 = {dataInMem_lo_hi_5, dataRegroupBySew_0_0};
  wire [15:0]      _GEN_67 = {dataRegroupBySew_5_0, dataRegroupBySew_4_0};
  wire [15:0]      dataInMem_hi_hi_21;
  assign dataInMem_hi_hi_21 = _GEN_67;
  wire [15:0]      dataInMem_hi_lo_23;
  assign dataInMem_hi_lo_23 = _GEN_67;
  wire [23:0]      dataInMem_hi_53 = {dataInMem_hi_hi_21, dataRegroupBySew_3_0};
  wire [23:0]      dataInMem_lo_38 = {dataInMem_lo_hi_6, dataRegroupBySew_0_1};
  wire [15:0]      _GEN_68 = {dataRegroupBySew_5_1, dataRegroupBySew_4_1};
  wire [15:0]      dataInMem_hi_hi_22;
  assign dataInMem_hi_hi_22 = _GEN_68;
  wire [15:0]      dataInMem_hi_lo_24;
  assign dataInMem_hi_lo_24 = _GEN_68;
  wire [23:0]      dataInMem_hi_54 = {dataInMem_hi_hi_22, dataRegroupBySew_3_1};
  wire [23:0]      dataInMem_lo_39 = {dataInMem_lo_hi_7, dataRegroupBySew_0_2};
  wire [15:0]      _GEN_69 = {dataRegroupBySew_5_2, dataRegroupBySew_4_2};
  wire [15:0]      dataInMem_hi_hi_23;
  assign dataInMem_hi_hi_23 = _GEN_69;
  wire [15:0]      dataInMem_hi_lo_25;
  assign dataInMem_hi_lo_25 = _GEN_69;
  wire [23:0]      dataInMem_hi_55 = {dataInMem_hi_hi_23, dataRegroupBySew_3_2};
  wire [23:0]      dataInMem_lo_40 = {dataInMem_lo_hi_8, dataRegroupBySew_0_3};
  wire [15:0]      _GEN_70 = {dataRegroupBySew_5_3, dataRegroupBySew_4_3};
  wire [15:0]      dataInMem_hi_hi_24;
  assign dataInMem_hi_hi_24 = _GEN_70;
  wire [15:0]      dataInMem_hi_lo_26;
  assign dataInMem_hi_lo_26 = _GEN_70;
  wire [23:0]      dataInMem_hi_56 = {dataInMem_hi_hi_24, dataRegroupBySew_3_3};
  wire [23:0]      dataInMem_lo_41 = {dataInMem_lo_hi_9, dataRegroupBySew_0_4};
  wire [15:0]      _GEN_71 = {dataRegroupBySew_5_4, dataRegroupBySew_4_4};
  wire [15:0]      dataInMem_hi_hi_25;
  assign dataInMem_hi_hi_25 = _GEN_71;
  wire [15:0]      dataInMem_hi_lo_27;
  assign dataInMem_hi_lo_27 = _GEN_71;
  wire [23:0]      dataInMem_hi_57 = {dataInMem_hi_hi_25, dataRegroupBySew_3_4};
  wire [23:0]      dataInMem_lo_42 = {dataInMem_lo_hi_10, dataRegroupBySew_0_5};
  wire [15:0]      _GEN_72 = {dataRegroupBySew_5_5, dataRegroupBySew_4_5};
  wire [15:0]      dataInMem_hi_hi_26;
  assign dataInMem_hi_hi_26 = _GEN_72;
  wire [15:0]      dataInMem_hi_lo_28;
  assign dataInMem_hi_lo_28 = _GEN_72;
  wire [23:0]      dataInMem_hi_58 = {dataInMem_hi_hi_26, dataRegroupBySew_3_5};
  wire [23:0]      dataInMem_lo_43 = {dataInMem_lo_hi_11, dataRegroupBySew_0_6};
  wire [15:0]      _GEN_73 = {dataRegroupBySew_5_6, dataRegroupBySew_4_6};
  wire [15:0]      dataInMem_hi_hi_27;
  assign dataInMem_hi_hi_27 = _GEN_73;
  wire [15:0]      dataInMem_hi_lo_29;
  assign dataInMem_hi_lo_29 = _GEN_73;
  wire [23:0]      dataInMem_hi_59 = {dataInMem_hi_hi_27, dataRegroupBySew_3_6};
  wire [23:0]      dataInMem_lo_44 = {dataInMem_lo_hi_12, dataRegroupBySew_0_7};
  wire [15:0]      _GEN_74 = {dataRegroupBySew_5_7, dataRegroupBySew_4_7};
  wire [15:0]      dataInMem_hi_hi_28;
  assign dataInMem_hi_hi_28 = _GEN_74;
  wire [15:0]      dataInMem_hi_lo_30;
  assign dataInMem_hi_lo_30 = _GEN_74;
  wire [23:0]      dataInMem_hi_60 = {dataInMem_hi_hi_28, dataRegroupBySew_3_7};
  wire [23:0]      dataInMem_lo_45 = {dataInMem_lo_hi_13, dataRegroupBySew_0_8};
  wire [15:0]      _GEN_75 = {dataRegroupBySew_5_8, dataRegroupBySew_4_8};
  wire [15:0]      dataInMem_hi_hi_29;
  assign dataInMem_hi_hi_29 = _GEN_75;
  wire [15:0]      dataInMem_hi_lo_31;
  assign dataInMem_hi_lo_31 = _GEN_75;
  wire [23:0]      dataInMem_hi_61 = {dataInMem_hi_hi_29, dataRegroupBySew_3_8};
  wire [23:0]      dataInMem_lo_46 = {dataInMem_lo_hi_14, dataRegroupBySew_0_9};
  wire [15:0]      _GEN_76 = {dataRegroupBySew_5_9, dataRegroupBySew_4_9};
  wire [15:0]      dataInMem_hi_hi_30;
  assign dataInMem_hi_hi_30 = _GEN_76;
  wire [15:0]      dataInMem_hi_lo_32;
  assign dataInMem_hi_lo_32 = _GEN_76;
  wire [23:0]      dataInMem_hi_62 = {dataInMem_hi_hi_30, dataRegroupBySew_3_9};
  wire [23:0]      dataInMem_lo_47 = {dataInMem_lo_hi_15, dataRegroupBySew_0_10};
  wire [15:0]      _GEN_77 = {dataRegroupBySew_5_10, dataRegroupBySew_4_10};
  wire [15:0]      dataInMem_hi_hi_31;
  assign dataInMem_hi_hi_31 = _GEN_77;
  wire [15:0]      dataInMem_hi_lo_33;
  assign dataInMem_hi_lo_33 = _GEN_77;
  wire [23:0]      dataInMem_hi_63 = {dataInMem_hi_hi_31, dataRegroupBySew_3_10};
  wire [23:0]      dataInMem_lo_48 = {dataInMem_lo_hi_16, dataRegroupBySew_0_11};
  wire [15:0]      _GEN_78 = {dataRegroupBySew_5_11, dataRegroupBySew_4_11};
  wire [15:0]      dataInMem_hi_hi_32;
  assign dataInMem_hi_hi_32 = _GEN_78;
  wire [15:0]      dataInMem_hi_lo_34;
  assign dataInMem_hi_lo_34 = _GEN_78;
  wire [23:0]      dataInMem_hi_64 = {dataInMem_hi_hi_32, dataRegroupBySew_3_11};
  wire [23:0]      dataInMem_lo_49 = {dataInMem_lo_hi_17, dataRegroupBySew_0_12};
  wire [15:0]      _GEN_79 = {dataRegroupBySew_5_12, dataRegroupBySew_4_12};
  wire [15:0]      dataInMem_hi_hi_33;
  assign dataInMem_hi_hi_33 = _GEN_79;
  wire [15:0]      dataInMem_hi_lo_35;
  assign dataInMem_hi_lo_35 = _GEN_79;
  wire [23:0]      dataInMem_hi_65 = {dataInMem_hi_hi_33, dataRegroupBySew_3_12};
  wire [23:0]      dataInMem_lo_50 = {dataInMem_lo_hi_18, dataRegroupBySew_0_13};
  wire [15:0]      _GEN_80 = {dataRegroupBySew_5_13, dataRegroupBySew_4_13};
  wire [15:0]      dataInMem_hi_hi_34;
  assign dataInMem_hi_hi_34 = _GEN_80;
  wire [15:0]      dataInMem_hi_lo_36;
  assign dataInMem_hi_lo_36 = _GEN_80;
  wire [23:0]      dataInMem_hi_66 = {dataInMem_hi_hi_34, dataRegroupBySew_3_13};
  wire [23:0]      dataInMem_lo_51 = {dataInMem_lo_hi_19, dataRegroupBySew_0_14};
  wire [15:0]      _GEN_81 = {dataRegroupBySew_5_14, dataRegroupBySew_4_14};
  wire [15:0]      dataInMem_hi_hi_35;
  assign dataInMem_hi_hi_35 = _GEN_81;
  wire [15:0]      dataInMem_hi_lo_37;
  assign dataInMem_hi_lo_37 = _GEN_81;
  wire [23:0]      dataInMem_hi_67 = {dataInMem_hi_hi_35, dataRegroupBySew_3_14};
  wire [23:0]      dataInMem_lo_52 = {dataInMem_lo_hi_20, dataRegroupBySew_0_15};
  wire [15:0]      _GEN_82 = {dataRegroupBySew_5_15, dataRegroupBySew_4_15};
  wire [15:0]      dataInMem_hi_hi_36;
  assign dataInMem_hi_hi_36 = _GEN_82;
  wire [15:0]      dataInMem_hi_lo_38;
  assign dataInMem_hi_lo_38 = _GEN_82;
  wire [23:0]      dataInMem_hi_68 = {dataInMem_hi_hi_36, dataRegroupBySew_3_15};
  wire [95:0]      dataInMem_lo_lo_lo_5 = {dataInMem_hi_54, dataInMem_lo_38, dataInMem_hi_53, dataInMem_lo_37};
  wire [95:0]      dataInMem_lo_lo_hi_5 = {dataInMem_hi_56, dataInMem_lo_40, dataInMem_hi_55, dataInMem_lo_39};
  wire [191:0]     dataInMem_lo_lo_5 = {dataInMem_lo_lo_hi_5, dataInMem_lo_lo_lo_5};
  wire [95:0]      dataInMem_lo_hi_lo_5 = {dataInMem_hi_58, dataInMem_lo_42, dataInMem_hi_57, dataInMem_lo_41};
  wire [95:0]      dataInMem_lo_hi_hi_5 = {dataInMem_hi_60, dataInMem_lo_44, dataInMem_hi_59, dataInMem_lo_43};
  wire [191:0]     dataInMem_lo_hi_21 = {dataInMem_lo_hi_hi_5, dataInMem_lo_hi_lo_5};
  wire [383:0]     dataInMem_lo_53 = {dataInMem_lo_hi_21, dataInMem_lo_lo_5};
  wire [95:0]      dataInMem_hi_lo_lo_5 = {dataInMem_hi_62, dataInMem_lo_46, dataInMem_hi_61, dataInMem_lo_45};
  wire [95:0]      dataInMem_hi_lo_hi_5 = {dataInMem_hi_64, dataInMem_lo_48, dataInMem_hi_63, dataInMem_lo_47};
  wire [191:0]     dataInMem_hi_lo_5 = {dataInMem_hi_lo_hi_5, dataInMem_hi_lo_lo_5};
  wire [95:0]      dataInMem_hi_hi_lo_5 = {dataInMem_hi_66, dataInMem_lo_50, dataInMem_hi_65, dataInMem_lo_49};
  wire [95:0]      dataInMem_hi_hi_hi_5 = {dataInMem_hi_68, dataInMem_lo_52, dataInMem_hi_67, dataInMem_lo_51};
  wire [191:0]     dataInMem_hi_hi_37 = {dataInMem_hi_hi_hi_5, dataInMem_hi_hi_lo_5};
  wire [383:0]     dataInMem_hi_69 = {dataInMem_hi_hi_37, dataInMem_hi_lo_5};
  wire [767:0]     dataInMem_5 = {dataInMem_hi_69, dataInMem_lo_53};
  wire [127:0]     regroupCacheLine_5_0 = dataInMem_5[127:0];
  wire [127:0]     regroupCacheLine_5_1 = dataInMem_5[255:128];
  wire [127:0]     regroupCacheLine_5_2 = dataInMem_5[383:256];
  wire [127:0]     regroupCacheLine_5_3 = dataInMem_5[511:384];
  wire [127:0]     regroupCacheLine_5_4 = dataInMem_5[639:512];
  wire [127:0]     regroupCacheLine_5_5 = dataInMem_5[767:640];
  wire [127:0]     res_40 = regroupCacheLine_5_0;
  wire [127:0]     res_41 = regroupCacheLine_5_1;
  wire [127:0]     res_42 = regroupCacheLine_5_2;
  wire [127:0]     res_43 = regroupCacheLine_5_3;
  wire [127:0]     res_44 = regroupCacheLine_5_4;
  wire [127:0]     res_45 = regroupCacheLine_5_5;
  wire [255:0]     lo_lo_5 = {res_41, res_40};
  wire [255:0]     lo_hi_5 = {res_43, res_42};
  wire [511:0]     lo_5 = {lo_hi_5, lo_lo_5};
  wire [255:0]     hi_lo_5 = {res_45, res_44};
  wire [511:0]     hi_5 = {256'h0, hi_lo_5};
  wire [1023:0]    regroupLoadData_0_5 = {hi_5, lo_5};
  wire [23:0]      dataInMem_lo_54 = {dataInMem_lo_hi_22, dataRegroupBySew_0_0};
  wire [15:0]      dataInMem_hi_hi_38 = {dataRegroupBySew_6_0, dataRegroupBySew_5_0};
  wire [31:0]      dataInMem_hi_70 = {dataInMem_hi_hi_38, dataInMem_hi_lo_6};
  wire [23:0]      dataInMem_lo_55 = {dataInMem_lo_hi_23, dataRegroupBySew_0_1};
  wire [15:0]      dataInMem_hi_hi_39 = {dataRegroupBySew_6_1, dataRegroupBySew_5_1};
  wire [31:0]      dataInMem_hi_71 = {dataInMem_hi_hi_39, dataInMem_hi_lo_7};
  wire [23:0]      dataInMem_lo_56 = {dataInMem_lo_hi_24, dataRegroupBySew_0_2};
  wire [15:0]      dataInMem_hi_hi_40 = {dataRegroupBySew_6_2, dataRegroupBySew_5_2};
  wire [31:0]      dataInMem_hi_72 = {dataInMem_hi_hi_40, dataInMem_hi_lo_8};
  wire [23:0]      dataInMem_lo_57 = {dataInMem_lo_hi_25, dataRegroupBySew_0_3};
  wire [15:0]      dataInMem_hi_hi_41 = {dataRegroupBySew_6_3, dataRegroupBySew_5_3};
  wire [31:0]      dataInMem_hi_73 = {dataInMem_hi_hi_41, dataInMem_hi_lo_9};
  wire [23:0]      dataInMem_lo_58 = {dataInMem_lo_hi_26, dataRegroupBySew_0_4};
  wire [15:0]      dataInMem_hi_hi_42 = {dataRegroupBySew_6_4, dataRegroupBySew_5_4};
  wire [31:0]      dataInMem_hi_74 = {dataInMem_hi_hi_42, dataInMem_hi_lo_10};
  wire [23:0]      dataInMem_lo_59 = {dataInMem_lo_hi_27, dataRegroupBySew_0_5};
  wire [15:0]      dataInMem_hi_hi_43 = {dataRegroupBySew_6_5, dataRegroupBySew_5_5};
  wire [31:0]      dataInMem_hi_75 = {dataInMem_hi_hi_43, dataInMem_hi_lo_11};
  wire [23:0]      dataInMem_lo_60 = {dataInMem_lo_hi_28, dataRegroupBySew_0_6};
  wire [15:0]      dataInMem_hi_hi_44 = {dataRegroupBySew_6_6, dataRegroupBySew_5_6};
  wire [31:0]      dataInMem_hi_76 = {dataInMem_hi_hi_44, dataInMem_hi_lo_12};
  wire [23:0]      dataInMem_lo_61 = {dataInMem_lo_hi_29, dataRegroupBySew_0_7};
  wire [15:0]      dataInMem_hi_hi_45 = {dataRegroupBySew_6_7, dataRegroupBySew_5_7};
  wire [31:0]      dataInMem_hi_77 = {dataInMem_hi_hi_45, dataInMem_hi_lo_13};
  wire [23:0]      dataInMem_lo_62 = {dataInMem_lo_hi_30, dataRegroupBySew_0_8};
  wire [15:0]      dataInMem_hi_hi_46 = {dataRegroupBySew_6_8, dataRegroupBySew_5_8};
  wire [31:0]      dataInMem_hi_78 = {dataInMem_hi_hi_46, dataInMem_hi_lo_14};
  wire [23:0]      dataInMem_lo_63 = {dataInMem_lo_hi_31, dataRegroupBySew_0_9};
  wire [15:0]      dataInMem_hi_hi_47 = {dataRegroupBySew_6_9, dataRegroupBySew_5_9};
  wire [31:0]      dataInMem_hi_79 = {dataInMem_hi_hi_47, dataInMem_hi_lo_15};
  wire [23:0]      dataInMem_lo_64 = {dataInMem_lo_hi_32, dataRegroupBySew_0_10};
  wire [15:0]      dataInMem_hi_hi_48 = {dataRegroupBySew_6_10, dataRegroupBySew_5_10};
  wire [31:0]      dataInMem_hi_80 = {dataInMem_hi_hi_48, dataInMem_hi_lo_16};
  wire [23:0]      dataInMem_lo_65 = {dataInMem_lo_hi_33, dataRegroupBySew_0_11};
  wire [15:0]      dataInMem_hi_hi_49 = {dataRegroupBySew_6_11, dataRegroupBySew_5_11};
  wire [31:0]      dataInMem_hi_81 = {dataInMem_hi_hi_49, dataInMem_hi_lo_17};
  wire [23:0]      dataInMem_lo_66 = {dataInMem_lo_hi_34, dataRegroupBySew_0_12};
  wire [15:0]      dataInMem_hi_hi_50 = {dataRegroupBySew_6_12, dataRegroupBySew_5_12};
  wire [31:0]      dataInMem_hi_82 = {dataInMem_hi_hi_50, dataInMem_hi_lo_18};
  wire [23:0]      dataInMem_lo_67 = {dataInMem_lo_hi_35, dataRegroupBySew_0_13};
  wire [15:0]      dataInMem_hi_hi_51 = {dataRegroupBySew_6_13, dataRegroupBySew_5_13};
  wire [31:0]      dataInMem_hi_83 = {dataInMem_hi_hi_51, dataInMem_hi_lo_19};
  wire [23:0]      dataInMem_lo_68 = {dataInMem_lo_hi_36, dataRegroupBySew_0_14};
  wire [15:0]      dataInMem_hi_hi_52 = {dataRegroupBySew_6_14, dataRegroupBySew_5_14};
  wire [31:0]      dataInMem_hi_84 = {dataInMem_hi_hi_52, dataInMem_hi_lo_20};
  wire [23:0]      dataInMem_lo_69 = {dataInMem_lo_hi_37, dataRegroupBySew_0_15};
  wire [15:0]      dataInMem_hi_hi_53 = {dataRegroupBySew_6_15, dataRegroupBySew_5_15};
  wire [31:0]      dataInMem_hi_85 = {dataInMem_hi_hi_53, dataInMem_hi_lo_21};
  wire [111:0]     dataInMem_lo_lo_lo_6 = {dataInMem_hi_71, dataInMem_lo_55, dataInMem_hi_70, dataInMem_lo_54};
  wire [111:0]     dataInMem_lo_lo_hi_6 = {dataInMem_hi_73, dataInMem_lo_57, dataInMem_hi_72, dataInMem_lo_56};
  wire [223:0]     dataInMem_lo_lo_6 = {dataInMem_lo_lo_hi_6, dataInMem_lo_lo_lo_6};
  wire [111:0]     dataInMem_lo_hi_lo_6 = {dataInMem_hi_75, dataInMem_lo_59, dataInMem_hi_74, dataInMem_lo_58};
  wire [111:0]     dataInMem_lo_hi_hi_6 = {dataInMem_hi_77, dataInMem_lo_61, dataInMem_hi_76, dataInMem_lo_60};
  wire [223:0]     dataInMem_lo_hi_38 = {dataInMem_lo_hi_hi_6, dataInMem_lo_hi_lo_6};
  wire [447:0]     dataInMem_lo_70 = {dataInMem_lo_hi_38, dataInMem_lo_lo_6};
  wire [111:0]     dataInMem_hi_lo_lo_6 = {dataInMem_hi_79, dataInMem_lo_63, dataInMem_hi_78, dataInMem_lo_62};
  wire [111:0]     dataInMem_hi_lo_hi_6 = {dataInMem_hi_81, dataInMem_lo_65, dataInMem_hi_80, dataInMem_lo_64};
  wire [223:0]     dataInMem_hi_lo_22 = {dataInMem_hi_lo_hi_6, dataInMem_hi_lo_lo_6};
  wire [111:0]     dataInMem_hi_hi_lo_6 = {dataInMem_hi_83, dataInMem_lo_67, dataInMem_hi_82, dataInMem_lo_66};
  wire [111:0]     dataInMem_hi_hi_hi_6 = {dataInMem_hi_85, dataInMem_lo_69, dataInMem_hi_84, dataInMem_lo_68};
  wire [223:0]     dataInMem_hi_hi_54 = {dataInMem_hi_hi_hi_6, dataInMem_hi_hi_lo_6};
  wire [447:0]     dataInMem_hi_86 = {dataInMem_hi_hi_54, dataInMem_hi_lo_22};
  wire [895:0]     dataInMem_6 = {dataInMem_hi_86, dataInMem_lo_70};
  wire [127:0]     regroupCacheLine_6_0 = dataInMem_6[127:0];
  wire [127:0]     regroupCacheLine_6_1 = dataInMem_6[255:128];
  wire [127:0]     regroupCacheLine_6_2 = dataInMem_6[383:256];
  wire [127:0]     regroupCacheLine_6_3 = dataInMem_6[511:384];
  wire [127:0]     regroupCacheLine_6_4 = dataInMem_6[639:512];
  wire [127:0]     regroupCacheLine_6_5 = dataInMem_6[767:640];
  wire [127:0]     regroupCacheLine_6_6 = dataInMem_6[895:768];
  wire [127:0]     res_48 = regroupCacheLine_6_0;
  wire [127:0]     res_49 = regroupCacheLine_6_1;
  wire [127:0]     res_50 = regroupCacheLine_6_2;
  wire [127:0]     res_51 = regroupCacheLine_6_3;
  wire [127:0]     res_52 = regroupCacheLine_6_4;
  wire [127:0]     res_53 = regroupCacheLine_6_5;
  wire [127:0]     res_54 = regroupCacheLine_6_6;
  wire [255:0]     lo_lo_6 = {res_49, res_48};
  wire [255:0]     lo_hi_6 = {res_51, res_50};
  wire [511:0]     lo_6 = {lo_hi_6, lo_lo_6};
  wire [255:0]     hi_lo_6 = {res_53, res_52};
  wire [255:0]     hi_hi_6 = {128'h0, res_54};
  wire [511:0]     hi_6 = {hi_hi_6, hi_lo_6};
  wire [1023:0]    regroupLoadData_0_6 = {hi_6, lo_6};
  wire [31:0]      dataInMem_lo_71 = {dataInMem_lo_hi_39, dataInMem_lo_lo_7};
  wire [15:0]      dataInMem_hi_hi_55 = {dataRegroupBySew_7_0, dataRegroupBySew_6_0};
  wire [31:0]      dataInMem_hi_87 = {dataInMem_hi_hi_55, dataInMem_hi_lo_23};
  wire [31:0]      dataInMem_lo_72 = {dataInMem_lo_hi_40, dataInMem_lo_lo_8};
  wire [15:0]      dataInMem_hi_hi_56 = {dataRegroupBySew_7_1, dataRegroupBySew_6_1};
  wire [31:0]      dataInMem_hi_88 = {dataInMem_hi_hi_56, dataInMem_hi_lo_24};
  wire [31:0]      dataInMem_lo_73 = {dataInMem_lo_hi_41, dataInMem_lo_lo_9};
  wire [15:0]      dataInMem_hi_hi_57 = {dataRegroupBySew_7_2, dataRegroupBySew_6_2};
  wire [31:0]      dataInMem_hi_89 = {dataInMem_hi_hi_57, dataInMem_hi_lo_25};
  wire [31:0]      dataInMem_lo_74 = {dataInMem_lo_hi_42, dataInMem_lo_lo_10};
  wire [15:0]      dataInMem_hi_hi_58 = {dataRegroupBySew_7_3, dataRegroupBySew_6_3};
  wire [31:0]      dataInMem_hi_90 = {dataInMem_hi_hi_58, dataInMem_hi_lo_26};
  wire [31:0]      dataInMem_lo_75 = {dataInMem_lo_hi_43, dataInMem_lo_lo_11};
  wire [15:0]      dataInMem_hi_hi_59 = {dataRegroupBySew_7_4, dataRegroupBySew_6_4};
  wire [31:0]      dataInMem_hi_91 = {dataInMem_hi_hi_59, dataInMem_hi_lo_27};
  wire [31:0]      dataInMem_lo_76 = {dataInMem_lo_hi_44, dataInMem_lo_lo_12};
  wire [15:0]      dataInMem_hi_hi_60 = {dataRegroupBySew_7_5, dataRegroupBySew_6_5};
  wire [31:0]      dataInMem_hi_92 = {dataInMem_hi_hi_60, dataInMem_hi_lo_28};
  wire [31:0]      dataInMem_lo_77 = {dataInMem_lo_hi_45, dataInMem_lo_lo_13};
  wire [15:0]      dataInMem_hi_hi_61 = {dataRegroupBySew_7_6, dataRegroupBySew_6_6};
  wire [31:0]      dataInMem_hi_93 = {dataInMem_hi_hi_61, dataInMem_hi_lo_29};
  wire [31:0]      dataInMem_lo_78 = {dataInMem_lo_hi_46, dataInMem_lo_lo_14};
  wire [15:0]      dataInMem_hi_hi_62 = {dataRegroupBySew_7_7, dataRegroupBySew_6_7};
  wire [31:0]      dataInMem_hi_94 = {dataInMem_hi_hi_62, dataInMem_hi_lo_30};
  wire [31:0]      dataInMem_lo_79 = {dataInMem_lo_hi_47, dataInMem_lo_lo_15};
  wire [15:0]      dataInMem_hi_hi_63 = {dataRegroupBySew_7_8, dataRegroupBySew_6_8};
  wire [31:0]      dataInMem_hi_95 = {dataInMem_hi_hi_63, dataInMem_hi_lo_31};
  wire [31:0]      dataInMem_lo_80 = {dataInMem_lo_hi_48, dataInMem_lo_lo_16};
  wire [15:0]      dataInMem_hi_hi_64 = {dataRegroupBySew_7_9, dataRegroupBySew_6_9};
  wire [31:0]      dataInMem_hi_96 = {dataInMem_hi_hi_64, dataInMem_hi_lo_32};
  wire [31:0]      dataInMem_lo_81 = {dataInMem_lo_hi_49, dataInMem_lo_lo_17};
  wire [15:0]      dataInMem_hi_hi_65 = {dataRegroupBySew_7_10, dataRegroupBySew_6_10};
  wire [31:0]      dataInMem_hi_97 = {dataInMem_hi_hi_65, dataInMem_hi_lo_33};
  wire [31:0]      dataInMem_lo_82 = {dataInMem_lo_hi_50, dataInMem_lo_lo_18};
  wire [15:0]      dataInMem_hi_hi_66 = {dataRegroupBySew_7_11, dataRegroupBySew_6_11};
  wire [31:0]      dataInMem_hi_98 = {dataInMem_hi_hi_66, dataInMem_hi_lo_34};
  wire [31:0]      dataInMem_lo_83 = {dataInMem_lo_hi_51, dataInMem_lo_lo_19};
  wire [15:0]      dataInMem_hi_hi_67 = {dataRegroupBySew_7_12, dataRegroupBySew_6_12};
  wire [31:0]      dataInMem_hi_99 = {dataInMem_hi_hi_67, dataInMem_hi_lo_35};
  wire [31:0]      dataInMem_lo_84 = {dataInMem_lo_hi_52, dataInMem_lo_lo_20};
  wire [15:0]      dataInMem_hi_hi_68 = {dataRegroupBySew_7_13, dataRegroupBySew_6_13};
  wire [31:0]      dataInMem_hi_100 = {dataInMem_hi_hi_68, dataInMem_hi_lo_36};
  wire [31:0]      dataInMem_lo_85 = {dataInMem_lo_hi_53, dataInMem_lo_lo_21};
  wire [15:0]      dataInMem_hi_hi_69 = {dataRegroupBySew_7_14, dataRegroupBySew_6_14};
  wire [31:0]      dataInMem_hi_101 = {dataInMem_hi_hi_69, dataInMem_hi_lo_37};
  wire [31:0]      dataInMem_lo_86 = {dataInMem_lo_hi_54, dataInMem_lo_lo_22};
  wire [15:0]      dataInMem_hi_hi_70 = {dataRegroupBySew_7_15, dataRegroupBySew_6_15};
  wire [31:0]      dataInMem_hi_102 = {dataInMem_hi_hi_70, dataInMem_hi_lo_38};
  wire [127:0]     dataInMem_lo_lo_lo_7 = {dataInMem_hi_88, dataInMem_lo_72, dataInMem_hi_87, dataInMem_lo_71};
  wire [127:0]     dataInMem_lo_lo_hi_7 = {dataInMem_hi_90, dataInMem_lo_74, dataInMem_hi_89, dataInMem_lo_73};
  wire [255:0]     dataInMem_lo_lo_23 = {dataInMem_lo_lo_hi_7, dataInMem_lo_lo_lo_7};
  wire [127:0]     dataInMem_lo_hi_lo_7 = {dataInMem_hi_92, dataInMem_lo_76, dataInMem_hi_91, dataInMem_lo_75};
  wire [127:0]     dataInMem_lo_hi_hi_7 = {dataInMem_hi_94, dataInMem_lo_78, dataInMem_hi_93, dataInMem_lo_77};
  wire [255:0]     dataInMem_lo_hi_55 = {dataInMem_lo_hi_hi_7, dataInMem_lo_hi_lo_7};
  wire [511:0]     dataInMem_lo_87 = {dataInMem_lo_hi_55, dataInMem_lo_lo_23};
  wire [127:0]     dataInMem_hi_lo_lo_7 = {dataInMem_hi_96, dataInMem_lo_80, dataInMem_hi_95, dataInMem_lo_79};
  wire [127:0]     dataInMem_hi_lo_hi_7 = {dataInMem_hi_98, dataInMem_lo_82, dataInMem_hi_97, dataInMem_lo_81};
  wire [255:0]     dataInMem_hi_lo_39 = {dataInMem_hi_lo_hi_7, dataInMem_hi_lo_lo_7};
  wire [127:0]     dataInMem_hi_hi_lo_7 = {dataInMem_hi_100, dataInMem_lo_84, dataInMem_hi_99, dataInMem_lo_83};
  wire [127:0]     dataInMem_hi_hi_hi_7 = {dataInMem_hi_102, dataInMem_lo_86, dataInMem_hi_101, dataInMem_lo_85};
  wire [255:0]     dataInMem_hi_hi_71 = {dataInMem_hi_hi_hi_7, dataInMem_hi_hi_lo_7};
  wire [511:0]     dataInMem_hi_103 = {dataInMem_hi_hi_71, dataInMem_hi_lo_39};
  wire [1023:0]    dataInMem_7 = {dataInMem_hi_103, dataInMem_lo_87};
  wire [127:0]     regroupCacheLine_7_0 = dataInMem_7[127:0];
  wire [127:0]     regroupCacheLine_7_1 = dataInMem_7[255:128];
  wire [127:0]     regroupCacheLine_7_2 = dataInMem_7[383:256];
  wire [127:0]     regroupCacheLine_7_3 = dataInMem_7[511:384];
  wire [127:0]     regroupCacheLine_7_4 = dataInMem_7[639:512];
  wire [127:0]     regroupCacheLine_7_5 = dataInMem_7[767:640];
  wire [127:0]     regroupCacheLine_7_6 = dataInMem_7[895:768];
  wire [127:0]     regroupCacheLine_7_7 = dataInMem_7[1023:896];
  wire [127:0]     res_56 = regroupCacheLine_7_0;
  wire [127:0]     res_57 = regroupCacheLine_7_1;
  wire [127:0]     res_58 = regroupCacheLine_7_2;
  wire [127:0]     res_59 = regroupCacheLine_7_3;
  wire [127:0]     res_60 = regroupCacheLine_7_4;
  wire [127:0]     res_61 = regroupCacheLine_7_5;
  wire [127:0]     res_62 = regroupCacheLine_7_6;
  wire [127:0]     res_63 = regroupCacheLine_7_7;
  wire [255:0]     lo_lo_7 = {res_57, res_56};
  wire [255:0]     lo_hi_7 = {res_59, res_58};
  wire [511:0]     lo_7 = {lo_hi_7, lo_lo_7};
  wire [255:0]     hi_lo_7 = {res_61, res_60};
  wire [255:0]     hi_hi_7 = {res_63, res_62};
  wire [511:0]     hi_7 = {hi_hi_7, hi_lo_7};
  wire [1023:0]    regroupLoadData_0_7 = {hi_7, lo_7};
  wire [15:0]      dataRegroupBySew_0_1_0 = bufferStageEnqueueData_0[15:0];
  wire [15:0]      dataRegroupBySew_0_1_1 = bufferStageEnqueueData_0[31:16];
  wire [15:0]      dataRegroupBySew_0_1_2 = bufferStageEnqueueData_0[47:32];
  wire [15:0]      dataRegroupBySew_0_1_3 = bufferStageEnqueueData_0[63:48];
  wire [15:0]      dataRegroupBySew_0_1_4 = bufferStageEnqueueData_0[79:64];
  wire [15:0]      dataRegroupBySew_0_1_5 = bufferStageEnqueueData_0[95:80];
  wire [15:0]      dataRegroupBySew_0_1_6 = bufferStageEnqueueData_0[111:96];
  wire [15:0]      dataRegroupBySew_0_1_7 = bufferStageEnqueueData_0[127:112];
  wire [15:0]      dataRegroupBySew_1_1_0 = bufferStageEnqueueData_1[15:0];
  wire [15:0]      dataRegroupBySew_1_1_1 = bufferStageEnqueueData_1[31:16];
  wire [15:0]      dataRegroupBySew_1_1_2 = bufferStageEnqueueData_1[47:32];
  wire [15:0]      dataRegroupBySew_1_1_3 = bufferStageEnqueueData_1[63:48];
  wire [15:0]      dataRegroupBySew_1_1_4 = bufferStageEnqueueData_1[79:64];
  wire [15:0]      dataRegroupBySew_1_1_5 = bufferStageEnqueueData_1[95:80];
  wire [15:0]      dataRegroupBySew_1_1_6 = bufferStageEnqueueData_1[111:96];
  wire [15:0]      dataRegroupBySew_1_1_7 = bufferStageEnqueueData_1[127:112];
  wire [15:0]      dataRegroupBySew_2_1_0 = bufferStageEnqueueData_2[15:0];
  wire [15:0]      dataRegroupBySew_2_1_1 = bufferStageEnqueueData_2[31:16];
  wire [15:0]      dataRegroupBySew_2_1_2 = bufferStageEnqueueData_2[47:32];
  wire [15:0]      dataRegroupBySew_2_1_3 = bufferStageEnqueueData_2[63:48];
  wire [15:0]      dataRegroupBySew_2_1_4 = bufferStageEnqueueData_2[79:64];
  wire [15:0]      dataRegroupBySew_2_1_5 = bufferStageEnqueueData_2[95:80];
  wire [15:0]      dataRegroupBySew_2_1_6 = bufferStageEnqueueData_2[111:96];
  wire [15:0]      dataRegroupBySew_2_1_7 = bufferStageEnqueueData_2[127:112];
  wire [15:0]      dataRegroupBySew_3_1_0 = bufferStageEnqueueData_3[15:0];
  wire [15:0]      dataRegroupBySew_3_1_1 = bufferStageEnqueueData_3[31:16];
  wire [15:0]      dataRegroupBySew_3_1_2 = bufferStageEnqueueData_3[47:32];
  wire [15:0]      dataRegroupBySew_3_1_3 = bufferStageEnqueueData_3[63:48];
  wire [15:0]      dataRegroupBySew_3_1_4 = bufferStageEnqueueData_3[79:64];
  wire [15:0]      dataRegroupBySew_3_1_5 = bufferStageEnqueueData_3[95:80];
  wire [15:0]      dataRegroupBySew_3_1_6 = bufferStageEnqueueData_3[111:96];
  wire [15:0]      dataRegroupBySew_3_1_7 = bufferStageEnqueueData_3[127:112];
  wire [15:0]      dataRegroupBySew_4_1_0 = bufferStageEnqueueData_4[15:0];
  wire [15:0]      dataRegroupBySew_4_1_1 = bufferStageEnqueueData_4[31:16];
  wire [15:0]      dataRegroupBySew_4_1_2 = bufferStageEnqueueData_4[47:32];
  wire [15:0]      dataRegroupBySew_4_1_3 = bufferStageEnqueueData_4[63:48];
  wire [15:0]      dataRegroupBySew_4_1_4 = bufferStageEnqueueData_4[79:64];
  wire [15:0]      dataRegroupBySew_4_1_5 = bufferStageEnqueueData_4[95:80];
  wire [15:0]      dataRegroupBySew_4_1_6 = bufferStageEnqueueData_4[111:96];
  wire [15:0]      dataRegroupBySew_4_1_7 = bufferStageEnqueueData_4[127:112];
  wire [15:0]      dataRegroupBySew_5_1_0 = bufferStageEnqueueData_5[15:0];
  wire [15:0]      dataRegroupBySew_5_1_1 = bufferStageEnqueueData_5[31:16];
  wire [15:0]      dataRegroupBySew_5_1_2 = bufferStageEnqueueData_5[47:32];
  wire [15:0]      dataRegroupBySew_5_1_3 = bufferStageEnqueueData_5[63:48];
  wire [15:0]      dataRegroupBySew_5_1_4 = bufferStageEnqueueData_5[79:64];
  wire [15:0]      dataRegroupBySew_5_1_5 = bufferStageEnqueueData_5[95:80];
  wire [15:0]      dataRegroupBySew_5_1_6 = bufferStageEnqueueData_5[111:96];
  wire [15:0]      dataRegroupBySew_5_1_7 = bufferStageEnqueueData_5[127:112];
  wire [15:0]      dataRegroupBySew_6_1_0 = bufferStageEnqueueData_6[15:0];
  wire [15:0]      dataRegroupBySew_6_1_1 = bufferStageEnqueueData_6[31:16];
  wire [15:0]      dataRegroupBySew_6_1_2 = bufferStageEnqueueData_6[47:32];
  wire [15:0]      dataRegroupBySew_6_1_3 = bufferStageEnqueueData_6[63:48];
  wire [15:0]      dataRegroupBySew_6_1_4 = bufferStageEnqueueData_6[79:64];
  wire [15:0]      dataRegroupBySew_6_1_5 = bufferStageEnqueueData_6[95:80];
  wire [15:0]      dataRegroupBySew_6_1_6 = bufferStageEnqueueData_6[111:96];
  wire [15:0]      dataRegroupBySew_6_1_7 = bufferStageEnqueueData_6[127:112];
  wire [15:0]      dataRegroupBySew_7_1_0 = bufferStageEnqueueData_7[15:0];
  wire [15:0]      dataRegroupBySew_7_1_1 = bufferStageEnqueueData_7[31:16];
  wire [15:0]      dataRegroupBySew_7_1_2 = bufferStageEnqueueData_7[47:32];
  wire [15:0]      dataRegroupBySew_7_1_3 = bufferStageEnqueueData_7[63:48];
  wire [15:0]      dataRegroupBySew_7_1_4 = bufferStageEnqueueData_7[79:64];
  wire [15:0]      dataRegroupBySew_7_1_5 = bufferStageEnqueueData_7[95:80];
  wire [15:0]      dataRegroupBySew_7_1_6 = bufferStageEnqueueData_7[111:96];
  wire [15:0]      dataRegroupBySew_7_1_7 = bufferStageEnqueueData_7[127:112];
  wire [31:0]      dataInMem_lo_lo_24 = {dataRegroupBySew_0_1_1, dataRegroupBySew_0_1_0};
  wire [31:0]      dataInMem_lo_hi_56 = {dataRegroupBySew_0_1_3, dataRegroupBySew_0_1_2};
  wire [63:0]      dataInMem_lo_88 = {dataInMem_lo_hi_56, dataInMem_lo_lo_24};
  wire [31:0]      dataInMem_hi_lo_40 = {dataRegroupBySew_0_1_5, dataRegroupBySew_0_1_4};
  wire [31:0]      dataInMem_hi_hi_72 = {dataRegroupBySew_0_1_7, dataRegroupBySew_0_1_6};
  wire [63:0]      dataInMem_hi_104 = {dataInMem_hi_hi_72, dataInMem_hi_lo_40};
  wire [127:0]     dataInMem_8 = {dataInMem_hi_104, dataInMem_lo_88};
  wire [127:0]     regroupCacheLine_8_0 = dataInMem_8;
  wire [127:0]     res_64 = regroupCacheLine_8_0;
  wire [255:0]     lo_lo_8 = {128'h0, res_64};
  wire [511:0]     lo_8 = {256'h0, lo_lo_8};
  wire [1023:0]    regroupLoadData_1_0 = {512'h0, lo_8};
  wire [63:0]      dataInMem_lo_lo_25 = {dataRegroupBySew_1_1_1, dataRegroupBySew_0_1_1, dataRegroupBySew_1_1_0, dataRegroupBySew_0_1_0};
  wire [63:0]      dataInMem_lo_hi_57 = {dataRegroupBySew_1_1_3, dataRegroupBySew_0_1_3, dataRegroupBySew_1_1_2, dataRegroupBySew_0_1_2};
  wire [127:0]     dataInMem_lo_89 = {dataInMem_lo_hi_57, dataInMem_lo_lo_25};
  wire [63:0]      dataInMem_hi_lo_41 = {dataRegroupBySew_1_1_5, dataRegroupBySew_0_1_5, dataRegroupBySew_1_1_4, dataRegroupBySew_0_1_4};
  wire [63:0]      dataInMem_hi_hi_73 = {dataRegroupBySew_1_1_7, dataRegroupBySew_0_1_7, dataRegroupBySew_1_1_6, dataRegroupBySew_0_1_6};
  wire [127:0]     dataInMem_hi_105 = {dataInMem_hi_hi_73, dataInMem_hi_lo_41};
  wire [255:0]     dataInMem_9 = {dataInMem_hi_105, dataInMem_lo_89};
  wire [127:0]     regroupCacheLine_9_0 = dataInMem_9[127:0];
  wire [127:0]     regroupCacheLine_9_1 = dataInMem_9[255:128];
  wire [127:0]     res_72 = regroupCacheLine_9_0;
  wire [127:0]     res_73 = regroupCacheLine_9_1;
  wire [255:0]     lo_lo_9 = {res_73, res_72};
  wire [511:0]     lo_9 = {256'h0, lo_lo_9};
  wire [1023:0]    regroupLoadData_1_1 = {512'h0, lo_9};
  wire [31:0]      _GEN_83 = {dataRegroupBySew_2_1_0, dataRegroupBySew_1_1_0};
  wire [31:0]      dataInMem_hi_106;
  assign dataInMem_hi_106 = _GEN_83;
  wire [31:0]      dataInMem_lo_hi_61;
  assign dataInMem_lo_hi_61 = _GEN_83;
  wire [31:0]      dataInMem_lo_hi_70;
  assign dataInMem_lo_hi_70 = _GEN_83;
  wire [31:0]      _GEN_84 = {dataRegroupBySew_2_1_1, dataRegroupBySew_1_1_1};
  wire [31:0]      dataInMem_hi_107;
  assign dataInMem_hi_107 = _GEN_84;
  wire [31:0]      dataInMem_lo_hi_62;
  assign dataInMem_lo_hi_62 = _GEN_84;
  wire [31:0]      dataInMem_lo_hi_71;
  assign dataInMem_lo_hi_71 = _GEN_84;
  wire [31:0]      _GEN_85 = {dataRegroupBySew_2_1_2, dataRegroupBySew_1_1_2};
  wire [31:0]      dataInMem_hi_108;
  assign dataInMem_hi_108 = _GEN_85;
  wire [31:0]      dataInMem_lo_hi_63;
  assign dataInMem_lo_hi_63 = _GEN_85;
  wire [31:0]      dataInMem_lo_hi_72;
  assign dataInMem_lo_hi_72 = _GEN_85;
  wire [31:0]      _GEN_86 = {dataRegroupBySew_2_1_3, dataRegroupBySew_1_1_3};
  wire [31:0]      dataInMem_hi_109;
  assign dataInMem_hi_109 = _GEN_86;
  wire [31:0]      dataInMem_lo_hi_64;
  assign dataInMem_lo_hi_64 = _GEN_86;
  wire [31:0]      dataInMem_lo_hi_73;
  assign dataInMem_lo_hi_73 = _GEN_86;
  wire [31:0]      _GEN_87 = {dataRegroupBySew_2_1_4, dataRegroupBySew_1_1_4};
  wire [31:0]      dataInMem_hi_110;
  assign dataInMem_hi_110 = _GEN_87;
  wire [31:0]      dataInMem_lo_hi_65;
  assign dataInMem_lo_hi_65 = _GEN_87;
  wire [31:0]      dataInMem_lo_hi_74;
  assign dataInMem_lo_hi_74 = _GEN_87;
  wire [31:0]      _GEN_88 = {dataRegroupBySew_2_1_5, dataRegroupBySew_1_1_5};
  wire [31:0]      dataInMem_hi_111;
  assign dataInMem_hi_111 = _GEN_88;
  wire [31:0]      dataInMem_lo_hi_66;
  assign dataInMem_lo_hi_66 = _GEN_88;
  wire [31:0]      dataInMem_lo_hi_75;
  assign dataInMem_lo_hi_75 = _GEN_88;
  wire [31:0]      _GEN_89 = {dataRegroupBySew_2_1_6, dataRegroupBySew_1_1_6};
  wire [31:0]      dataInMem_hi_112;
  assign dataInMem_hi_112 = _GEN_89;
  wire [31:0]      dataInMem_lo_hi_67;
  assign dataInMem_lo_hi_67 = _GEN_89;
  wire [31:0]      dataInMem_lo_hi_76;
  assign dataInMem_lo_hi_76 = _GEN_89;
  wire [31:0]      _GEN_90 = {dataRegroupBySew_2_1_7, dataRegroupBySew_1_1_7};
  wire [31:0]      dataInMem_hi_113;
  assign dataInMem_hi_113 = _GEN_90;
  wire [31:0]      dataInMem_lo_hi_68;
  assign dataInMem_lo_hi_68 = _GEN_90;
  wire [31:0]      dataInMem_lo_hi_77;
  assign dataInMem_lo_hi_77 = _GEN_90;
  wire [95:0]      dataInMem_lo_lo_26 = {dataInMem_hi_107, dataRegroupBySew_0_1_1, dataInMem_hi_106, dataRegroupBySew_0_1_0};
  wire [95:0]      dataInMem_lo_hi_58 = {dataInMem_hi_109, dataRegroupBySew_0_1_3, dataInMem_hi_108, dataRegroupBySew_0_1_2};
  wire [191:0]     dataInMem_lo_90 = {dataInMem_lo_hi_58, dataInMem_lo_lo_26};
  wire [95:0]      dataInMem_hi_lo_42 = {dataInMem_hi_111, dataRegroupBySew_0_1_5, dataInMem_hi_110, dataRegroupBySew_0_1_4};
  wire [95:0]      dataInMem_hi_hi_74 = {dataInMem_hi_113, dataRegroupBySew_0_1_7, dataInMem_hi_112, dataRegroupBySew_0_1_6};
  wire [191:0]     dataInMem_hi_114 = {dataInMem_hi_hi_74, dataInMem_hi_lo_42};
  wire [383:0]     dataInMem_10 = {dataInMem_hi_114, dataInMem_lo_90};
  wire [127:0]     regroupCacheLine_10_0 = dataInMem_10[127:0];
  wire [127:0]     regroupCacheLine_10_1 = dataInMem_10[255:128];
  wire [127:0]     regroupCacheLine_10_2 = dataInMem_10[383:256];
  wire [127:0]     res_80 = regroupCacheLine_10_0;
  wire [127:0]     res_81 = regroupCacheLine_10_1;
  wire [127:0]     res_82 = regroupCacheLine_10_2;
  wire [255:0]     lo_lo_10 = {res_81, res_80};
  wire [255:0]     lo_hi_10 = {128'h0, res_82};
  wire [511:0]     lo_10 = {lo_hi_10, lo_lo_10};
  wire [1023:0]    regroupLoadData_1_2 = {512'h0, lo_10};
  wire [31:0]      _GEN_91 = {dataRegroupBySew_1_1_0, dataRegroupBySew_0_1_0};
  wire [31:0]      dataInMem_lo_91;
  assign dataInMem_lo_91 = _GEN_91;
  wire [31:0]      dataInMem_lo_100;
  assign dataInMem_lo_100 = _GEN_91;
  wire [31:0]      dataInMem_lo_lo_31;
  assign dataInMem_lo_lo_31 = _GEN_91;
  wire [31:0]      _GEN_92 = {dataRegroupBySew_3_1_0, dataRegroupBySew_2_1_0};
  wire [31:0]      dataInMem_hi_115;
  assign dataInMem_hi_115 = _GEN_92;
  wire [31:0]      dataInMem_lo_hi_79;
  assign dataInMem_lo_hi_79 = _GEN_92;
  wire [31:0]      _GEN_93 = {dataRegroupBySew_1_1_1, dataRegroupBySew_0_1_1};
  wire [31:0]      dataInMem_lo_92;
  assign dataInMem_lo_92 = _GEN_93;
  wire [31:0]      dataInMem_lo_101;
  assign dataInMem_lo_101 = _GEN_93;
  wire [31:0]      dataInMem_lo_lo_32;
  assign dataInMem_lo_lo_32 = _GEN_93;
  wire [31:0]      _GEN_94 = {dataRegroupBySew_3_1_1, dataRegroupBySew_2_1_1};
  wire [31:0]      dataInMem_hi_116;
  assign dataInMem_hi_116 = _GEN_94;
  wire [31:0]      dataInMem_lo_hi_80;
  assign dataInMem_lo_hi_80 = _GEN_94;
  wire [31:0]      _GEN_95 = {dataRegroupBySew_1_1_2, dataRegroupBySew_0_1_2};
  wire [31:0]      dataInMem_lo_93;
  assign dataInMem_lo_93 = _GEN_95;
  wire [31:0]      dataInMem_lo_102;
  assign dataInMem_lo_102 = _GEN_95;
  wire [31:0]      dataInMem_lo_lo_33;
  assign dataInMem_lo_lo_33 = _GEN_95;
  wire [31:0]      _GEN_96 = {dataRegroupBySew_3_1_2, dataRegroupBySew_2_1_2};
  wire [31:0]      dataInMem_hi_117;
  assign dataInMem_hi_117 = _GEN_96;
  wire [31:0]      dataInMem_lo_hi_81;
  assign dataInMem_lo_hi_81 = _GEN_96;
  wire [31:0]      _GEN_97 = {dataRegroupBySew_1_1_3, dataRegroupBySew_0_1_3};
  wire [31:0]      dataInMem_lo_94;
  assign dataInMem_lo_94 = _GEN_97;
  wire [31:0]      dataInMem_lo_103;
  assign dataInMem_lo_103 = _GEN_97;
  wire [31:0]      dataInMem_lo_lo_34;
  assign dataInMem_lo_lo_34 = _GEN_97;
  wire [31:0]      _GEN_98 = {dataRegroupBySew_3_1_3, dataRegroupBySew_2_1_3};
  wire [31:0]      dataInMem_hi_118;
  assign dataInMem_hi_118 = _GEN_98;
  wire [31:0]      dataInMem_lo_hi_82;
  assign dataInMem_lo_hi_82 = _GEN_98;
  wire [31:0]      _GEN_99 = {dataRegroupBySew_1_1_4, dataRegroupBySew_0_1_4};
  wire [31:0]      dataInMem_lo_95;
  assign dataInMem_lo_95 = _GEN_99;
  wire [31:0]      dataInMem_lo_104;
  assign dataInMem_lo_104 = _GEN_99;
  wire [31:0]      dataInMem_lo_lo_35;
  assign dataInMem_lo_lo_35 = _GEN_99;
  wire [31:0]      _GEN_100 = {dataRegroupBySew_3_1_4, dataRegroupBySew_2_1_4};
  wire [31:0]      dataInMem_hi_119;
  assign dataInMem_hi_119 = _GEN_100;
  wire [31:0]      dataInMem_lo_hi_83;
  assign dataInMem_lo_hi_83 = _GEN_100;
  wire [31:0]      _GEN_101 = {dataRegroupBySew_1_1_5, dataRegroupBySew_0_1_5};
  wire [31:0]      dataInMem_lo_96;
  assign dataInMem_lo_96 = _GEN_101;
  wire [31:0]      dataInMem_lo_105;
  assign dataInMem_lo_105 = _GEN_101;
  wire [31:0]      dataInMem_lo_lo_36;
  assign dataInMem_lo_lo_36 = _GEN_101;
  wire [31:0]      _GEN_102 = {dataRegroupBySew_3_1_5, dataRegroupBySew_2_1_5};
  wire [31:0]      dataInMem_hi_120;
  assign dataInMem_hi_120 = _GEN_102;
  wire [31:0]      dataInMem_lo_hi_84;
  assign dataInMem_lo_hi_84 = _GEN_102;
  wire [31:0]      _GEN_103 = {dataRegroupBySew_1_1_6, dataRegroupBySew_0_1_6};
  wire [31:0]      dataInMem_lo_97;
  assign dataInMem_lo_97 = _GEN_103;
  wire [31:0]      dataInMem_lo_106;
  assign dataInMem_lo_106 = _GEN_103;
  wire [31:0]      dataInMem_lo_lo_37;
  assign dataInMem_lo_lo_37 = _GEN_103;
  wire [31:0]      _GEN_104 = {dataRegroupBySew_3_1_6, dataRegroupBySew_2_1_6};
  wire [31:0]      dataInMem_hi_121;
  assign dataInMem_hi_121 = _GEN_104;
  wire [31:0]      dataInMem_lo_hi_85;
  assign dataInMem_lo_hi_85 = _GEN_104;
  wire [31:0]      _GEN_105 = {dataRegroupBySew_1_1_7, dataRegroupBySew_0_1_7};
  wire [31:0]      dataInMem_lo_98;
  assign dataInMem_lo_98 = _GEN_105;
  wire [31:0]      dataInMem_lo_107;
  assign dataInMem_lo_107 = _GEN_105;
  wire [31:0]      dataInMem_lo_lo_38;
  assign dataInMem_lo_lo_38 = _GEN_105;
  wire [31:0]      _GEN_106 = {dataRegroupBySew_3_1_7, dataRegroupBySew_2_1_7};
  wire [31:0]      dataInMem_hi_122;
  assign dataInMem_hi_122 = _GEN_106;
  wire [31:0]      dataInMem_lo_hi_86;
  assign dataInMem_lo_hi_86 = _GEN_106;
  wire [127:0]     dataInMem_lo_lo_27 = {dataInMem_hi_116, dataInMem_lo_92, dataInMem_hi_115, dataInMem_lo_91};
  wire [127:0]     dataInMem_lo_hi_59 = {dataInMem_hi_118, dataInMem_lo_94, dataInMem_hi_117, dataInMem_lo_93};
  wire [255:0]     dataInMem_lo_99 = {dataInMem_lo_hi_59, dataInMem_lo_lo_27};
  wire [127:0]     dataInMem_hi_lo_43 = {dataInMem_hi_120, dataInMem_lo_96, dataInMem_hi_119, dataInMem_lo_95};
  wire [127:0]     dataInMem_hi_hi_75 = {dataInMem_hi_122, dataInMem_lo_98, dataInMem_hi_121, dataInMem_lo_97};
  wire [255:0]     dataInMem_hi_123 = {dataInMem_hi_hi_75, dataInMem_hi_lo_43};
  wire [511:0]     dataInMem_11 = {dataInMem_hi_123, dataInMem_lo_99};
  wire [127:0]     regroupCacheLine_11_0 = dataInMem_11[127:0];
  wire [127:0]     regroupCacheLine_11_1 = dataInMem_11[255:128];
  wire [127:0]     regroupCacheLine_11_2 = dataInMem_11[383:256];
  wire [127:0]     regroupCacheLine_11_3 = dataInMem_11[511:384];
  wire [127:0]     res_88 = regroupCacheLine_11_0;
  wire [127:0]     res_89 = regroupCacheLine_11_1;
  wire [127:0]     res_90 = regroupCacheLine_11_2;
  wire [127:0]     res_91 = regroupCacheLine_11_3;
  wire [255:0]     lo_lo_11 = {res_89, res_88};
  wire [255:0]     lo_hi_11 = {res_91, res_90};
  wire [511:0]     lo_11 = {lo_hi_11, lo_lo_11};
  wire [1023:0]    regroupLoadData_1_3 = {512'h0, lo_11};
  wire [31:0]      _GEN_107 = {dataRegroupBySew_4_1_0, dataRegroupBySew_3_1_0};
  wire [31:0]      dataInMem_hi_hi_76;
  assign dataInMem_hi_hi_76 = _GEN_107;
  wire [31:0]      dataInMem_hi_lo_46;
  assign dataInMem_hi_lo_46 = _GEN_107;
  wire [47:0]      dataInMem_hi_124 = {dataInMem_hi_hi_76, dataRegroupBySew_2_1_0};
  wire [31:0]      _GEN_108 = {dataRegroupBySew_4_1_1, dataRegroupBySew_3_1_1};
  wire [31:0]      dataInMem_hi_hi_77;
  assign dataInMem_hi_hi_77 = _GEN_108;
  wire [31:0]      dataInMem_hi_lo_47;
  assign dataInMem_hi_lo_47 = _GEN_108;
  wire [47:0]      dataInMem_hi_125 = {dataInMem_hi_hi_77, dataRegroupBySew_2_1_1};
  wire [31:0]      _GEN_109 = {dataRegroupBySew_4_1_2, dataRegroupBySew_3_1_2};
  wire [31:0]      dataInMem_hi_hi_78;
  assign dataInMem_hi_hi_78 = _GEN_109;
  wire [31:0]      dataInMem_hi_lo_48;
  assign dataInMem_hi_lo_48 = _GEN_109;
  wire [47:0]      dataInMem_hi_126 = {dataInMem_hi_hi_78, dataRegroupBySew_2_1_2};
  wire [31:0]      _GEN_110 = {dataRegroupBySew_4_1_3, dataRegroupBySew_3_1_3};
  wire [31:0]      dataInMem_hi_hi_79;
  assign dataInMem_hi_hi_79 = _GEN_110;
  wire [31:0]      dataInMem_hi_lo_49;
  assign dataInMem_hi_lo_49 = _GEN_110;
  wire [47:0]      dataInMem_hi_127 = {dataInMem_hi_hi_79, dataRegroupBySew_2_1_3};
  wire [31:0]      _GEN_111 = {dataRegroupBySew_4_1_4, dataRegroupBySew_3_1_4};
  wire [31:0]      dataInMem_hi_hi_80;
  assign dataInMem_hi_hi_80 = _GEN_111;
  wire [31:0]      dataInMem_hi_lo_50;
  assign dataInMem_hi_lo_50 = _GEN_111;
  wire [47:0]      dataInMem_hi_128 = {dataInMem_hi_hi_80, dataRegroupBySew_2_1_4};
  wire [31:0]      _GEN_112 = {dataRegroupBySew_4_1_5, dataRegroupBySew_3_1_5};
  wire [31:0]      dataInMem_hi_hi_81;
  assign dataInMem_hi_hi_81 = _GEN_112;
  wire [31:0]      dataInMem_hi_lo_51;
  assign dataInMem_hi_lo_51 = _GEN_112;
  wire [47:0]      dataInMem_hi_129 = {dataInMem_hi_hi_81, dataRegroupBySew_2_1_5};
  wire [31:0]      _GEN_113 = {dataRegroupBySew_4_1_6, dataRegroupBySew_3_1_6};
  wire [31:0]      dataInMem_hi_hi_82;
  assign dataInMem_hi_hi_82 = _GEN_113;
  wire [31:0]      dataInMem_hi_lo_52;
  assign dataInMem_hi_lo_52 = _GEN_113;
  wire [47:0]      dataInMem_hi_130 = {dataInMem_hi_hi_82, dataRegroupBySew_2_1_6};
  wire [31:0]      _GEN_114 = {dataRegroupBySew_4_1_7, dataRegroupBySew_3_1_7};
  wire [31:0]      dataInMem_hi_hi_83;
  assign dataInMem_hi_hi_83 = _GEN_114;
  wire [31:0]      dataInMem_hi_lo_53;
  assign dataInMem_hi_lo_53 = _GEN_114;
  wire [47:0]      dataInMem_hi_131 = {dataInMem_hi_hi_83, dataRegroupBySew_2_1_7};
  wire [159:0]     dataInMem_lo_lo_28 = {dataInMem_hi_125, dataInMem_lo_101, dataInMem_hi_124, dataInMem_lo_100};
  wire [159:0]     dataInMem_lo_hi_60 = {dataInMem_hi_127, dataInMem_lo_103, dataInMem_hi_126, dataInMem_lo_102};
  wire [319:0]     dataInMem_lo_108 = {dataInMem_lo_hi_60, dataInMem_lo_lo_28};
  wire [159:0]     dataInMem_hi_lo_44 = {dataInMem_hi_129, dataInMem_lo_105, dataInMem_hi_128, dataInMem_lo_104};
  wire [159:0]     dataInMem_hi_hi_84 = {dataInMem_hi_131, dataInMem_lo_107, dataInMem_hi_130, dataInMem_lo_106};
  wire [319:0]     dataInMem_hi_132 = {dataInMem_hi_hi_84, dataInMem_hi_lo_44};
  wire [639:0]     dataInMem_12 = {dataInMem_hi_132, dataInMem_lo_108};
  wire [127:0]     regroupCacheLine_12_0 = dataInMem_12[127:0];
  wire [127:0]     regroupCacheLine_12_1 = dataInMem_12[255:128];
  wire [127:0]     regroupCacheLine_12_2 = dataInMem_12[383:256];
  wire [127:0]     regroupCacheLine_12_3 = dataInMem_12[511:384];
  wire [127:0]     regroupCacheLine_12_4 = dataInMem_12[639:512];
  wire [127:0]     res_96 = regroupCacheLine_12_0;
  wire [127:0]     res_97 = regroupCacheLine_12_1;
  wire [127:0]     res_98 = regroupCacheLine_12_2;
  wire [127:0]     res_99 = regroupCacheLine_12_3;
  wire [127:0]     res_100 = regroupCacheLine_12_4;
  wire [255:0]     lo_lo_12 = {res_97, res_96};
  wire [255:0]     lo_hi_12 = {res_99, res_98};
  wire [511:0]     lo_12 = {lo_hi_12, lo_lo_12};
  wire [255:0]     hi_lo_12 = {128'h0, res_100};
  wire [511:0]     hi_12 = {256'h0, hi_lo_12};
  wire [1023:0]    regroupLoadData_1_4 = {hi_12, lo_12};
  wire [47:0]      dataInMem_lo_109 = {dataInMem_lo_hi_61, dataRegroupBySew_0_1_0};
  wire [31:0]      _GEN_115 = {dataRegroupBySew_5_1_0, dataRegroupBySew_4_1_0};
  wire [31:0]      dataInMem_hi_hi_85;
  assign dataInMem_hi_hi_85 = _GEN_115;
  wire [31:0]      dataInMem_hi_lo_55;
  assign dataInMem_hi_lo_55 = _GEN_115;
  wire [47:0]      dataInMem_hi_133 = {dataInMem_hi_hi_85, dataRegroupBySew_3_1_0};
  wire [47:0]      dataInMem_lo_110 = {dataInMem_lo_hi_62, dataRegroupBySew_0_1_1};
  wire [31:0]      _GEN_116 = {dataRegroupBySew_5_1_1, dataRegroupBySew_4_1_1};
  wire [31:0]      dataInMem_hi_hi_86;
  assign dataInMem_hi_hi_86 = _GEN_116;
  wire [31:0]      dataInMem_hi_lo_56;
  assign dataInMem_hi_lo_56 = _GEN_116;
  wire [47:0]      dataInMem_hi_134 = {dataInMem_hi_hi_86, dataRegroupBySew_3_1_1};
  wire [47:0]      dataInMem_lo_111 = {dataInMem_lo_hi_63, dataRegroupBySew_0_1_2};
  wire [31:0]      _GEN_117 = {dataRegroupBySew_5_1_2, dataRegroupBySew_4_1_2};
  wire [31:0]      dataInMem_hi_hi_87;
  assign dataInMem_hi_hi_87 = _GEN_117;
  wire [31:0]      dataInMem_hi_lo_57;
  assign dataInMem_hi_lo_57 = _GEN_117;
  wire [47:0]      dataInMem_hi_135 = {dataInMem_hi_hi_87, dataRegroupBySew_3_1_2};
  wire [47:0]      dataInMem_lo_112 = {dataInMem_lo_hi_64, dataRegroupBySew_0_1_3};
  wire [31:0]      _GEN_118 = {dataRegroupBySew_5_1_3, dataRegroupBySew_4_1_3};
  wire [31:0]      dataInMem_hi_hi_88;
  assign dataInMem_hi_hi_88 = _GEN_118;
  wire [31:0]      dataInMem_hi_lo_58;
  assign dataInMem_hi_lo_58 = _GEN_118;
  wire [47:0]      dataInMem_hi_136 = {dataInMem_hi_hi_88, dataRegroupBySew_3_1_3};
  wire [47:0]      dataInMem_lo_113 = {dataInMem_lo_hi_65, dataRegroupBySew_0_1_4};
  wire [31:0]      _GEN_119 = {dataRegroupBySew_5_1_4, dataRegroupBySew_4_1_4};
  wire [31:0]      dataInMem_hi_hi_89;
  assign dataInMem_hi_hi_89 = _GEN_119;
  wire [31:0]      dataInMem_hi_lo_59;
  assign dataInMem_hi_lo_59 = _GEN_119;
  wire [47:0]      dataInMem_hi_137 = {dataInMem_hi_hi_89, dataRegroupBySew_3_1_4};
  wire [47:0]      dataInMem_lo_114 = {dataInMem_lo_hi_66, dataRegroupBySew_0_1_5};
  wire [31:0]      _GEN_120 = {dataRegroupBySew_5_1_5, dataRegroupBySew_4_1_5};
  wire [31:0]      dataInMem_hi_hi_90;
  assign dataInMem_hi_hi_90 = _GEN_120;
  wire [31:0]      dataInMem_hi_lo_60;
  assign dataInMem_hi_lo_60 = _GEN_120;
  wire [47:0]      dataInMem_hi_138 = {dataInMem_hi_hi_90, dataRegroupBySew_3_1_5};
  wire [47:0]      dataInMem_lo_115 = {dataInMem_lo_hi_67, dataRegroupBySew_0_1_6};
  wire [31:0]      _GEN_121 = {dataRegroupBySew_5_1_6, dataRegroupBySew_4_1_6};
  wire [31:0]      dataInMem_hi_hi_91;
  assign dataInMem_hi_hi_91 = _GEN_121;
  wire [31:0]      dataInMem_hi_lo_61;
  assign dataInMem_hi_lo_61 = _GEN_121;
  wire [47:0]      dataInMem_hi_139 = {dataInMem_hi_hi_91, dataRegroupBySew_3_1_6};
  wire [47:0]      dataInMem_lo_116 = {dataInMem_lo_hi_68, dataRegroupBySew_0_1_7};
  wire [31:0]      _GEN_122 = {dataRegroupBySew_5_1_7, dataRegroupBySew_4_1_7};
  wire [31:0]      dataInMem_hi_hi_92;
  assign dataInMem_hi_hi_92 = _GEN_122;
  wire [31:0]      dataInMem_hi_lo_62;
  assign dataInMem_hi_lo_62 = _GEN_122;
  wire [47:0]      dataInMem_hi_140 = {dataInMem_hi_hi_92, dataRegroupBySew_3_1_7};
  wire [191:0]     dataInMem_lo_lo_29 = {dataInMem_hi_134, dataInMem_lo_110, dataInMem_hi_133, dataInMem_lo_109};
  wire [191:0]     dataInMem_lo_hi_69 = {dataInMem_hi_136, dataInMem_lo_112, dataInMem_hi_135, dataInMem_lo_111};
  wire [383:0]     dataInMem_lo_117 = {dataInMem_lo_hi_69, dataInMem_lo_lo_29};
  wire [191:0]     dataInMem_hi_lo_45 = {dataInMem_hi_138, dataInMem_lo_114, dataInMem_hi_137, dataInMem_lo_113};
  wire [191:0]     dataInMem_hi_hi_93 = {dataInMem_hi_140, dataInMem_lo_116, dataInMem_hi_139, dataInMem_lo_115};
  wire [383:0]     dataInMem_hi_141 = {dataInMem_hi_hi_93, dataInMem_hi_lo_45};
  wire [767:0]     dataInMem_13 = {dataInMem_hi_141, dataInMem_lo_117};
  wire [127:0]     regroupCacheLine_13_0 = dataInMem_13[127:0];
  wire [127:0]     regroupCacheLine_13_1 = dataInMem_13[255:128];
  wire [127:0]     regroupCacheLine_13_2 = dataInMem_13[383:256];
  wire [127:0]     regroupCacheLine_13_3 = dataInMem_13[511:384];
  wire [127:0]     regroupCacheLine_13_4 = dataInMem_13[639:512];
  wire [127:0]     regroupCacheLine_13_5 = dataInMem_13[767:640];
  wire [127:0]     res_104 = regroupCacheLine_13_0;
  wire [127:0]     res_105 = regroupCacheLine_13_1;
  wire [127:0]     res_106 = regroupCacheLine_13_2;
  wire [127:0]     res_107 = regroupCacheLine_13_3;
  wire [127:0]     res_108 = regroupCacheLine_13_4;
  wire [127:0]     res_109 = regroupCacheLine_13_5;
  wire [255:0]     lo_lo_13 = {res_105, res_104};
  wire [255:0]     lo_hi_13 = {res_107, res_106};
  wire [511:0]     lo_13 = {lo_hi_13, lo_lo_13};
  wire [255:0]     hi_lo_13 = {res_109, res_108};
  wire [511:0]     hi_13 = {256'h0, hi_lo_13};
  wire [1023:0]    regroupLoadData_1_5 = {hi_13, lo_13};
  wire [47:0]      dataInMem_lo_118 = {dataInMem_lo_hi_70, dataRegroupBySew_0_1_0};
  wire [31:0]      dataInMem_hi_hi_94 = {dataRegroupBySew_6_1_0, dataRegroupBySew_5_1_0};
  wire [63:0]      dataInMem_hi_142 = {dataInMem_hi_hi_94, dataInMem_hi_lo_46};
  wire [47:0]      dataInMem_lo_119 = {dataInMem_lo_hi_71, dataRegroupBySew_0_1_1};
  wire [31:0]      dataInMem_hi_hi_95 = {dataRegroupBySew_6_1_1, dataRegroupBySew_5_1_1};
  wire [63:0]      dataInMem_hi_143 = {dataInMem_hi_hi_95, dataInMem_hi_lo_47};
  wire [47:0]      dataInMem_lo_120 = {dataInMem_lo_hi_72, dataRegroupBySew_0_1_2};
  wire [31:0]      dataInMem_hi_hi_96 = {dataRegroupBySew_6_1_2, dataRegroupBySew_5_1_2};
  wire [63:0]      dataInMem_hi_144 = {dataInMem_hi_hi_96, dataInMem_hi_lo_48};
  wire [47:0]      dataInMem_lo_121 = {dataInMem_lo_hi_73, dataRegroupBySew_0_1_3};
  wire [31:0]      dataInMem_hi_hi_97 = {dataRegroupBySew_6_1_3, dataRegroupBySew_5_1_3};
  wire [63:0]      dataInMem_hi_145 = {dataInMem_hi_hi_97, dataInMem_hi_lo_49};
  wire [47:0]      dataInMem_lo_122 = {dataInMem_lo_hi_74, dataRegroupBySew_0_1_4};
  wire [31:0]      dataInMem_hi_hi_98 = {dataRegroupBySew_6_1_4, dataRegroupBySew_5_1_4};
  wire [63:0]      dataInMem_hi_146 = {dataInMem_hi_hi_98, dataInMem_hi_lo_50};
  wire [47:0]      dataInMem_lo_123 = {dataInMem_lo_hi_75, dataRegroupBySew_0_1_5};
  wire [31:0]      dataInMem_hi_hi_99 = {dataRegroupBySew_6_1_5, dataRegroupBySew_5_1_5};
  wire [63:0]      dataInMem_hi_147 = {dataInMem_hi_hi_99, dataInMem_hi_lo_51};
  wire [47:0]      dataInMem_lo_124 = {dataInMem_lo_hi_76, dataRegroupBySew_0_1_6};
  wire [31:0]      dataInMem_hi_hi_100 = {dataRegroupBySew_6_1_6, dataRegroupBySew_5_1_6};
  wire [63:0]      dataInMem_hi_148 = {dataInMem_hi_hi_100, dataInMem_hi_lo_52};
  wire [47:0]      dataInMem_lo_125 = {dataInMem_lo_hi_77, dataRegroupBySew_0_1_7};
  wire [31:0]      dataInMem_hi_hi_101 = {dataRegroupBySew_6_1_7, dataRegroupBySew_5_1_7};
  wire [63:0]      dataInMem_hi_149 = {dataInMem_hi_hi_101, dataInMem_hi_lo_53};
  wire [223:0]     dataInMem_lo_lo_30 = {dataInMem_hi_143, dataInMem_lo_119, dataInMem_hi_142, dataInMem_lo_118};
  wire [223:0]     dataInMem_lo_hi_78 = {dataInMem_hi_145, dataInMem_lo_121, dataInMem_hi_144, dataInMem_lo_120};
  wire [447:0]     dataInMem_lo_126 = {dataInMem_lo_hi_78, dataInMem_lo_lo_30};
  wire [223:0]     dataInMem_hi_lo_54 = {dataInMem_hi_147, dataInMem_lo_123, dataInMem_hi_146, dataInMem_lo_122};
  wire [223:0]     dataInMem_hi_hi_102 = {dataInMem_hi_149, dataInMem_lo_125, dataInMem_hi_148, dataInMem_lo_124};
  wire [447:0]     dataInMem_hi_150 = {dataInMem_hi_hi_102, dataInMem_hi_lo_54};
  wire [895:0]     dataInMem_14 = {dataInMem_hi_150, dataInMem_lo_126};
  wire [127:0]     regroupCacheLine_14_0 = dataInMem_14[127:0];
  wire [127:0]     regroupCacheLine_14_1 = dataInMem_14[255:128];
  wire [127:0]     regroupCacheLine_14_2 = dataInMem_14[383:256];
  wire [127:0]     regroupCacheLine_14_3 = dataInMem_14[511:384];
  wire [127:0]     regroupCacheLine_14_4 = dataInMem_14[639:512];
  wire [127:0]     regroupCacheLine_14_5 = dataInMem_14[767:640];
  wire [127:0]     regroupCacheLine_14_6 = dataInMem_14[895:768];
  wire [127:0]     res_112 = regroupCacheLine_14_0;
  wire [127:0]     res_113 = regroupCacheLine_14_1;
  wire [127:0]     res_114 = regroupCacheLine_14_2;
  wire [127:0]     res_115 = regroupCacheLine_14_3;
  wire [127:0]     res_116 = regroupCacheLine_14_4;
  wire [127:0]     res_117 = regroupCacheLine_14_5;
  wire [127:0]     res_118 = regroupCacheLine_14_6;
  wire [255:0]     lo_lo_14 = {res_113, res_112};
  wire [255:0]     lo_hi_14 = {res_115, res_114};
  wire [511:0]     lo_14 = {lo_hi_14, lo_lo_14};
  wire [255:0]     hi_lo_14 = {res_117, res_116};
  wire [255:0]     hi_hi_14 = {128'h0, res_118};
  wire [511:0]     hi_14 = {hi_hi_14, hi_lo_14};
  wire [1023:0]    regroupLoadData_1_6 = {hi_14, lo_14};
  wire [63:0]      dataInMem_lo_127 = {dataInMem_lo_hi_79, dataInMem_lo_lo_31};
  wire [31:0]      dataInMem_hi_hi_103 = {dataRegroupBySew_7_1_0, dataRegroupBySew_6_1_0};
  wire [63:0]      dataInMem_hi_151 = {dataInMem_hi_hi_103, dataInMem_hi_lo_55};
  wire [63:0]      dataInMem_lo_128 = {dataInMem_lo_hi_80, dataInMem_lo_lo_32};
  wire [31:0]      dataInMem_hi_hi_104 = {dataRegroupBySew_7_1_1, dataRegroupBySew_6_1_1};
  wire [63:0]      dataInMem_hi_152 = {dataInMem_hi_hi_104, dataInMem_hi_lo_56};
  wire [63:0]      dataInMem_lo_129 = {dataInMem_lo_hi_81, dataInMem_lo_lo_33};
  wire [31:0]      dataInMem_hi_hi_105 = {dataRegroupBySew_7_1_2, dataRegroupBySew_6_1_2};
  wire [63:0]      dataInMem_hi_153 = {dataInMem_hi_hi_105, dataInMem_hi_lo_57};
  wire [63:0]      dataInMem_lo_130 = {dataInMem_lo_hi_82, dataInMem_lo_lo_34};
  wire [31:0]      dataInMem_hi_hi_106 = {dataRegroupBySew_7_1_3, dataRegroupBySew_6_1_3};
  wire [63:0]      dataInMem_hi_154 = {dataInMem_hi_hi_106, dataInMem_hi_lo_58};
  wire [63:0]      dataInMem_lo_131 = {dataInMem_lo_hi_83, dataInMem_lo_lo_35};
  wire [31:0]      dataInMem_hi_hi_107 = {dataRegroupBySew_7_1_4, dataRegroupBySew_6_1_4};
  wire [63:0]      dataInMem_hi_155 = {dataInMem_hi_hi_107, dataInMem_hi_lo_59};
  wire [63:0]      dataInMem_lo_132 = {dataInMem_lo_hi_84, dataInMem_lo_lo_36};
  wire [31:0]      dataInMem_hi_hi_108 = {dataRegroupBySew_7_1_5, dataRegroupBySew_6_1_5};
  wire [63:0]      dataInMem_hi_156 = {dataInMem_hi_hi_108, dataInMem_hi_lo_60};
  wire [63:0]      dataInMem_lo_133 = {dataInMem_lo_hi_85, dataInMem_lo_lo_37};
  wire [31:0]      dataInMem_hi_hi_109 = {dataRegroupBySew_7_1_6, dataRegroupBySew_6_1_6};
  wire [63:0]      dataInMem_hi_157 = {dataInMem_hi_hi_109, dataInMem_hi_lo_61};
  wire [63:0]      dataInMem_lo_134 = {dataInMem_lo_hi_86, dataInMem_lo_lo_38};
  wire [31:0]      dataInMem_hi_hi_110 = {dataRegroupBySew_7_1_7, dataRegroupBySew_6_1_7};
  wire [63:0]      dataInMem_hi_158 = {dataInMem_hi_hi_110, dataInMem_hi_lo_62};
  wire [255:0]     dataInMem_lo_lo_39 = {dataInMem_hi_152, dataInMem_lo_128, dataInMem_hi_151, dataInMem_lo_127};
  wire [255:0]     dataInMem_lo_hi_87 = {dataInMem_hi_154, dataInMem_lo_130, dataInMem_hi_153, dataInMem_lo_129};
  wire [511:0]     dataInMem_lo_135 = {dataInMem_lo_hi_87, dataInMem_lo_lo_39};
  wire [255:0]     dataInMem_hi_lo_63 = {dataInMem_hi_156, dataInMem_lo_132, dataInMem_hi_155, dataInMem_lo_131};
  wire [255:0]     dataInMem_hi_hi_111 = {dataInMem_hi_158, dataInMem_lo_134, dataInMem_hi_157, dataInMem_lo_133};
  wire [511:0]     dataInMem_hi_159 = {dataInMem_hi_hi_111, dataInMem_hi_lo_63};
  wire [1023:0]    dataInMem_15 = {dataInMem_hi_159, dataInMem_lo_135};
  wire [127:0]     regroupCacheLine_15_0 = dataInMem_15[127:0];
  wire [127:0]     regroupCacheLine_15_1 = dataInMem_15[255:128];
  wire [127:0]     regroupCacheLine_15_2 = dataInMem_15[383:256];
  wire [127:0]     regroupCacheLine_15_3 = dataInMem_15[511:384];
  wire [127:0]     regroupCacheLine_15_4 = dataInMem_15[639:512];
  wire [127:0]     regroupCacheLine_15_5 = dataInMem_15[767:640];
  wire [127:0]     regroupCacheLine_15_6 = dataInMem_15[895:768];
  wire [127:0]     regroupCacheLine_15_7 = dataInMem_15[1023:896];
  wire [127:0]     res_120 = regroupCacheLine_15_0;
  wire [127:0]     res_121 = regroupCacheLine_15_1;
  wire [127:0]     res_122 = regroupCacheLine_15_2;
  wire [127:0]     res_123 = regroupCacheLine_15_3;
  wire [127:0]     res_124 = regroupCacheLine_15_4;
  wire [127:0]     res_125 = regroupCacheLine_15_5;
  wire [127:0]     res_126 = regroupCacheLine_15_6;
  wire [127:0]     res_127 = regroupCacheLine_15_7;
  wire [255:0]     lo_lo_15 = {res_121, res_120};
  wire [255:0]     lo_hi_15 = {res_123, res_122};
  wire [511:0]     lo_15 = {lo_hi_15, lo_lo_15};
  wire [255:0]     hi_lo_15 = {res_125, res_124};
  wire [255:0]     hi_hi_15 = {res_127, res_126};
  wire [511:0]     hi_15 = {hi_hi_15, hi_lo_15};
  wire [1023:0]    regroupLoadData_1_7 = {hi_15, lo_15};
  wire [31:0]      dataRegroupBySew_0_2_0 = bufferStageEnqueueData_0[31:0];
  wire [31:0]      dataRegroupBySew_0_2_1 = bufferStageEnqueueData_0[63:32];
  wire [31:0]      dataRegroupBySew_0_2_2 = bufferStageEnqueueData_0[95:64];
  wire [31:0]      dataRegroupBySew_0_2_3 = bufferStageEnqueueData_0[127:96];
  wire [31:0]      dataRegroupBySew_1_2_0 = bufferStageEnqueueData_1[31:0];
  wire [31:0]      dataRegroupBySew_1_2_1 = bufferStageEnqueueData_1[63:32];
  wire [31:0]      dataRegroupBySew_1_2_2 = bufferStageEnqueueData_1[95:64];
  wire [31:0]      dataRegroupBySew_1_2_3 = bufferStageEnqueueData_1[127:96];
  wire [31:0]      dataRegroupBySew_2_2_0 = bufferStageEnqueueData_2[31:0];
  wire [31:0]      dataRegroupBySew_2_2_1 = bufferStageEnqueueData_2[63:32];
  wire [31:0]      dataRegroupBySew_2_2_2 = bufferStageEnqueueData_2[95:64];
  wire [31:0]      dataRegroupBySew_2_2_3 = bufferStageEnqueueData_2[127:96];
  wire [31:0]      dataRegroupBySew_3_2_0 = bufferStageEnqueueData_3[31:0];
  wire [31:0]      dataRegroupBySew_3_2_1 = bufferStageEnqueueData_3[63:32];
  wire [31:0]      dataRegroupBySew_3_2_2 = bufferStageEnqueueData_3[95:64];
  wire [31:0]      dataRegroupBySew_3_2_3 = bufferStageEnqueueData_3[127:96];
  wire [31:0]      dataRegroupBySew_4_2_0 = bufferStageEnqueueData_4[31:0];
  wire [31:0]      dataRegroupBySew_4_2_1 = bufferStageEnqueueData_4[63:32];
  wire [31:0]      dataRegroupBySew_4_2_2 = bufferStageEnqueueData_4[95:64];
  wire [31:0]      dataRegroupBySew_4_2_3 = bufferStageEnqueueData_4[127:96];
  wire [31:0]      dataRegroupBySew_5_2_0 = bufferStageEnqueueData_5[31:0];
  wire [31:0]      dataRegroupBySew_5_2_1 = bufferStageEnqueueData_5[63:32];
  wire [31:0]      dataRegroupBySew_5_2_2 = bufferStageEnqueueData_5[95:64];
  wire [31:0]      dataRegroupBySew_5_2_3 = bufferStageEnqueueData_5[127:96];
  wire [31:0]      dataRegroupBySew_6_2_0 = bufferStageEnqueueData_6[31:0];
  wire [31:0]      dataRegroupBySew_6_2_1 = bufferStageEnqueueData_6[63:32];
  wire [31:0]      dataRegroupBySew_6_2_2 = bufferStageEnqueueData_6[95:64];
  wire [31:0]      dataRegroupBySew_6_2_3 = bufferStageEnqueueData_6[127:96];
  wire [31:0]      dataRegroupBySew_7_2_0 = bufferStageEnqueueData_7[31:0];
  wire [31:0]      dataRegroupBySew_7_2_1 = bufferStageEnqueueData_7[63:32];
  wire [31:0]      dataRegroupBySew_7_2_2 = bufferStageEnqueueData_7[95:64];
  wire [31:0]      dataRegroupBySew_7_2_3 = bufferStageEnqueueData_7[127:96];
  wire [63:0]      dataInMem_lo_136 = {dataRegroupBySew_0_2_1, dataRegroupBySew_0_2_0};
  wire [63:0]      dataInMem_hi_160 = {dataRegroupBySew_0_2_3, dataRegroupBySew_0_2_2};
  wire [127:0]     dataInMem_16 = {dataInMem_hi_160, dataInMem_lo_136};
  wire [127:0]     regroupCacheLine_16_0 = dataInMem_16;
  wire [127:0]     res_128 = regroupCacheLine_16_0;
  wire [255:0]     lo_lo_16 = {128'h0, res_128};
  wire [511:0]     lo_16 = {256'h0, lo_lo_16};
  wire [1023:0]    regroupLoadData_2_0 = {512'h0, lo_16};
  wire [127:0]     dataInMem_lo_137 = {dataRegroupBySew_1_2_1, dataRegroupBySew_0_2_1, dataRegroupBySew_1_2_0, dataRegroupBySew_0_2_0};
  wire [127:0]     dataInMem_hi_161 = {dataRegroupBySew_1_2_3, dataRegroupBySew_0_2_3, dataRegroupBySew_1_2_2, dataRegroupBySew_0_2_2};
  wire [255:0]     dataInMem_17 = {dataInMem_hi_161, dataInMem_lo_137};
  wire [127:0]     regroupCacheLine_17_0 = dataInMem_17[127:0];
  wire [127:0]     regroupCacheLine_17_1 = dataInMem_17[255:128];
  wire [127:0]     res_136 = regroupCacheLine_17_0;
  wire [127:0]     res_137 = regroupCacheLine_17_1;
  wire [255:0]     lo_lo_17 = {res_137, res_136};
  wire [511:0]     lo_17 = {256'h0, lo_lo_17};
  wire [1023:0]    regroupLoadData_2_1 = {512'h0, lo_17};
  wire [63:0]      _GEN_123 = {dataRegroupBySew_2_2_0, dataRegroupBySew_1_2_0};
  wire [63:0]      dataInMem_hi_162;
  assign dataInMem_hi_162 = _GEN_123;
  wire [63:0]      dataInMem_lo_hi_88;
  assign dataInMem_lo_hi_88 = _GEN_123;
  wire [63:0]      dataInMem_lo_hi_92;
  assign dataInMem_lo_hi_92 = _GEN_123;
  wire [63:0]      _GEN_124 = {dataRegroupBySew_2_2_1, dataRegroupBySew_1_2_1};
  wire [63:0]      dataInMem_hi_163;
  assign dataInMem_hi_163 = _GEN_124;
  wire [63:0]      dataInMem_lo_hi_89;
  assign dataInMem_lo_hi_89 = _GEN_124;
  wire [63:0]      dataInMem_lo_hi_93;
  assign dataInMem_lo_hi_93 = _GEN_124;
  wire [63:0]      _GEN_125 = {dataRegroupBySew_2_2_2, dataRegroupBySew_1_2_2};
  wire [63:0]      dataInMem_hi_164;
  assign dataInMem_hi_164 = _GEN_125;
  wire [63:0]      dataInMem_lo_hi_90;
  assign dataInMem_lo_hi_90 = _GEN_125;
  wire [63:0]      dataInMem_lo_hi_94;
  assign dataInMem_lo_hi_94 = _GEN_125;
  wire [63:0]      _GEN_126 = {dataRegroupBySew_2_2_3, dataRegroupBySew_1_2_3};
  wire [63:0]      dataInMem_hi_165;
  assign dataInMem_hi_165 = _GEN_126;
  wire [63:0]      dataInMem_lo_hi_91;
  assign dataInMem_lo_hi_91 = _GEN_126;
  wire [63:0]      dataInMem_lo_hi_95;
  assign dataInMem_lo_hi_95 = _GEN_126;
  wire [191:0]     dataInMem_lo_138 = {dataInMem_hi_163, dataRegroupBySew_0_2_1, dataInMem_hi_162, dataRegroupBySew_0_2_0};
  wire [191:0]     dataInMem_hi_166 = {dataInMem_hi_165, dataRegroupBySew_0_2_3, dataInMem_hi_164, dataRegroupBySew_0_2_2};
  wire [383:0]     dataInMem_18 = {dataInMem_hi_166, dataInMem_lo_138};
  wire [127:0]     regroupCacheLine_18_0 = dataInMem_18[127:0];
  wire [127:0]     regroupCacheLine_18_1 = dataInMem_18[255:128];
  wire [127:0]     regroupCacheLine_18_2 = dataInMem_18[383:256];
  wire [127:0]     res_144 = regroupCacheLine_18_0;
  wire [127:0]     res_145 = regroupCacheLine_18_1;
  wire [127:0]     res_146 = regroupCacheLine_18_2;
  wire [255:0]     lo_lo_18 = {res_145, res_144};
  wire [255:0]     lo_hi_18 = {128'h0, res_146};
  wire [511:0]     lo_18 = {lo_hi_18, lo_lo_18};
  wire [1023:0]    regroupLoadData_2_2 = {512'h0, lo_18};
  wire [63:0]      _GEN_127 = {dataRegroupBySew_1_2_0, dataRegroupBySew_0_2_0};
  wire [63:0]      dataInMem_lo_139;
  assign dataInMem_lo_139 = _GEN_127;
  wire [63:0]      dataInMem_lo_144;
  assign dataInMem_lo_144 = _GEN_127;
  wire [63:0]      dataInMem_lo_lo_40;
  assign dataInMem_lo_lo_40 = _GEN_127;
  wire [63:0]      _GEN_128 = {dataRegroupBySew_3_2_0, dataRegroupBySew_2_2_0};
  wire [63:0]      dataInMem_hi_167;
  assign dataInMem_hi_167 = _GEN_128;
  wire [63:0]      dataInMem_lo_hi_96;
  assign dataInMem_lo_hi_96 = _GEN_128;
  wire [63:0]      _GEN_129 = {dataRegroupBySew_1_2_1, dataRegroupBySew_0_2_1};
  wire [63:0]      dataInMem_lo_140;
  assign dataInMem_lo_140 = _GEN_129;
  wire [63:0]      dataInMem_lo_145;
  assign dataInMem_lo_145 = _GEN_129;
  wire [63:0]      dataInMem_lo_lo_41;
  assign dataInMem_lo_lo_41 = _GEN_129;
  wire [63:0]      _GEN_130 = {dataRegroupBySew_3_2_1, dataRegroupBySew_2_2_1};
  wire [63:0]      dataInMem_hi_168;
  assign dataInMem_hi_168 = _GEN_130;
  wire [63:0]      dataInMem_lo_hi_97;
  assign dataInMem_lo_hi_97 = _GEN_130;
  wire [63:0]      _GEN_131 = {dataRegroupBySew_1_2_2, dataRegroupBySew_0_2_2};
  wire [63:0]      dataInMem_lo_141;
  assign dataInMem_lo_141 = _GEN_131;
  wire [63:0]      dataInMem_lo_146;
  assign dataInMem_lo_146 = _GEN_131;
  wire [63:0]      dataInMem_lo_lo_42;
  assign dataInMem_lo_lo_42 = _GEN_131;
  wire [63:0]      _GEN_132 = {dataRegroupBySew_3_2_2, dataRegroupBySew_2_2_2};
  wire [63:0]      dataInMem_hi_169;
  assign dataInMem_hi_169 = _GEN_132;
  wire [63:0]      dataInMem_lo_hi_98;
  assign dataInMem_lo_hi_98 = _GEN_132;
  wire [63:0]      _GEN_133 = {dataRegroupBySew_1_2_3, dataRegroupBySew_0_2_3};
  wire [63:0]      dataInMem_lo_142;
  assign dataInMem_lo_142 = _GEN_133;
  wire [63:0]      dataInMem_lo_147;
  assign dataInMem_lo_147 = _GEN_133;
  wire [63:0]      dataInMem_lo_lo_43;
  assign dataInMem_lo_lo_43 = _GEN_133;
  wire [63:0]      _GEN_134 = {dataRegroupBySew_3_2_3, dataRegroupBySew_2_2_3};
  wire [63:0]      dataInMem_hi_170;
  assign dataInMem_hi_170 = _GEN_134;
  wire [63:0]      dataInMem_lo_hi_99;
  assign dataInMem_lo_hi_99 = _GEN_134;
  wire [255:0]     dataInMem_lo_143 = {dataInMem_hi_168, dataInMem_lo_140, dataInMem_hi_167, dataInMem_lo_139};
  wire [255:0]     dataInMem_hi_171 = {dataInMem_hi_170, dataInMem_lo_142, dataInMem_hi_169, dataInMem_lo_141};
  wire [511:0]     dataInMem_19 = {dataInMem_hi_171, dataInMem_lo_143};
  wire [127:0]     regroupCacheLine_19_0 = dataInMem_19[127:0];
  wire [127:0]     regroupCacheLine_19_1 = dataInMem_19[255:128];
  wire [127:0]     regroupCacheLine_19_2 = dataInMem_19[383:256];
  wire [127:0]     regroupCacheLine_19_3 = dataInMem_19[511:384];
  wire [127:0]     res_152 = regroupCacheLine_19_0;
  wire [127:0]     res_153 = regroupCacheLine_19_1;
  wire [127:0]     res_154 = regroupCacheLine_19_2;
  wire [127:0]     res_155 = regroupCacheLine_19_3;
  wire [255:0]     lo_lo_19 = {res_153, res_152};
  wire [255:0]     lo_hi_19 = {res_155, res_154};
  wire [511:0]     lo_19 = {lo_hi_19, lo_lo_19};
  wire [1023:0]    regroupLoadData_2_3 = {512'h0, lo_19};
  wire [63:0]      _GEN_135 = {dataRegroupBySew_4_2_0, dataRegroupBySew_3_2_0};
  wire [63:0]      dataInMem_hi_hi_112;
  assign dataInMem_hi_hi_112 = _GEN_135;
  wire [63:0]      dataInMem_hi_lo_64;
  assign dataInMem_hi_lo_64 = _GEN_135;
  wire [95:0]      dataInMem_hi_172 = {dataInMem_hi_hi_112, dataRegroupBySew_2_2_0};
  wire [63:0]      _GEN_136 = {dataRegroupBySew_4_2_1, dataRegroupBySew_3_2_1};
  wire [63:0]      dataInMem_hi_hi_113;
  assign dataInMem_hi_hi_113 = _GEN_136;
  wire [63:0]      dataInMem_hi_lo_65;
  assign dataInMem_hi_lo_65 = _GEN_136;
  wire [95:0]      dataInMem_hi_173 = {dataInMem_hi_hi_113, dataRegroupBySew_2_2_1};
  wire [63:0]      _GEN_137 = {dataRegroupBySew_4_2_2, dataRegroupBySew_3_2_2};
  wire [63:0]      dataInMem_hi_hi_114;
  assign dataInMem_hi_hi_114 = _GEN_137;
  wire [63:0]      dataInMem_hi_lo_66;
  assign dataInMem_hi_lo_66 = _GEN_137;
  wire [95:0]      dataInMem_hi_174 = {dataInMem_hi_hi_114, dataRegroupBySew_2_2_2};
  wire [63:0]      _GEN_138 = {dataRegroupBySew_4_2_3, dataRegroupBySew_3_2_3};
  wire [63:0]      dataInMem_hi_hi_115;
  assign dataInMem_hi_hi_115 = _GEN_138;
  wire [63:0]      dataInMem_hi_lo_67;
  assign dataInMem_hi_lo_67 = _GEN_138;
  wire [95:0]      dataInMem_hi_175 = {dataInMem_hi_hi_115, dataRegroupBySew_2_2_3};
  wire [319:0]     dataInMem_lo_148 = {dataInMem_hi_173, dataInMem_lo_145, dataInMem_hi_172, dataInMem_lo_144};
  wire [319:0]     dataInMem_hi_176 = {dataInMem_hi_175, dataInMem_lo_147, dataInMem_hi_174, dataInMem_lo_146};
  wire [639:0]     dataInMem_20 = {dataInMem_hi_176, dataInMem_lo_148};
  wire [127:0]     regroupCacheLine_20_0 = dataInMem_20[127:0];
  wire [127:0]     regroupCacheLine_20_1 = dataInMem_20[255:128];
  wire [127:0]     regroupCacheLine_20_2 = dataInMem_20[383:256];
  wire [127:0]     regroupCacheLine_20_3 = dataInMem_20[511:384];
  wire [127:0]     regroupCacheLine_20_4 = dataInMem_20[639:512];
  wire [127:0]     res_160 = regroupCacheLine_20_0;
  wire [127:0]     res_161 = regroupCacheLine_20_1;
  wire [127:0]     res_162 = regroupCacheLine_20_2;
  wire [127:0]     res_163 = regroupCacheLine_20_3;
  wire [127:0]     res_164 = regroupCacheLine_20_4;
  wire [255:0]     lo_lo_20 = {res_161, res_160};
  wire [255:0]     lo_hi_20 = {res_163, res_162};
  wire [511:0]     lo_20 = {lo_hi_20, lo_lo_20};
  wire [255:0]     hi_lo_20 = {128'h0, res_164};
  wire [511:0]     hi_20 = {256'h0, hi_lo_20};
  wire [1023:0]    regroupLoadData_2_4 = {hi_20, lo_20};
  wire [95:0]      dataInMem_lo_149 = {dataInMem_lo_hi_88, dataRegroupBySew_0_2_0};
  wire [63:0]      _GEN_139 = {dataRegroupBySew_5_2_0, dataRegroupBySew_4_2_0};
  wire [63:0]      dataInMem_hi_hi_116;
  assign dataInMem_hi_hi_116 = _GEN_139;
  wire [63:0]      dataInMem_hi_lo_68;
  assign dataInMem_hi_lo_68 = _GEN_139;
  wire [95:0]      dataInMem_hi_177 = {dataInMem_hi_hi_116, dataRegroupBySew_3_2_0};
  wire [95:0]      dataInMem_lo_150 = {dataInMem_lo_hi_89, dataRegroupBySew_0_2_1};
  wire [63:0]      _GEN_140 = {dataRegroupBySew_5_2_1, dataRegroupBySew_4_2_1};
  wire [63:0]      dataInMem_hi_hi_117;
  assign dataInMem_hi_hi_117 = _GEN_140;
  wire [63:0]      dataInMem_hi_lo_69;
  assign dataInMem_hi_lo_69 = _GEN_140;
  wire [95:0]      dataInMem_hi_178 = {dataInMem_hi_hi_117, dataRegroupBySew_3_2_1};
  wire [95:0]      dataInMem_lo_151 = {dataInMem_lo_hi_90, dataRegroupBySew_0_2_2};
  wire [63:0]      _GEN_141 = {dataRegroupBySew_5_2_2, dataRegroupBySew_4_2_2};
  wire [63:0]      dataInMem_hi_hi_118;
  assign dataInMem_hi_hi_118 = _GEN_141;
  wire [63:0]      dataInMem_hi_lo_70;
  assign dataInMem_hi_lo_70 = _GEN_141;
  wire [95:0]      dataInMem_hi_179 = {dataInMem_hi_hi_118, dataRegroupBySew_3_2_2};
  wire [95:0]      dataInMem_lo_152 = {dataInMem_lo_hi_91, dataRegroupBySew_0_2_3};
  wire [63:0]      _GEN_142 = {dataRegroupBySew_5_2_3, dataRegroupBySew_4_2_3};
  wire [63:0]      dataInMem_hi_hi_119;
  assign dataInMem_hi_hi_119 = _GEN_142;
  wire [63:0]      dataInMem_hi_lo_71;
  assign dataInMem_hi_lo_71 = _GEN_142;
  wire [95:0]      dataInMem_hi_180 = {dataInMem_hi_hi_119, dataRegroupBySew_3_2_3};
  wire [383:0]     dataInMem_lo_153 = {dataInMem_hi_178, dataInMem_lo_150, dataInMem_hi_177, dataInMem_lo_149};
  wire [383:0]     dataInMem_hi_181 = {dataInMem_hi_180, dataInMem_lo_152, dataInMem_hi_179, dataInMem_lo_151};
  wire [767:0]     dataInMem_21 = {dataInMem_hi_181, dataInMem_lo_153};
  wire [127:0]     regroupCacheLine_21_0 = dataInMem_21[127:0];
  wire [127:0]     regroupCacheLine_21_1 = dataInMem_21[255:128];
  wire [127:0]     regroupCacheLine_21_2 = dataInMem_21[383:256];
  wire [127:0]     regroupCacheLine_21_3 = dataInMem_21[511:384];
  wire [127:0]     regroupCacheLine_21_4 = dataInMem_21[639:512];
  wire [127:0]     regroupCacheLine_21_5 = dataInMem_21[767:640];
  wire [127:0]     res_168 = regroupCacheLine_21_0;
  wire [127:0]     res_169 = regroupCacheLine_21_1;
  wire [127:0]     res_170 = regroupCacheLine_21_2;
  wire [127:0]     res_171 = regroupCacheLine_21_3;
  wire [127:0]     res_172 = regroupCacheLine_21_4;
  wire [127:0]     res_173 = regroupCacheLine_21_5;
  wire [255:0]     lo_lo_21 = {res_169, res_168};
  wire [255:0]     lo_hi_21 = {res_171, res_170};
  wire [511:0]     lo_21 = {lo_hi_21, lo_lo_21};
  wire [255:0]     hi_lo_21 = {res_173, res_172};
  wire [511:0]     hi_21 = {256'h0, hi_lo_21};
  wire [1023:0]    regroupLoadData_2_5 = {hi_21, lo_21};
  wire [95:0]      dataInMem_lo_154 = {dataInMem_lo_hi_92, dataRegroupBySew_0_2_0};
  wire [63:0]      dataInMem_hi_hi_120 = {dataRegroupBySew_6_2_0, dataRegroupBySew_5_2_0};
  wire [127:0]     dataInMem_hi_182 = {dataInMem_hi_hi_120, dataInMem_hi_lo_64};
  wire [95:0]      dataInMem_lo_155 = {dataInMem_lo_hi_93, dataRegroupBySew_0_2_1};
  wire [63:0]      dataInMem_hi_hi_121 = {dataRegroupBySew_6_2_1, dataRegroupBySew_5_2_1};
  wire [127:0]     dataInMem_hi_183 = {dataInMem_hi_hi_121, dataInMem_hi_lo_65};
  wire [95:0]      dataInMem_lo_156 = {dataInMem_lo_hi_94, dataRegroupBySew_0_2_2};
  wire [63:0]      dataInMem_hi_hi_122 = {dataRegroupBySew_6_2_2, dataRegroupBySew_5_2_2};
  wire [127:0]     dataInMem_hi_184 = {dataInMem_hi_hi_122, dataInMem_hi_lo_66};
  wire [95:0]      dataInMem_lo_157 = {dataInMem_lo_hi_95, dataRegroupBySew_0_2_3};
  wire [63:0]      dataInMem_hi_hi_123 = {dataRegroupBySew_6_2_3, dataRegroupBySew_5_2_3};
  wire [127:0]     dataInMem_hi_185 = {dataInMem_hi_hi_123, dataInMem_hi_lo_67};
  wire [447:0]     dataInMem_lo_158 = {dataInMem_hi_183, dataInMem_lo_155, dataInMem_hi_182, dataInMem_lo_154};
  wire [447:0]     dataInMem_hi_186 = {dataInMem_hi_185, dataInMem_lo_157, dataInMem_hi_184, dataInMem_lo_156};
  wire [895:0]     dataInMem_22 = {dataInMem_hi_186, dataInMem_lo_158};
  wire [127:0]     regroupCacheLine_22_0 = dataInMem_22[127:0];
  wire [127:0]     regroupCacheLine_22_1 = dataInMem_22[255:128];
  wire [127:0]     regroupCacheLine_22_2 = dataInMem_22[383:256];
  wire [127:0]     regroupCacheLine_22_3 = dataInMem_22[511:384];
  wire [127:0]     regroupCacheLine_22_4 = dataInMem_22[639:512];
  wire [127:0]     regroupCacheLine_22_5 = dataInMem_22[767:640];
  wire [127:0]     regroupCacheLine_22_6 = dataInMem_22[895:768];
  wire [127:0]     res_176 = regroupCacheLine_22_0;
  wire [127:0]     res_177 = regroupCacheLine_22_1;
  wire [127:0]     res_178 = regroupCacheLine_22_2;
  wire [127:0]     res_179 = regroupCacheLine_22_3;
  wire [127:0]     res_180 = regroupCacheLine_22_4;
  wire [127:0]     res_181 = regroupCacheLine_22_5;
  wire [127:0]     res_182 = regroupCacheLine_22_6;
  wire [255:0]     lo_lo_22 = {res_177, res_176};
  wire [255:0]     lo_hi_22 = {res_179, res_178};
  wire [511:0]     lo_22 = {lo_hi_22, lo_lo_22};
  wire [255:0]     hi_lo_22 = {res_181, res_180};
  wire [255:0]     hi_hi_22 = {128'h0, res_182};
  wire [511:0]     hi_22 = {hi_hi_22, hi_lo_22};
  wire [1023:0]    regroupLoadData_2_6 = {hi_22, lo_22};
  wire [127:0]     dataInMem_lo_159 = {dataInMem_lo_hi_96, dataInMem_lo_lo_40};
  wire [63:0]      dataInMem_hi_hi_124 = {dataRegroupBySew_7_2_0, dataRegroupBySew_6_2_0};
  wire [127:0]     dataInMem_hi_187 = {dataInMem_hi_hi_124, dataInMem_hi_lo_68};
  wire [127:0]     dataInMem_lo_160 = {dataInMem_lo_hi_97, dataInMem_lo_lo_41};
  wire [63:0]      dataInMem_hi_hi_125 = {dataRegroupBySew_7_2_1, dataRegroupBySew_6_2_1};
  wire [127:0]     dataInMem_hi_188 = {dataInMem_hi_hi_125, dataInMem_hi_lo_69};
  wire [127:0]     dataInMem_lo_161 = {dataInMem_lo_hi_98, dataInMem_lo_lo_42};
  wire [63:0]      dataInMem_hi_hi_126 = {dataRegroupBySew_7_2_2, dataRegroupBySew_6_2_2};
  wire [127:0]     dataInMem_hi_189 = {dataInMem_hi_hi_126, dataInMem_hi_lo_70};
  wire [127:0]     dataInMem_lo_162 = {dataInMem_lo_hi_99, dataInMem_lo_lo_43};
  wire [63:0]      dataInMem_hi_hi_127 = {dataRegroupBySew_7_2_3, dataRegroupBySew_6_2_3};
  wire [127:0]     dataInMem_hi_190 = {dataInMem_hi_hi_127, dataInMem_hi_lo_71};
  wire [511:0]     dataInMem_lo_163 = {dataInMem_hi_188, dataInMem_lo_160, dataInMem_hi_187, dataInMem_lo_159};
  wire [511:0]     dataInMem_hi_191 = {dataInMem_hi_190, dataInMem_lo_162, dataInMem_hi_189, dataInMem_lo_161};
  wire [1023:0]    dataInMem_23 = {dataInMem_hi_191, dataInMem_lo_163};
  wire [127:0]     regroupCacheLine_23_0 = dataInMem_23[127:0];
  wire [127:0]     regroupCacheLine_23_1 = dataInMem_23[255:128];
  wire [127:0]     regroupCacheLine_23_2 = dataInMem_23[383:256];
  wire [127:0]     regroupCacheLine_23_3 = dataInMem_23[511:384];
  wire [127:0]     regroupCacheLine_23_4 = dataInMem_23[639:512];
  wire [127:0]     regroupCacheLine_23_5 = dataInMem_23[767:640];
  wire [127:0]     regroupCacheLine_23_6 = dataInMem_23[895:768];
  wire [127:0]     regroupCacheLine_23_7 = dataInMem_23[1023:896];
  wire [127:0]     res_184 = regroupCacheLine_23_0;
  wire [127:0]     res_185 = regroupCacheLine_23_1;
  wire [127:0]     res_186 = regroupCacheLine_23_2;
  wire [127:0]     res_187 = regroupCacheLine_23_3;
  wire [127:0]     res_188 = regroupCacheLine_23_4;
  wire [127:0]     res_189 = regroupCacheLine_23_5;
  wire [127:0]     res_190 = regroupCacheLine_23_6;
  wire [127:0]     res_191 = regroupCacheLine_23_7;
  wire [255:0]     lo_lo_23 = {res_185, res_184};
  wire [255:0]     lo_hi_23 = {res_187, res_186};
  wire [511:0]     lo_23 = {lo_hi_23, lo_lo_23};
  wire [255:0]     hi_lo_23 = {res_189, res_188};
  wire [255:0]     hi_hi_23 = {res_191, res_190};
  wire [511:0]     hi_23 = {hi_hi_23, hi_lo_23};
  wire [1023:0]    regroupLoadData_2_7 = {hi_23, lo_23};
  wire             _GEN_143 = lsuRequest_valid | accessBufferDequeueFire;
  wire             _GEN_144 = isLastDataGroup & ~isLastMaskGroup;
  wire             _maskSelect_valid_output = _GEN_143 & _GEN_144;
  wire [7:0][15:0] _GEN_145 = {{maskForBufferData_7}, {maskForBufferData_6}, {maskForBufferData_5}, {maskForBufferData_4}, {maskForBufferData_3}, {maskForBufferData_2}, {maskForBufferData_1}, {maskForBufferData_0}};
  wire [15:0]      _GEN_146 = _GEN_145[cacheLineIndexInBuffer];
  wire             needSendTail = {7'h0, bufferBaseCacheLineIndex} == cacheLineNumberReg;
  assign memRequest_valid_0 = (bufferValid | canSendTail & needSendTail) & addressQueueFree;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo = {cacheLineTemp[8], cacheLineTemp[0]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi = {cacheLineTemp[24], cacheLineTemp[16]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo = {memRequest_bits_data_lo_lo_lo_hi, memRequest_bits_data_lo_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo = {cacheLineTemp[40], cacheLineTemp[32]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi = {cacheLineTemp[56], cacheLineTemp[48]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi = {memRequest_bits_data_lo_lo_hi_hi, memRequest_bits_data_lo_lo_hi_lo};
  wire [7:0]       memRequest_bits_data_lo_lo = {memRequest_bits_data_lo_lo_hi, memRequest_bits_data_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo = {cacheLineTemp[72], cacheLineTemp[64]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi = {cacheLineTemp[88], cacheLineTemp[80]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo = {memRequest_bits_data_lo_hi_lo_hi, memRequest_bits_data_lo_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo = {cacheLineTemp[104], cacheLineTemp[96]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi = {cacheLineTemp[120], cacheLineTemp[112]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi = {memRequest_bits_data_lo_hi_hi_hi, memRequest_bits_data_lo_hi_hi_lo};
  wire [7:0]       memRequest_bits_data_lo_hi = {memRequest_bits_data_lo_hi_hi, memRequest_bits_data_lo_hi_lo};
  wire [15:0]      memRequest_bits_data_lo = {memRequest_bits_data_lo_hi, memRequest_bits_data_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo = {dataBuffer_0[8], dataBuffer_0[0]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi = {dataBuffer_0[24], dataBuffer_0[16]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo = {memRequest_bits_data_hi_lo_lo_hi, memRequest_bits_data_hi_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo = {dataBuffer_0[40], dataBuffer_0[32]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi = {dataBuffer_0[56], dataBuffer_0[48]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi = {memRequest_bits_data_hi_lo_hi_hi, memRequest_bits_data_hi_lo_hi_lo};
  wire [7:0]       memRequest_bits_data_hi_lo = {memRequest_bits_data_hi_lo_hi, memRequest_bits_data_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo = {dataBuffer_0[72], dataBuffer_0[64]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi = {dataBuffer_0[88], dataBuffer_0[80]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo = {memRequest_bits_data_hi_hi_lo_hi, memRequest_bits_data_hi_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo = {dataBuffer_0[104], dataBuffer_0[96]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi = {dataBuffer_0[120], dataBuffer_0[112]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi = {memRequest_bits_data_hi_hi_hi_hi, memRequest_bits_data_hi_hi_hi_lo};
  wire [7:0]       memRequest_bits_data_hi_hi = {memRequest_bits_data_hi_hi_hi, memRequest_bits_data_hi_hi_lo};
  wire [15:0]      memRequest_bits_data_hi = {memRequest_bits_data_hi_hi, memRequest_bits_data_hi_lo};
  wire [46:0]      _GEN_147 = {43'h0, initOffset};
  wire [46:0]      _memRequest_bits_data_T_258 = {15'h0, memRequest_bits_data_hi, memRequest_bits_data_lo} << _GEN_147;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_1 = {cacheLineTemp[9], cacheLineTemp[1]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_1 = {cacheLineTemp[25], cacheLineTemp[17]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_1 = {memRequest_bits_data_lo_lo_lo_hi_1, memRequest_bits_data_lo_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_1 = {cacheLineTemp[41], cacheLineTemp[33]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_1 = {cacheLineTemp[57], cacheLineTemp[49]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_1 = {memRequest_bits_data_lo_lo_hi_hi_1, memRequest_bits_data_lo_lo_hi_lo_1};
  wire [7:0]       memRequest_bits_data_lo_lo_1 = {memRequest_bits_data_lo_lo_hi_1, memRequest_bits_data_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_1 = {cacheLineTemp[73], cacheLineTemp[65]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_1 = {cacheLineTemp[89], cacheLineTemp[81]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_1 = {memRequest_bits_data_lo_hi_lo_hi_1, memRequest_bits_data_lo_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_1 = {cacheLineTemp[105], cacheLineTemp[97]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_1 = {cacheLineTemp[121], cacheLineTemp[113]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_1 = {memRequest_bits_data_lo_hi_hi_hi_1, memRequest_bits_data_lo_hi_hi_lo_1};
  wire [7:0]       memRequest_bits_data_lo_hi_1 = {memRequest_bits_data_lo_hi_hi_1, memRequest_bits_data_lo_hi_lo_1};
  wire [15:0]      memRequest_bits_data_lo_1 = {memRequest_bits_data_lo_hi_1, memRequest_bits_data_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_1 = {dataBuffer_0[9], dataBuffer_0[1]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_1 = {dataBuffer_0[25], dataBuffer_0[17]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_1 = {memRequest_bits_data_hi_lo_lo_hi_1, memRequest_bits_data_hi_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_1 = {dataBuffer_0[41], dataBuffer_0[33]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_1 = {dataBuffer_0[57], dataBuffer_0[49]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_1 = {memRequest_bits_data_hi_lo_hi_hi_1, memRequest_bits_data_hi_lo_hi_lo_1};
  wire [7:0]       memRequest_bits_data_hi_lo_1 = {memRequest_bits_data_hi_lo_hi_1, memRequest_bits_data_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_1 = {dataBuffer_0[73], dataBuffer_0[65]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_1 = {dataBuffer_0[89], dataBuffer_0[81]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_1 = {memRequest_bits_data_hi_hi_lo_hi_1, memRequest_bits_data_hi_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_1 = {dataBuffer_0[105], dataBuffer_0[97]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_1 = {dataBuffer_0[121], dataBuffer_0[113]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_1 = {memRequest_bits_data_hi_hi_hi_hi_1, memRequest_bits_data_hi_hi_hi_lo_1};
  wire [7:0]       memRequest_bits_data_hi_hi_1 = {memRequest_bits_data_hi_hi_hi_1, memRequest_bits_data_hi_hi_lo_1};
  wire [15:0]      memRequest_bits_data_hi_1 = {memRequest_bits_data_hi_hi_1, memRequest_bits_data_hi_lo_1};
  wire [46:0]      _memRequest_bits_data_T_307 = {15'h0, memRequest_bits_data_hi_1, memRequest_bits_data_lo_1} << _GEN_147;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_2 = {cacheLineTemp[10], cacheLineTemp[2]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_2 = {cacheLineTemp[26], cacheLineTemp[18]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_2 = {memRequest_bits_data_lo_lo_lo_hi_2, memRequest_bits_data_lo_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_2 = {cacheLineTemp[42], cacheLineTemp[34]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_2 = {cacheLineTemp[58], cacheLineTemp[50]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_2 = {memRequest_bits_data_lo_lo_hi_hi_2, memRequest_bits_data_lo_lo_hi_lo_2};
  wire [7:0]       memRequest_bits_data_lo_lo_2 = {memRequest_bits_data_lo_lo_hi_2, memRequest_bits_data_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_2 = {cacheLineTemp[74], cacheLineTemp[66]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_2 = {cacheLineTemp[90], cacheLineTemp[82]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_2 = {memRequest_bits_data_lo_hi_lo_hi_2, memRequest_bits_data_lo_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_2 = {cacheLineTemp[106], cacheLineTemp[98]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_2 = {cacheLineTemp[122], cacheLineTemp[114]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_2 = {memRequest_bits_data_lo_hi_hi_hi_2, memRequest_bits_data_lo_hi_hi_lo_2};
  wire [7:0]       memRequest_bits_data_lo_hi_2 = {memRequest_bits_data_lo_hi_hi_2, memRequest_bits_data_lo_hi_lo_2};
  wire [15:0]      memRequest_bits_data_lo_2 = {memRequest_bits_data_lo_hi_2, memRequest_bits_data_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_2 = {dataBuffer_0[10], dataBuffer_0[2]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_2 = {dataBuffer_0[26], dataBuffer_0[18]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_2 = {memRequest_bits_data_hi_lo_lo_hi_2, memRequest_bits_data_hi_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_2 = {dataBuffer_0[42], dataBuffer_0[34]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_2 = {dataBuffer_0[58], dataBuffer_0[50]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_2 = {memRequest_bits_data_hi_lo_hi_hi_2, memRequest_bits_data_hi_lo_hi_lo_2};
  wire [7:0]       memRequest_bits_data_hi_lo_2 = {memRequest_bits_data_hi_lo_hi_2, memRequest_bits_data_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_2 = {dataBuffer_0[74], dataBuffer_0[66]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_2 = {dataBuffer_0[90], dataBuffer_0[82]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_2 = {memRequest_bits_data_hi_hi_lo_hi_2, memRequest_bits_data_hi_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_2 = {dataBuffer_0[106], dataBuffer_0[98]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_2 = {dataBuffer_0[122], dataBuffer_0[114]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_2 = {memRequest_bits_data_hi_hi_hi_hi_2, memRequest_bits_data_hi_hi_hi_lo_2};
  wire [7:0]       memRequest_bits_data_hi_hi_2 = {memRequest_bits_data_hi_hi_hi_2, memRequest_bits_data_hi_hi_lo_2};
  wire [15:0]      memRequest_bits_data_hi_2 = {memRequest_bits_data_hi_hi_2, memRequest_bits_data_hi_lo_2};
  wire [46:0]      _memRequest_bits_data_T_356 = {15'h0, memRequest_bits_data_hi_2, memRequest_bits_data_lo_2} << _GEN_147;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_3 = {cacheLineTemp[11], cacheLineTemp[3]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_3 = {cacheLineTemp[27], cacheLineTemp[19]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_3 = {memRequest_bits_data_lo_lo_lo_hi_3, memRequest_bits_data_lo_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_3 = {cacheLineTemp[43], cacheLineTemp[35]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_3 = {cacheLineTemp[59], cacheLineTemp[51]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_3 = {memRequest_bits_data_lo_lo_hi_hi_3, memRequest_bits_data_lo_lo_hi_lo_3};
  wire [7:0]       memRequest_bits_data_lo_lo_3 = {memRequest_bits_data_lo_lo_hi_3, memRequest_bits_data_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_3 = {cacheLineTemp[75], cacheLineTemp[67]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_3 = {cacheLineTemp[91], cacheLineTemp[83]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_3 = {memRequest_bits_data_lo_hi_lo_hi_3, memRequest_bits_data_lo_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_3 = {cacheLineTemp[107], cacheLineTemp[99]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_3 = {cacheLineTemp[123], cacheLineTemp[115]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_3 = {memRequest_bits_data_lo_hi_hi_hi_3, memRequest_bits_data_lo_hi_hi_lo_3};
  wire [7:0]       memRequest_bits_data_lo_hi_3 = {memRequest_bits_data_lo_hi_hi_3, memRequest_bits_data_lo_hi_lo_3};
  wire [15:0]      memRequest_bits_data_lo_3 = {memRequest_bits_data_lo_hi_3, memRequest_bits_data_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_3 = {dataBuffer_0[11], dataBuffer_0[3]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_3 = {dataBuffer_0[27], dataBuffer_0[19]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_3 = {memRequest_bits_data_hi_lo_lo_hi_3, memRequest_bits_data_hi_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_3 = {dataBuffer_0[43], dataBuffer_0[35]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_3 = {dataBuffer_0[59], dataBuffer_0[51]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_3 = {memRequest_bits_data_hi_lo_hi_hi_3, memRequest_bits_data_hi_lo_hi_lo_3};
  wire [7:0]       memRequest_bits_data_hi_lo_3 = {memRequest_bits_data_hi_lo_hi_3, memRequest_bits_data_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_3 = {dataBuffer_0[75], dataBuffer_0[67]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_3 = {dataBuffer_0[91], dataBuffer_0[83]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_3 = {memRequest_bits_data_hi_hi_lo_hi_3, memRequest_bits_data_hi_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_3 = {dataBuffer_0[107], dataBuffer_0[99]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_3 = {dataBuffer_0[123], dataBuffer_0[115]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_3 = {memRequest_bits_data_hi_hi_hi_hi_3, memRequest_bits_data_hi_hi_hi_lo_3};
  wire [7:0]       memRequest_bits_data_hi_hi_3 = {memRequest_bits_data_hi_hi_hi_3, memRequest_bits_data_hi_hi_lo_3};
  wire [15:0]      memRequest_bits_data_hi_3 = {memRequest_bits_data_hi_hi_3, memRequest_bits_data_hi_lo_3};
  wire [46:0]      _memRequest_bits_data_T_405 = {15'h0, memRequest_bits_data_hi_3, memRequest_bits_data_lo_3} << _GEN_147;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_4 = {cacheLineTemp[12], cacheLineTemp[4]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_4 = {cacheLineTemp[28], cacheLineTemp[20]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_4 = {memRequest_bits_data_lo_lo_lo_hi_4, memRequest_bits_data_lo_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_4 = {cacheLineTemp[44], cacheLineTemp[36]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_4 = {cacheLineTemp[60], cacheLineTemp[52]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_4 = {memRequest_bits_data_lo_lo_hi_hi_4, memRequest_bits_data_lo_lo_hi_lo_4};
  wire [7:0]       memRequest_bits_data_lo_lo_4 = {memRequest_bits_data_lo_lo_hi_4, memRequest_bits_data_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_4 = {cacheLineTemp[76], cacheLineTemp[68]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_4 = {cacheLineTemp[92], cacheLineTemp[84]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_4 = {memRequest_bits_data_lo_hi_lo_hi_4, memRequest_bits_data_lo_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_4 = {cacheLineTemp[108], cacheLineTemp[100]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_4 = {cacheLineTemp[124], cacheLineTemp[116]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_4 = {memRequest_bits_data_lo_hi_hi_hi_4, memRequest_bits_data_lo_hi_hi_lo_4};
  wire [7:0]       memRequest_bits_data_lo_hi_4 = {memRequest_bits_data_lo_hi_hi_4, memRequest_bits_data_lo_hi_lo_4};
  wire [15:0]      memRequest_bits_data_lo_4 = {memRequest_bits_data_lo_hi_4, memRequest_bits_data_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_4 = {dataBuffer_0[12], dataBuffer_0[4]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_4 = {dataBuffer_0[28], dataBuffer_0[20]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_4 = {memRequest_bits_data_hi_lo_lo_hi_4, memRequest_bits_data_hi_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_4 = {dataBuffer_0[44], dataBuffer_0[36]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_4 = {dataBuffer_0[60], dataBuffer_0[52]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_4 = {memRequest_bits_data_hi_lo_hi_hi_4, memRequest_bits_data_hi_lo_hi_lo_4};
  wire [7:0]       memRequest_bits_data_hi_lo_4 = {memRequest_bits_data_hi_lo_hi_4, memRequest_bits_data_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_4 = {dataBuffer_0[76], dataBuffer_0[68]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_4 = {dataBuffer_0[92], dataBuffer_0[84]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_4 = {memRequest_bits_data_hi_hi_lo_hi_4, memRequest_bits_data_hi_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_4 = {dataBuffer_0[108], dataBuffer_0[100]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_4 = {dataBuffer_0[124], dataBuffer_0[116]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_4 = {memRequest_bits_data_hi_hi_hi_hi_4, memRequest_bits_data_hi_hi_hi_lo_4};
  wire [7:0]       memRequest_bits_data_hi_hi_4 = {memRequest_bits_data_hi_hi_hi_4, memRequest_bits_data_hi_hi_lo_4};
  wire [15:0]      memRequest_bits_data_hi_4 = {memRequest_bits_data_hi_hi_4, memRequest_bits_data_hi_lo_4};
  wire [46:0]      _memRequest_bits_data_T_454 = {15'h0, memRequest_bits_data_hi_4, memRequest_bits_data_lo_4} << _GEN_147;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_5 = {cacheLineTemp[13], cacheLineTemp[5]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_5 = {cacheLineTemp[29], cacheLineTemp[21]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_5 = {memRequest_bits_data_lo_lo_lo_hi_5, memRequest_bits_data_lo_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_5 = {cacheLineTemp[45], cacheLineTemp[37]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_5 = {cacheLineTemp[61], cacheLineTemp[53]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_5 = {memRequest_bits_data_lo_lo_hi_hi_5, memRequest_bits_data_lo_lo_hi_lo_5};
  wire [7:0]       memRequest_bits_data_lo_lo_5 = {memRequest_bits_data_lo_lo_hi_5, memRequest_bits_data_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_5 = {cacheLineTemp[77], cacheLineTemp[69]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_5 = {cacheLineTemp[93], cacheLineTemp[85]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_5 = {memRequest_bits_data_lo_hi_lo_hi_5, memRequest_bits_data_lo_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_5 = {cacheLineTemp[109], cacheLineTemp[101]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_5 = {cacheLineTemp[125], cacheLineTemp[117]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_5 = {memRequest_bits_data_lo_hi_hi_hi_5, memRequest_bits_data_lo_hi_hi_lo_5};
  wire [7:0]       memRequest_bits_data_lo_hi_5 = {memRequest_bits_data_lo_hi_hi_5, memRequest_bits_data_lo_hi_lo_5};
  wire [15:0]      memRequest_bits_data_lo_5 = {memRequest_bits_data_lo_hi_5, memRequest_bits_data_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_5 = {dataBuffer_0[13], dataBuffer_0[5]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_5 = {dataBuffer_0[29], dataBuffer_0[21]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_5 = {memRequest_bits_data_hi_lo_lo_hi_5, memRequest_bits_data_hi_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_5 = {dataBuffer_0[45], dataBuffer_0[37]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_5 = {dataBuffer_0[61], dataBuffer_0[53]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_5 = {memRequest_bits_data_hi_lo_hi_hi_5, memRequest_bits_data_hi_lo_hi_lo_5};
  wire [7:0]       memRequest_bits_data_hi_lo_5 = {memRequest_bits_data_hi_lo_hi_5, memRequest_bits_data_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_5 = {dataBuffer_0[77], dataBuffer_0[69]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_5 = {dataBuffer_0[93], dataBuffer_0[85]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_5 = {memRequest_bits_data_hi_hi_lo_hi_5, memRequest_bits_data_hi_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_5 = {dataBuffer_0[109], dataBuffer_0[101]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_5 = {dataBuffer_0[125], dataBuffer_0[117]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_5 = {memRequest_bits_data_hi_hi_hi_hi_5, memRequest_bits_data_hi_hi_hi_lo_5};
  wire [7:0]       memRequest_bits_data_hi_hi_5 = {memRequest_bits_data_hi_hi_hi_5, memRequest_bits_data_hi_hi_lo_5};
  wire [15:0]      memRequest_bits_data_hi_5 = {memRequest_bits_data_hi_hi_5, memRequest_bits_data_hi_lo_5};
  wire [46:0]      _memRequest_bits_data_T_503 = {15'h0, memRequest_bits_data_hi_5, memRequest_bits_data_lo_5} << _GEN_147;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_6 = {cacheLineTemp[14], cacheLineTemp[6]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_6 = {cacheLineTemp[30], cacheLineTemp[22]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_6 = {memRequest_bits_data_lo_lo_lo_hi_6, memRequest_bits_data_lo_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_6 = {cacheLineTemp[46], cacheLineTemp[38]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_6 = {cacheLineTemp[62], cacheLineTemp[54]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_6 = {memRequest_bits_data_lo_lo_hi_hi_6, memRequest_bits_data_lo_lo_hi_lo_6};
  wire [7:0]       memRequest_bits_data_lo_lo_6 = {memRequest_bits_data_lo_lo_hi_6, memRequest_bits_data_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_6 = {cacheLineTemp[78], cacheLineTemp[70]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_6 = {cacheLineTemp[94], cacheLineTemp[86]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_6 = {memRequest_bits_data_lo_hi_lo_hi_6, memRequest_bits_data_lo_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_6 = {cacheLineTemp[110], cacheLineTemp[102]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_6 = {cacheLineTemp[126], cacheLineTemp[118]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_6 = {memRequest_bits_data_lo_hi_hi_hi_6, memRequest_bits_data_lo_hi_hi_lo_6};
  wire [7:0]       memRequest_bits_data_lo_hi_6 = {memRequest_bits_data_lo_hi_hi_6, memRequest_bits_data_lo_hi_lo_6};
  wire [15:0]      memRequest_bits_data_lo_6 = {memRequest_bits_data_lo_hi_6, memRequest_bits_data_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_6 = {dataBuffer_0[14], dataBuffer_0[6]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_6 = {dataBuffer_0[30], dataBuffer_0[22]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_6 = {memRequest_bits_data_hi_lo_lo_hi_6, memRequest_bits_data_hi_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_6 = {dataBuffer_0[46], dataBuffer_0[38]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_6 = {dataBuffer_0[62], dataBuffer_0[54]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_6 = {memRequest_bits_data_hi_lo_hi_hi_6, memRequest_bits_data_hi_lo_hi_lo_6};
  wire [7:0]       memRequest_bits_data_hi_lo_6 = {memRequest_bits_data_hi_lo_hi_6, memRequest_bits_data_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_6 = {dataBuffer_0[78], dataBuffer_0[70]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_6 = {dataBuffer_0[94], dataBuffer_0[86]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_6 = {memRequest_bits_data_hi_hi_lo_hi_6, memRequest_bits_data_hi_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_6 = {dataBuffer_0[110], dataBuffer_0[102]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_6 = {dataBuffer_0[126], dataBuffer_0[118]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_6 = {memRequest_bits_data_hi_hi_hi_hi_6, memRequest_bits_data_hi_hi_hi_lo_6};
  wire [7:0]       memRequest_bits_data_hi_hi_6 = {memRequest_bits_data_hi_hi_hi_6, memRequest_bits_data_hi_hi_lo_6};
  wire [15:0]      memRequest_bits_data_hi_6 = {memRequest_bits_data_hi_hi_6, memRequest_bits_data_hi_lo_6};
  wire [46:0]      _memRequest_bits_data_T_552 = {15'h0, memRequest_bits_data_hi_6, memRequest_bits_data_lo_6} << _GEN_147;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_7 = {cacheLineTemp[15], cacheLineTemp[7]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_7 = {cacheLineTemp[31], cacheLineTemp[23]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_7 = {memRequest_bits_data_lo_lo_lo_hi_7, memRequest_bits_data_lo_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_7 = {cacheLineTemp[47], cacheLineTemp[39]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_7 = {cacheLineTemp[63], cacheLineTemp[55]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_7 = {memRequest_bits_data_lo_lo_hi_hi_7, memRequest_bits_data_lo_lo_hi_lo_7};
  wire [7:0]       memRequest_bits_data_lo_lo_7 = {memRequest_bits_data_lo_lo_hi_7, memRequest_bits_data_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_7 = {cacheLineTemp[79], cacheLineTemp[71]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_7 = {cacheLineTemp[95], cacheLineTemp[87]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_7 = {memRequest_bits_data_lo_hi_lo_hi_7, memRequest_bits_data_lo_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_7 = {cacheLineTemp[111], cacheLineTemp[103]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_7 = {cacheLineTemp[127], cacheLineTemp[119]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_7 = {memRequest_bits_data_lo_hi_hi_hi_7, memRequest_bits_data_lo_hi_hi_lo_7};
  wire [7:0]       memRequest_bits_data_lo_hi_7 = {memRequest_bits_data_lo_hi_hi_7, memRequest_bits_data_lo_hi_lo_7};
  wire [15:0]      memRequest_bits_data_lo_7 = {memRequest_bits_data_lo_hi_7, memRequest_bits_data_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_7 = {dataBuffer_0[15], dataBuffer_0[7]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_7 = {dataBuffer_0[31], dataBuffer_0[23]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_7 = {memRequest_bits_data_hi_lo_lo_hi_7, memRequest_bits_data_hi_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_7 = {dataBuffer_0[47], dataBuffer_0[39]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_7 = {dataBuffer_0[63], dataBuffer_0[55]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_7 = {memRequest_bits_data_hi_lo_hi_hi_7, memRequest_bits_data_hi_lo_hi_lo_7};
  wire [7:0]       memRequest_bits_data_hi_lo_7 = {memRequest_bits_data_hi_lo_hi_7, memRequest_bits_data_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_7 = {dataBuffer_0[79], dataBuffer_0[71]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_7 = {dataBuffer_0[95], dataBuffer_0[87]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_7 = {memRequest_bits_data_hi_hi_lo_hi_7, memRequest_bits_data_hi_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_7 = {dataBuffer_0[111], dataBuffer_0[103]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_7 = {dataBuffer_0[127], dataBuffer_0[119]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_7 = {memRequest_bits_data_hi_hi_hi_hi_7, memRequest_bits_data_hi_hi_hi_lo_7};
  wire [7:0]       memRequest_bits_data_hi_hi_7 = {memRequest_bits_data_hi_hi_hi_7, memRequest_bits_data_hi_hi_lo_7};
  wire [15:0]      memRequest_bits_data_hi_7 = {memRequest_bits_data_hi_hi_7, memRequest_bits_data_hi_lo_7};
  wire [46:0]      _memRequest_bits_data_T_601 = {15'h0, memRequest_bits_data_hi_7, memRequest_bits_data_lo_7} << _GEN_147;
  wire [1:0]       memRequest_bits_data_lo_lo_8 = {_memRequest_bits_data_T_307[0], _memRequest_bits_data_T_258[0]};
  wire [1:0]       memRequest_bits_data_lo_hi_8 = {_memRequest_bits_data_T_405[0], _memRequest_bits_data_T_356[0]};
  wire [3:0]       memRequest_bits_data_lo_8 = {memRequest_bits_data_lo_hi_8, memRequest_bits_data_lo_lo_8};
  wire [1:0]       memRequest_bits_data_hi_lo_8 = {_memRequest_bits_data_T_503[0], _memRequest_bits_data_T_454[0]};
  wire [1:0]       memRequest_bits_data_hi_hi_8 = {_memRequest_bits_data_T_601[0], _memRequest_bits_data_T_552[0]};
  wire [3:0]       memRequest_bits_data_hi_8 = {memRequest_bits_data_hi_hi_8, memRequest_bits_data_hi_lo_8};
  wire [1:0]       memRequest_bits_data_lo_lo_9 = {_memRequest_bits_data_T_307[1], _memRequest_bits_data_T_258[1]};
  wire [1:0]       memRequest_bits_data_lo_hi_9 = {_memRequest_bits_data_T_405[1], _memRequest_bits_data_T_356[1]};
  wire [3:0]       memRequest_bits_data_lo_9 = {memRequest_bits_data_lo_hi_9, memRequest_bits_data_lo_lo_9};
  wire [1:0]       memRequest_bits_data_hi_lo_9 = {_memRequest_bits_data_T_503[1], _memRequest_bits_data_T_454[1]};
  wire [1:0]       memRequest_bits_data_hi_hi_9 = {_memRequest_bits_data_T_601[1], _memRequest_bits_data_T_552[1]};
  wire [3:0]       memRequest_bits_data_hi_9 = {memRequest_bits_data_hi_hi_9, memRequest_bits_data_hi_lo_9};
  wire [1:0]       memRequest_bits_data_lo_lo_10 = {_memRequest_bits_data_T_307[2], _memRequest_bits_data_T_258[2]};
  wire [1:0]       memRequest_bits_data_lo_hi_10 = {_memRequest_bits_data_T_405[2], _memRequest_bits_data_T_356[2]};
  wire [3:0]       memRequest_bits_data_lo_10 = {memRequest_bits_data_lo_hi_10, memRequest_bits_data_lo_lo_10};
  wire [1:0]       memRequest_bits_data_hi_lo_10 = {_memRequest_bits_data_T_503[2], _memRequest_bits_data_T_454[2]};
  wire [1:0]       memRequest_bits_data_hi_hi_10 = {_memRequest_bits_data_T_601[2], _memRequest_bits_data_T_552[2]};
  wire [3:0]       memRequest_bits_data_hi_10 = {memRequest_bits_data_hi_hi_10, memRequest_bits_data_hi_lo_10};
  wire [1:0]       memRequest_bits_data_lo_lo_11 = {_memRequest_bits_data_T_307[3], _memRequest_bits_data_T_258[3]};
  wire [1:0]       memRequest_bits_data_lo_hi_11 = {_memRequest_bits_data_T_405[3], _memRequest_bits_data_T_356[3]};
  wire [3:0]       memRequest_bits_data_lo_11 = {memRequest_bits_data_lo_hi_11, memRequest_bits_data_lo_lo_11};
  wire [1:0]       memRequest_bits_data_hi_lo_11 = {_memRequest_bits_data_T_503[3], _memRequest_bits_data_T_454[3]};
  wire [1:0]       memRequest_bits_data_hi_hi_11 = {_memRequest_bits_data_T_601[3], _memRequest_bits_data_T_552[3]};
  wire [3:0]       memRequest_bits_data_hi_11 = {memRequest_bits_data_hi_hi_11, memRequest_bits_data_hi_lo_11};
  wire [1:0]       memRequest_bits_data_lo_lo_12 = {_memRequest_bits_data_T_307[4], _memRequest_bits_data_T_258[4]};
  wire [1:0]       memRequest_bits_data_lo_hi_12 = {_memRequest_bits_data_T_405[4], _memRequest_bits_data_T_356[4]};
  wire [3:0]       memRequest_bits_data_lo_12 = {memRequest_bits_data_lo_hi_12, memRequest_bits_data_lo_lo_12};
  wire [1:0]       memRequest_bits_data_hi_lo_12 = {_memRequest_bits_data_T_503[4], _memRequest_bits_data_T_454[4]};
  wire [1:0]       memRequest_bits_data_hi_hi_12 = {_memRequest_bits_data_T_601[4], _memRequest_bits_data_T_552[4]};
  wire [3:0]       memRequest_bits_data_hi_12 = {memRequest_bits_data_hi_hi_12, memRequest_bits_data_hi_lo_12};
  wire [1:0]       memRequest_bits_data_lo_lo_13 = {_memRequest_bits_data_T_307[5], _memRequest_bits_data_T_258[5]};
  wire [1:0]       memRequest_bits_data_lo_hi_13 = {_memRequest_bits_data_T_405[5], _memRequest_bits_data_T_356[5]};
  wire [3:0]       memRequest_bits_data_lo_13 = {memRequest_bits_data_lo_hi_13, memRequest_bits_data_lo_lo_13};
  wire [1:0]       memRequest_bits_data_hi_lo_13 = {_memRequest_bits_data_T_503[5], _memRequest_bits_data_T_454[5]};
  wire [1:0]       memRequest_bits_data_hi_hi_13 = {_memRequest_bits_data_T_601[5], _memRequest_bits_data_T_552[5]};
  wire [3:0]       memRequest_bits_data_hi_13 = {memRequest_bits_data_hi_hi_13, memRequest_bits_data_hi_lo_13};
  wire [1:0]       memRequest_bits_data_lo_lo_14 = {_memRequest_bits_data_T_307[6], _memRequest_bits_data_T_258[6]};
  wire [1:0]       memRequest_bits_data_lo_hi_14 = {_memRequest_bits_data_T_405[6], _memRequest_bits_data_T_356[6]};
  wire [3:0]       memRequest_bits_data_lo_14 = {memRequest_bits_data_lo_hi_14, memRequest_bits_data_lo_lo_14};
  wire [1:0]       memRequest_bits_data_hi_lo_14 = {_memRequest_bits_data_T_503[6], _memRequest_bits_data_T_454[6]};
  wire [1:0]       memRequest_bits_data_hi_hi_14 = {_memRequest_bits_data_T_601[6], _memRequest_bits_data_T_552[6]};
  wire [3:0]       memRequest_bits_data_hi_14 = {memRequest_bits_data_hi_hi_14, memRequest_bits_data_hi_lo_14};
  wire [1:0]       memRequest_bits_data_lo_lo_15 = {_memRequest_bits_data_T_307[7], _memRequest_bits_data_T_258[7]};
  wire [1:0]       memRequest_bits_data_lo_hi_15 = {_memRequest_bits_data_T_405[7], _memRequest_bits_data_T_356[7]};
  wire [3:0]       memRequest_bits_data_lo_15 = {memRequest_bits_data_lo_hi_15, memRequest_bits_data_lo_lo_15};
  wire [1:0]       memRequest_bits_data_hi_lo_15 = {_memRequest_bits_data_T_503[7], _memRequest_bits_data_T_454[7]};
  wire [1:0]       memRequest_bits_data_hi_hi_15 = {_memRequest_bits_data_T_601[7], _memRequest_bits_data_T_552[7]};
  wire [3:0]       memRequest_bits_data_hi_15 = {memRequest_bits_data_hi_hi_15, memRequest_bits_data_hi_lo_15};
  wire [1:0]       memRequest_bits_data_lo_lo_16 = {_memRequest_bits_data_T_307[8], _memRequest_bits_data_T_258[8]};
  wire [1:0]       memRequest_bits_data_lo_hi_16 = {_memRequest_bits_data_T_405[8], _memRequest_bits_data_T_356[8]};
  wire [3:0]       memRequest_bits_data_lo_16 = {memRequest_bits_data_lo_hi_16, memRequest_bits_data_lo_lo_16};
  wire [1:0]       memRequest_bits_data_hi_lo_16 = {_memRequest_bits_data_T_503[8], _memRequest_bits_data_T_454[8]};
  wire [1:0]       memRequest_bits_data_hi_hi_16 = {_memRequest_bits_data_T_601[8], _memRequest_bits_data_T_552[8]};
  wire [3:0]       memRequest_bits_data_hi_16 = {memRequest_bits_data_hi_hi_16, memRequest_bits_data_hi_lo_16};
  wire [1:0]       memRequest_bits_data_lo_lo_17 = {_memRequest_bits_data_T_307[9], _memRequest_bits_data_T_258[9]};
  wire [1:0]       memRequest_bits_data_lo_hi_17 = {_memRequest_bits_data_T_405[9], _memRequest_bits_data_T_356[9]};
  wire [3:0]       memRequest_bits_data_lo_17 = {memRequest_bits_data_lo_hi_17, memRequest_bits_data_lo_lo_17};
  wire [1:0]       memRequest_bits_data_hi_lo_17 = {_memRequest_bits_data_T_503[9], _memRequest_bits_data_T_454[9]};
  wire [1:0]       memRequest_bits_data_hi_hi_17 = {_memRequest_bits_data_T_601[9], _memRequest_bits_data_T_552[9]};
  wire [3:0]       memRequest_bits_data_hi_17 = {memRequest_bits_data_hi_hi_17, memRequest_bits_data_hi_lo_17};
  wire [1:0]       memRequest_bits_data_lo_lo_18 = {_memRequest_bits_data_T_307[10], _memRequest_bits_data_T_258[10]};
  wire [1:0]       memRequest_bits_data_lo_hi_18 = {_memRequest_bits_data_T_405[10], _memRequest_bits_data_T_356[10]};
  wire [3:0]       memRequest_bits_data_lo_18 = {memRequest_bits_data_lo_hi_18, memRequest_bits_data_lo_lo_18};
  wire [1:0]       memRequest_bits_data_hi_lo_18 = {_memRequest_bits_data_T_503[10], _memRequest_bits_data_T_454[10]};
  wire [1:0]       memRequest_bits_data_hi_hi_18 = {_memRequest_bits_data_T_601[10], _memRequest_bits_data_T_552[10]};
  wire [3:0]       memRequest_bits_data_hi_18 = {memRequest_bits_data_hi_hi_18, memRequest_bits_data_hi_lo_18};
  wire [1:0]       memRequest_bits_data_lo_lo_19 = {_memRequest_bits_data_T_307[11], _memRequest_bits_data_T_258[11]};
  wire [1:0]       memRequest_bits_data_lo_hi_19 = {_memRequest_bits_data_T_405[11], _memRequest_bits_data_T_356[11]};
  wire [3:0]       memRequest_bits_data_lo_19 = {memRequest_bits_data_lo_hi_19, memRequest_bits_data_lo_lo_19};
  wire [1:0]       memRequest_bits_data_hi_lo_19 = {_memRequest_bits_data_T_503[11], _memRequest_bits_data_T_454[11]};
  wire [1:0]       memRequest_bits_data_hi_hi_19 = {_memRequest_bits_data_T_601[11], _memRequest_bits_data_T_552[11]};
  wire [3:0]       memRequest_bits_data_hi_19 = {memRequest_bits_data_hi_hi_19, memRequest_bits_data_hi_lo_19};
  wire [1:0]       memRequest_bits_data_lo_lo_20 = {_memRequest_bits_data_T_307[12], _memRequest_bits_data_T_258[12]};
  wire [1:0]       memRequest_bits_data_lo_hi_20 = {_memRequest_bits_data_T_405[12], _memRequest_bits_data_T_356[12]};
  wire [3:0]       memRequest_bits_data_lo_20 = {memRequest_bits_data_lo_hi_20, memRequest_bits_data_lo_lo_20};
  wire [1:0]       memRequest_bits_data_hi_lo_20 = {_memRequest_bits_data_T_503[12], _memRequest_bits_data_T_454[12]};
  wire [1:0]       memRequest_bits_data_hi_hi_20 = {_memRequest_bits_data_T_601[12], _memRequest_bits_data_T_552[12]};
  wire [3:0]       memRequest_bits_data_hi_20 = {memRequest_bits_data_hi_hi_20, memRequest_bits_data_hi_lo_20};
  wire [1:0]       memRequest_bits_data_lo_lo_21 = {_memRequest_bits_data_T_307[13], _memRequest_bits_data_T_258[13]};
  wire [1:0]       memRequest_bits_data_lo_hi_21 = {_memRequest_bits_data_T_405[13], _memRequest_bits_data_T_356[13]};
  wire [3:0]       memRequest_bits_data_lo_21 = {memRequest_bits_data_lo_hi_21, memRequest_bits_data_lo_lo_21};
  wire [1:0]       memRequest_bits_data_hi_lo_21 = {_memRequest_bits_data_T_503[13], _memRequest_bits_data_T_454[13]};
  wire [1:0]       memRequest_bits_data_hi_hi_21 = {_memRequest_bits_data_T_601[13], _memRequest_bits_data_T_552[13]};
  wire [3:0]       memRequest_bits_data_hi_21 = {memRequest_bits_data_hi_hi_21, memRequest_bits_data_hi_lo_21};
  wire [1:0]       memRequest_bits_data_lo_lo_22 = {_memRequest_bits_data_T_307[14], _memRequest_bits_data_T_258[14]};
  wire [1:0]       memRequest_bits_data_lo_hi_22 = {_memRequest_bits_data_T_405[14], _memRequest_bits_data_T_356[14]};
  wire [3:0]       memRequest_bits_data_lo_22 = {memRequest_bits_data_lo_hi_22, memRequest_bits_data_lo_lo_22};
  wire [1:0]       memRequest_bits_data_hi_lo_22 = {_memRequest_bits_data_T_503[14], _memRequest_bits_data_T_454[14]};
  wire [1:0]       memRequest_bits_data_hi_hi_22 = {_memRequest_bits_data_T_601[14], _memRequest_bits_data_T_552[14]};
  wire [3:0]       memRequest_bits_data_hi_22 = {memRequest_bits_data_hi_hi_22, memRequest_bits_data_hi_lo_22};
  wire [1:0]       memRequest_bits_data_lo_lo_23 = {_memRequest_bits_data_T_307[15], _memRequest_bits_data_T_258[15]};
  wire [1:0]       memRequest_bits_data_lo_hi_23 = {_memRequest_bits_data_T_405[15], _memRequest_bits_data_T_356[15]};
  wire [3:0]       memRequest_bits_data_lo_23 = {memRequest_bits_data_lo_hi_23, memRequest_bits_data_lo_lo_23};
  wire [1:0]       memRequest_bits_data_hi_lo_23 = {_memRequest_bits_data_T_503[15], _memRequest_bits_data_T_454[15]};
  wire [1:0]       memRequest_bits_data_hi_hi_23 = {_memRequest_bits_data_T_601[15], _memRequest_bits_data_T_552[15]};
  wire [3:0]       memRequest_bits_data_hi_23 = {memRequest_bits_data_hi_hi_23, memRequest_bits_data_hi_lo_23};
  wire [1:0]       memRequest_bits_data_lo_lo_24 = {_memRequest_bits_data_T_307[16], _memRequest_bits_data_T_258[16]};
  wire [1:0]       memRequest_bits_data_lo_hi_24 = {_memRequest_bits_data_T_405[16], _memRequest_bits_data_T_356[16]};
  wire [3:0]       memRequest_bits_data_lo_24 = {memRequest_bits_data_lo_hi_24, memRequest_bits_data_lo_lo_24};
  wire [1:0]       memRequest_bits_data_hi_lo_24 = {_memRequest_bits_data_T_503[16], _memRequest_bits_data_T_454[16]};
  wire [1:0]       memRequest_bits_data_hi_hi_24 = {_memRequest_bits_data_T_601[16], _memRequest_bits_data_T_552[16]};
  wire [3:0]       memRequest_bits_data_hi_24 = {memRequest_bits_data_hi_hi_24, memRequest_bits_data_hi_lo_24};
  wire [1:0]       memRequest_bits_data_lo_lo_25 = {_memRequest_bits_data_T_307[17], _memRequest_bits_data_T_258[17]};
  wire [1:0]       memRequest_bits_data_lo_hi_25 = {_memRequest_bits_data_T_405[17], _memRequest_bits_data_T_356[17]};
  wire [3:0]       memRequest_bits_data_lo_25 = {memRequest_bits_data_lo_hi_25, memRequest_bits_data_lo_lo_25};
  wire [1:0]       memRequest_bits_data_hi_lo_25 = {_memRequest_bits_data_T_503[17], _memRequest_bits_data_T_454[17]};
  wire [1:0]       memRequest_bits_data_hi_hi_25 = {_memRequest_bits_data_T_601[17], _memRequest_bits_data_T_552[17]};
  wire [3:0]       memRequest_bits_data_hi_25 = {memRequest_bits_data_hi_hi_25, memRequest_bits_data_hi_lo_25};
  wire [1:0]       memRequest_bits_data_lo_lo_26 = {_memRequest_bits_data_T_307[18], _memRequest_bits_data_T_258[18]};
  wire [1:0]       memRequest_bits_data_lo_hi_26 = {_memRequest_bits_data_T_405[18], _memRequest_bits_data_T_356[18]};
  wire [3:0]       memRequest_bits_data_lo_26 = {memRequest_bits_data_lo_hi_26, memRequest_bits_data_lo_lo_26};
  wire [1:0]       memRequest_bits_data_hi_lo_26 = {_memRequest_bits_data_T_503[18], _memRequest_bits_data_T_454[18]};
  wire [1:0]       memRequest_bits_data_hi_hi_26 = {_memRequest_bits_data_T_601[18], _memRequest_bits_data_T_552[18]};
  wire [3:0]       memRequest_bits_data_hi_26 = {memRequest_bits_data_hi_hi_26, memRequest_bits_data_hi_lo_26};
  wire [1:0]       memRequest_bits_data_lo_lo_27 = {_memRequest_bits_data_T_307[19], _memRequest_bits_data_T_258[19]};
  wire [1:0]       memRequest_bits_data_lo_hi_27 = {_memRequest_bits_data_T_405[19], _memRequest_bits_data_T_356[19]};
  wire [3:0]       memRequest_bits_data_lo_27 = {memRequest_bits_data_lo_hi_27, memRequest_bits_data_lo_lo_27};
  wire [1:0]       memRequest_bits_data_hi_lo_27 = {_memRequest_bits_data_T_503[19], _memRequest_bits_data_T_454[19]};
  wire [1:0]       memRequest_bits_data_hi_hi_27 = {_memRequest_bits_data_T_601[19], _memRequest_bits_data_T_552[19]};
  wire [3:0]       memRequest_bits_data_hi_27 = {memRequest_bits_data_hi_hi_27, memRequest_bits_data_hi_lo_27};
  wire [1:0]       memRequest_bits_data_lo_lo_28 = {_memRequest_bits_data_T_307[20], _memRequest_bits_data_T_258[20]};
  wire [1:0]       memRequest_bits_data_lo_hi_28 = {_memRequest_bits_data_T_405[20], _memRequest_bits_data_T_356[20]};
  wire [3:0]       memRequest_bits_data_lo_28 = {memRequest_bits_data_lo_hi_28, memRequest_bits_data_lo_lo_28};
  wire [1:0]       memRequest_bits_data_hi_lo_28 = {_memRequest_bits_data_T_503[20], _memRequest_bits_data_T_454[20]};
  wire [1:0]       memRequest_bits_data_hi_hi_28 = {_memRequest_bits_data_T_601[20], _memRequest_bits_data_T_552[20]};
  wire [3:0]       memRequest_bits_data_hi_28 = {memRequest_bits_data_hi_hi_28, memRequest_bits_data_hi_lo_28};
  wire [1:0]       memRequest_bits_data_lo_lo_29 = {_memRequest_bits_data_T_307[21], _memRequest_bits_data_T_258[21]};
  wire [1:0]       memRequest_bits_data_lo_hi_29 = {_memRequest_bits_data_T_405[21], _memRequest_bits_data_T_356[21]};
  wire [3:0]       memRequest_bits_data_lo_29 = {memRequest_bits_data_lo_hi_29, memRequest_bits_data_lo_lo_29};
  wire [1:0]       memRequest_bits_data_hi_lo_29 = {_memRequest_bits_data_T_503[21], _memRequest_bits_data_T_454[21]};
  wire [1:0]       memRequest_bits_data_hi_hi_29 = {_memRequest_bits_data_T_601[21], _memRequest_bits_data_T_552[21]};
  wire [3:0]       memRequest_bits_data_hi_29 = {memRequest_bits_data_hi_hi_29, memRequest_bits_data_hi_lo_29};
  wire [1:0]       memRequest_bits_data_lo_lo_30 = {_memRequest_bits_data_T_307[22], _memRequest_bits_data_T_258[22]};
  wire [1:0]       memRequest_bits_data_lo_hi_30 = {_memRequest_bits_data_T_405[22], _memRequest_bits_data_T_356[22]};
  wire [3:0]       memRequest_bits_data_lo_30 = {memRequest_bits_data_lo_hi_30, memRequest_bits_data_lo_lo_30};
  wire [1:0]       memRequest_bits_data_hi_lo_30 = {_memRequest_bits_data_T_503[22], _memRequest_bits_data_T_454[22]};
  wire [1:0]       memRequest_bits_data_hi_hi_30 = {_memRequest_bits_data_T_601[22], _memRequest_bits_data_T_552[22]};
  wire [3:0]       memRequest_bits_data_hi_30 = {memRequest_bits_data_hi_hi_30, memRequest_bits_data_hi_lo_30};
  wire [1:0]       memRequest_bits_data_lo_lo_31 = {_memRequest_bits_data_T_307[23], _memRequest_bits_data_T_258[23]};
  wire [1:0]       memRequest_bits_data_lo_hi_31 = {_memRequest_bits_data_T_405[23], _memRequest_bits_data_T_356[23]};
  wire [3:0]       memRequest_bits_data_lo_31 = {memRequest_bits_data_lo_hi_31, memRequest_bits_data_lo_lo_31};
  wire [1:0]       memRequest_bits_data_hi_lo_31 = {_memRequest_bits_data_T_503[23], _memRequest_bits_data_T_454[23]};
  wire [1:0]       memRequest_bits_data_hi_hi_31 = {_memRequest_bits_data_T_601[23], _memRequest_bits_data_T_552[23]};
  wire [3:0]       memRequest_bits_data_hi_31 = {memRequest_bits_data_hi_hi_31, memRequest_bits_data_hi_lo_31};
  wire [1:0]       memRequest_bits_data_lo_lo_32 = {_memRequest_bits_data_T_307[24], _memRequest_bits_data_T_258[24]};
  wire [1:0]       memRequest_bits_data_lo_hi_32 = {_memRequest_bits_data_T_405[24], _memRequest_bits_data_T_356[24]};
  wire [3:0]       memRequest_bits_data_lo_32 = {memRequest_bits_data_lo_hi_32, memRequest_bits_data_lo_lo_32};
  wire [1:0]       memRequest_bits_data_hi_lo_32 = {_memRequest_bits_data_T_503[24], _memRequest_bits_data_T_454[24]};
  wire [1:0]       memRequest_bits_data_hi_hi_32 = {_memRequest_bits_data_T_601[24], _memRequest_bits_data_T_552[24]};
  wire [3:0]       memRequest_bits_data_hi_32 = {memRequest_bits_data_hi_hi_32, memRequest_bits_data_hi_lo_32};
  wire [1:0]       memRequest_bits_data_lo_lo_33 = {_memRequest_bits_data_T_307[25], _memRequest_bits_data_T_258[25]};
  wire [1:0]       memRequest_bits_data_lo_hi_33 = {_memRequest_bits_data_T_405[25], _memRequest_bits_data_T_356[25]};
  wire [3:0]       memRequest_bits_data_lo_33 = {memRequest_bits_data_lo_hi_33, memRequest_bits_data_lo_lo_33};
  wire [1:0]       memRequest_bits_data_hi_lo_33 = {_memRequest_bits_data_T_503[25], _memRequest_bits_data_T_454[25]};
  wire [1:0]       memRequest_bits_data_hi_hi_33 = {_memRequest_bits_data_T_601[25], _memRequest_bits_data_T_552[25]};
  wire [3:0]       memRequest_bits_data_hi_33 = {memRequest_bits_data_hi_hi_33, memRequest_bits_data_hi_lo_33};
  wire [1:0]       memRequest_bits_data_lo_lo_34 = {_memRequest_bits_data_T_307[26], _memRequest_bits_data_T_258[26]};
  wire [1:0]       memRequest_bits_data_lo_hi_34 = {_memRequest_bits_data_T_405[26], _memRequest_bits_data_T_356[26]};
  wire [3:0]       memRequest_bits_data_lo_34 = {memRequest_bits_data_lo_hi_34, memRequest_bits_data_lo_lo_34};
  wire [1:0]       memRequest_bits_data_hi_lo_34 = {_memRequest_bits_data_T_503[26], _memRequest_bits_data_T_454[26]};
  wire [1:0]       memRequest_bits_data_hi_hi_34 = {_memRequest_bits_data_T_601[26], _memRequest_bits_data_T_552[26]};
  wire [3:0]       memRequest_bits_data_hi_34 = {memRequest_bits_data_hi_hi_34, memRequest_bits_data_hi_lo_34};
  wire [1:0]       memRequest_bits_data_lo_lo_35 = {_memRequest_bits_data_T_307[27], _memRequest_bits_data_T_258[27]};
  wire [1:0]       memRequest_bits_data_lo_hi_35 = {_memRequest_bits_data_T_405[27], _memRequest_bits_data_T_356[27]};
  wire [3:0]       memRequest_bits_data_lo_35 = {memRequest_bits_data_lo_hi_35, memRequest_bits_data_lo_lo_35};
  wire [1:0]       memRequest_bits_data_hi_lo_35 = {_memRequest_bits_data_T_503[27], _memRequest_bits_data_T_454[27]};
  wire [1:0]       memRequest_bits_data_hi_hi_35 = {_memRequest_bits_data_T_601[27], _memRequest_bits_data_T_552[27]};
  wire [3:0]       memRequest_bits_data_hi_35 = {memRequest_bits_data_hi_hi_35, memRequest_bits_data_hi_lo_35};
  wire [1:0]       memRequest_bits_data_lo_lo_36 = {_memRequest_bits_data_T_307[28], _memRequest_bits_data_T_258[28]};
  wire [1:0]       memRequest_bits_data_lo_hi_36 = {_memRequest_bits_data_T_405[28], _memRequest_bits_data_T_356[28]};
  wire [3:0]       memRequest_bits_data_lo_36 = {memRequest_bits_data_lo_hi_36, memRequest_bits_data_lo_lo_36};
  wire [1:0]       memRequest_bits_data_hi_lo_36 = {_memRequest_bits_data_T_503[28], _memRequest_bits_data_T_454[28]};
  wire [1:0]       memRequest_bits_data_hi_hi_36 = {_memRequest_bits_data_T_601[28], _memRequest_bits_data_T_552[28]};
  wire [3:0]       memRequest_bits_data_hi_36 = {memRequest_bits_data_hi_hi_36, memRequest_bits_data_hi_lo_36};
  wire [1:0]       memRequest_bits_data_lo_lo_37 = {_memRequest_bits_data_T_307[29], _memRequest_bits_data_T_258[29]};
  wire [1:0]       memRequest_bits_data_lo_hi_37 = {_memRequest_bits_data_T_405[29], _memRequest_bits_data_T_356[29]};
  wire [3:0]       memRequest_bits_data_lo_37 = {memRequest_bits_data_lo_hi_37, memRequest_bits_data_lo_lo_37};
  wire [1:0]       memRequest_bits_data_hi_lo_37 = {_memRequest_bits_data_T_503[29], _memRequest_bits_data_T_454[29]};
  wire [1:0]       memRequest_bits_data_hi_hi_37 = {_memRequest_bits_data_T_601[29], _memRequest_bits_data_T_552[29]};
  wire [3:0]       memRequest_bits_data_hi_37 = {memRequest_bits_data_hi_hi_37, memRequest_bits_data_hi_lo_37};
  wire [1:0]       memRequest_bits_data_lo_lo_38 = {_memRequest_bits_data_T_307[30], _memRequest_bits_data_T_258[30]};
  wire [1:0]       memRequest_bits_data_lo_hi_38 = {_memRequest_bits_data_T_405[30], _memRequest_bits_data_T_356[30]};
  wire [3:0]       memRequest_bits_data_lo_38 = {memRequest_bits_data_lo_hi_38, memRequest_bits_data_lo_lo_38};
  wire [1:0]       memRequest_bits_data_hi_lo_38 = {_memRequest_bits_data_T_503[30], _memRequest_bits_data_T_454[30]};
  wire [1:0]       memRequest_bits_data_hi_hi_38 = {_memRequest_bits_data_T_601[30], _memRequest_bits_data_T_552[30]};
  wire [3:0]       memRequest_bits_data_hi_38 = {memRequest_bits_data_hi_hi_38, memRequest_bits_data_hi_lo_38};
  wire [1:0]       memRequest_bits_data_lo_lo_39 = {_memRequest_bits_data_T_307[31], _memRequest_bits_data_T_258[31]};
  wire [1:0]       memRequest_bits_data_lo_hi_39 = {_memRequest_bits_data_T_405[31], _memRequest_bits_data_T_356[31]};
  wire [3:0]       memRequest_bits_data_lo_39 = {memRequest_bits_data_lo_hi_39, memRequest_bits_data_lo_lo_39};
  wire [1:0]       memRequest_bits_data_hi_lo_39 = {_memRequest_bits_data_T_503[31], _memRequest_bits_data_T_454[31]};
  wire [1:0]       memRequest_bits_data_hi_hi_39 = {_memRequest_bits_data_T_601[31], _memRequest_bits_data_T_552[31]};
  wire [3:0]       memRequest_bits_data_hi_39 = {memRequest_bits_data_hi_hi_39, memRequest_bits_data_hi_lo_39};
  wire [1:0]       memRequest_bits_data_lo_lo_40 = {_memRequest_bits_data_T_307[32], _memRequest_bits_data_T_258[32]};
  wire [1:0]       memRequest_bits_data_lo_hi_40 = {_memRequest_bits_data_T_405[32], _memRequest_bits_data_T_356[32]};
  wire [3:0]       memRequest_bits_data_lo_40 = {memRequest_bits_data_lo_hi_40, memRequest_bits_data_lo_lo_40};
  wire [1:0]       memRequest_bits_data_hi_lo_40 = {_memRequest_bits_data_T_503[32], _memRequest_bits_data_T_454[32]};
  wire [1:0]       memRequest_bits_data_hi_hi_40 = {_memRequest_bits_data_T_601[32], _memRequest_bits_data_T_552[32]};
  wire [3:0]       memRequest_bits_data_hi_40 = {memRequest_bits_data_hi_hi_40, memRequest_bits_data_hi_lo_40};
  wire [1:0]       memRequest_bits_data_lo_lo_41 = {_memRequest_bits_data_T_307[33], _memRequest_bits_data_T_258[33]};
  wire [1:0]       memRequest_bits_data_lo_hi_41 = {_memRequest_bits_data_T_405[33], _memRequest_bits_data_T_356[33]};
  wire [3:0]       memRequest_bits_data_lo_41 = {memRequest_bits_data_lo_hi_41, memRequest_bits_data_lo_lo_41};
  wire [1:0]       memRequest_bits_data_hi_lo_41 = {_memRequest_bits_data_T_503[33], _memRequest_bits_data_T_454[33]};
  wire [1:0]       memRequest_bits_data_hi_hi_41 = {_memRequest_bits_data_T_601[33], _memRequest_bits_data_T_552[33]};
  wire [3:0]       memRequest_bits_data_hi_41 = {memRequest_bits_data_hi_hi_41, memRequest_bits_data_hi_lo_41};
  wire [1:0]       memRequest_bits_data_lo_lo_42 = {_memRequest_bits_data_T_307[34], _memRequest_bits_data_T_258[34]};
  wire [1:0]       memRequest_bits_data_lo_hi_42 = {_memRequest_bits_data_T_405[34], _memRequest_bits_data_T_356[34]};
  wire [3:0]       memRequest_bits_data_lo_42 = {memRequest_bits_data_lo_hi_42, memRequest_bits_data_lo_lo_42};
  wire [1:0]       memRequest_bits_data_hi_lo_42 = {_memRequest_bits_data_T_503[34], _memRequest_bits_data_T_454[34]};
  wire [1:0]       memRequest_bits_data_hi_hi_42 = {_memRequest_bits_data_T_601[34], _memRequest_bits_data_T_552[34]};
  wire [3:0]       memRequest_bits_data_hi_42 = {memRequest_bits_data_hi_hi_42, memRequest_bits_data_hi_lo_42};
  wire [1:0]       memRequest_bits_data_lo_lo_43 = {_memRequest_bits_data_T_307[35], _memRequest_bits_data_T_258[35]};
  wire [1:0]       memRequest_bits_data_lo_hi_43 = {_memRequest_bits_data_T_405[35], _memRequest_bits_data_T_356[35]};
  wire [3:0]       memRequest_bits_data_lo_43 = {memRequest_bits_data_lo_hi_43, memRequest_bits_data_lo_lo_43};
  wire [1:0]       memRequest_bits_data_hi_lo_43 = {_memRequest_bits_data_T_503[35], _memRequest_bits_data_T_454[35]};
  wire [1:0]       memRequest_bits_data_hi_hi_43 = {_memRequest_bits_data_T_601[35], _memRequest_bits_data_T_552[35]};
  wire [3:0]       memRequest_bits_data_hi_43 = {memRequest_bits_data_hi_hi_43, memRequest_bits_data_hi_lo_43};
  wire [1:0]       memRequest_bits_data_lo_lo_44 = {_memRequest_bits_data_T_307[36], _memRequest_bits_data_T_258[36]};
  wire [1:0]       memRequest_bits_data_lo_hi_44 = {_memRequest_bits_data_T_405[36], _memRequest_bits_data_T_356[36]};
  wire [3:0]       memRequest_bits_data_lo_44 = {memRequest_bits_data_lo_hi_44, memRequest_bits_data_lo_lo_44};
  wire [1:0]       memRequest_bits_data_hi_lo_44 = {_memRequest_bits_data_T_503[36], _memRequest_bits_data_T_454[36]};
  wire [1:0]       memRequest_bits_data_hi_hi_44 = {_memRequest_bits_data_T_601[36], _memRequest_bits_data_T_552[36]};
  wire [3:0]       memRequest_bits_data_hi_44 = {memRequest_bits_data_hi_hi_44, memRequest_bits_data_hi_lo_44};
  wire [1:0]       memRequest_bits_data_lo_lo_45 = {_memRequest_bits_data_T_307[37], _memRequest_bits_data_T_258[37]};
  wire [1:0]       memRequest_bits_data_lo_hi_45 = {_memRequest_bits_data_T_405[37], _memRequest_bits_data_T_356[37]};
  wire [3:0]       memRequest_bits_data_lo_45 = {memRequest_bits_data_lo_hi_45, memRequest_bits_data_lo_lo_45};
  wire [1:0]       memRequest_bits_data_hi_lo_45 = {_memRequest_bits_data_T_503[37], _memRequest_bits_data_T_454[37]};
  wire [1:0]       memRequest_bits_data_hi_hi_45 = {_memRequest_bits_data_T_601[37], _memRequest_bits_data_T_552[37]};
  wire [3:0]       memRequest_bits_data_hi_45 = {memRequest_bits_data_hi_hi_45, memRequest_bits_data_hi_lo_45};
  wire [1:0]       memRequest_bits_data_lo_lo_46 = {_memRequest_bits_data_T_307[38], _memRequest_bits_data_T_258[38]};
  wire [1:0]       memRequest_bits_data_lo_hi_46 = {_memRequest_bits_data_T_405[38], _memRequest_bits_data_T_356[38]};
  wire [3:0]       memRequest_bits_data_lo_46 = {memRequest_bits_data_lo_hi_46, memRequest_bits_data_lo_lo_46};
  wire [1:0]       memRequest_bits_data_hi_lo_46 = {_memRequest_bits_data_T_503[38], _memRequest_bits_data_T_454[38]};
  wire [1:0]       memRequest_bits_data_hi_hi_46 = {_memRequest_bits_data_T_601[38], _memRequest_bits_data_T_552[38]};
  wire [3:0]       memRequest_bits_data_hi_46 = {memRequest_bits_data_hi_hi_46, memRequest_bits_data_hi_lo_46};
  wire [1:0]       memRequest_bits_data_lo_lo_47 = {_memRequest_bits_data_T_307[39], _memRequest_bits_data_T_258[39]};
  wire [1:0]       memRequest_bits_data_lo_hi_47 = {_memRequest_bits_data_T_405[39], _memRequest_bits_data_T_356[39]};
  wire [3:0]       memRequest_bits_data_lo_47 = {memRequest_bits_data_lo_hi_47, memRequest_bits_data_lo_lo_47};
  wire [1:0]       memRequest_bits_data_hi_lo_47 = {_memRequest_bits_data_T_503[39], _memRequest_bits_data_T_454[39]};
  wire [1:0]       memRequest_bits_data_hi_hi_47 = {_memRequest_bits_data_T_601[39], _memRequest_bits_data_T_552[39]};
  wire [3:0]       memRequest_bits_data_hi_47 = {memRequest_bits_data_hi_hi_47, memRequest_bits_data_hi_lo_47};
  wire [1:0]       memRequest_bits_data_lo_lo_48 = {_memRequest_bits_data_T_307[40], _memRequest_bits_data_T_258[40]};
  wire [1:0]       memRequest_bits_data_lo_hi_48 = {_memRequest_bits_data_T_405[40], _memRequest_bits_data_T_356[40]};
  wire [3:0]       memRequest_bits_data_lo_48 = {memRequest_bits_data_lo_hi_48, memRequest_bits_data_lo_lo_48};
  wire [1:0]       memRequest_bits_data_hi_lo_48 = {_memRequest_bits_data_T_503[40], _memRequest_bits_data_T_454[40]};
  wire [1:0]       memRequest_bits_data_hi_hi_48 = {_memRequest_bits_data_T_601[40], _memRequest_bits_data_T_552[40]};
  wire [3:0]       memRequest_bits_data_hi_48 = {memRequest_bits_data_hi_hi_48, memRequest_bits_data_hi_lo_48};
  wire [1:0]       memRequest_bits_data_lo_lo_49 = {_memRequest_bits_data_T_307[41], _memRequest_bits_data_T_258[41]};
  wire [1:0]       memRequest_bits_data_lo_hi_49 = {_memRequest_bits_data_T_405[41], _memRequest_bits_data_T_356[41]};
  wire [3:0]       memRequest_bits_data_lo_49 = {memRequest_bits_data_lo_hi_49, memRequest_bits_data_lo_lo_49};
  wire [1:0]       memRequest_bits_data_hi_lo_49 = {_memRequest_bits_data_T_503[41], _memRequest_bits_data_T_454[41]};
  wire [1:0]       memRequest_bits_data_hi_hi_49 = {_memRequest_bits_data_T_601[41], _memRequest_bits_data_T_552[41]};
  wire [3:0]       memRequest_bits_data_hi_49 = {memRequest_bits_data_hi_hi_49, memRequest_bits_data_hi_lo_49};
  wire [1:0]       memRequest_bits_data_lo_lo_50 = {_memRequest_bits_data_T_307[42], _memRequest_bits_data_T_258[42]};
  wire [1:0]       memRequest_bits_data_lo_hi_50 = {_memRequest_bits_data_T_405[42], _memRequest_bits_data_T_356[42]};
  wire [3:0]       memRequest_bits_data_lo_50 = {memRequest_bits_data_lo_hi_50, memRequest_bits_data_lo_lo_50};
  wire [1:0]       memRequest_bits_data_hi_lo_50 = {_memRequest_bits_data_T_503[42], _memRequest_bits_data_T_454[42]};
  wire [1:0]       memRequest_bits_data_hi_hi_50 = {_memRequest_bits_data_T_601[42], _memRequest_bits_data_T_552[42]};
  wire [3:0]       memRequest_bits_data_hi_50 = {memRequest_bits_data_hi_hi_50, memRequest_bits_data_hi_lo_50};
  wire [1:0]       memRequest_bits_data_lo_lo_51 = {_memRequest_bits_data_T_307[43], _memRequest_bits_data_T_258[43]};
  wire [1:0]       memRequest_bits_data_lo_hi_51 = {_memRequest_bits_data_T_405[43], _memRequest_bits_data_T_356[43]};
  wire [3:0]       memRequest_bits_data_lo_51 = {memRequest_bits_data_lo_hi_51, memRequest_bits_data_lo_lo_51};
  wire [1:0]       memRequest_bits_data_hi_lo_51 = {_memRequest_bits_data_T_503[43], _memRequest_bits_data_T_454[43]};
  wire [1:0]       memRequest_bits_data_hi_hi_51 = {_memRequest_bits_data_T_601[43], _memRequest_bits_data_T_552[43]};
  wire [3:0]       memRequest_bits_data_hi_51 = {memRequest_bits_data_hi_hi_51, memRequest_bits_data_hi_lo_51};
  wire [1:0]       memRequest_bits_data_lo_lo_52 = {_memRequest_bits_data_T_307[44], _memRequest_bits_data_T_258[44]};
  wire [1:0]       memRequest_bits_data_lo_hi_52 = {_memRequest_bits_data_T_405[44], _memRequest_bits_data_T_356[44]};
  wire [3:0]       memRequest_bits_data_lo_52 = {memRequest_bits_data_lo_hi_52, memRequest_bits_data_lo_lo_52};
  wire [1:0]       memRequest_bits_data_hi_lo_52 = {_memRequest_bits_data_T_503[44], _memRequest_bits_data_T_454[44]};
  wire [1:0]       memRequest_bits_data_hi_hi_52 = {_memRequest_bits_data_T_601[44], _memRequest_bits_data_T_552[44]};
  wire [3:0]       memRequest_bits_data_hi_52 = {memRequest_bits_data_hi_hi_52, memRequest_bits_data_hi_lo_52};
  wire [1:0]       memRequest_bits_data_lo_lo_53 = {_memRequest_bits_data_T_307[45], _memRequest_bits_data_T_258[45]};
  wire [1:0]       memRequest_bits_data_lo_hi_53 = {_memRequest_bits_data_T_405[45], _memRequest_bits_data_T_356[45]};
  wire [3:0]       memRequest_bits_data_lo_53 = {memRequest_bits_data_lo_hi_53, memRequest_bits_data_lo_lo_53};
  wire [1:0]       memRequest_bits_data_hi_lo_53 = {_memRequest_bits_data_T_503[45], _memRequest_bits_data_T_454[45]};
  wire [1:0]       memRequest_bits_data_hi_hi_53 = {_memRequest_bits_data_T_601[45], _memRequest_bits_data_T_552[45]};
  wire [3:0]       memRequest_bits_data_hi_53 = {memRequest_bits_data_hi_hi_53, memRequest_bits_data_hi_lo_53};
  wire [1:0]       memRequest_bits_data_lo_lo_54 = {_memRequest_bits_data_T_307[46], _memRequest_bits_data_T_258[46]};
  wire [1:0]       memRequest_bits_data_lo_hi_54 = {_memRequest_bits_data_T_405[46], _memRequest_bits_data_T_356[46]};
  wire [3:0]       memRequest_bits_data_lo_54 = {memRequest_bits_data_lo_hi_54, memRequest_bits_data_lo_lo_54};
  wire [1:0]       memRequest_bits_data_hi_lo_54 = {_memRequest_bits_data_T_503[46], _memRequest_bits_data_T_454[46]};
  wire [1:0]       memRequest_bits_data_hi_hi_54 = {_memRequest_bits_data_T_601[46], _memRequest_bits_data_T_552[46]};
  wire [3:0]       memRequest_bits_data_hi_54 = {memRequest_bits_data_hi_hi_54, memRequest_bits_data_hi_lo_54};
  wire [15:0]      memRequest_bits_data_lo_lo_lo_lo_8 = {memRequest_bits_data_hi_9, memRequest_bits_data_lo_9, memRequest_bits_data_hi_8, memRequest_bits_data_lo_8};
  wire [15:0]      memRequest_bits_data_lo_lo_lo_hi_hi = {memRequest_bits_data_hi_12, memRequest_bits_data_lo_12, memRequest_bits_data_hi_11, memRequest_bits_data_lo_11};
  wire [23:0]      memRequest_bits_data_lo_lo_lo_hi_8 = {memRequest_bits_data_lo_lo_lo_hi_hi, memRequest_bits_data_hi_10, memRequest_bits_data_lo_10};
  wire [39:0]      memRequest_bits_data_lo_lo_lo_8 = {memRequest_bits_data_lo_lo_lo_hi_8, memRequest_bits_data_lo_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_lo_hi_lo_hi = {memRequest_bits_data_hi_15, memRequest_bits_data_lo_15, memRequest_bits_data_hi_14, memRequest_bits_data_lo_14};
  wire [23:0]      memRequest_bits_data_lo_lo_hi_lo_8 = {memRequest_bits_data_lo_lo_hi_lo_hi, memRequest_bits_data_hi_13, memRequest_bits_data_lo_13};
  wire [15:0]      memRequest_bits_data_lo_lo_hi_hi_hi = {memRequest_bits_data_hi_18, memRequest_bits_data_lo_18, memRequest_bits_data_hi_17, memRequest_bits_data_lo_17};
  wire [23:0]      memRequest_bits_data_lo_lo_hi_hi_8 = {memRequest_bits_data_lo_lo_hi_hi_hi, memRequest_bits_data_hi_16, memRequest_bits_data_lo_16};
  wire [47:0]      memRequest_bits_data_lo_lo_hi_8 = {memRequest_bits_data_lo_lo_hi_hi_8, memRequest_bits_data_lo_lo_hi_lo_8};
  wire [87:0]      memRequest_bits_data_lo_lo_55 = {memRequest_bits_data_lo_lo_hi_8, memRequest_bits_data_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_hi_lo_lo_hi = {memRequest_bits_data_hi_21, memRequest_bits_data_lo_21, memRequest_bits_data_hi_20, memRequest_bits_data_lo_20};
  wire [23:0]      memRequest_bits_data_lo_hi_lo_lo_8 = {memRequest_bits_data_lo_hi_lo_lo_hi, memRequest_bits_data_hi_19, memRequest_bits_data_lo_19};
  wire [15:0]      memRequest_bits_data_lo_hi_lo_hi_hi = {memRequest_bits_data_hi_24, memRequest_bits_data_lo_24, memRequest_bits_data_hi_23, memRequest_bits_data_lo_23};
  wire [23:0]      memRequest_bits_data_lo_hi_lo_hi_8 = {memRequest_bits_data_lo_hi_lo_hi_hi, memRequest_bits_data_hi_22, memRequest_bits_data_lo_22};
  wire [47:0]      memRequest_bits_data_lo_hi_lo_8 = {memRequest_bits_data_lo_hi_lo_hi_8, memRequest_bits_data_lo_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_hi_hi_lo_hi = {memRequest_bits_data_hi_27, memRequest_bits_data_lo_27, memRequest_bits_data_hi_26, memRequest_bits_data_lo_26};
  wire [23:0]      memRequest_bits_data_lo_hi_hi_lo_8 = {memRequest_bits_data_lo_hi_hi_lo_hi, memRequest_bits_data_hi_25, memRequest_bits_data_lo_25};
  wire [15:0]      memRequest_bits_data_lo_hi_hi_hi_hi = {memRequest_bits_data_hi_30, memRequest_bits_data_lo_30, memRequest_bits_data_hi_29, memRequest_bits_data_lo_29};
  wire [23:0]      memRequest_bits_data_lo_hi_hi_hi_8 = {memRequest_bits_data_lo_hi_hi_hi_hi, memRequest_bits_data_hi_28, memRequest_bits_data_lo_28};
  wire [47:0]      memRequest_bits_data_lo_hi_hi_8 = {memRequest_bits_data_lo_hi_hi_hi_8, memRequest_bits_data_lo_hi_hi_lo_8};
  wire [95:0]      memRequest_bits_data_lo_hi_55 = {memRequest_bits_data_lo_hi_hi_8, memRequest_bits_data_lo_hi_lo_8};
  wire [183:0]     memRequest_bits_data_lo_55 = {memRequest_bits_data_lo_hi_55, memRequest_bits_data_lo_lo_55};
  wire [15:0]      memRequest_bits_data_hi_lo_lo_lo_hi = {memRequest_bits_data_hi_33, memRequest_bits_data_lo_33, memRequest_bits_data_hi_32, memRequest_bits_data_lo_32};
  wire [23:0]      memRequest_bits_data_hi_lo_lo_lo_8 = {memRequest_bits_data_hi_lo_lo_lo_hi, memRequest_bits_data_hi_31, memRequest_bits_data_lo_31};
  wire [15:0]      memRequest_bits_data_hi_lo_lo_hi_hi = {memRequest_bits_data_hi_36, memRequest_bits_data_lo_36, memRequest_bits_data_hi_35, memRequest_bits_data_lo_35};
  wire [23:0]      memRequest_bits_data_hi_lo_lo_hi_8 = {memRequest_bits_data_hi_lo_lo_hi_hi, memRequest_bits_data_hi_34, memRequest_bits_data_lo_34};
  wire [47:0]      memRequest_bits_data_hi_lo_lo_8 = {memRequest_bits_data_hi_lo_lo_hi_8, memRequest_bits_data_hi_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_lo_hi_lo_hi = {memRequest_bits_data_hi_39, memRequest_bits_data_lo_39, memRequest_bits_data_hi_38, memRequest_bits_data_lo_38};
  wire [23:0]      memRequest_bits_data_hi_lo_hi_lo_8 = {memRequest_bits_data_hi_lo_hi_lo_hi, memRequest_bits_data_hi_37, memRequest_bits_data_lo_37};
  wire [15:0]      memRequest_bits_data_hi_lo_hi_hi_hi = {memRequest_bits_data_hi_42, memRequest_bits_data_lo_42, memRequest_bits_data_hi_41, memRequest_bits_data_lo_41};
  wire [23:0]      memRequest_bits_data_hi_lo_hi_hi_8 = {memRequest_bits_data_hi_lo_hi_hi_hi, memRequest_bits_data_hi_40, memRequest_bits_data_lo_40};
  wire [47:0]      memRequest_bits_data_hi_lo_hi_8 = {memRequest_bits_data_hi_lo_hi_hi_8, memRequest_bits_data_hi_lo_hi_lo_8};
  wire [95:0]      memRequest_bits_data_hi_lo_55 = {memRequest_bits_data_hi_lo_hi_8, memRequest_bits_data_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_hi_lo_lo_hi = {memRequest_bits_data_hi_45, memRequest_bits_data_lo_45, memRequest_bits_data_hi_44, memRequest_bits_data_lo_44};
  wire [23:0]      memRequest_bits_data_hi_hi_lo_lo_8 = {memRequest_bits_data_hi_hi_lo_lo_hi, memRequest_bits_data_hi_43, memRequest_bits_data_lo_43};
  wire [15:0]      memRequest_bits_data_hi_hi_lo_hi_hi = {memRequest_bits_data_hi_48, memRequest_bits_data_lo_48, memRequest_bits_data_hi_47, memRequest_bits_data_lo_47};
  wire [23:0]      memRequest_bits_data_hi_hi_lo_hi_8 = {memRequest_bits_data_hi_hi_lo_hi_hi, memRequest_bits_data_hi_46, memRequest_bits_data_lo_46};
  wire [47:0]      memRequest_bits_data_hi_hi_lo_8 = {memRequest_bits_data_hi_hi_lo_hi_8, memRequest_bits_data_hi_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_hi_hi_lo_hi = {memRequest_bits_data_hi_51, memRequest_bits_data_lo_51, memRequest_bits_data_hi_50, memRequest_bits_data_lo_50};
  wire [23:0]      memRequest_bits_data_hi_hi_hi_lo_8 = {memRequest_bits_data_hi_hi_hi_lo_hi, memRequest_bits_data_hi_49, memRequest_bits_data_lo_49};
  wire [15:0]      memRequest_bits_data_hi_hi_hi_hi_hi = {memRequest_bits_data_hi_54, memRequest_bits_data_lo_54, memRequest_bits_data_hi_53, memRequest_bits_data_lo_53};
  wire [23:0]      memRequest_bits_data_hi_hi_hi_hi_8 = {memRequest_bits_data_hi_hi_hi_hi_hi, memRequest_bits_data_hi_52, memRequest_bits_data_lo_52};
  wire [47:0]      memRequest_bits_data_hi_hi_hi_8 = {memRequest_bits_data_hi_hi_hi_hi_8, memRequest_bits_data_hi_hi_hi_lo_8};
  wire [95:0]      memRequest_bits_data_hi_hi_55 = {memRequest_bits_data_hi_hi_hi_8, memRequest_bits_data_hi_hi_lo_8};
  wire [191:0]     memRequest_bits_data_hi_55 = {memRequest_bits_data_hi_hi_55, memRequest_bits_data_hi_lo_55};
  wire [127:0]     memRequest_bits_data_0 = {memRequest_bits_data_hi_55[71:0], memRequest_bits_data_lo_55[183:128]};
  wire [15:0]      selectMaskForTail = bufferValid ? _GEN_146 : 16'h0;
  wire [46:0]      _memRequest_bits_mask_T_1 = {15'h0, selectMaskForTail, maskTemp} << _GEN_147;
  wire [15:0]      memRequest_bits_mask_0 = _memRequest_bits_mask_T_1[31:16];
  assign alignedDequeueAddress = {lsuRequestReg_rs1Data[31:4] + {19'h0, bufferBaseCacheLineIndex}, 4'h0};
  wire [31:0]      memRequest_bits_address_0 = alignedDequeueAddress;
  wire [31:0]      addressQueue_enq_bits = alignedDequeueAddress;
  assign addressQueueFree = addressQueue_enq_ready;
  wire             addressQueue_deq_valid;
  assign addressQueue_deq_valid = ~_addressQueue_fifo_empty;
  assign addressQueue_enq_ready = ~_addressQueue_fifo_full;
  wire             _status_idle_output = ~bufferValid & ~readStageValid & readQueueClear & ~bufferFull & ~addressQueue_deq_valid;
  reg              idleNext;
  wire [31:0]      addressQueue_deq_bits;
  always @(posedge clock) begin
    if (reset) begin
      lsuRequestReg_instructionInformation_nf <= 3'h0;
      lsuRequestReg_instructionInformation_mew <= 1'h0;
      lsuRequestReg_instructionInformation_mop <= 2'h0;
      lsuRequestReg_instructionInformation_lumop <= 5'h0;
      lsuRequestReg_instructionInformation_eew <= 2'h0;
      lsuRequestReg_instructionInformation_vs3 <= 5'h0;
      lsuRequestReg_instructionInformation_isStore <= 1'h0;
      lsuRequestReg_instructionInformation_maskedLoadStore <= 1'h0;
      lsuRequestReg_rs1Data <= 32'h0;
      lsuRequestReg_rs2Data <= 32'h0;
      lsuRequestReg_instructionIndex <= 3'h0;
      csrInterfaceReg_vl <= 13'h0;
      csrInterfaceReg_vStart <= 13'h0;
      csrInterfaceReg_vlmul <= 3'h0;
      csrInterfaceReg_vSew <= 2'h0;
      csrInterfaceReg_vxrm <= 2'h0;
      csrInterfaceReg_vta <= 1'h0;
      csrInterfaceReg_vma <= 1'h0;
      requestFireNext <= 1'h0;
      dataEEW <= 2'h0;
      maskReg <= 16'h0;
      needAmend <= 1'h0;
      lastMaskAmendReg <= 15'h0;
      maskGroupCounter <= 8'h0;
      maskCounterInGroup <= 2'h0;
      isLastMaskGroup <= 1'h0;
      accessData_0 <= 128'h0;
      accessData_1 <= 128'h0;
      accessData_2 <= 128'h0;
      accessData_3 <= 128'h0;
      accessData_4 <= 128'h0;
      accessData_5 <= 128'h0;
      accessData_6 <= 128'h0;
      accessData_7 <= 128'h0;
      accessPtr <= 3'h0;
      dataGroup <= 8'h0;
      dataBuffer_0 <= 128'h0;
      dataBuffer_1 <= 128'h0;
      dataBuffer_2 <= 128'h0;
      dataBuffer_3 <= 128'h0;
      dataBuffer_4 <= 128'h0;
      dataBuffer_5 <= 128'h0;
      dataBuffer_6 <= 128'h0;
      dataBuffer_7 <= 128'h0;
      bufferBaseCacheLineIndex <= 9'h0;
      cacheLineIndexInBuffer <= 3'h0;
      segmentInstructionIndexInterval <= 4'h0;
      lastWriteVrfIndexReg <= 16'h0;
      lastCacheNeedPush <= 1'h0;
      cacheLineNumberReg <= 16'h0;
      lastDataGroupReg <= 12'h0;
      hazardCheck <= 1'h0;
      readStageValid_segPtr <= 3'h0;
      readStageValid_readCount <= 8'h0;
      readStageValid_stageValid <= 1'h0;
      readStageValid_readCounter <= 4'h0;
      readStageValid_segPtr_1 <= 3'h0;
      readStageValid_readCount_1 <= 8'h0;
      readStageValid_stageValid_1 <= 1'h0;
      readStageValid_readCounter_1 <= 4'h0;
      readStageValid_segPtr_2 <= 3'h0;
      readStageValid_readCount_2 <= 8'h0;
      readStageValid_stageValid_2 <= 1'h0;
      readStageValid_readCounter_2 <= 4'h0;
      readStageValid_segPtr_3 <= 3'h0;
      readStageValid_readCount_3 <= 8'h0;
      readStageValid_stageValid_3 <= 1'h0;
      readStageValid_readCounter_3 <= 4'h0;
      bufferFull <= 1'h0;
      bufferValid <= 1'h0;
      maskForBufferData_0 <= 16'h0;
      maskForBufferData_1 <= 16'h0;
      maskForBufferData_2 <= 16'h0;
      maskForBufferData_3 <= 16'h0;
      maskForBufferData_4 <= 16'h0;
      maskForBufferData_5 <= 16'h0;
      maskForBufferData_6 <= 16'h0;
      maskForBufferData_7 <= 16'h0;
      lastDataGroupInDataBuffer <= 1'h0;
      cacheLineTemp <= 128'h0;
      maskTemp <= 16'h0;
      canSendTail <= 1'h0;
      idleNext <= 1'h1;
    end
    else begin
      if (lsuRequest_valid) begin
        lsuRequestReg_instructionInformation_nf <= nfCorrection;
        lsuRequestReg_instructionInformation_mew <= ~invalidInstruction & lsuRequest_bits_instructionInformation_mew;
        lsuRequestReg_instructionInformation_mop <= invalidInstruction ? 2'h0 : lsuRequest_bits_instructionInformation_mop;
        lsuRequestReg_instructionInformation_lumop <= invalidInstruction ? 5'h0 : lsuRequest_bits_instructionInformation_lumop;
        lsuRequestReg_instructionInformation_eew <= invalidInstruction ? 2'h0 : lsuRequest_bits_instructionInformation_eew;
        lsuRequestReg_instructionInformation_vs3 <= invalidInstruction ? 5'h0 : lsuRequest_bits_instructionInformation_vs3;
        lsuRequestReg_instructionInformation_isStore <= ~invalidInstruction & lsuRequest_bits_instructionInformation_isStore;
        lsuRequestReg_instructionInformation_maskedLoadStore <= ~invalidInstruction & lsuRequest_bits_instructionInformation_maskedLoadStore;
        lsuRequestReg_rs1Data <= invalidInstruction ? 32'h0 : lsuRequest_bits_rs1Data;
        lsuRequestReg_rs2Data <= invalidInstruction ? 32'h0 : lsuRequest_bits_rs2Data;
        lsuRequestReg_instructionIndex <= lsuRequest_bits_instructionIndex;
        csrInterfaceReg_vl <= csrInterface_vl;
        csrInterfaceReg_vStart <= csrInterface_vStart;
        csrInterfaceReg_vlmul <= csrInterface_vlmul;
        csrInterfaceReg_vSew <= csrInterface_vSew;
        csrInterfaceReg_vxrm <= csrInterface_vxrm;
        csrInterfaceReg_vta <= csrInterface_vta;
        csrInterfaceReg_vma <= csrInterface_vma;
        dataEEW <= lsuRequest_bits_instructionInformation_eew;
        needAmend <= |(csrInterface_vl[3:0]);
        lastMaskAmendReg <= lastMaskAmend;
        segmentInstructionIndexInterval <= csrInterface_vlmul[2] ? 4'h1 : 4'h1 << csrInterface_vlmul[1:0];
        lastWriteVrfIndexReg <= lastWriteVrfIndex;
        lastCacheNeedPush <= lastCacheLineIndex == lastWriteVrfIndex;
        cacheLineNumberReg <= lastCacheLineIndex;
        lastDataGroupReg <= lastDataGroupForInstruction;
      end
      requestFireNext <= lsuRequest_valid;
      if (_maskSelect_valid_output | lsuRequest_valid) begin
        maskReg <= maskAmend;
        isLastMaskGroup <= lsuRequest_valid ? csrInterface_vl[12:4] == 9'h0 : {1'h0, _maskSelect_bits_output} == csrInterfaceReg_vl[12:4];
      end
      if (_GEN_143 & (_GEN_144 | lsuRequest_valid))
        maskGroupCounter <= _maskSelect_bits_output;
      if (_GEN_143) begin
        maskCounterInGroup <= isLastDataGroup | lsuRequest_valid ? 2'h0 : nextMaskCount;
        dataGroup <= nextDataGroup;
      end
      if (accessBufferDequeueFire | accessBufferEnqueueFire | requestFireNext) begin
        accessData_0 <= accessDataUpdate_0;
        accessData_1 <= accessDataUpdate_1;
        accessData_2 <= accessDataUpdate_2;
        accessData_3 <= accessDataUpdate_3;
        accessData_4 <= accessDataUpdate_4;
        accessData_5 <= accessDataUpdate_5;
        accessData_6 <= accessDataUpdate_6;
        accessData_7 <= accessDataUpdate_7;
        accessPtr <= accessBufferDequeueFire | lastPtr | requestFireNext ? lsuRequestReg_instructionInformation_nf - {2'h0, accessBufferEnqueueFire & ~lastPtr} : accessPtr - 3'h1;
      end
      if (accessBufferDequeueFire) begin
        automatic logic [1023:0] _GEN_148 =
          (dataEEWOH[0]
             ? (_fillBySeg_T[0] ? regroupLoadData_0_0 : 1024'h0) | (_fillBySeg_T[1] ? regroupLoadData_0_1 : 1024'h0) | (_fillBySeg_T[2] ? regroupLoadData_0_2 : 1024'h0) | (_fillBySeg_T[3] ? regroupLoadData_0_3 : 1024'h0)
               | (_fillBySeg_T[4] ? regroupLoadData_0_4 : 1024'h0) | (_fillBySeg_T[5] ? regroupLoadData_0_5 : 1024'h0) | (_fillBySeg_T[6] ? regroupLoadData_0_6 : 1024'h0) | (_fillBySeg_T[7] ? regroupLoadData_0_7 : 1024'h0)
             : 1024'h0)
          | (dataEEWOH[1]
               ? (_fillBySeg_T[0] ? regroupLoadData_1_0 : 1024'h0) | (_fillBySeg_T[1] ? regroupLoadData_1_1 : 1024'h0) | (_fillBySeg_T[2] ? regroupLoadData_1_2 : 1024'h0) | (_fillBySeg_T[3] ? regroupLoadData_1_3 : 1024'h0)
                 | (_fillBySeg_T[4] ? regroupLoadData_1_4 : 1024'h0) | (_fillBySeg_T[5] ? regroupLoadData_1_5 : 1024'h0) | (_fillBySeg_T[6] ? regroupLoadData_1_6 : 1024'h0) | (_fillBySeg_T[7] ? regroupLoadData_1_7 : 1024'h0)
               : 1024'h0)
          | (dataEEWOH[2]
               ? (_fillBySeg_T[0] ? regroupLoadData_2_0 : 1024'h0) | (_fillBySeg_T[1] ? regroupLoadData_2_1 : 1024'h0) | (_fillBySeg_T[2] ? regroupLoadData_2_2 : 1024'h0) | (_fillBySeg_T[3] ? regroupLoadData_2_3 : 1024'h0)
                 | (_fillBySeg_T[4] ? regroupLoadData_2_4 : 1024'h0) | (_fillBySeg_T[5] ? regroupLoadData_2_5 : 1024'h0) | (_fillBySeg_T[6] ? regroupLoadData_2_6 : 1024'h0) | (_fillBySeg_T[7] ? regroupLoadData_2_7 : 1024'h0)
               : 1024'h0);
        dataBuffer_0 <= _GEN_148[127:0];
        dataBuffer_1 <= _GEN_148[255:128];
        dataBuffer_2 <= _GEN_148[383:256];
        dataBuffer_3 <= _GEN_148[511:384];
        dataBuffer_4 <= _GEN_148[639:512];
        dataBuffer_5 <= _GEN_148[767:640];
        dataBuffer_6 <= _GEN_148[895:768];
        dataBuffer_7 <= _GEN_148[1023:896];
        maskForBufferData_0 <= fillBySeg[15:0];
        maskForBufferData_1 <= fillBySeg[31:16];
        maskForBufferData_2 <= fillBySeg[47:32];
        maskForBufferData_3 <= fillBySeg[63:48];
        maskForBufferData_4 <= fillBySeg[79:64];
        maskForBufferData_5 <= fillBySeg[95:80];
        maskForBufferData_6 <= fillBySeg[111:96];
        maskForBufferData_7 <= fillBySeg[127:112];
        lastDataGroupInDataBuffer <= isLastRead;
      end
      else if (alignedDequeueFire) begin
        dataBuffer_0 <= dataBuffer_1;
        dataBuffer_1 <= dataBuffer_2;
        dataBuffer_2 <= dataBuffer_3;
        dataBuffer_3 <= dataBuffer_4;
        dataBuffer_4 <= dataBuffer_5;
        dataBuffer_5 <= dataBuffer_6;
        dataBuffer_6 <= dataBuffer_7;
        dataBuffer_7 <= 128'h0;
      end
      if (lsuRequest_valid | alignedDequeueFire) begin
        bufferBaseCacheLineIndex <= lsuRequest_valid ? 9'h0 : bufferBaseCacheLineIndex + 9'h1;
        maskTemp <= lsuRequest_valid ? 16'h0 : _GEN_146;
        canSendTail <= ~lsuRequest_valid & bufferValid & isLastCacheLineInBuffer & lastDataGroupInDataBuffer;
      end
      if (accessBufferDequeueFire | alignedDequeueFire)
        cacheLineIndexInBuffer <= accessBufferDequeueFire ? 3'h0 : cacheLineIndexInBuffer + 3'h1;
      hazardCheck <= ~lsuRequest_valid;
      if (lsuRequest_valid | _readStageValid_T_11)
        readStageValid_segPtr <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_11 & readStageValid_lastReadPtr)
        readStageValid_readCount <= readStageValid_nextReadCount;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup & readStageValid_lastReadPtr & _readStageValid_T_11)
        readStageValid_stageValid <= lsuRequest_valid;
      if (_readStageValid_T_11 ^ vrfReadQueueVec_0_deq_ready & vrfReadQueueVec_0_deq_valid)
        readStageValid_readCounter <= readStageValid_readCounter + readStageValid_counterChange;
      if (lsuRequest_valid | _readStageValid_T_30)
        readStageValid_segPtr_1 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_1 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_1 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_30 & readStageValid_lastReadPtr_1)
        readStageValid_readCount_1 <= readStageValid_nextReadCount_1;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_1 & readStageValid_lastReadPtr_1 & _readStageValid_T_30)
        readStageValid_stageValid_1 <= lsuRequest_valid;
      if (_readStageValid_T_30 ^ vrfReadQueueVec_1_deq_ready & vrfReadQueueVec_1_deq_valid)
        readStageValid_readCounter_1 <= readStageValid_readCounter_1 + readStageValid_counterChange_1;
      if (lsuRequest_valid | _readStageValid_T_49)
        readStageValid_segPtr_2 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_2 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_2 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_49 & readStageValid_lastReadPtr_2)
        readStageValid_readCount_2 <= readStageValid_nextReadCount_2;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_2 & readStageValid_lastReadPtr_2 & _readStageValid_T_49)
        readStageValid_stageValid_2 <= lsuRequest_valid;
      if (_readStageValid_T_49 ^ vrfReadQueueVec_2_deq_ready & vrfReadQueueVec_2_deq_valid)
        readStageValid_readCounter_2 <= readStageValid_readCounter_2 + readStageValid_counterChange_2;
      if (lsuRequest_valid | _readStageValid_T_68)
        readStageValid_segPtr_3 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_3 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_3 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_68 & readStageValid_lastReadPtr_3)
        readStageValid_readCount_3 <= readStageValid_nextReadCount_3;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_3 & readStageValid_lastReadPtr_3 & _readStageValid_T_68)
        readStageValid_stageValid_3 <= lsuRequest_valid;
      if (_readStageValid_T_68 ^ vrfReadQueueVec_3_deq_ready & vrfReadQueueVec_3_deq_valid)
        readStageValid_readCounter_3 <= readStageValid_readCounter_3 + readStageValid_counterChange_3;
      if (lastPtrEnq ^ accessBufferDequeueFire)
        bufferFull <= lastPtrEnq;
      if (accessBufferDequeueFire ^ bufferWillClear)
        bufferValid <= accessBufferDequeueFire;
      if (alignedDequeueFire)
        cacheLineTemp <= dataBuffer_0;
      idleNext <= _status_idle_output;
    end
    invalidInstructionNext <= invalidInstruction & lsuRequest_valid;
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:82];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [6:0] i = 7'h0; i < 7'h53; i += 7'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        lsuRequestReg_instructionInformation_nf = _RANDOM[7'h0][2:0];
        lsuRequestReg_instructionInformation_mew = _RANDOM[7'h0][3];
        lsuRequestReg_instructionInformation_mop = _RANDOM[7'h0][5:4];
        lsuRequestReg_instructionInformation_lumop = _RANDOM[7'h0][10:6];
        lsuRequestReg_instructionInformation_eew = _RANDOM[7'h0][12:11];
        lsuRequestReg_instructionInformation_vs3 = _RANDOM[7'h0][17:13];
        lsuRequestReg_instructionInformation_isStore = _RANDOM[7'h0][18];
        lsuRequestReg_instructionInformation_maskedLoadStore = _RANDOM[7'h0][19];
        lsuRequestReg_rs1Data = {_RANDOM[7'h0][31:20], _RANDOM[7'h1][19:0]};
        lsuRequestReg_rs2Data = {_RANDOM[7'h1][31:20], _RANDOM[7'h2][19:0]};
        lsuRequestReg_instructionIndex = _RANDOM[7'h2][22:20];
        csrInterfaceReg_vl = {_RANDOM[7'h2][31:23], _RANDOM[7'h3][3:0]};
        csrInterfaceReg_vStart = _RANDOM[7'h3][16:4];
        csrInterfaceReg_vlmul = _RANDOM[7'h3][19:17];
        csrInterfaceReg_vSew = _RANDOM[7'h3][21:20];
        csrInterfaceReg_vxrm = _RANDOM[7'h3][23:22];
        csrInterfaceReg_vta = _RANDOM[7'h3][24];
        csrInterfaceReg_vma = _RANDOM[7'h3][25];
        requestFireNext = _RANDOM[7'h3][26];
        dataEEW = _RANDOM[7'h3][28:27];
        maskReg = {_RANDOM[7'h3][31:29], _RANDOM[7'h4][12:0]};
        needAmend = _RANDOM[7'h4][13];
        lastMaskAmendReg = _RANDOM[7'h4][28:14];
        maskGroupCounter = {_RANDOM[7'h4][31:29], _RANDOM[7'h5][4:0]};
        maskCounterInGroup = _RANDOM[7'h5][6:5];
        isLastMaskGroup = _RANDOM[7'h5][23];
        accessData_0 = {_RANDOM[7'h5][31:24], _RANDOM[7'h6], _RANDOM[7'h7], _RANDOM[7'h8], _RANDOM[7'h9][23:0]};
        accessData_1 = {_RANDOM[7'h9][31:24], _RANDOM[7'hA], _RANDOM[7'hB], _RANDOM[7'hC], _RANDOM[7'hD][23:0]};
        accessData_2 = {_RANDOM[7'hD][31:24], _RANDOM[7'hE], _RANDOM[7'hF], _RANDOM[7'h10], _RANDOM[7'h11][23:0]};
        accessData_3 = {_RANDOM[7'h11][31:24], _RANDOM[7'h12], _RANDOM[7'h13], _RANDOM[7'h14], _RANDOM[7'h15][23:0]};
        accessData_4 = {_RANDOM[7'h15][31:24], _RANDOM[7'h16], _RANDOM[7'h17], _RANDOM[7'h18], _RANDOM[7'h19][23:0]};
        accessData_5 = {_RANDOM[7'h19][31:24], _RANDOM[7'h1A], _RANDOM[7'h1B], _RANDOM[7'h1C], _RANDOM[7'h1D][23:0]};
        accessData_6 = {_RANDOM[7'h1D][31:24], _RANDOM[7'h1E], _RANDOM[7'h1F], _RANDOM[7'h20], _RANDOM[7'h21][23:0]};
        accessData_7 = {_RANDOM[7'h21][31:24], _RANDOM[7'h22], _RANDOM[7'h23], _RANDOM[7'h24], _RANDOM[7'h25][23:0]};
        accessPtr = _RANDOM[7'h25][26:24];
        dataGroup = {_RANDOM[7'h25][31], _RANDOM[7'h26][6:0]};
        dataBuffer_0 = {_RANDOM[7'h26][31:7], _RANDOM[7'h27], _RANDOM[7'h28], _RANDOM[7'h29], _RANDOM[7'h2A][6:0]};
        dataBuffer_1 = {_RANDOM[7'h2A][31:7], _RANDOM[7'h2B], _RANDOM[7'h2C], _RANDOM[7'h2D], _RANDOM[7'h2E][6:0]};
        dataBuffer_2 = {_RANDOM[7'h2E][31:7], _RANDOM[7'h2F], _RANDOM[7'h30], _RANDOM[7'h31], _RANDOM[7'h32][6:0]};
        dataBuffer_3 = {_RANDOM[7'h32][31:7], _RANDOM[7'h33], _RANDOM[7'h34], _RANDOM[7'h35], _RANDOM[7'h36][6:0]};
        dataBuffer_4 = {_RANDOM[7'h36][31:7], _RANDOM[7'h37], _RANDOM[7'h38], _RANDOM[7'h39], _RANDOM[7'h3A][6:0]};
        dataBuffer_5 = {_RANDOM[7'h3A][31:7], _RANDOM[7'h3B], _RANDOM[7'h3C], _RANDOM[7'h3D], _RANDOM[7'h3E][6:0]};
        dataBuffer_6 = {_RANDOM[7'h3E][31:7], _RANDOM[7'h3F], _RANDOM[7'h40], _RANDOM[7'h41], _RANDOM[7'h42][6:0]};
        dataBuffer_7 = {_RANDOM[7'h42][31:7], _RANDOM[7'h43], _RANDOM[7'h44], _RANDOM[7'h45], _RANDOM[7'h46][6:0]};
        bufferBaseCacheLineIndex = _RANDOM[7'h46][15:7];
        cacheLineIndexInBuffer = _RANDOM[7'h46][18:16];
        invalidInstructionNext = _RANDOM[7'h46][19];
        segmentInstructionIndexInterval = _RANDOM[7'h46][23:20];
        lastWriteVrfIndexReg = {_RANDOM[7'h46][31:24], _RANDOM[7'h47][7:0]};
        lastCacheNeedPush = _RANDOM[7'h47][8];
        cacheLineNumberReg = _RANDOM[7'h47][24:9];
        lastDataGroupReg = {_RANDOM[7'h47][31:25], _RANDOM[7'h48][4:0]};
        hazardCheck = _RANDOM[7'h48][5];
        readStageValid_segPtr = _RANDOM[7'h48][8:6];
        readStageValid_readCount = _RANDOM[7'h48][16:9];
        readStageValid_stageValid = _RANDOM[7'h48][17];
        readStageValid_readCounter = _RANDOM[7'h48][21:18];
        readStageValid_segPtr_1 = _RANDOM[7'h48][24:22];
        readStageValid_readCount_1 = {_RANDOM[7'h48][31:25], _RANDOM[7'h49][0]};
        readStageValid_stageValid_1 = _RANDOM[7'h49][1];
        readStageValid_readCounter_1 = _RANDOM[7'h49][5:2];
        readStageValid_segPtr_2 = _RANDOM[7'h49][8:6];
        readStageValid_readCount_2 = _RANDOM[7'h49][16:9];
        readStageValid_stageValid_2 = _RANDOM[7'h49][17];
        readStageValid_readCounter_2 = _RANDOM[7'h49][21:18];
        readStageValid_segPtr_3 = _RANDOM[7'h49][24:22];
        readStageValid_readCount_3 = {_RANDOM[7'h49][31:25], _RANDOM[7'h4A][0]};
        readStageValid_stageValid_3 = _RANDOM[7'h4A][1];
        readStageValid_readCounter_3 = _RANDOM[7'h4A][5:2];
        bufferFull = _RANDOM[7'h4A][6];
        bufferValid = _RANDOM[7'h4A][7];
        maskForBufferData_0 = _RANDOM[7'h4A][23:8];
        maskForBufferData_1 = {_RANDOM[7'h4A][31:24], _RANDOM[7'h4B][7:0]};
        maskForBufferData_2 = _RANDOM[7'h4B][23:8];
        maskForBufferData_3 = {_RANDOM[7'h4B][31:24], _RANDOM[7'h4C][7:0]};
        maskForBufferData_4 = _RANDOM[7'h4C][23:8];
        maskForBufferData_5 = {_RANDOM[7'h4C][31:24], _RANDOM[7'h4D][7:0]};
        maskForBufferData_6 = _RANDOM[7'h4D][23:8];
        maskForBufferData_7 = {_RANDOM[7'h4D][31:24], _RANDOM[7'h4E][7:0]};
        lastDataGroupInDataBuffer = _RANDOM[7'h4E][8];
        cacheLineTemp = {_RANDOM[7'h4E][31:9], _RANDOM[7'h4F], _RANDOM[7'h50], _RANDOM[7'h51], _RANDOM[7'h52][8:0]};
        maskTemp = _RANDOM[7'h52][24:9];
        canSendTail = _RANDOM[7'h52][25];
        idleNext = _RANDOM[7'h52][26];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  wire             vrfReadQueueVec_0_empty;
  assign vrfReadQueueVec_0_empty = _vrfReadQueueVec_fifo_empty;
  wire             vrfReadQueueVec_0_full;
  assign vrfReadQueueVec_0_full = _vrfReadQueueVec_fifo_full;
  wire             vrfReadQueueVec_1_empty;
  assign vrfReadQueueVec_1_empty = _vrfReadQueueVec_fifo_1_empty;
  wire             vrfReadQueueVec_1_full;
  assign vrfReadQueueVec_1_full = _vrfReadQueueVec_fifo_1_full;
  wire             vrfReadQueueVec_2_empty;
  assign vrfReadQueueVec_2_empty = _vrfReadQueueVec_fifo_2_empty;
  wire             vrfReadQueueVec_2_full;
  assign vrfReadQueueVec_2_full = _vrfReadQueueVec_fifo_2_full;
  wire             vrfReadQueueVec_3_empty;
  assign vrfReadQueueVec_3_empty = _vrfReadQueueVec_fifo_3_empty;
  wire             vrfReadQueueVec_3_full;
  assign vrfReadQueueVec_3_full = _vrfReadQueueVec_fifo_3_full;
  wire             addressQueue_empty;
  assign addressQueue_empty = _addressQueue_fifo_empty;
  wire             addressQueue_full;
  assign addressQueue_full = _addressQueue_fifo_full;
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_0_enq_ready & vrfReadQueueVec_0_enq_valid & ~(_vrfReadQueueVec_fifo_empty & vrfReadQueueVec_0_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_0_deq_ready & ~_vrfReadQueueVec_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_0_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_empty),
    .almost_empty (vrfReadQueueVec_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_0_almostFull),
    .full         (_vrfReadQueueVec_fifo_full),
    .error        (_vrfReadQueueVec_fifo_error),
    .data_out     (_vrfReadQueueVec_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_1_enq_ready & vrfReadQueueVec_1_enq_valid & ~(_vrfReadQueueVec_fifo_1_empty & vrfReadQueueVec_1_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_1_deq_ready & ~_vrfReadQueueVec_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_1_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_1_empty),
    .almost_empty (vrfReadQueueVec_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_1_almostFull),
    .full         (_vrfReadQueueVec_fifo_1_full),
    .error        (_vrfReadQueueVec_fifo_1_error),
    .data_out     (_vrfReadQueueVec_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_2_enq_ready & vrfReadQueueVec_2_enq_valid & ~(_vrfReadQueueVec_fifo_2_empty & vrfReadQueueVec_2_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_2_deq_ready & ~_vrfReadQueueVec_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_2_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_2_empty),
    .almost_empty (vrfReadQueueVec_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_2_almostFull),
    .full         (_vrfReadQueueVec_fifo_2_full),
    .error        (_vrfReadQueueVec_fifo_2_error),
    .data_out     (_vrfReadQueueVec_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_3_enq_ready & vrfReadQueueVec_3_enq_valid & ~(_vrfReadQueueVec_fifo_3_empty & vrfReadQueueVec_3_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_3_deq_ready & ~_vrfReadQueueVec_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_3_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_3_empty),
    .almost_empty (vrfReadQueueVec_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_3_almostFull),
    .full         (_vrfReadQueueVec_fifo_3_full),
    .error        (_vrfReadQueueVec_fifo_3_error),
    .data_out     (_vrfReadQueueVec_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) addressQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(addressQueue_enq_ready & addressQueue_enq_valid)),
    .pop_req_n    (~(addressQueue_deq_ready & ~_addressQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (addressQueue_enq_bits),
    .empty        (_addressQueue_fifo_empty),
    .almost_empty (addressQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (addressQueue_almostFull),
    .full         (_addressQueue_fifo_full),
    .error        (_addressQueue_fifo_error),
    .data_out     (addressQueue_deq_bits)
  );
  assign maskSelect_valid = _maskSelect_valid_output;
  assign maskSelect_bits = _maskSelect_bits_output;
  assign memRequest_valid = memRequest_valid_0;
  assign memRequest_bits_data = memRequest_bits_data_0;
  assign memRequest_bits_mask = memRequest_bits_mask_0;
  assign memRequest_bits_index = memRequest_bits_index_0;
  assign memRequest_bits_address = memRequest_bits_address_0;
  assign status_idle = _status_idle_output;
  assign status_last = ~idleNext & _status_idle_output | invalidInstructionNext;
  assign status_instructionIndex = lsuRequestReg_instructionIndex;
  assign status_changeMaskGroup = _maskSelect_valid_output & ~lsuRequest_valid;
  assign status_startAddress = addressQueue_deq_valid ? addressQueue_deq_bits : alignedDequeueAddress;
  assign status_endAddress = {lsuRequestReg_rs1Data[31:4] + {12'h0, cacheLineNumberReg}, 4'h0};
  assign vrfReadDataPorts_0_valid = vrfReadDataPorts_0_valid_0;
  assign vrfReadDataPorts_0_bits_vs = vrfReadDataPorts_0_bits_vs_0;
  assign vrfReadDataPorts_0_bits_offset = vrfReadDataPorts_0_bits_offset_0;
  assign vrfReadDataPorts_0_bits_instructionIndex = vrfReadDataPorts_0_bits_instructionIndex_0;
  assign vrfReadDataPorts_1_valid = vrfReadDataPorts_1_valid_0;
  assign vrfReadDataPorts_1_bits_vs = vrfReadDataPorts_1_bits_vs_0;
  assign vrfReadDataPorts_1_bits_offset = vrfReadDataPorts_1_bits_offset_0;
  assign vrfReadDataPorts_1_bits_instructionIndex = vrfReadDataPorts_1_bits_instructionIndex_0;
  assign vrfReadDataPorts_2_valid = vrfReadDataPorts_2_valid_0;
  assign vrfReadDataPorts_2_bits_vs = vrfReadDataPorts_2_bits_vs_0;
  assign vrfReadDataPorts_2_bits_offset = vrfReadDataPorts_2_bits_offset_0;
  assign vrfReadDataPorts_2_bits_instructionIndex = vrfReadDataPorts_2_bits_instructionIndex_0;
  assign vrfReadDataPorts_3_valid = vrfReadDataPorts_3_valid_0;
  assign vrfReadDataPorts_3_bits_vs = vrfReadDataPorts_3_bits_vs_0;
  assign vrfReadDataPorts_3_bits_offset = vrfReadDataPorts_3_bits_offset_0;
  assign vrfReadDataPorts_3_bits_instructionIndex = vrfReadDataPorts_3_bits_instructionIndex_0;
endmodule

