
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module T1(
  input          indexedLoadStorePort_aw_ready,
  output         indexedLoadStorePort_aw_valid,
  output [1:0]   indexedLoadStorePort_aw_bits_id,
  output [31:0]  indexedLoadStorePort_aw_bits_addr,
  output [7:0]   indexedLoadStorePort_aw_bits_len,
  output [2:0]   indexedLoadStorePort_aw_bits_size,
  output [1:0]   indexedLoadStorePort_aw_bits_burst,
  output         indexedLoadStorePort_aw_bits_lock,
  output [3:0]   indexedLoadStorePort_aw_bits_cache,
  output [2:0]   indexedLoadStorePort_aw_bits_prot,
  output [3:0]   indexedLoadStorePort_aw_bits_qos,
                 indexedLoadStorePort_aw_bits_region,
  input          indexedLoadStorePort_w_ready,
  output         indexedLoadStorePort_w_valid,
  output [31:0]  indexedLoadStorePort_w_bits_data,
  output [3:0]   indexedLoadStorePort_w_bits_strb,
  output         indexedLoadStorePort_w_bits_last,
                 indexedLoadStorePort_b_ready,
  input          indexedLoadStorePort_b_valid,
  input  [1:0]   indexedLoadStorePort_b_bits_id,
                 indexedLoadStorePort_b_bits_resp,
  input          indexedLoadStorePort_ar_ready,
  output         indexedLoadStorePort_ar_valid,
  output [1:0]   indexedLoadStorePort_ar_bits_id,
  output [31:0]  indexedLoadStorePort_ar_bits_addr,
  output [7:0]   indexedLoadStorePort_ar_bits_len,
  output [2:0]   indexedLoadStorePort_ar_bits_size,
  output [1:0]   indexedLoadStorePort_ar_bits_burst,
  output         indexedLoadStorePort_ar_bits_lock,
  output [3:0]   indexedLoadStorePort_ar_bits_cache,
  output [2:0]   indexedLoadStorePort_ar_bits_prot,
  output [3:0]   indexedLoadStorePort_ar_bits_qos,
                 indexedLoadStorePort_ar_bits_region,
  output         indexedLoadStorePort_r_ready,
  input          indexedLoadStorePort_r_valid,
  input  [1:0]   indexedLoadStorePort_r_bits_id,
  input  [31:0]  indexedLoadStorePort_r_bits_data,
  input  [1:0]   indexedLoadStorePort_r_bits_resp,
  input          indexedLoadStorePort_r_bits_last,
                 highBandwidthLoadStorePort_aw_ready,
  output         highBandwidthLoadStorePort_aw_valid,
  output [1:0]   highBandwidthLoadStorePort_aw_bits_id,
  output [31:0]  highBandwidthLoadStorePort_aw_bits_addr,
  output [7:0]   highBandwidthLoadStorePort_aw_bits_len,
  output [2:0]   highBandwidthLoadStorePort_aw_bits_size,
  output [1:0]   highBandwidthLoadStorePort_aw_bits_burst,
  output         highBandwidthLoadStorePort_aw_bits_lock,
  output [3:0]   highBandwidthLoadStorePort_aw_bits_cache,
  output [2:0]   highBandwidthLoadStorePort_aw_bits_prot,
  output [3:0]   highBandwidthLoadStorePort_aw_bits_qos,
                 highBandwidthLoadStorePort_aw_bits_region,
  input          highBandwidthLoadStorePort_w_ready,
  output         highBandwidthLoadStorePort_w_valid,
  output [255:0] highBandwidthLoadStorePort_w_bits_data,
  output [31:0]  highBandwidthLoadStorePort_w_bits_strb,
  output         highBandwidthLoadStorePort_w_bits_last,
                 highBandwidthLoadStorePort_b_ready,
  input          highBandwidthLoadStorePort_b_valid,
  input  [1:0]   highBandwidthLoadStorePort_b_bits_id,
                 highBandwidthLoadStorePort_b_bits_resp,
  input          highBandwidthLoadStorePort_ar_ready,
  output         highBandwidthLoadStorePort_ar_valid,
  output [1:0]   highBandwidthLoadStorePort_ar_bits_id,
  output [31:0]  highBandwidthLoadStorePort_ar_bits_addr,
  output [7:0]   highBandwidthLoadStorePort_ar_bits_len,
  output [2:0]   highBandwidthLoadStorePort_ar_bits_size,
  output [1:0]   highBandwidthLoadStorePort_ar_bits_burst,
  output         highBandwidthLoadStorePort_ar_bits_lock,
  output [3:0]   highBandwidthLoadStorePort_ar_bits_cache,
  output [2:0]   highBandwidthLoadStorePort_ar_bits_prot,
  output [3:0]   highBandwidthLoadStorePort_ar_bits_qos,
                 highBandwidthLoadStorePort_ar_bits_region,
  output         highBandwidthLoadStorePort_r_ready,
  input          highBandwidthLoadStorePort_r_valid,
  input  [1:0]   highBandwidthLoadStorePort_r_bits_id,
  input  [255:0] highBandwidthLoadStorePort_r_bits_data,
  input  [1:0]   highBandwidthLoadStorePort_r_bits_resp,
  input          highBandwidthLoadStorePort_r_bits_last,
  output         retire_rd_valid,
  output [4:0]   retire_rd_bits_rdAddress,
  output [31:0]  retire_rd_bits_rdData,
  output         retire_rd_bits_isFp,
                 retire_csr_valid,
  output [31:0]  retire_csr_bits_vxsat,
                 retire_csr_bits_fflag,
  output         retire_mem_valid,
                 issue_ready,
  input          issue_valid,
  input  [31:0]  issue_bits_instruction,
                 issue_bits_rs1Data,
                 issue_bits_rs2Data,
                 issue_bits_vtype,
                 issue_bits_vl,
                 issue_bits_vstart,
                 issue_bits_vcsr,
  input          reset,
                 clock
);

  wire         _sinkVec_queue_fifo_31_empty;
  wire         _sinkVec_queue_fifo_31_full;
  wire         _sinkVec_queue_fifo_31_error;
  wire [47:0]  _sinkVec_queue_fifo_31_data_out;
  wire         _sinkVec_queue_fifo_30_empty;
  wire         _sinkVec_queue_fifo_30_full;
  wire         _sinkVec_queue_fifo_30_error;
  wire [47:0]  _sinkVec_queue_fifo_30_data_out;
  wire         _sinkVec_queue_fifo_29_empty;
  wire         _sinkVec_queue_fifo_29_full;
  wire         _sinkVec_queue_fifo_29_error;
  wire [12:0]  _sinkVec_queue_fifo_29_data_out;
  wire         _sinkVec_queue_fifo_28_empty;
  wire         _sinkVec_queue_fifo_28_full;
  wire         _sinkVec_queue_fifo_28_error;
  wire [12:0]  _sinkVec_queue_fifo_28_data_out;
  wire         _laneVec_7_readBusPort_0_enqRelease;
  wire         _laneVec_7_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_7_readBusPort_0_deq_bits_data;
  wire         _laneVec_7_readBusPort_1_enqRelease;
  wire         _laneVec_7_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_7_readBusPort_1_deq_bits_data;
  wire         _laneVec_7_writeBusPort_0_enqRelease;
  wire         _laneVec_7_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_7_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_7_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_7_writeBusPort_0_deq_bits_instructionIndex;
  wire [6:0]   _laneVec_7_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_7_writeBusPort_1_enqRelease;
  wire         _laneVec_7_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_7_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_7_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_7_writeBusPort_1_deq_bits_instructionIndex;
  wire [6:0]   _laneVec_7_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_7_laneRequest_ready;
  wire         _laneVec_7_maskUnitRequest_valid;
  wire [31:0]  _laneVec_7_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_7_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_7_maskUnitRequest_bits_index;
  wire         _laneVec_7_maskUnitRequest_bits_ffo;
  wire         _laneVec_7_maskRequestToLSU;
  wire [31:0]  _laneVec_7_vrfReadDataChannel;
  wire [7:0]   _laneVec_7_instructionFinished;
  wire [7:0]   _laneVec_7_vxsatReport;
  wire         _laneVec_7_v0Update_valid;
  wire [31:0]  _laneVec_7_v0Update_bits_data;
  wire [2:0]   _laneVec_7_v0Update_bits_offset;
  wire [3:0]   _laneVec_7_v0Update_bits_mask;
  wire [5:0]   _laneVec_7_maskSelect;
  wire [1:0]   _laneVec_7_maskSelectSew;
  wire         _sinkVec_queue_fifo_27_empty;
  wire         _sinkVec_queue_fifo_27_full;
  wire         _sinkVec_queue_fifo_27_error;
  wire [47:0]  _sinkVec_queue_fifo_27_data_out;
  wire         _sinkVec_queue_fifo_26_empty;
  wire         _sinkVec_queue_fifo_26_full;
  wire         _sinkVec_queue_fifo_26_error;
  wire [47:0]  _sinkVec_queue_fifo_26_data_out;
  wire         _sinkVec_queue_fifo_25_empty;
  wire         _sinkVec_queue_fifo_25_full;
  wire         _sinkVec_queue_fifo_25_error;
  wire [12:0]  _sinkVec_queue_fifo_25_data_out;
  wire         _sinkVec_queue_fifo_24_empty;
  wire         _sinkVec_queue_fifo_24_full;
  wire         _sinkVec_queue_fifo_24_error;
  wire [12:0]  _sinkVec_queue_fifo_24_data_out;
  wire         _laneVec_6_readBusPort_0_enqRelease;
  wire         _laneVec_6_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_6_readBusPort_0_deq_bits_data;
  wire         _laneVec_6_readBusPort_1_enqRelease;
  wire         _laneVec_6_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_6_readBusPort_1_deq_bits_data;
  wire         _laneVec_6_writeBusPort_0_enqRelease;
  wire         _laneVec_6_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_6_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_6_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_6_writeBusPort_0_deq_bits_instructionIndex;
  wire [6:0]   _laneVec_6_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_6_writeBusPort_1_enqRelease;
  wire         _laneVec_6_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_6_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_6_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_6_writeBusPort_1_deq_bits_instructionIndex;
  wire [6:0]   _laneVec_6_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_6_laneRequest_ready;
  wire         _laneVec_6_maskUnitRequest_valid;
  wire [31:0]  _laneVec_6_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_6_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_6_maskUnitRequest_bits_index;
  wire         _laneVec_6_maskUnitRequest_bits_ffo;
  wire         _laneVec_6_maskRequestToLSU;
  wire [31:0]  _laneVec_6_vrfReadDataChannel;
  wire [7:0]   _laneVec_6_instructionFinished;
  wire [7:0]   _laneVec_6_vxsatReport;
  wire         _laneVec_6_v0Update_valid;
  wire [31:0]  _laneVec_6_v0Update_bits_data;
  wire [2:0]   _laneVec_6_v0Update_bits_offset;
  wire [3:0]   _laneVec_6_v0Update_bits_mask;
  wire [5:0]   _laneVec_6_maskSelect;
  wire [1:0]   _laneVec_6_maskSelectSew;
  wire         _sinkVec_queue_fifo_23_empty;
  wire         _sinkVec_queue_fifo_23_full;
  wire         _sinkVec_queue_fifo_23_error;
  wire [47:0]  _sinkVec_queue_fifo_23_data_out;
  wire         _sinkVec_queue_fifo_22_empty;
  wire         _sinkVec_queue_fifo_22_full;
  wire         _sinkVec_queue_fifo_22_error;
  wire [47:0]  _sinkVec_queue_fifo_22_data_out;
  wire         _sinkVec_queue_fifo_21_empty;
  wire         _sinkVec_queue_fifo_21_full;
  wire         _sinkVec_queue_fifo_21_error;
  wire [12:0]  _sinkVec_queue_fifo_21_data_out;
  wire         _sinkVec_queue_fifo_20_empty;
  wire         _sinkVec_queue_fifo_20_full;
  wire         _sinkVec_queue_fifo_20_error;
  wire [12:0]  _sinkVec_queue_fifo_20_data_out;
  wire         _laneVec_5_readBusPort_0_enqRelease;
  wire         _laneVec_5_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_5_readBusPort_0_deq_bits_data;
  wire         _laneVec_5_readBusPort_1_enqRelease;
  wire         _laneVec_5_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_5_readBusPort_1_deq_bits_data;
  wire         _laneVec_5_writeBusPort_0_enqRelease;
  wire         _laneVec_5_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_5_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_5_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_5_writeBusPort_0_deq_bits_instructionIndex;
  wire [6:0]   _laneVec_5_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_5_writeBusPort_1_enqRelease;
  wire         _laneVec_5_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_5_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_5_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_5_writeBusPort_1_deq_bits_instructionIndex;
  wire [6:0]   _laneVec_5_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_5_laneRequest_ready;
  wire         _laneVec_5_maskUnitRequest_valid;
  wire [31:0]  _laneVec_5_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_5_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_5_maskUnitRequest_bits_index;
  wire         _laneVec_5_maskUnitRequest_bits_ffo;
  wire         _laneVec_5_maskRequestToLSU;
  wire [31:0]  _laneVec_5_vrfReadDataChannel;
  wire [7:0]   _laneVec_5_instructionFinished;
  wire [7:0]   _laneVec_5_vxsatReport;
  wire         _laneVec_5_v0Update_valid;
  wire [31:0]  _laneVec_5_v0Update_bits_data;
  wire [2:0]   _laneVec_5_v0Update_bits_offset;
  wire [3:0]   _laneVec_5_v0Update_bits_mask;
  wire [5:0]   _laneVec_5_maskSelect;
  wire [1:0]   _laneVec_5_maskSelectSew;
  wire         _sinkVec_queue_fifo_19_empty;
  wire         _sinkVec_queue_fifo_19_full;
  wire         _sinkVec_queue_fifo_19_error;
  wire [47:0]  _sinkVec_queue_fifo_19_data_out;
  wire         _sinkVec_queue_fifo_18_empty;
  wire         _sinkVec_queue_fifo_18_full;
  wire         _sinkVec_queue_fifo_18_error;
  wire [47:0]  _sinkVec_queue_fifo_18_data_out;
  wire         _sinkVec_queue_fifo_17_empty;
  wire         _sinkVec_queue_fifo_17_full;
  wire         _sinkVec_queue_fifo_17_error;
  wire [12:0]  _sinkVec_queue_fifo_17_data_out;
  wire         _sinkVec_queue_fifo_16_empty;
  wire         _sinkVec_queue_fifo_16_full;
  wire         _sinkVec_queue_fifo_16_error;
  wire [12:0]  _sinkVec_queue_fifo_16_data_out;
  wire         _laneVec_4_readBusPort_0_enqRelease;
  wire         _laneVec_4_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_4_readBusPort_0_deq_bits_data;
  wire         _laneVec_4_readBusPort_1_enqRelease;
  wire         _laneVec_4_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_4_readBusPort_1_deq_bits_data;
  wire         _laneVec_4_writeBusPort_0_enqRelease;
  wire         _laneVec_4_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_4_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_4_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_4_writeBusPort_0_deq_bits_instructionIndex;
  wire [6:0]   _laneVec_4_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_4_writeBusPort_1_enqRelease;
  wire         _laneVec_4_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_4_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_4_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_4_writeBusPort_1_deq_bits_instructionIndex;
  wire [6:0]   _laneVec_4_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_4_laneRequest_ready;
  wire         _laneVec_4_maskUnitRequest_valid;
  wire [31:0]  _laneVec_4_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_4_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_4_maskUnitRequest_bits_index;
  wire         _laneVec_4_maskUnitRequest_bits_ffo;
  wire         _laneVec_4_maskRequestToLSU;
  wire [31:0]  _laneVec_4_vrfReadDataChannel;
  wire [7:0]   _laneVec_4_instructionFinished;
  wire [7:0]   _laneVec_4_vxsatReport;
  wire         _laneVec_4_v0Update_valid;
  wire [31:0]  _laneVec_4_v0Update_bits_data;
  wire [2:0]   _laneVec_4_v0Update_bits_offset;
  wire [3:0]   _laneVec_4_v0Update_bits_mask;
  wire [5:0]   _laneVec_4_maskSelect;
  wire [1:0]   _laneVec_4_maskSelectSew;
  wire         _sinkVec_queue_fifo_15_empty;
  wire         _sinkVec_queue_fifo_15_full;
  wire         _sinkVec_queue_fifo_15_error;
  wire [47:0]  _sinkVec_queue_fifo_15_data_out;
  wire         _sinkVec_queue_fifo_14_empty;
  wire         _sinkVec_queue_fifo_14_full;
  wire         _sinkVec_queue_fifo_14_error;
  wire [47:0]  _sinkVec_queue_fifo_14_data_out;
  wire         _sinkVec_queue_fifo_13_empty;
  wire         _sinkVec_queue_fifo_13_full;
  wire         _sinkVec_queue_fifo_13_error;
  wire [12:0]  _sinkVec_queue_fifo_13_data_out;
  wire         _sinkVec_queue_fifo_12_empty;
  wire         _sinkVec_queue_fifo_12_full;
  wire         _sinkVec_queue_fifo_12_error;
  wire [12:0]  _sinkVec_queue_fifo_12_data_out;
  wire         _laneVec_3_readBusPort_0_enqRelease;
  wire         _laneVec_3_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_3_readBusPort_0_deq_bits_data;
  wire         _laneVec_3_readBusPort_1_enqRelease;
  wire         _laneVec_3_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_3_readBusPort_1_deq_bits_data;
  wire         _laneVec_3_writeBusPort_0_enqRelease;
  wire         _laneVec_3_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_3_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_3_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_3_writeBusPort_0_deq_bits_instructionIndex;
  wire [6:0]   _laneVec_3_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_3_writeBusPort_1_enqRelease;
  wire         _laneVec_3_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_3_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_3_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_3_writeBusPort_1_deq_bits_instructionIndex;
  wire [6:0]   _laneVec_3_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_3_laneRequest_ready;
  wire         _laneVec_3_maskUnitRequest_valid;
  wire [31:0]  _laneVec_3_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_3_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_3_maskUnitRequest_bits_index;
  wire         _laneVec_3_maskUnitRequest_bits_ffo;
  wire         _laneVec_3_maskRequestToLSU;
  wire [31:0]  _laneVec_3_vrfReadDataChannel;
  wire [7:0]   _laneVec_3_instructionFinished;
  wire [7:0]   _laneVec_3_vxsatReport;
  wire         _laneVec_3_v0Update_valid;
  wire [31:0]  _laneVec_3_v0Update_bits_data;
  wire [2:0]   _laneVec_3_v0Update_bits_offset;
  wire [3:0]   _laneVec_3_v0Update_bits_mask;
  wire [5:0]   _laneVec_3_maskSelect;
  wire [1:0]   _laneVec_3_maskSelectSew;
  wire         _sinkVec_queue_fifo_11_empty;
  wire         _sinkVec_queue_fifo_11_full;
  wire         _sinkVec_queue_fifo_11_error;
  wire [47:0]  _sinkVec_queue_fifo_11_data_out;
  wire         _sinkVec_queue_fifo_10_empty;
  wire         _sinkVec_queue_fifo_10_full;
  wire         _sinkVec_queue_fifo_10_error;
  wire [47:0]  _sinkVec_queue_fifo_10_data_out;
  wire         _sinkVec_queue_fifo_9_empty;
  wire         _sinkVec_queue_fifo_9_full;
  wire         _sinkVec_queue_fifo_9_error;
  wire [12:0]  _sinkVec_queue_fifo_9_data_out;
  wire         _sinkVec_queue_fifo_8_empty;
  wire         _sinkVec_queue_fifo_8_full;
  wire         _sinkVec_queue_fifo_8_error;
  wire [12:0]  _sinkVec_queue_fifo_8_data_out;
  wire         _laneVec_2_readBusPort_0_enqRelease;
  wire         _laneVec_2_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_2_readBusPort_0_deq_bits_data;
  wire         _laneVec_2_readBusPort_1_enqRelease;
  wire         _laneVec_2_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_2_readBusPort_1_deq_bits_data;
  wire         _laneVec_2_writeBusPort_0_enqRelease;
  wire         _laneVec_2_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_2_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_2_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_2_writeBusPort_0_deq_bits_instructionIndex;
  wire [6:0]   _laneVec_2_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_2_writeBusPort_1_enqRelease;
  wire         _laneVec_2_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_2_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_2_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_2_writeBusPort_1_deq_bits_instructionIndex;
  wire [6:0]   _laneVec_2_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_2_laneRequest_ready;
  wire         _laneVec_2_maskUnitRequest_valid;
  wire [31:0]  _laneVec_2_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_2_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_2_maskUnitRequest_bits_index;
  wire         _laneVec_2_maskUnitRequest_bits_ffo;
  wire         _laneVec_2_maskRequestToLSU;
  wire [31:0]  _laneVec_2_vrfReadDataChannel;
  wire [7:0]   _laneVec_2_instructionFinished;
  wire [7:0]   _laneVec_2_vxsatReport;
  wire         _laneVec_2_v0Update_valid;
  wire [31:0]  _laneVec_2_v0Update_bits_data;
  wire [2:0]   _laneVec_2_v0Update_bits_offset;
  wire [3:0]   _laneVec_2_v0Update_bits_mask;
  wire [5:0]   _laneVec_2_maskSelect;
  wire [1:0]   _laneVec_2_maskSelectSew;
  wire         _sinkVec_queue_fifo_7_empty;
  wire         _sinkVec_queue_fifo_7_full;
  wire         _sinkVec_queue_fifo_7_error;
  wire [47:0]  _sinkVec_queue_fifo_7_data_out;
  wire         _sinkVec_queue_fifo_6_empty;
  wire         _sinkVec_queue_fifo_6_full;
  wire         _sinkVec_queue_fifo_6_error;
  wire [47:0]  _sinkVec_queue_fifo_6_data_out;
  wire         _sinkVec_queue_fifo_5_empty;
  wire         _sinkVec_queue_fifo_5_full;
  wire         _sinkVec_queue_fifo_5_error;
  wire [12:0]  _sinkVec_queue_fifo_5_data_out;
  wire         _sinkVec_queue_fifo_4_empty;
  wire         _sinkVec_queue_fifo_4_full;
  wire         _sinkVec_queue_fifo_4_error;
  wire [12:0]  _sinkVec_queue_fifo_4_data_out;
  wire         _laneVec_1_readBusPort_0_enqRelease;
  wire         _laneVec_1_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_1_readBusPort_0_deq_bits_data;
  wire         _laneVec_1_readBusPort_1_enqRelease;
  wire         _laneVec_1_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_1_readBusPort_1_deq_bits_data;
  wire         _laneVec_1_writeBusPort_0_enqRelease;
  wire         _laneVec_1_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_1_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_1_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_1_writeBusPort_0_deq_bits_instructionIndex;
  wire [6:0]   _laneVec_1_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_1_writeBusPort_1_enqRelease;
  wire         _laneVec_1_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_1_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_1_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_1_writeBusPort_1_deq_bits_instructionIndex;
  wire [6:0]   _laneVec_1_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_1_laneRequest_ready;
  wire         _laneVec_1_maskUnitRequest_valid;
  wire [31:0]  _laneVec_1_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_1_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_1_maskUnitRequest_bits_index;
  wire         _laneVec_1_maskUnitRequest_bits_ffo;
  wire         _laneVec_1_maskRequestToLSU;
  wire [31:0]  _laneVec_1_vrfReadDataChannel;
  wire [7:0]   _laneVec_1_instructionFinished;
  wire [7:0]   _laneVec_1_vxsatReport;
  wire         _laneVec_1_v0Update_valid;
  wire [31:0]  _laneVec_1_v0Update_bits_data;
  wire [2:0]   _laneVec_1_v0Update_bits_offset;
  wire [3:0]   _laneVec_1_v0Update_bits_mask;
  wire [5:0]   _laneVec_1_maskSelect;
  wire [1:0]   _laneVec_1_maskSelectSew;
  wire         _sinkVec_queue_fifo_3_empty;
  wire         _sinkVec_queue_fifo_3_full;
  wire         _sinkVec_queue_fifo_3_error;
  wire [47:0]  _sinkVec_queue_fifo_3_data_out;
  wire         _sinkVec_queue_fifo_2_empty;
  wire         _sinkVec_queue_fifo_2_full;
  wire         _sinkVec_queue_fifo_2_error;
  wire [47:0]  _sinkVec_queue_fifo_2_data_out;
  wire         _sinkVec_queue_fifo_1_empty;
  wire         _sinkVec_queue_fifo_1_full;
  wire         _sinkVec_queue_fifo_1_error;
  wire [12:0]  _sinkVec_queue_fifo_1_data_out;
  wire         _sinkVec_queue_fifo_empty;
  wire         _sinkVec_queue_fifo_full;
  wire         _sinkVec_queue_fifo_error;
  wire [12:0]  _sinkVec_queue_fifo_data_out;
  wire         _laneVec_0_readBusPort_0_enqRelease;
  wire         _laneVec_0_readBusPort_0_deq_valid;
  wire [31:0]  _laneVec_0_readBusPort_0_deq_bits_data;
  wire         _laneVec_0_readBusPort_1_enqRelease;
  wire         _laneVec_0_readBusPort_1_deq_valid;
  wire [31:0]  _laneVec_0_readBusPort_1_deq_bits_data;
  wire         _laneVec_0_writeBusPort_0_enqRelease;
  wire         _laneVec_0_writeBusPort_0_deq_valid;
  wire [31:0]  _laneVec_0_writeBusPort_0_deq_bits_data;
  wire [1:0]   _laneVec_0_writeBusPort_0_deq_bits_mask;
  wire [2:0]   _laneVec_0_writeBusPort_0_deq_bits_instructionIndex;
  wire [6:0]   _laneVec_0_writeBusPort_0_deq_bits_counter;
  wire         _laneVec_0_writeBusPort_1_enqRelease;
  wire         _laneVec_0_writeBusPort_1_deq_valid;
  wire [31:0]  _laneVec_0_writeBusPort_1_deq_bits_data;
  wire [1:0]   _laneVec_0_writeBusPort_1_deq_bits_mask;
  wire [2:0]   _laneVec_0_writeBusPort_1_deq_bits_instructionIndex;
  wire [6:0]   _laneVec_0_writeBusPort_1_deq_bits_counter;
  wire         _laneVec_0_laneRequest_ready;
  wire         _laneVec_0_maskUnitRequest_valid;
  wire [31:0]  _laneVec_0_maskUnitRequest_bits_source1;
  wire [31:0]  _laneVec_0_maskUnitRequest_bits_source2;
  wire [2:0]   _laneVec_0_maskUnitRequest_bits_index;
  wire         _laneVec_0_maskUnitRequest_bits_ffo;
  wire         _laneVec_0_maskRequestToLSU;
  wire [31:0]  _laneVec_0_vrfReadDataChannel;
  wire [7:0]   _laneVec_0_instructionFinished;
  wire [7:0]   _laneVec_0_vxsatReport;
  wire         _laneVec_0_v0Update_valid;
  wire [31:0]  _laneVec_0_v0Update_bits_data;
  wire [2:0]   _laneVec_0_v0Update_bits_offset;
  wire [3:0]   _laneVec_0_v0Update_bits_mask;
  wire [5:0]   _laneVec_0_maskSelect;
  wire [1:0]   _laneVec_0_maskSelectSew;
  wire         _queue_fifo_7_empty;
  wire         _queue_fifo_7_full;
  wire         _queue_fifo_7_error;
  wire [144:0] _queue_fifo_7_data_out;
  wire         _queue_fifo_6_empty;
  wire         _queue_fifo_6_full;
  wire         _queue_fifo_6_error;
  wire [144:0] _queue_fifo_6_data_out;
  wire         _queue_fifo_5_empty;
  wire         _queue_fifo_5_full;
  wire         _queue_fifo_5_error;
  wire [144:0] _queue_fifo_5_data_out;
  wire         _queue_fifo_4_empty;
  wire         _queue_fifo_4_full;
  wire         _queue_fifo_4_error;
  wire [144:0] _queue_fifo_4_data_out;
  wire         _queue_fifo_3_empty;
  wire         _queue_fifo_3_full;
  wire         _queue_fifo_3_error;
  wire [144:0] _queue_fifo_3_data_out;
  wire         _queue_fifo_2_empty;
  wire         _queue_fifo_2_full;
  wire         _queue_fifo_2_error;
  wire [144:0] _queue_fifo_2_data_out;
  wire         _queue_fifo_1_empty;
  wire         _queue_fifo_1_full;
  wire         _queue_fifo_1_error;
  wire [144:0] _queue_fifo_1_data_out;
  wire         _queue_fifo_empty;
  wire         _queue_fifo_full;
  wire         _queue_fifo_error;
  wire [144:0] _queue_fifo_data_out;
  wire         _tokenManager_issueAllow;
  wire [7:0]   _tokenManager_v0WriteValid;
  wire         _maskUnit_exeResp_0_valid;
  wire [3:0]   _maskUnit_exeResp_0_bits_mask;
  wire [2:0]   _maskUnit_exeResp_0_bits_instructionIndex;
  wire         _maskUnit_exeResp_1_valid;
  wire [3:0]   _maskUnit_exeResp_1_bits_mask;
  wire [2:0]   _maskUnit_exeResp_1_bits_instructionIndex;
  wire         _maskUnit_exeResp_2_valid;
  wire [3:0]   _maskUnit_exeResp_2_bits_mask;
  wire [2:0]   _maskUnit_exeResp_2_bits_instructionIndex;
  wire         _maskUnit_exeResp_3_valid;
  wire [3:0]   _maskUnit_exeResp_3_bits_mask;
  wire [2:0]   _maskUnit_exeResp_3_bits_instructionIndex;
  wire         _maskUnit_exeResp_4_valid;
  wire [3:0]   _maskUnit_exeResp_4_bits_mask;
  wire [2:0]   _maskUnit_exeResp_4_bits_instructionIndex;
  wire         _maskUnit_exeResp_5_valid;
  wire [3:0]   _maskUnit_exeResp_5_bits_mask;
  wire [2:0]   _maskUnit_exeResp_5_bits_instructionIndex;
  wire         _maskUnit_exeResp_6_valid;
  wire [3:0]   _maskUnit_exeResp_6_bits_mask;
  wire [2:0]   _maskUnit_exeResp_6_bits_instructionIndex;
  wire         _maskUnit_exeResp_7_valid;
  wire [3:0]   _maskUnit_exeResp_7_bits_mask;
  wire [2:0]   _maskUnit_exeResp_7_bits_instructionIndex;
  wire         _maskUnit_tokenIO_0_maskRequestRelease;
  wire         _maskUnit_tokenIO_1_maskRequestRelease;
  wire         _maskUnit_tokenIO_2_maskRequestRelease;
  wire         _maskUnit_tokenIO_3_maskRequestRelease;
  wire         _maskUnit_tokenIO_4_maskRequestRelease;
  wire         _maskUnit_tokenIO_5_maskRequestRelease;
  wire         _maskUnit_tokenIO_6_maskRequestRelease;
  wire         _maskUnit_tokenIO_7_maskRequestRelease;
  wire [7:0]   _maskUnit_lastReport;
  wire [31:0]  _maskUnit_laneMaskInput_0;
  wire [31:0]  _maskUnit_laneMaskInput_1;
  wire [31:0]  _maskUnit_laneMaskInput_2;
  wire [31:0]  _maskUnit_laneMaskInput_3;
  wire [31:0]  _maskUnit_laneMaskInput_4;
  wire [31:0]  _maskUnit_laneMaskInput_5;
  wire [31:0]  _maskUnit_laneMaskInput_6;
  wire [31:0]  _maskUnit_laneMaskInput_7;
  wire         _maskUnit_gatherData_valid;
  wire [31:0]  _maskUnit_gatherData_bits;
  wire         _decode_decodeResult_specialSlot;
  wire [4:0]   _decode_decodeResult_topUop;
  wire         _decode_decodeResult_popCount;
  wire         _decode_decodeResult_ffo;
  wire         _decode_decodeResult_average;
  wire         _decode_decodeResult_reverse;
  wire         _decode_decodeResult_dontNeedExecuteInLane;
  wire         _decode_decodeResult_scheduler;
  wire         _decode_decodeResult_sReadVD;
  wire         _decode_decodeResult_vtype;
  wire         _decode_decodeResult_sWrite;
  wire         _decode_decodeResult_crossRead;
  wire         _decode_decodeResult_crossWrite;
  wire         _decode_decodeResult_maskUnit;
  wire         _decode_decodeResult_special;
  wire         _decode_decodeResult_saturate;
  wire         _decode_decodeResult_vwmacc;
  wire         _decode_decodeResult_readOnly;
  wire         _decode_decodeResult_maskSource;
  wire         _decode_decodeResult_maskDestination;
  wire         _decode_decodeResult_maskLogic;
  wire [3:0]   _decode_decodeResult_uop;
  wire         _decode_decodeResult_iota;
  wire         _decode_decodeResult_mv;
  wire         _decode_decodeResult_extend;
  wire         _decode_decodeResult_unOrderWrite;
  wire         _decode_decodeResult_compress;
  wire         _decode_decodeResult_gather16;
  wire         _decode_decodeResult_gather;
  wire         _decode_decodeResult_slid;
  wire         _decode_decodeResult_targetRd;
  wire         _decode_decodeResult_widenReduce;
  wire         _decode_decodeResult_red;
  wire         _decode_decodeResult_nr;
  wire         _decode_decodeResult_itype;
  wire         _decode_decodeResult_unsigned1;
  wire         _decode_decodeResult_unsigned0;
  wire         _decode_decodeResult_other;
  wire         _decode_decodeResult_multiCycle;
  wire         _decode_decodeResult_divider;
  wire         _decode_decodeResult_multiplier;
  wire         _decode_decodeResult_shift;
  wire         _decode_decodeResult_adder;
  wire         _decode_decodeResult_logic;
  wire         _lsu_request_ready;
  wire         _lsu_vrfWritePort_0_valid;
  wire [4:0]   _lsu_vrfWritePort_0_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_0_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_0_bits_instructionIndex;
  wire         _lsu_vrfWritePort_1_valid;
  wire [4:0]   _lsu_vrfWritePort_1_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_1_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_1_bits_instructionIndex;
  wire         _lsu_vrfWritePort_2_valid;
  wire [4:0]   _lsu_vrfWritePort_2_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_2_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_2_bits_instructionIndex;
  wire         _lsu_vrfWritePort_3_valid;
  wire [4:0]   _lsu_vrfWritePort_3_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_3_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_3_bits_instructionIndex;
  wire         _lsu_vrfWritePort_4_valid;
  wire [4:0]   _lsu_vrfWritePort_4_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_4_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_4_bits_instructionIndex;
  wire         _lsu_vrfWritePort_5_valid;
  wire [4:0]   _lsu_vrfWritePort_5_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_5_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_5_bits_instructionIndex;
  wire         _lsu_vrfWritePort_6_valid;
  wire [4:0]   _lsu_vrfWritePort_6_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_6_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_6_bits_instructionIndex;
  wire         _lsu_vrfWritePort_7_valid;
  wire [4:0]   _lsu_vrfWritePort_7_bits_vd;
  wire [3:0]   _lsu_vrfWritePort_7_bits_mask;
  wire [2:0]   _lsu_vrfWritePort_7_bits_instructionIndex;
  wire [7:0]   _lsu_dataInWriteQueue_0;
  wire [7:0]   _lsu_dataInWriteQueue_1;
  wire [7:0]   _lsu_dataInWriteQueue_2;
  wire [7:0]   _lsu_dataInWriteQueue_3;
  wire [7:0]   _lsu_dataInWriteQueue_4;
  wire [7:0]   _lsu_dataInWriteQueue_5;
  wire [7:0]   _lsu_dataInWriteQueue_6;
  wire [7:0]   _lsu_dataInWriteQueue_7;
  wire [7:0]   _lsu_lastReport;
  wire [7:0]   _lsu_tokenIO_offsetGroupRelease;
  wire         sinkVec_queue_31_almostFull;
  wire         sinkVec_queue_31_almostEmpty;
  wire         sinkVec_queue_30_almostFull;
  wire         sinkVec_queue_30_almostEmpty;
  wire         sinkVec_queue_29_almostFull;
  wire         sinkVec_queue_29_almostEmpty;
  wire         sinkVec_queue_28_almostFull;
  wire         sinkVec_queue_28_almostEmpty;
  wire         sinkVec_queue_27_almostFull;
  wire         sinkVec_queue_27_almostEmpty;
  wire         sinkVec_queue_26_almostFull;
  wire         sinkVec_queue_26_almostEmpty;
  wire         sinkVec_queue_25_almostFull;
  wire         sinkVec_queue_25_almostEmpty;
  wire         sinkVec_queue_24_almostFull;
  wire         sinkVec_queue_24_almostEmpty;
  wire         sinkVec_queue_23_almostFull;
  wire         sinkVec_queue_23_almostEmpty;
  wire         sinkVec_queue_22_almostFull;
  wire         sinkVec_queue_22_almostEmpty;
  wire         sinkVec_queue_21_almostFull;
  wire         sinkVec_queue_21_almostEmpty;
  wire         sinkVec_queue_20_almostFull;
  wire         sinkVec_queue_20_almostEmpty;
  wire         sinkVec_queue_19_almostFull;
  wire         sinkVec_queue_19_almostEmpty;
  wire         sinkVec_queue_18_almostFull;
  wire         sinkVec_queue_18_almostEmpty;
  wire         sinkVec_queue_17_almostFull;
  wire         sinkVec_queue_17_almostEmpty;
  wire         sinkVec_queue_16_almostFull;
  wire         sinkVec_queue_16_almostEmpty;
  wire         sinkVec_queue_15_almostFull;
  wire         sinkVec_queue_15_almostEmpty;
  wire         sinkVec_queue_14_almostFull;
  wire         sinkVec_queue_14_almostEmpty;
  wire         sinkVec_queue_13_almostFull;
  wire         sinkVec_queue_13_almostEmpty;
  wire         sinkVec_queue_12_almostFull;
  wire         sinkVec_queue_12_almostEmpty;
  wire         sinkVec_queue_11_almostFull;
  wire         sinkVec_queue_11_almostEmpty;
  wire         sinkVec_queue_10_almostFull;
  wire         sinkVec_queue_10_almostEmpty;
  wire         sinkVec_queue_9_almostFull;
  wire         sinkVec_queue_9_almostEmpty;
  wire         sinkVec_queue_8_almostFull;
  wire         sinkVec_queue_8_almostEmpty;
  wire         sinkVec_queue_7_almostFull;
  wire         sinkVec_queue_7_almostEmpty;
  wire         sinkVec_queue_6_almostFull;
  wire         sinkVec_queue_6_almostEmpty;
  wire         sinkVec_queue_5_almostFull;
  wire         sinkVec_queue_5_almostEmpty;
  wire         sinkVec_queue_4_almostFull;
  wire         sinkVec_queue_4_almostEmpty;
  wire         sinkVec_queue_3_almostFull;
  wire         sinkVec_queue_3_almostEmpty;
  wire         sinkVec_queue_2_almostFull;
  wire         sinkVec_queue_2_almostEmpty;
  wire         sinkVec_queue_1_almostFull;
  wire         sinkVec_queue_1_almostEmpty;
  wire         sinkVec_queue_almostFull;
  wire         sinkVec_queue_almostEmpty;
  wire         queue_7_almostFull;
  wire         queue_7_almostEmpty;
  wire         queue_6_almostFull;
  wire         queue_6_almostEmpty;
  wire         queue_5_almostFull;
  wire         queue_5_almostEmpty;
  wire         queue_4_almostFull;
  wire         queue_4_almostEmpty;
  wire         queue_3_almostFull;
  wire         queue_3_almostEmpty;
  wire         queue_2_almostFull;
  wire         queue_2_almostEmpty;
  wire         queue_1_almostFull;
  wire         queue_1_almostEmpty;
  wire         queue_almostFull;
  wire         queue_almostEmpty;
  wire [31:0]  retire_rd_bits_rdData_0;
  wire         highBandwidthLoadStorePort_r_ready_0;
  wire [31:0]  highBandwidthLoadStorePort_ar_bits_addr_0;
  wire         highBandwidthLoadStorePort_ar_valid_0;
  wire [31:0]  highBandwidthLoadStorePort_w_bits_strb_0;
  wire [255:0] highBandwidthLoadStorePort_w_bits_data_0;
  wire         highBandwidthLoadStorePort_w_valid_0;
  wire [31:0]  highBandwidthLoadStorePort_aw_bits_addr_0;
  wire [1:0]   highBandwidthLoadStorePort_aw_bits_id_0;
  wire         highBandwidthLoadStorePort_aw_valid_0;
  wire         indexedLoadStorePort_r_ready_0;
  wire [31:0]  indexedLoadStorePort_ar_bits_addr_0;
  wire         indexedLoadStorePort_ar_valid_0;
  wire [3:0]   indexedLoadStorePort_w_bits_strb_0;
  wire [31:0]  indexedLoadStorePort_w_bits_data_0;
  wire         indexedLoadStorePort_w_valid_0;
  wire [2:0]   indexedLoadStorePort_aw_bits_size_0;
  wire [31:0]  indexedLoadStorePort_aw_bits_addr_0;
  wire [1:0]   indexedLoadStorePort_aw_bits_id_0;
  wire         indexedLoadStorePort_aw_valid_0;
  wire [2:0]   x22_7_1_bits_instructionIndex;
  wire         x22_7_1_bits_last;
  wire [31:0]  x22_7_1_bits_data;
  wire [3:0]   x22_7_1_bits_mask;
  wire [2:0]   x22_7_1_bits_offset;
  wire [4:0]   x22_7_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_31_bits_instructionIndex;
  wire         sinkVec_sinkWire_31_bits_last;
  wire [31:0]  sinkVec_sinkWire_31_bits_data;
  wire [3:0]   sinkVec_sinkWire_31_bits_mask;
  wire [2:0]   sinkVec_sinkWire_31_bits_offset;
  wire [4:0]   sinkVec_sinkWire_31_bits_vd;
  wire         sinkVec_sinkWire_31_valid;
  wire         sinkVec_sinkWire_31_ready;
  wire [2:0]   x22_7_0_bits_instructionIndex;
  wire [31:0]  x22_7_0_bits_data;
  wire [3:0]   x22_7_0_bits_mask;
  wire [2:0]   x22_7_0_bits_offset;
  wire [4:0]   x22_7_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_30_bits_instructionIndex;
  wire         sinkVec_sinkWire_30_bits_last;
  wire [31:0]  sinkVec_sinkWire_30_bits_data;
  wire [3:0]   sinkVec_sinkWire_30_bits_mask;
  wire [2:0]   sinkVec_sinkWire_30_bits_offset;
  wire [4:0]   sinkVec_sinkWire_30_bits_vd;
  wire         sinkVec_sinkWire_30_valid;
  wire         sinkVec_sinkWire_30_ready;
  wire [2:0]   x13_7_1_bits_instructionIndex;
  wire [2:0]   x13_7_1_bits_offset;
  wire [4:0]   x13_7_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_29_bits_instructionIndex;
  wire [2:0]   sinkVec_sinkWire_29_bits_offset;
  wire [1:0]   sinkVec_sinkWire_29_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_29_bits_vs;
  wire         sinkVec_sinkWire_29_valid;
  wire         sinkVec_sinkWire_29_ready;
  wire [2:0]   x13_7_0_bits_instructionIndex;
  wire [2:0]   x13_7_0_bits_offset;
  wire [4:0]   x13_7_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_28_bits_instructionIndex;
  wire [2:0]   sinkVec_sinkWire_28_bits_offset;
  wire [1:0]   sinkVec_sinkWire_28_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_28_bits_vs;
  wire         sinkVec_sinkWire_28_valid;
  wire         sinkVec_sinkWire_28_ready;
  wire [2:0]   x22_6_1_bits_instructionIndex;
  wire         x22_6_1_bits_last;
  wire [31:0]  x22_6_1_bits_data;
  wire [3:0]   x22_6_1_bits_mask;
  wire [2:0]   x22_6_1_bits_offset;
  wire [4:0]   x22_6_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_27_bits_instructionIndex;
  wire         sinkVec_sinkWire_27_bits_last;
  wire [31:0]  sinkVec_sinkWire_27_bits_data;
  wire [3:0]   sinkVec_sinkWire_27_bits_mask;
  wire [2:0]   sinkVec_sinkWire_27_bits_offset;
  wire [4:0]   sinkVec_sinkWire_27_bits_vd;
  wire         sinkVec_sinkWire_27_valid;
  wire         sinkVec_sinkWire_27_ready;
  wire [2:0]   x22_6_0_bits_instructionIndex;
  wire [31:0]  x22_6_0_bits_data;
  wire [3:0]   x22_6_0_bits_mask;
  wire [2:0]   x22_6_0_bits_offset;
  wire [4:0]   x22_6_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_26_bits_instructionIndex;
  wire         sinkVec_sinkWire_26_bits_last;
  wire [31:0]  sinkVec_sinkWire_26_bits_data;
  wire [3:0]   sinkVec_sinkWire_26_bits_mask;
  wire [2:0]   sinkVec_sinkWire_26_bits_offset;
  wire [4:0]   sinkVec_sinkWire_26_bits_vd;
  wire         sinkVec_sinkWire_26_valid;
  wire         sinkVec_sinkWire_26_ready;
  wire [2:0]   x13_6_1_bits_instructionIndex;
  wire [2:0]   x13_6_1_bits_offset;
  wire [4:0]   x13_6_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_25_bits_instructionIndex;
  wire [2:0]   sinkVec_sinkWire_25_bits_offset;
  wire [1:0]   sinkVec_sinkWire_25_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_25_bits_vs;
  wire         sinkVec_sinkWire_25_valid;
  wire         sinkVec_sinkWire_25_ready;
  wire [2:0]   x13_6_0_bits_instructionIndex;
  wire [2:0]   x13_6_0_bits_offset;
  wire [4:0]   x13_6_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_24_bits_instructionIndex;
  wire [2:0]   sinkVec_sinkWire_24_bits_offset;
  wire [1:0]   sinkVec_sinkWire_24_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_24_bits_vs;
  wire         sinkVec_sinkWire_24_valid;
  wire         sinkVec_sinkWire_24_ready;
  wire [2:0]   x22_5_1_bits_instructionIndex;
  wire         x22_5_1_bits_last;
  wire [31:0]  x22_5_1_bits_data;
  wire [3:0]   x22_5_1_bits_mask;
  wire [2:0]   x22_5_1_bits_offset;
  wire [4:0]   x22_5_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_23_bits_instructionIndex;
  wire         sinkVec_sinkWire_23_bits_last;
  wire [31:0]  sinkVec_sinkWire_23_bits_data;
  wire [3:0]   sinkVec_sinkWire_23_bits_mask;
  wire [2:0]   sinkVec_sinkWire_23_bits_offset;
  wire [4:0]   sinkVec_sinkWire_23_bits_vd;
  wire         sinkVec_sinkWire_23_valid;
  wire         sinkVec_sinkWire_23_ready;
  wire [2:0]   x22_5_0_bits_instructionIndex;
  wire [31:0]  x22_5_0_bits_data;
  wire [3:0]   x22_5_0_bits_mask;
  wire [2:0]   x22_5_0_bits_offset;
  wire [4:0]   x22_5_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_22_bits_instructionIndex;
  wire         sinkVec_sinkWire_22_bits_last;
  wire [31:0]  sinkVec_sinkWire_22_bits_data;
  wire [3:0]   sinkVec_sinkWire_22_bits_mask;
  wire [2:0]   sinkVec_sinkWire_22_bits_offset;
  wire [4:0]   sinkVec_sinkWire_22_bits_vd;
  wire         sinkVec_sinkWire_22_valid;
  wire         sinkVec_sinkWire_22_ready;
  wire [2:0]   x13_5_1_bits_instructionIndex;
  wire [2:0]   x13_5_1_bits_offset;
  wire [4:0]   x13_5_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_21_bits_instructionIndex;
  wire [2:0]   sinkVec_sinkWire_21_bits_offset;
  wire [1:0]   sinkVec_sinkWire_21_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_21_bits_vs;
  wire         sinkVec_sinkWire_21_valid;
  wire         sinkVec_sinkWire_21_ready;
  wire [2:0]   x13_5_0_bits_instructionIndex;
  wire [2:0]   x13_5_0_bits_offset;
  wire [4:0]   x13_5_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_20_bits_instructionIndex;
  wire [2:0]   sinkVec_sinkWire_20_bits_offset;
  wire [1:0]   sinkVec_sinkWire_20_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_20_bits_vs;
  wire         sinkVec_sinkWire_20_valid;
  wire         sinkVec_sinkWire_20_ready;
  wire [2:0]   x22_4_1_bits_instructionIndex;
  wire         x22_4_1_bits_last;
  wire [31:0]  x22_4_1_bits_data;
  wire [3:0]   x22_4_1_bits_mask;
  wire [2:0]   x22_4_1_bits_offset;
  wire [4:0]   x22_4_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_19_bits_instructionIndex;
  wire         sinkVec_sinkWire_19_bits_last;
  wire [31:0]  sinkVec_sinkWire_19_bits_data;
  wire [3:0]   sinkVec_sinkWire_19_bits_mask;
  wire [2:0]   sinkVec_sinkWire_19_bits_offset;
  wire [4:0]   sinkVec_sinkWire_19_bits_vd;
  wire         sinkVec_sinkWire_19_valid;
  wire         sinkVec_sinkWire_19_ready;
  wire [2:0]   x22_4_0_bits_instructionIndex;
  wire [31:0]  x22_4_0_bits_data;
  wire [3:0]   x22_4_0_bits_mask;
  wire [2:0]   x22_4_0_bits_offset;
  wire [4:0]   x22_4_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_18_bits_instructionIndex;
  wire         sinkVec_sinkWire_18_bits_last;
  wire [31:0]  sinkVec_sinkWire_18_bits_data;
  wire [3:0]   sinkVec_sinkWire_18_bits_mask;
  wire [2:0]   sinkVec_sinkWire_18_bits_offset;
  wire [4:0]   sinkVec_sinkWire_18_bits_vd;
  wire         sinkVec_sinkWire_18_valid;
  wire         sinkVec_sinkWire_18_ready;
  wire [2:0]   x13_4_1_bits_instructionIndex;
  wire [2:0]   x13_4_1_bits_offset;
  wire [4:0]   x13_4_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_17_bits_instructionIndex;
  wire [2:0]   sinkVec_sinkWire_17_bits_offset;
  wire [1:0]   sinkVec_sinkWire_17_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_17_bits_vs;
  wire         sinkVec_sinkWire_17_valid;
  wire         sinkVec_sinkWire_17_ready;
  wire [2:0]   x13_4_0_bits_instructionIndex;
  wire [2:0]   x13_4_0_bits_offset;
  wire [4:0]   x13_4_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_16_bits_instructionIndex;
  wire [2:0]   sinkVec_sinkWire_16_bits_offset;
  wire [1:0]   sinkVec_sinkWire_16_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_16_bits_vs;
  wire         sinkVec_sinkWire_16_valid;
  wire         sinkVec_sinkWire_16_ready;
  wire [2:0]   x22_3_1_bits_instructionIndex;
  wire         x22_3_1_bits_last;
  wire [31:0]  x22_3_1_bits_data;
  wire [3:0]   x22_3_1_bits_mask;
  wire [2:0]   x22_3_1_bits_offset;
  wire [4:0]   x22_3_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_15_bits_instructionIndex;
  wire         sinkVec_sinkWire_15_bits_last;
  wire [31:0]  sinkVec_sinkWire_15_bits_data;
  wire [3:0]   sinkVec_sinkWire_15_bits_mask;
  wire [2:0]   sinkVec_sinkWire_15_bits_offset;
  wire [4:0]   sinkVec_sinkWire_15_bits_vd;
  wire         sinkVec_sinkWire_15_valid;
  wire         sinkVec_sinkWire_15_ready;
  wire [2:0]   x22_3_0_bits_instructionIndex;
  wire [31:0]  x22_3_0_bits_data;
  wire [3:0]   x22_3_0_bits_mask;
  wire [2:0]   x22_3_0_bits_offset;
  wire [4:0]   x22_3_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_14_bits_instructionIndex;
  wire         sinkVec_sinkWire_14_bits_last;
  wire [31:0]  sinkVec_sinkWire_14_bits_data;
  wire [3:0]   sinkVec_sinkWire_14_bits_mask;
  wire [2:0]   sinkVec_sinkWire_14_bits_offset;
  wire [4:0]   sinkVec_sinkWire_14_bits_vd;
  wire         sinkVec_sinkWire_14_valid;
  wire         sinkVec_sinkWire_14_ready;
  wire [2:0]   x13_3_1_bits_instructionIndex;
  wire [2:0]   x13_3_1_bits_offset;
  wire [4:0]   x13_3_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_13_bits_instructionIndex;
  wire [2:0]   sinkVec_sinkWire_13_bits_offset;
  wire [1:0]   sinkVec_sinkWire_13_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_13_bits_vs;
  wire         sinkVec_sinkWire_13_valid;
  wire         sinkVec_sinkWire_13_ready;
  wire [2:0]   x13_3_0_bits_instructionIndex;
  wire [2:0]   x13_3_0_bits_offset;
  wire [4:0]   x13_3_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_12_bits_instructionIndex;
  wire [2:0]   sinkVec_sinkWire_12_bits_offset;
  wire [1:0]   sinkVec_sinkWire_12_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_12_bits_vs;
  wire         sinkVec_sinkWire_12_valid;
  wire         sinkVec_sinkWire_12_ready;
  wire [2:0]   x22_2_1_bits_instructionIndex;
  wire         x22_2_1_bits_last;
  wire [31:0]  x22_2_1_bits_data;
  wire [3:0]   x22_2_1_bits_mask;
  wire [2:0]   x22_2_1_bits_offset;
  wire [4:0]   x22_2_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_11_bits_instructionIndex;
  wire         sinkVec_sinkWire_11_bits_last;
  wire [31:0]  sinkVec_sinkWire_11_bits_data;
  wire [3:0]   sinkVec_sinkWire_11_bits_mask;
  wire [2:0]   sinkVec_sinkWire_11_bits_offset;
  wire [4:0]   sinkVec_sinkWire_11_bits_vd;
  wire         sinkVec_sinkWire_11_valid;
  wire         sinkVec_sinkWire_11_ready;
  wire [2:0]   x22_2_0_bits_instructionIndex;
  wire [31:0]  x22_2_0_bits_data;
  wire [3:0]   x22_2_0_bits_mask;
  wire [2:0]   x22_2_0_bits_offset;
  wire [4:0]   x22_2_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_10_bits_instructionIndex;
  wire         sinkVec_sinkWire_10_bits_last;
  wire [31:0]  sinkVec_sinkWire_10_bits_data;
  wire [3:0]   sinkVec_sinkWire_10_bits_mask;
  wire [2:0]   sinkVec_sinkWire_10_bits_offset;
  wire [4:0]   sinkVec_sinkWire_10_bits_vd;
  wire         sinkVec_sinkWire_10_valid;
  wire         sinkVec_sinkWire_10_ready;
  wire [2:0]   x13_2_1_bits_instructionIndex;
  wire [2:0]   x13_2_1_bits_offset;
  wire [4:0]   x13_2_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_9_bits_instructionIndex;
  wire [2:0]   sinkVec_sinkWire_9_bits_offset;
  wire [1:0]   sinkVec_sinkWire_9_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_9_bits_vs;
  wire         sinkVec_sinkWire_9_valid;
  wire         sinkVec_sinkWire_9_ready;
  wire [2:0]   x13_2_0_bits_instructionIndex;
  wire [2:0]   x13_2_0_bits_offset;
  wire [4:0]   x13_2_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_8_bits_instructionIndex;
  wire [2:0]   sinkVec_sinkWire_8_bits_offset;
  wire [1:0]   sinkVec_sinkWire_8_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_8_bits_vs;
  wire         sinkVec_sinkWire_8_valid;
  wire         sinkVec_sinkWire_8_ready;
  wire [2:0]   x22_1_1_bits_instructionIndex;
  wire         x22_1_1_bits_last;
  wire [31:0]  x22_1_1_bits_data;
  wire [3:0]   x22_1_1_bits_mask;
  wire [2:0]   x22_1_1_bits_offset;
  wire [4:0]   x22_1_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_7_bits_instructionIndex;
  wire         sinkVec_sinkWire_7_bits_last;
  wire [31:0]  sinkVec_sinkWire_7_bits_data;
  wire [3:0]   sinkVec_sinkWire_7_bits_mask;
  wire [2:0]   sinkVec_sinkWire_7_bits_offset;
  wire [4:0]   sinkVec_sinkWire_7_bits_vd;
  wire         sinkVec_sinkWire_7_valid;
  wire         sinkVec_sinkWire_7_ready;
  wire [2:0]   x22_1_0_bits_instructionIndex;
  wire [31:0]  x22_1_0_bits_data;
  wire [3:0]   x22_1_0_bits_mask;
  wire [2:0]   x22_1_0_bits_offset;
  wire [4:0]   x22_1_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_6_bits_instructionIndex;
  wire         sinkVec_sinkWire_6_bits_last;
  wire [31:0]  sinkVec_sinkWire_6_bits_data;
  wire [3:0]   sinkVec_sinkWire_6_bits_mask;
  wire [2:0]   sinkVec_sinkWire_6_bits_offset;
  wire [4:0]   sinkVec_sinkWire_6_bits_vd;
  wire         sinkVec_sinkWire_6_valid;
  wire         sinkVec_sinkWire_6_ready;
  wire [2:0]   x13_1_1_bits_instructionIndex;
  wire [2:0]   x13_1_1_bits_offset;
  wire [4:0]   x13_1_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_5_bits_instructionIndex;
  wire [2:0]   sinkVec_sinkWire_5_bits_offset;
  wire [1:0]   sinkVec_sinkWire_5_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_5_bits_vs;
  wire         sinkVec_sinkWire_5_valid;
  wire         sinkVec_sinkWire_5_ready;
  wire [2:0]   x13_1_0_bits_instructionIndex;
  wire [2:0]   x13_1_0_bits_offset;
  wire [4:0]   x13_1_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_4_bits_instructionIndex;
  wire [2:0]   sinkVec_sinkWire_4_bits_offset;
  wire [1:0]   sinkVec_sinkWire_4_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_4_bits_vs;
  wire         sinkVec_sinkWire_4_valid;
  wire         sinkVec_sinkWire_4_ready;
  wire [2:0]   x22_1_bits_instructionIndex;
  wire         x22_1_bits_last;
  wire [31:0]  x22_1_bits_data;
  wire [3:0]   x22_1_bits_mask;
  wire [2:0]   x22_1_bits_offset;
  wire [4:0]   x22_1_bits_vd;
  wire [2:0]   sinkVec_sinkWire_3_bits_instructionIndex;
  wire         sinkVec_sinkWire_3_bits_last;
  wire [31:0]  sinkVec_sinkWire_3_bits_data;
  wire [3:0]   sinkVec_sinkWire_3_bits_mask;
  wire [2:0]   sinkVec_sinkWire_3_bits_offset;
  wire [4:0]   sinkVec_sinkWire_3_bits_vd;
  wire         sinkVec_sinkWire_3_valid;
  wire         sinkVec_sinkWire_3_ready;
  wire [2:0]   x22_0_bits_instructionIndex;
  wire [31:0]  x22_0_bits_data;
  wire [3:0]   x22_0_bits_mask;
  wire [2:0]   x22_0_bits_offset;
  wire [4:0]   x22_0_bits_vd;
  wire [2:0]   sinkVec_sinkWire_2_bits_instructionIndex;
  wire         sinkVec_sinkWire_2_bits_last;
  wire [31:0]  sinkVec_sinkWire_2_bits_data;
  wire [3:0]   sinkVec_sinkWire_2_bits_mask;
  wire [2:0]   sinkVec_sinkWire_2_bits_offset;
  wire [4:0]   sinkVec_sinkWire_2_bits_vd;
  wire         sinkVec_sinkWire_2_valid;
  wire         sinkVec_sinkWire_2_ready;
  wire [2:0]   x13_1_bits_instructionIndex;
  wire [2:0]   x13_1_bits_offset;
  wire [4:0]   x13_1_bits_vs;
  wire [2:0]   sinkVec_sinkWire_1_bits_instructionIndex;
  wire [2:0]   sinkVec_sinkWire_1_bits_offset;
  wire [1:0]   sinkVec_sinkWire_1_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_1_bits_vs;
  wire         sinkVec_sinkWire_1_valid;
  wire         sinkVec_sinkWire_1_ready;
  wire [2:0]   x13_0_bits_instructionIndex;
  wire [2:0]   x13_0_bits_offset;
  wire [4:0]   x13_0_bits_vs;
  wire [2:0]   sinkVec_sinkWire_bits_instructionIndex;
  wire [2:0]   sinkVec_sinkWire_bits_offset;
  wire [1:0]   sinkVec_sinkWire_bits_readSource;
  wire [4:0]   sinkVec_sinkWire_bits_vs;
  wire         sinkVec_sinkWire_valid;
  wire         sinkVec_sinkWire_ready;
  wire [1:0]   laneRequestSourceWire_7_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_7_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_7_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_7_bits_segment;
  wire [1:0]   laneRequestSourceWire_7_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_7_bits_vd;
  wire [4:0]   laneRequestSourceWire_7_bits_vs1;
  wire         laneRequestSourceWire_7_bits_issueInst;
  wire         laneRequestSinkWire_7_ready;
  wire [1:0]   laneRequestSourceWire_6_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_6_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_6_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_6_bits_segment;
  wire [1:0]   laneRequestSourceWire_6_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_6_bits_vd;
  wire [4:0]   laneRequestSourceWire_6_bits_vs1;
  wire         laneRequestSourceWire_6_bits_issueInst;
  wire         laneRequestSinkWire_6_ready;
  wire [1:0]   laneRequestSourceWire_5_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_5_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_5_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_5_bits_segment;
  wire [1:0]   laneRequestSourceWire_5_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_5_bits_vd;
  wire [4:0]   laneRequestSourceWire_5_bits_vs1;
  wire         laneRequestSourceWire_5_bits_issueInst;
  wire         laneRequestSinkWire_5_ready;
  wire [1:0]   laneRequestSourceWire_4_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_4_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_4_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_4_bits_segment;
  wire [1:0]   laneRequestSourceWire_4_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_4_bits_vd;
  wire [4:0]   laneRequestSourceWire_4_bits_vs1;
  wire         laneRequestSourceWire_4_bits_issueInst;
  wire         laneRequestSinkWire_4_ready;
  wire [1:0]   laneRequestSourceWire_3_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_3_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_3_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_3_bits_segment;
  wire [1:0]   laneRequestSourceWire_3_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_3_bits_vd;
  wire [4:0]   laneRequestSourceWire_3_bits_vs1;
  wire         laneRequestSourceWire_3_bits_issueInst;
  wire         laneRequestSinkWire_3_ready;
  wire [1:0]   laneRequestSourceWire_2_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_2_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_2_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_2_bits_segment;
  wire [1:0]   laneRequestSourceWire_2_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_2_bits_vd;
  wire [4:0]   laneRequestSourceWire_2_bits_vs1;
  wire         laneRequestSourceWire_2_bits_issueInst;
  wire         laneRequestSinkWire_2_ready;
  wire [1:0]   laneRequestSourceWire_1_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_1_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_1_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_1_bits_segment;
  wire [1:0]   laneRequestSourceWire_1_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_1_bits_vd;
  wire [4:0]   laneRequestSourceWire_1_bits_vs1;
  wire         laneRequestSourceWire_1_bits_issueInst;
  wire         laneRequestSinkWire_1_ready;
  wire [1:0]   laneRequestSourceWire_0_bits_csrInterface_vSew;
  wire [11:0]  laneRequestSourceWire_0_bits_csrInterface_vl;
  wire [31:0]  laneRequestSourceWire_0_bits_readFromScalar;
  wire [2:0]   laneRequestSourceWire_0_bits_segment;
  wire [1:0]   laneRequestSourceWire_0_bits_loadStoreEEW;
  wire [4:0]   laneRequestSourceWire_0_bits_vd;
  wire [4:0]   laneRequestSourceWire_0_bits_vs1;
  wire         laneRequestSourceWire_0_bits_issueInst;
  wire         laneRequestSinkWire_0_ready;
  wire [1:0]   requestRegCSR_vxrm;
  wire [11:0]  requestRegCSR_vStart;
  wire         requestRegCSR_vma;
  wire         requestRegCSR_vta;
  wire [2:0]   requestRegCSR_vlmul;
  wire         indexedLoadStorePort_aw_ready_0 = indexedLoadStorePort_aw_ready;
  wire         indexedLoadStorePort_w_ready_0 = indexedLoadStorePort_w_ready;
  wire         indexedLoadStorePort_b_valid_0 = indexedLoadStorePort_b_valid;
  wire [1:0]   indexedLoadStorePort_b_bits_id_0 = indexedLoadStorePort_b_bits_id;
  wire [1:0]   indexedLoadStorePort_b_bits_resp_0 = indexedLoadStorePort_b_bits_resp;
  wire         indexedLoadStorePort_ar_ready_0 = indexedLoadStorePort_ar_ready;
  wire         indexedLoadStorePort_r_valid_0 = indexedLoadStorePort_r_valid;
  wire [1:0]   indexedLoadStorePort_r_bits_id_0 = indexedLoadStorePort_r_bits_id;
  wire [31:0]  indexedLoadStorePort_r_bits_data_0 = indexedLoadStorePort_r_bits_data;
  wire [1:0]   indexedLoadStorePort_r_bits_resp_0 = indexedLoadStorePort_r_bits_resp;
  wire         indexedLoadStorePort_r_bits_last_0 = indexedLoadStorePort_r_bits_last;
  wire         highBandwidthLoadStorePort_aw_ready_0 = highBandwidthLoadStorePort_aw_ready;
  wire         highBandwidthLoadStorePort_w_ready_0 = highBandwidthLoadStorePort_w_ready;
  wire         highBandwidthLoadStorePort_b_valid_0 = highBandwidthLoadStorePort_b_valid;
  wire [1:0]   highBandwidthLoadStorePort_b_bits_id_0 = highBandwidthLoadStorePort_b_bits_id;
  wire [1:0]   highBandwidthLoadStorePort_b_bits_resp_0 = highBandwidthLoadStorePort_b_bits_resp;
  wire         highBandwidthLoadStorePort_ar_ready_0 = highBandwidthLoadStorePort_ar_ready;
  wire         highBandwidthLoadStorePort_r_valid_0 = highBandwidthLoadStorePort_r_valid;
  wire [1:0]   highBandwidthLoadStorePort_r_bits_id_0 = highBandwidthLoadStorePort_r_bits_id;
  wire [255:0] highBandwidthLoadStorePort_r_bits_data_0 = highBandwidthLoadStorePort_r_bits_data;
  wire [1:0]   highBandwidthLoadStorePort_r_bits_resp_0 = highBandwidthLoadStorePort_r_bits_resp;
  wire         highBandwidthLoadStorePort_r_bits_last_0 = highBandwidthLoadStorePort_r_bits_last;
  wire         issue_valid_0 = issue_valid;
  wire [31:0]  issue_bits_instruction_0 = issue_bits_instruction;
  wire [31:0]  issue_bits_rs1Data_0 = issue_bits_rs1Data;
  wire [31:0]  issue_bits_rs2Data_0 = issue_bits_rs2Data;
  wire [31:0]  issue_bits_vtype_0 = issue_bits_vtype;
  wire [31:0]  issue_bits_vl_0 = issue_bits_vl;
  wire [31:0]  issue_bits_vstart_0 = issue_bits_vstart;
  wire [31:0]  issue_bits_vcsr_0 = issue_bits_vcsr;
  wire [7:0]   indexedLoadStorePort_aw_bits_len_0 = 8'h0;
  wire [7:0]   indexedLoadStorePort_ar_bits_len_0 = 8'h0;
  wire [7:0]   highBandwidthLoadStorePort_aw_bits_len_0 = 8'h0;
  wire [7:0]   highBandwidthLoadStorePort_ar_bits_len_0 = 8'h0;
  wire [1:0]   indexedLoadStorePort_ar_bits_id_0 = 2'h0;
  wire [1:0]   highBandwidthLoadStorePort_ar_bits_id_0 = 2'h0;
  wire [1:0]   indexedLoadStorePort_aw_bits_burst_0 = 2'h1;
  wire [1:0]   indexedLoadStorePort_ar_bits_burst_0 = 2'h1;
  wire [1:0]   highBandwidthLoadStorePort_aw_bits_burst_0 = 2'h1;
  wire [1:0]   highBandwidthLoadStorePort_ar_bits_burst_0 = 2'h1;
  wire [3:0]   indexedLoadStorePort_aw_bits_cache_0 = 4'h0;
  wire [3:0]   indexedLoadStorePort_aw_bits_qos_0 = 4'h0;
  wire [3:0]   indexedLoadStorePort_aw_bits_region_0 = 4'h0;
  wire [3:0]   indexedLoadStorePort_ar_bits_cache_0 = 4'h0;
  wire [3:0]   indexedLoadStorePort_ar_bits_qos_0 = 4'h0;
  wire [3:0]   indexedLoadStorePort_ar_bits_region_0 = 4'h0;
  wire [3:0]   highBandwidthLoadStorePort_aw_bits_cache_0 = 4'h0;
  wire [3:0]   highBandwidthLoadStorePort_aw_bits_qos_0 = 4'h0;
  wire [3:0]   highBandwidthLoadStorePort_aw_bits_region_0 = 4'h0;
  wire [3:0]   highBandwidthLoadStorePort_ar_bits_cache_0 = 4'h0;
  wire [3:0]   highBandwidthLoadStorePort_ar_bits_qos_0 = 4'h0;
  wire [3:0]   highBandwidthLoadStorePort_ar_bits_region_0 = 4'h0;
  wire [31:0]  retire_csr_bits_fflag_0 = 32'h0;
  wire [2:0]   indexedLoadStorePort_aw_bits_prot_0 = 3'h0;
  wire [2:0]   indexedLoadStorePort_ar_bits_prot_0 = 3'h0;
  wire [2:0]   highBandwidthLoadStorePort_aw_bits_prot_0 = 3'h0;
  wire [2:0]   highBandwidthLoadStorePort_ar_bits_prot_0 = 3'h0;
  wire [2:0]   indexedLoadStorePort_ar_bits_size_0 = 3'h2;
  wire [2:0]   highBandwidthLoadStorePort_aw_bits_size_0 = 3'h5;
  wire [2:0]   highBandwidthLoadStorePort_ar_bits_size_0 = 3'h5;
  wire [1:0]   x13_0_bits_readSource = 2'h2;
  wire [1:0]   x13_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_1_bits_readSource = 2'h2;
  wire [1:0]   x13_1_0_bits_readSource = 2'h2;
  wire [1:0]   x13_1_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_4_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_5_bits_readSource = 2'h2;
  wire [1:0]   x13_2_0_bits_readSource = 2'h2;
  wire [1:0]   x13_2_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_8_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_9_bits_readSource = 2'h2;
  wire [1:0]   x13_3_0_bits_readSource = 2'h2;
  wire [1:0]   x13_3_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_12_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_13_bits_readSource = 2'h2;
  wire [1:0]   x13_4_0_bits_readSource = 2'h2;
  wire [1:0]   x13_4_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_16_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_17_bits_readSource = 2'h2;
  wire [1:0]   x13_5_0_bits_readSource = 2'h2;
  wire [1:0]   x13_5_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_20_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_21_bits_readSource = 2'h2;
  wire [1:0]   x13_6_0_bits_readSource = 2'h2;
  wire [1:0]   x13_6_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_24_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_25_bits_readSource = 2'h2;
  wire [1:0]   x13_7_0_bits_readSource = 2'h2;
  wire [1:0]   x13_7_1_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_28_bits_readSource = 2'h2;
  wire [1:0]   sinkVec_validSource_29_bits_readSource = 2'h2;
  wire [1:0]   lo_lo = 2'h3;
  wire [1:0]   lo_hi = 2'h3;
  wire [1:0]   hi_lo = 2'h3;
  wire [1:0]   hi_hi = 2'h3;
  wire [1:0]   lo_lo_1 = 2'h3;
  wire [1:0]   lo_hi_1 = 2'h3;
  wire [1:0]   hi_lo_1 = 2'h3;
  wire [1:0]   hi_hi_1 = 2'h3;
  wire [3:0]   lo = 4'hF;
  wire [3:0]   hi = 4'hF;
  wire [3:0]   lo_1 = 4'hF;
  wire [3:0]   hi_1 = 4'hF;
  wire         indexedLoadStorePort_w_bits_last_0 = 1'h1;
  wire         indexedLoadStorePort_b_ready_0 = 1'h1;
  wire         highBandwidthLoadStorePort_w_bits_last_0 = 1'h1;
  wire         highBandwidthLoadStorePort_b_ready_0 = 1'h1;
  wire [2:0]   vSewOHForMask = 3'h1;
  wire         indexedLoadStorePort_aw_bits_lock_0 = 1'h0;
  wire         indexedLoadStorePort_ar_bits_lock_0 = 1'h0;
  wire         highBandwidthLoadStorePort_aw_bits_lock_0 = 1'h0;
  wire         highBandwidthLoadStorePort_ar_bits_lock_0 = 1'h0;
  wire         retire_rd_bits_isFp_0 = 1'h0;
  wire         retire_csr_valid_0 = 1'h0;
  wire         x22_0_bits_last = 1'h0;
  wire         sinkVec_queue_2_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_2_bits_last = 1'h0;
  wire         sinkVec_validSink_2_bits_last = 1'h0;
  wire         x22_1_0_bits_last = 1'h0;
  wire         sinkVec_queue_6_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_6_bits_last = 1'h0;
  wire         sinkVec_validSink_6_bits_last = 1'h0;
  wire         x22_2_0_bits_last = 1'h0;
  wire         sinkVec_queue_10_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_10_bits_last = 1'h0;
  wire         sinkVec_validSink_10_bits_last = 1'h0;
  wire         x22_3_0_bits_last = 1'h0;
  wire         sinkVec_queue_14_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_14_bits_last = 1'h0;
  wire         sinkVec_validSink_14_bits_last = 1'h0;
  wire         x22_4_0_bits_last = 1'h0;
  wire         sinkVec_queue_18_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_18_bits_last = 1'h0;
  wire         sinkVec_validSink_18_bits_last = 1'h0;
  wire         x22_5_0_bits_last = 1'h0;
  wire         sinkVec_queue_22_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_22_bits_last = 1'h0;
  wire         sinkVec_validSink_22_bits_last = 1'h0;
  wire         x22_6_0_bits_last = 1'h0;
  wire         sinkVec_queue_26_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_26_bits_last = 1'h0;
  wire         sinkVec_validSink_26_bits_last = 1'h0;
  wire         x22_7_0_bits_last = 1'h0;
  wire         sinkVec_queue_30_enq_bits_last = 1'h0;
  wire         sinkVec_validSource_30_bits_last = 1'h0;
  wire         sinkVec_validSink_30_bits_last = 1'h0;
  reg  [2:0]   instructionCounter;
  wire [2:0]   nextInstructionCounter = instructionCounter + 3'h1;
  wire         issue_ready_0;
  wire         _probeWire_issue_valid_T = issue_ready_0 & issue_valid_0;
  reg  [2:0]   responseCounter;
  wire [2:0]   nextResponseCounter = responseCounter + 3'h1;
  reg          requestReg_valid;
  wire         requestRegDequeue_valid = requestReg_valid;
  reg  [31:0]  requestReg_bits_issue_instruction;
  wire [31:0]  requestRegDequeue_bits_instruction = requestReg_bits_issue_instruction;
  reg  [31:0]  requestReg_bits_issue_rs1Data;
  wire [31:0]  requestRegDequeue_bits_rs1Data = requestReg_bits_issue_rs1Data;
  reg  [31:0]  requestReg_bits_issue_rs2Data;
  wire [31:0]  requestRegDequeue_bits_rs2Data = requestReg_bits_issue_rs2Data;
  reg  [31:0]  requestReg_bits_issue_vtype;
  wire [31:0]  requestRegDequeue_bits_vtype = requestReg_bits_issue_vtype;
  reg  [31:0]  requestReg_bits_issue_vl;
  wire [31:0]  requestRegDequeue_bits_vl = requestReg_bits_issue_vl;
  reg  [31:0]  requestReg_bits_issue_vstart;
  wire [31:0]  requestRegDequeue_bits_vstart = requestReg_bits_issue_vstart;
  reg  [31:0]  requestReg_bits_issue_vcsr;
  wire [31:0]  requestRegDequeue_bits_vcsr = requestReg_bits_issue_vcsr;
  reg          requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_0_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_1_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_2_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_3_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_4_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_5_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_6_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  wire         laneRequestSourceWire_7_bits_decodeResult_specialSlot = requestReg_bits_decodeResult_specialSlot;
  reg  [4:0]   requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_0_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_1_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_2_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_3_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_4_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_5_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_6_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  wire [4:0]   laneRequestSourceWire_7_bits_decodeResult_topUop = requestReg_bits_decodeResult_topUop;
  reg          requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_0_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_1_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_2_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_3_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_4_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_5_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_6_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  wire         laneRequestSourceWire_7_bits_decodeResult_popCount = requestReg_bits_decodeResult_popCount;
  reg          requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_0_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_1_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_2_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_3_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_4_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_5_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_6_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  wire         laneRequestSourceWire_7_bits_decodeResult_ffo = requestReg_bits_decodeResult_ffo;
  reg          requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_0_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_1_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_2_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_3_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_4_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_5_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_6_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  wire         laneRequestSourceWire_7_bits_decodeResult_average = requestReg_bits_decodeResult_average;
  reg          requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_0_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_1_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_2_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_3_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_4_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_5_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_6_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  wire         laneRequestSourceWire_7_bits_decodeResult_reverse = requestReg_bits_decodeResult_reverse;
  reg          requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_0_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_1_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_2_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_3_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_4_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_5_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_6_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSourceWire_7_bits_decodeResult_dontNeedExecuteInLane = requestReg_bits_decodeResult_dontNeedExecuteInLane;
  reg          requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_0_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_1_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_2_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_3_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_4_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_5_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_6_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  wire         laneRequestSourceWire_7_bits_decodeResult_scheduler = requestReg_bits_decodeResult_scheduler;
  reg          requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_0_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_1_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_2_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_3_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_4_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_5_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_6_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  wire         laneRequestSourceWire_7_bits_decodeResult_sReadVD = requestReg_bits_decodeResult_sReadVD;
  reg          requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_0_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_1_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_2_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_3_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_4_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_5_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_6_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  wire         laneRequestSourceWire_7_bits_decodeResult_vtype = requestReg_bits_decodeResult_vtype;
  reg          requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_0_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_1_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_2_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_3_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_4_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_5_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_6_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  wire         laneRequestSourceWire_7_bits_decodeResult_sWrite = requestReg_bits_decodeResult_sWrite;
  reg          requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_0_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_1_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_2_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_3_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_4_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_5_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_6_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  wire         laneRequestSourceWire_7_bits_decodeResult_crossRead = requestReg_bits_decodeResult_crossRead;
  reg          requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_0_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_1_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_2_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_3_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_4_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_5_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_6_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  wire         laneRequestSourceWire_7_bits_decodeResult_crossWrite = requestReg_bits_decodeResult_crossWrite;
  reg          requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_0_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_1_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_2_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_3_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_4_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_5_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_6_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  wire         laneRequestSourceWire_7_bits_decodeResult_maskUnit = requestReg_bits_decodeResult_maskUnit;
  reg          requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_0_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_1_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_2_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_3_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_4_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_5_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_6_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  wire         laneRequestSourceWire_7_bits_decodeResult_special = requestReg_bits_decodeResult_special;
  reg          requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_0_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_1_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_2_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_3_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_4_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_5_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_6_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  wire         laneRequestSourceWire_7_bits_decodeResult_saturate = requestReg_bits_decodeResult_saturate;
  reg          requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_0_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_1_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_2_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_3_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_4_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_5_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_6_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  wire         laneRequestSourceWire_7_bits_decodeResult_vwmacc = requestReg_bits_decodeResult_vwmacc;
  reg          requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_0_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_1_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_2_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_3_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_4_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_5_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_6_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  wire         laneRequestSourceWire_7_bits_decodeResult_readOnly = requestReg_bits_decodeResult_readOnly;
  reg          requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_0_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_1_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_2_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_3_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_4_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_5_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_6_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  wire         laneRequestSourceWire_7_bits_decodeResult_maskSource = requestReg_bits_decodeResult_maskSource;
  reg          requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_0_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_1_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_2_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_3_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_4_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_5_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_6_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  wire         laneRequestSourceWire_7_bits_decodeResult_maskDestination = requestReg_bits_decodeResult_maskDestination;
  reg          requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_0_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_1_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_2_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_3_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_4_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_5_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_6_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  wire         laneRequestSourceWire_7_bits_decodeResult_maskLogic = requestReg_bits_decodeResult_maskLogic;
  reg  [3:0]   requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_0_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_1_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_2_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_3_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_4_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_5_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_6_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  wire [3:0]   laneRequestSourceWire_7_bits_decodeResult_uop = requestReg_bits_decodeResult_uop;
  reg          requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_0_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_1_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_2_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_3_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_4_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_5_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_6_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  wire         laneRequestSourceWire_7_bits_decodeResult_iota = requestReg_bits_decodeResult_iota;
  reg          requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_0_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_1_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_2_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_3_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_4_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_5_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_6_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  wire         laneRequestSourceWire_7_bits_decodeResult_mv = requestReg_bits_decodeResult_mv;
  reg          requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_0_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_1_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_2_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_3_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_4_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_5_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_6_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  wire         laneRequestSourceWire_7_bits_decodeResult_extend = requestReg_bits_decodeResult_extend;
  reg          requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_0_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_1_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_2_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_3_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_4_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_5_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_6_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  wire         laneRequestSourceWire_7_bits_decodeResult_unOrderWrite = requestReg_bits_decodeResult_unOrderWrite;
  reg          requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_0_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_1_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_2_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_3_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_4_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_5_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_6_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  wire         laneRequestSourceWire_7_bits_decodeResult_compress = requestReg_bits_decodeResult_compress;
  reg          requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_0_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_1_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_2_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_3_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_4_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_5_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_6_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  wire         laneRequestSourceWire_7_bits_decodeResult_gather16 = requestReg_bits_decodeResult_gather16;
  reg          requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_0_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_1_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_2_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_3_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_4_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_5_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_6_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  wire         laneRequestSourceWire_7_bits_decodeResult_gather = requestReg_bits_decodeResult_gather;
  reg          requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_0_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_1_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_2_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_3_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_4_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_5_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_6_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  wire         laneRequestSourceWire_7_bits_decodeResult_slid = requestReg_bits_decodeResult_slid;
  reg          requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_0_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_1_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_2_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_3_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_4_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_5_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_6_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  wire         laneRequestSourceWire_7_bits_decodeResult_targetRd = requestReg_bits_decodeResult_targetRd;
  reg          requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_0_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_1_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_2_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_3_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_4_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_5_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_6_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  wire         laneRequestSourceWire_7_bits_decodeResult_widenReduce = requestReg_bits_decodeResult_widenReduce;
  reg          requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_0_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_1_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_2_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_3_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_4_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_5_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_6_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  wire         laneRequestSourceWire_7_bits_decodeResult_red = requestReg_bits_decodeResult_red;
  reg          requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_0_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_1_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_2_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_3_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_4_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_5_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_6_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  wire         laneRequestSourceWire_7_bits_decodeResult_nr = requestReg_bits_decodeResult_nr;
  reg          requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_0_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_1_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_2_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_3_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_4_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_5_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_6_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  wire         laneRequestSourceWire_7_bits_decodeResult_itype = requestReg_bits_decodeResult_itype;
  reg          requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_0_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_1_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_2_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_3_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_4_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_5_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_6_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  wire         laneRequestSourceWire_7_bits_decodeResult_unsigned1 = requestReg_bits_decodeResult_unsigned1;
  reg          requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_0_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_1_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_2_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_3_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_4_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_5_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_6_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  wire         laneRequestSourceWire_7_bits_decodeResult_unsigned0 = requestReg_bits_decodeResult_unsigned0;
  reg          requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_0_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_1_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_2_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_3_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_4_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_5_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_6_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  wire         laneRequestSourceWire_7_bits_decodeResult_other = requestReg_bits_decodeResult_other;
  reg          requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_0_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_1_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_2_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_3_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_4_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_5_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_6_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  wire         laneRequestSourceWire_7_bits_decodeResult_multiCycle = requestReg_bits_decodeResult_multiCycle;
  reg          requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_0_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_1_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_2_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_3_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_4_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_5_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_6_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  wire         laneRequestSourceWire_7_bits_decodeResult_divider = requestReg_bits_decodeResult_divider;
  reg          requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_0_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_1_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_2_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_3_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_4_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_5_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_6_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  wire         laneRequestSourceWire_7_bits_decodeResult_multiplier = requestReg_bits_decodeResult_multiplier;
  reg          requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_0_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_1_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_2_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_3_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_4_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_5_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_6_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  wire         laneRequestSourceWire_7_bits_decodeResult_shift = requestReg_bits_decodeResult_shift;
  reg          requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_0_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_1_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_2_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_3_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_4_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_5_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_6_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  wire         laneRequestSourceWire_7_bits_decodeResult_adder = requestReg_bits_decodeResult_adder;
  reg          requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_0_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_1_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_2_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_3_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_4_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_5_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_6_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  wire         laneRequestSourceWire_7_bits_decodeResult_logic = requestReg_bits_decodeResult_logic;
  reg  [2:0]   requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_0_bits_instructionIndex = requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_1_bits_instructionIndex = requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_2_bits_instructionIndex = requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_3_bits_instructionIndex = requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_4_bits_instructionIndex = requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_5_bits_instructionIndex = requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_6_bits_instructionIndex = requestReg_bits_instructionIndex;
  wire [2:0]   laneRequestSourceWire_7_bits_instructionIndex = requestReg_bits_instructionIndex;
  reg          requestReg_bits_vdIsV0;
  reg  [11:0]  requestReg_bits_writeByte;
  wire [11:0]  laneRequestSourceWire_0_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [11:0]  laneRequestSourceWire_1_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [11:0]  laneRequestSourceWire_2_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [11:0]  laneRequestSourceWire_3_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [11:0]  laneRequestSourceWire_4_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [11:0]  laneRequestSourceWire_5_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [11:0]  laneRequestSourceWire_6_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [11:0]  laneRequestSourceWire_7_bits_csrInterface_vStart = requestRegCSR_vStart;
  wire [2:0]   laneRequestSourceWire_0_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [2:0]   laneRequestSourceWire_1_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [2:0]   laneRequestSourceWire_2_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [2:0]   laneRequestSourceWire_3_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [2:0]   laneRequestSourceWire_4_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [2:0]   laneRequestSourceWire_5_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [2:0]   laneRequestSourceWire_6_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [2:0]   laneRequestSourceWire_7_bits_csrInterface_vlmul = requestRegCSR_vlmul;
  wire [1:0]   laneRequestSourceWire_0_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire [1:0]   laneRequestSourceWire_1_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire [1:0]   laneRequestSourceWire_2_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire [1:0]   laneRequestSourceWire_3_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire [1:0]   laneRequestSourceWire_4_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire [1:0]   laneRequestSourceWire_5_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire [1:0]   laneRequestSourceWire_6_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire [1:0]   laneRequestSourceWire_7_bits_csrInterface_vxrm = requestRegCSR_vxrm;
  wire         laneRequestSourceWire_0_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_1_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_2_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_3_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_4_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_5_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_6_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_7_bits_csrInterface_vta = requestRegCSR_vta;
  wire         laneRequestSourceWire_0_bits_csrInterface_vma = requestRegCSR_vma;
  wire         laneRequestSourceWire_1_bits_csrInterface_vma = requestRegCSR_vma;
  wire         laneRequestSourceWire_2_bits_csrInterface_vma = requestRegCSR_vma;
  wire         laneRequestSourceWire_3_bits_csrInterface_vma = requestRegCSR_vma;
  wire         laneRequestSourceWire_4_bits_csrInterface_vma = requestRegCSR_vma;
  wire         laneRequestSourceWire_5_bits_csrInterface_vma = requestRegCSR_vma;
  wire         laneRequestSourceWire_6_bits_csrInterface_vma = requestRegCSR_vma;
  wire         laneRequestSourceWire_7_bits_csrInterface_vma = requestRegCSR_vma;
  assign requestRegCSR_vlmul = requestReg_bits_issue_vtype[2:0];
  wire [1:0]   requestRegCSR_vSew = requestReg_bits_issue_vtype[4:3];
  assign requestRegCSR_vta = requestReg_bits_issue_vtype[6];
  assign requestRegCSR_vma = requestReg_bits_issue_vtype[7];
  wire [11:0]  requestRegCSR_vl = requestReg_bits_issue_vl[11:0];
  assign requestRegCSR_vStart = requestReg_bits_issue_vstart[11:0];
  assign requestRegCSR_vxrm = requestReg_bits_issue_vcsr[2:1];
  wire         requestRegDequeue_ready;
  wire         maskUnit_gatherData_ready = requestRegDequeue_ready & requestRegDequeue_valid;
  wire         laneRequestSourceWire_0_valid;
  assign laneRequestSourceWire_0_valid = maskUnit_gatherData_ready;
  wire         laneRequestSourceWire_1_valid;
  assign laneRequestSourceWire_1_valid = maskUnit_gatherData_ready;
  wire         laneRequestSourceWire_2_valid;
  assign laneRequestSourceWire_2_valid = maskUnit_gatherData_ready;
  wire         laneRequestSourceWire_3_valid;
  assign laneRequestSourceWire_3_valid = maskUnit_gatherData_ready;
  wire         laneRequestSourceWire_4_valid;
  assign laneRequestSourceWire_4_valid = maskUnit_gatherData_ready;
  wire         laneRequestSourceWire_5_valid;
  assign laneRequestSourceWire_5_valid = maskUnit_gatherData_ready;
  wire         laneRequestSourceWire_6_valid;
  assign laneRequestSourceWire_6_valid = maskUnit_gatherData_ready;
  wire         laneRequestSourceWire_7_valid;
  assign laneRequestSourceWire_7_valid = maskUnit_gatherData_ready;
  assign issue_ready_0 = ~requestReg_valid | requestRegDequeue_ready;
  wire         isLoadStoreType = ~(requestRegDequeue_bits_instruction[6]) & requestRegDequeue_valid;
  wire         laneRequestSourceWire_0_bits_loadStore = isLoadStoreType;
  wire         laneRequestSourceWire_1_bits_loadStore = isLoadStoreType;
  wire         laneRequestSourceWire_2_bits_loadStore = isLoadStoreType;
  wire         laneRequestSourceWire_3_bits_loadStore = isLoadStoreType;
  wire         laneRequestSourceWire_4_bits_loadStore = isLoadStoreType;
  wire         laneRequestSourceWire_5_bits_loadStore = isLoadStoreType;
  wire         laneRequestSourceWire_6_bits_loadStore = isLoadStoreType;
  wire         laneRequestSourceWire_7_bits_loadStore = isLoadStoreType;
  wire         isStoreType = ~(requestRegDequeue_bits_instruction[6]) & requestRegDequeue_bits_instruction[5];
  wire         laneRequestSourceWire_0_bits_store = isStoreType;
  wire         laneRequestSourceWire_1_bits_store = isStoreType;
  wire         laneRequestSourceWire_2_bits_store = isStoreType;
  wire         laneRequestSourceWire_3_bits_store = isStoreType;
  wire         laneRequestSourceWire_4_bits_store = isStoreType;
  wire         laneRequestSourceWire_5_bits_store = isStoreType;
  wire         laneRequestSourceWire_6_bits_store = isStoreType;
  wire         laneRequestSourceWire_7_bits_store = isStoreType;
  wire         maskType = ~(requestRegDequeue_bits_instruction[25]);
  wire         laneRequestSourceWire_0_bits_mask = maskType;
  wire         laneRequestSourceWire_1_bits_mask = maskType;
  wire         laneRequestSourceWire_2_bits_mask = maskType;
  wire         laneRequestSourceWire_3_bits_mask = maskType;
  wire         laneRequestSourceWire_4_bits_mask = maskType;
  wire         laneRequestSourceWire_5_bits_mask = maskType;
  wire         laneRequestSourceWire_6_bits_mask = maskType;
  wire         laneRequestSourceWire_7_bits_mask = maskType;
  wire [4:0]   laneRequestSourceWire_0_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire [4:0]   laneRequestSourceWire_1_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire [4:0]   laneRequestSourceWire_2_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire [4:0]   laneRequestSourceWire_3_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire [4:0]   laneRequestSourceWire_4_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire [4:0]   laneRequestSourceWire_5_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire [4:0]   laneRequestSourceWire_6_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire [4:0]   laneRequestSourceWire_7_bits_vs2 = requestRegDequeue_bits_instruction[24:20];
  wire         lsWholeReg = isLoadStoreType & requestRegDequeue_bits_instruction[27:26] == 2'h0 & requestRegDequeue_bits_instruction[24:20] == 5'h8;
  wire         laneRequestSourceWire_0_bits_lsWholeReg = lsWholeReg;
  wire         laneRequestSourceWire_1_bits_lsWholeReg = lsWholeReg;
  wire         laneRequestSourceWire_2_bits_lsWholeReg = lsWholeReg;
  wire         laneRequestSourceWire_3_bits_lsWholeReg = lsWholeReg;
  wire         laneRequestSourceWire_4_bits_lsWholeReg = lsWholeReg;
  wire         laneRequestSourceWire_5_bits_lsWholeReg = lsWholeReg;
  wire         laneRequestSourceWire_6_bits_lsWholeReg = lsWholeReg;
  wire         laneRequestSourceWire_7_bits_lsWholeReg = lsWholeReg;
  wire         maskUnitInstruction = requestReg_bits_decodeResult_slid | requestReg_bits_decodeResult_mv;
  wire         skipLastFromLane = isStoreType | maskUnitInstruction | requestReg_bits_decodeResult_readOnly;
  wire         instructionValid = requestReg_bits_issue_vl > requestReg_bits_issue_vstart;
  wire         noOffsetReadLoadStore = isLoadStoreType & ~(requestRegDequeue_bits_instruction[26]);
  wire [7:0]   vSew1H = 8'h1 << requestReg_bits_issue_vtype[5:3];
  wire [31:0]  source1Extend =
    (vSew1H[0] ? {{24{requestRegDequeue_bits_rs1Data[7] & ~requestReg_bits_decodeResult_unsigned0}}, requestRegDequeue_bits_rs1Data[7:0]} : 32'h0)
    | (vSew1H[1] ? {{16{requestRegDequeue_bits_rs1Data[15] & ~requestReg_bits_decodeResult_unsigned0}}, requestRegDequeue_bits_rs1Data[15:0]} : 32'h0) | (vSew1H[2] ? requestRegDequeue_bits_rs1Data : 32'h0);
  wire         src1IsSInt;
  assign src1IsSInt = ~requestReg_bits_decodeResult_unsigned0;
  wire [4:0]   imm = requestReg_bits_issue_instruction[19:15];
  wire [31:0]  immSignExtend = {{16{imm[4] & (vSew1H[2] | src1IsSInt)}}, {8{imm[4] & (vSew1H[1] | vSew1H[2] | src1IsSInt)}}, {3{imm[4]}}, imm};
  wire         slotCommit_3;
  wire [3:0]   vxsatReportVec_0;
  wire [3:0]   vxsatReportVec_1;
  wire [3:0]   vxsatReportVec_2;
  wire [3:0]   vxsatReportVec_3;
  wire [3:0]   vxsatReportVec_4;
  wire [3:0]   vxsatReportVec_5;
  wire [3:0]   vxsatReportVec_6;
  wire [3:0]   vxsatReportVec_7;
  wire [3:0]   vxsatReport = vxsatReportVec_0 | vxsatReportVec_1 | vxsatReportVec_2 | vxsatReportVec_3 | vxsatReportVec_4 | vxsatReportVec_5 | vxsatReportVec_6 | vxsatReportVec_7;
  wire         specialInstruction = requestReg_bits_decodeResult_special | requestReg_bits_vdIsV0;
  wire         laneRequestSourceWire_0_bits_special = specialInstruction;
  wire         laneRequestSourceWire_1_bits_special = specialInstruction;
  wire         laneRequestSourceWire_2_bits_special = specialInstruction;
  wire         laneRequestSourceWire_3_bits_special = specialInstruction;
  wire         laneRequestSourceWire_4_bits_special = specialInstruction;
  wire         laneRequestSourceWire_5_bits_special = specialInstruction;
  wire         laneRequestSourceWire_6_bits_special = specialInstruction;
  wire         laneRequestSourceWire_7_bits_special = specialInstruction;
  wire [7:0]   dataInWritePipeVec_0;
  wire [7:0]   dataInWritePipeVec_1;
  wire [7:0]   dataInWritePipeVec_2;
  wire [7:0]   dataInWritePipeVec_3;
  wire [7:0]   dataInWritePipeVec_4;
  wire [7:0]   dataInWritePipeVec_5;
  wire [7:0]   dataInWritePipeVec_6;
  wire [7:0]   dataInWritePipeVec_7;
  wire [7:0]   dataInWritePipe = dataInWritePipeVec_0 | dataInWritePipeVec_1 | dataInWritePipeVec_2 | dataInWritePipeVec_3 | dataInWritePipeVec_4 | dataInWritePipeVec_5 | dataInWritePipeVec_6 | dataInWritePipeVec_7;
  wire         gatherNeedRead = requestRegDequeue_valid & requestReg_bits_decodeResult_gather & ~requestReg_bits_decodeResult_vtype;
  reg  [2:0]   slots_0_record_instructionIndex;
  reg          slots_0_record_isLoadStore;
  reg          slots_0_record_maskType;
  reg          slots_0_state_wLast;
  reg          slots_0_state_idle;
  reg          slots_0_state_wMaskUnitLast;
  reg          slots_0_state_wVRFWrite;
  reg          slots_0_state_sCommit;
  reg          slots_0_endTag_0;
  reg          slots_0_endTag_1;
  reg          slots_0_endTag_2;
  reg          slots_0_endTag_3;
  reg          slots_0_endTag_4;
  reg          slots_0_endTag_5;
  reg          slots_0_endTag_6;
  reg          slots_0_endTag_7;
  reg          slots_0_endTag_8;
  reg          slots_0_vxsat;
  wire [1:0]   slots_laneAndLSUFinish_lo_lo = {slots_0_endTag_1, slots_0_endTag_0};
  wire [1:0]   slots_laneAndLSUFinish_lo_hi = {slots_0_endTag_3, slots_0_endTag_2};
  wire [3:0]   slots_laneAndLSUFinish_lo = {slots_laneAndLSUFinish_lo_hi, slots_laneAndLSUFinish_lo_lo};
  wire [1:0]   slots_laneAndLSUFinish_hi_lo = {slots_0_endTag_5, slots_0_endTag_4};
  wire [1:0]   slots_laneAndLSUFinish_hi_hi_hi = {slots_0_endTag_8, slots_0_endTag_7};
  wire [2:0]   slots_laneAndLSUFinish_hi_hi = {slots_laneAndLSUFinish_hi_hi_hi, slots_0_endTag_6};
  wire [4:0]   slots_laneAndLSUFinish_hi = {slots_laneAndLSUFinish_hi_hi, slots_laneAndLSUFinish_hi_lo};
  wire         slots_laneAndLSUFinish = &{slots_laneAndLSUFinish_hi, slots_laneAndLSUFinish_lo};
  wire [7:0]   _GEN = {5'h0, slots_0_record_instructionIndex};
  wire         slots_v0WriteFinish = (8'h1 << _GEN & _tokenManager_v0WriteValid) == 8'h0;
  wire         slots_lsuFinished = |(8'h1 << _GEN & _lsu_lastReport);
  wire [7:0]   _slots_vxsatUpdate_T_1 = 8'h1 << _GEN;
  wire         slots_vxsatUpdate = |(_slots_vxsatUpdate_T_1[3:0] & vxsatReport);
  wire         slots_dataInWritePipeCheck = |(8'h1 << _GEN & dataInWritePipe);
  reg  [2:0]   slots_1_record_instructionIndex;
  reg          slots_1_record_isLoadStore;
  reg          slots_1_record_maskType;
  reg          slots_1_state_wLast;
  reg          slots_1_state_idle;
  reg          slots_1_state_wMaskUnitLast;
  reg          slots_1_state_wVRFWrite;
  reg          slots_1_state_sCommit;
  reg          slots_1_endTag_0;
  reg          slots_1_endTag_1;
  reg          slots_1_endTag_2;
  reg          slots_1_endTag_3;
  reg          slots_1_endTag_4;
  reg          slots_1_endTag_5;
  reg          slots_1_endTag_6;
  reg          slots_1_endTag_7;
  reg          slots_1_endTag_8;
  reg          slots_1_vxsat;
  wire [1:0]   slots_laneAndLSUFinish_lo_lo_1 = {slots_1_endTag_1, slots_1_endTag_0};
  wire [1:0]   slots_laneAndLSUFinish_lo_hi_1 = {slots_1_endTag_3, slots_1_endTag_2};
  wire [3:0]   slots_laneAndLSUFinish_lo_1 = {slots_laneAndLSUFinish_lo_hi_1, slots_laneAndLSUFinish_lo_lo_1};
  wire [1:0]   slots_laneAndLSUFinish_hi_lo_1 = {slots_1_endTag_5, slots_1_endTag_4};
  wire [1:0]   slots_laneAndLSUFinish_hi_hi_hi_1 = {slots_1_endTag_8, slots_1_endTag_7};
  wire [2:0]   slots_laneAndLSUFinish_hi_hi_1 = {slots_laneAndLSUFinish_hi_hi_hi_1, slots_1_endTag_6};
  wire [4:0]   slots_laneAndLSUFinish_hi_1 = {slots_laneAndLSUFinish_hi_hi_1, slots_laneAndLSUFinish_hi_lo_1};
  wire         slots_laneAndLSUFinish_1 = &{slots_laneAndLSUFinish_hi_1, slots_laneAndLSUFinish_lo_1};
  wire [7:0]   _GEN_0 = {5'h0, slots_1_record_instructionIndex};
  wire         slots_v0WriteFinish_1 = (8'h1 << _GEN_0 & _tokenManager_v0WriteValid) == 8'h0;
  wire         slots_lsuFinished_1 = |(8'h1 << _GEN_0 & _lsu_lastReport);
  wire [7:0]   _slots_vxsatUpdate_T_4 = 8'h1 << _GEN_0;
  wire         slots_vxsatUpdate_1 = |(_slots_vxsatUpdate_T_4[3:0] & vxsatReport);
  wire         slots_dataInWritePipeCheck_1 = |(8'h1 << _GEN_0 & dataInWritePipe);
  reg  [2:0]   slots_2_record_instructionIndex;
  reg          slots_2_record_isLoadStore;
  reg          slots_2_record_maskType;
  reg          slots_2_state_wLast;
  reg          slots_2_state_idle;
  reg          slots_2_state_wMaskUnitLast;
  reg          slots_2_state_wVRFWrite;
  reg          slots_2_state_sCommit;
  reg          slots_2_endTag_0;
  reg          slots_2_endTag_1;
  reg          slots_2_endTag_2;
  reg          slots_2_endTag_3;
  reg          slots_2_endTag_4;
  reg          slots_2_endTag_5;
  reg          slots_2_endTag_6;
  reg          slots_2_endTag_7;
  reg          slots_2_endTag_8;
  reg          slots_2_vxsat;
  wire [1:0]   slots_laneAndLSUFinish_lo_lo_2 = {slots_2_endTag_1, slots_2_endTag_0};
  wire [1:0]   slots_laneAndLSUFinish_lo_hi_2 = {slots_2_endTag_3, slots_2_endTag_2};
  wire [3:0]   slots_laneAndLSUFinish_lo_2 = {slots_laneAndLSUFinish_lo_hi_2, slots_laneAndLSUFinish_lo_lo_2};
  wire [1:0]   slots_laneAndLSUFinish_hi_lo_2 = {slots_2_endTag_5, slots_2_endTag_4};
  wire [1:0]   slots_laneAndLSUFinish_hi_hi_hi_2 = {slots_2_endTag_8, slots_2_endTag_7};
  wire [2:0]   slots_laneAndLSUFinish_hi_hi_2 = {slots_laneAndLSUFinish_hi_hi_hi_2, slots_2_endTag_6};
  wire [4:0]   slots_laneAndLSUFinish_hi_2 = {slots_laneAndLSUFinish_hi_hi_2, slots_laneAndLSUFinish_hi_lo_2};
  wire         slots_laneAndLSUFinish_2 = &{slots_laneAndLSUFinish_hi_2, slots_laneAndLSUFinish_lo_2};
  wire [7:0]   _GEN_1 = {5'h0, slots_2_record_instructionIndex};
  wire         slots_v0WriteFinish_2 = (8'h1 << _GEN_1 & _tokenManager_v0WriteValid) == 8'h0;
  wire         slots_lsuFinished_2 = |(8'h1 << _GEN_1 & _lsu_lastReport);
  wire [7:0]   _slots_vxsatUpdate_T_7 = 8'h1 << _GEN_1;
  wire         slots_vxsatUpdate_2 = |(_slots_vxsatUpdate_T_7[3:0] & vxsatReport);
  wire         slots_dataInWritePipeCheck_2 = |(8'h1 << _GEN_1 & dataInWritePipe);
  reg  [2:0]   slots_3_record_instructionIndex;
  reg          slots_3_record_isLoadStore;
  reg          slots_3_record_maskType;
  reg          slots_3_state_wLast;
  reg          slots_3_state_idle;
  reg          slots_3_state_wMaskUnitLast;
  reg          slots_3_state_wVRFWrite;
  reg          slots_3_state_sCommit;
  reg          slots_3_endTag_0;
  reg          slots_3_endTag_1;
  reg          slots_3_endTag_2;
  reg          slots_3_endTag_3;
  reg          slots_3_endTag_4;
  reg          slots_3_endTag_5;
  reg          slots_3_endTag_6;
  reg          slots_3_endTag_7;
  reg          slots_3_endTag_8;
  reg          slots_3_vxsat;
  wire [1:0]   slots_laneAndLSUFinish_lo_lo_3 = {slots_3_endTag_1, slots_3_endTag_0};
  wire [1:0]   slots_laneAndLSUFinish_lo_hi_3 = {slots_3_endTag_3, slots_3_endTag_2};
  wire [3:0]   slots_laneAndLSUFinish_lo_3 = {slots_laneAndLSUFinish_lo_hi_3, slots_laneAndLSUFinish_lo_lo_3};
  wire [1:0]   slots_laneAndLSUFinish_hi_lo_3 = {slots_3_endTag_5, slots_3_endTag_4};
  wire [1:0]   slots_laneAndLSUFinish_hi_hi_hi_3 = {slots_3_endTag_8, slots_3_endTag_7};
  wire [2:0]   slots_laneAndLSUFinish_hi_hi_3 = {slots_laneAndLSUFinish_hi_hi_hi_3, slots_3_endTag_6};
  wire [4:0]   slots_laneAndLSUFinish_hi_3 = {slots_laneAndLSUFinish_hi_hi_3, slots_laneAndLSUFinish_hi_lo_3};
  wire         slots_laneAndLSUFinish_3 = &{slots_laneAndLSUFinish_hi_3, slots_laneAndLSUFinish_lo_3};
  wire [7:0]   _GEN_2 = {5'h0, slots_3_record_instructionIndex};
  wire         slots_v0WriteFinish_3 = (8'h1 << _GEN_2 & _tokenManager_v0WriteValid) == 8'h0;
  wire         slots_lsuFinished_3 = |(8'h1 << _GEN_2 & _lsu_lastReport);
  wire [7:0]   _slots_vxsatUpdate_T_10 = 8'h1 << _GEN_2;
  wire         slots_vxsatUpdate_3 = |(_slots_vxsatUpdate_T_10[3:0] & vxsatReport);
  wire         slots_dataInWritePipeCheck_3 = |(8'h1 << _GEN_2 & dataInWritePipe);
  reg          slots_writeRD;
  reg  [4:0]   slots_vd;
  wire [4:0]   retire_rd_bits_rdAddress_0 = slots_vd;
  wire         lastSlotCommit;
  wire         retire_rd_valid_0 = lastSlotCommit & slots_writeRD;
  wire         tokenCheck;
  wire [2:0]   validSource_bits_instructionIndex = laneRequestSourceWire_0_bits_instructionIndex;
  wire         validSource_bits_decodeResult_specialSlot = laneRequestSourceWire_0_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_bits_decodeResult_topUop = laneRequestSourceWire_0_bits_decodeResult_topUop;
  wire         validSource_bits_decodeResult_popCount = laneRequestSourceWire_0_bits_decodeResult_popCount;
  wire         validSource_bits_decodeResult_ffo = laneRequestSourceWire_0_bits_decodeResult_ffo;
  wire         validSource_bits_decodeResult_average = laneRequestSourceWire_0_bits_decodeResult_average;
  wire         validSource_bits_decodeResult_reverse = laneRequestSourceWire_0_bits_decodeResult_reverse;
  wire         validSource_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_0_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_bits_decodeResult_scheduler = laneRequestSourceWire_0_bits_decodeResult_scheduler;
  wire         validSource_bits_decodeResult_sReadVD = laneRequestSourceWire_0_bits_decodeResult_sReadVD;
  wire         validSource_bits_decodeResult_vtype = laneRequestSourceWire_0_bits_decodeResult_vtype;
  wire         validSource_bits_decodeResult_sWrite = laneRequestSourceWire_0_bits_decodeResult_sWrite;
  wire         validSource_bits_decodeResult_crossRead = laneRequestSourceWire_0_bits_decodeResult_crossRead;
  wire         validSource_bits_decodeResult_crossWrite = laneRequestSourceWire_0_bits_decodeResult_crossWrite;
  wire         validSource_bits_decodeResult_maskUnit = laneRequestSourceWire_0_bits_decodeResult_maskUnit;
  wire         validSource_bits_decodeResult_special = laneRequestSourceWire_0_bits_decodeResult_special;
  wire         validSource_bits_decodeResult_saturate = laneRequestSourceWire_0_bits_decodeResult_saturate;
  wire         validSource_bits_decodeResult_vwmacc = laneRequestSourceWire_0_bits_decodeResult_vwmacc;
  wire         validSource_bits_decodeResult_readOnly = laneRequestSourceWire_0_bits_decodeResult_readOnly;
  wire         validSource_bits_decodeResult_maskSource = laneRequestSourceWire_0_bits_decodeResult_maskSource;
  wire         validSource_bits_decodeResult_maskDestination = laneRequestSourceWire_0_bits_decodeResult_maskDestination;
  wire         validSource_bits_decodeResult_maskLogic = laneRequestSourceWire_0_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_bits_decodeResult_uop = laneRequestSourceWire_0_bits_decodeResult_uop;
  wire         validSource_bits_decodeResult_iota = laneRequestSourceWire_0_bits_decodeResult_iota;
  wire         validSource_bits_decodeResult_mv = laneRequestSourceWire_0_bits_decodeResult_mv;
  wire         validSource_bits_decodeResult_extend = laneRequestSourceWire_0_bits_decodeResult_extend;
  wire         validSource_bits_decodeResult_unOrderWrite = laneRequestSourceWire_0_bits_decodeResult_unOrderWrite;
  wire         validSource_bits_decodeResult_compress = laneRequestSourceWire_0_bits_decodeResult_compress;
  wire         validSource_bits_decodeResult_gather16 = laneRequestSourceWire_0_bits_decodeResult_gather16;
  wire         validSource_bits_decodeResult_gather = laneRequestSourceWire_0_bits_decodeResult_gather;
  wire         validSource_bits_decodeResult_slid = laneRequestSourceWire_0_bits_decodeResult_slid;
  wire         validSource_bits_decodeResult_targetRd = laneRequestSourceWire_0_bits_decodeResult_targetRd;
  wire         validSource_bits_decodeResult_widenReduce = laneRequestSourceWire_0_bits_decodeResult_widenReduce;
  wire         validSource_bits_decodeResult_red = laneRequestSourceWire_0_bits_decodeResult_red;
  wire         validSource_bits_decodeResult_nr = laneRequestSourceWire_0_bits_decodeResult_nr;
  wire         validSource_bits_decodeResult_itype = laneRequestSourceWire_0_bits_decodeResult_itype;
  wire         validSource_bits_decodeResult_unsigned1 = laneRequestSourceWire_0_bits_decodeResult_unsigned1;
  wire         validSource_bits_decodeResult_unsigned0 = laneRequestSourceWire_0_bits_decodeResult_unsigned0;
  wire         validSource_bits_decodeResult_other = laneRequestSourceWire_0_bits_decodeResult_other;
  wire         validSource_bits_decodeResult_multiCycle = laneRequestSourceWire_0_bits_decodeResult_multiCycle;
  wire         validSource_bits_decodeResult_divider = laneRequestSourceWire_0_bits_decodeResult_divider;
  wire         validSource_bits_decodeResult_multiplier = laneRequestSourceWire_0_bits_decodeResult_multiplier;
  wire         validSource_bits_decodeResult_shift = laneRequestSourceWire_0_bits_decodeResult_shift;
  wire         validSource_bits_decodeResult_adder = laneRequestSourceWire_0_bits_decodeResult_adder;
  wire         validSource_bits_decodeResult_logic = laneRequestSourceWire_0_bits_decodeResult_logic;
  wire         validSource_bits_loadStore = laneRequestSourceWire_0_bits_loadStore;
  wire         validSource_bits_issueInst = laneRequestSourceWire_0_bits_issueInst;
  wire         validSource_bits_store = laneRequestSourceWire_0_bits_store;
  wire         validSource_bits_special = laneRequestSourceWire_0_bits_special;
  wire         validSource_bits_lsWholeReg = laneRequestSourceWire_0_bits_lsWholeReg;
  wire [4:0]   validSource_bits_vs1 = laneRequestSourceWire_0_bits_vs1;
  wire [4:0]   validSource_bits_vs2 = laneRequestSourceWire_0_bits_vs2;
  wire [4:0]   validSource_bits_vd = laneRequestSourceWire_0_bits_vd;
  wire [1:0]   validSource_bits_loadStoreEEW = laneRequestSourceWire_0_bits_loadStoreEEW;
  wire         validSource_bits_mask = laneRequestSourceWire_0_bits_mask;
  wire [2:0]   validSource_bits_segment = laneRequestSourceWire_0_bits_segment;
  wire [31:0]  source1Select;
  wire [31:0]  validSource_bits_readFromScalar = laneRequestSourceWire_0_bits_readFromScalar;
  wire [11:0]  validSource_bits_csrInterface_vl = laneRequestSourceWire_0_bits_csrInterface_vl;
  wire [11:0]  validSource_bits_csrInterface_vStart = laneRequestSourceWire_0_bits_csrInterface_vStart;
  wire [2:0]   validSource_bits_csrInterface_vlmul = laneRequestSourceWire_0_bits_csrInterface_vlmul;
  wire [1:0]   validSource_bits_csrInterface_vSew = laneRequestSourceWire_0_bits_csrInterface_vSew;
  wire [1:0]   validSource_bits_csrInterface_vxrm = laneRequestSourceWire_0_bits_csrInterface_vxrm;
  wire         validSource_bits_csrInterface_vta = laneRequestSourceWire_0_bits_csrInterface_vta;
  wire         validSource_bits_csrInterface_vma = laneRequestSourceWire_0_bits_csrInterface_vma;
  wire         tokenCheck_1;
  wire [2:0]   validSource_1_bits_instructionIndex = laneRequestSourceWire_1_bits_instructionIndex;
  wire         validSource_1_bits_decodeResult_specialSlot = laneRequestSourceWire_1_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_1_bits_decodeResult_topUop = laneRequestSourceWire_1_bits_decodeResult_topUop;
  wire         validSource_1_bits_decodeResult_popCount = laneRequestSourceWire_1_bits_decodeResult_popCount;
  wire         validSource_1_bits_decodeResult_ffo = laneRequestSourceWire_1_bits_decodeResult_ffo;
  wire         validSource_1_bits_decodeResult_average = laneRequestSourceWire_1_bits_decodeResult_average;
  wire         validSource_1_bits_decodeResult_reverse = laneRequestSourceWire_1_bits_decodeResult_reverse;
  wire         validSource_1_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_1_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_1_bits_decodeResult_scheduler = laneRequestSourceWire_1_bits_decodeResult_scheduler;
  wire         validSource_1_bits_decodeResult_sReadVD = laneRequestSourceWire_1_bits_decodeResult_sReadVD;
  wire         validSource_1_bits_decodeResult_vtype = laneRequestSourceWire_1_bits_decodeResult_vtype;
  wire         validSource_1_bits_decodeResult_sWrite = laneRequestSourceWire_1_bits_decodeResult_sWrite;
  wire         validSource_1_bits_decodeResult_crossRead = laneRequestSourceWire_1_bits_decodeResult_crossRead;
  wire         validSource_1_bits_decodeResult_crossWrite = laneRequestSourceWire_1_bits_decodeResult_crossWrite;
  wire         validSource_1_bits_decodeResult_maskUnit = laneRequestSourceWire_1_bits_decodeResult_maskUnit;
  wire         validSource_1_bits_decodeResult_special = laneRequestSourceWire_1_bits_decodeResult_special;
  wire         validSource_1_bits_decodeResult_saturate = laneRequestSourceWire_1_bits_decodeResult_saturate;
  wire         validSource_1_bits_decodeResult_vwmacc = laneRequestSourceWire_1_bits_decodeResult_vwmacc;
  wire         validSource_1_bits_decodeResult_readOnly = laneRequestSourceWire_1_bits_decodeResult_readOnly;
  wire         validSource_1_bits_decodeResult_maskSource = laneRequestSourceWire_1_bits_decodeResult_maskSource;
  wire         validSource_1_bits_decodeResult_maskDestination = laneRequestSourceWire_1_bits_decodeResult_maskDestination;
  wire         validSource_1_bits_decodeResult_maskLogic = laneRequestSourceWire_1_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_1_bits_decodeResult_uop = laneRequestSourceWire_1_bits_decodeResult_uop;
  wire         validSource_1_bits_decodeResult_iota = laneRequestSourceWire_1_bits_decodeResult_iota;
  wire         validSource_1_bits_decodeResult_mv = laneRequestSourceWire_1_bits_decodeResult_mv;
  wire         validSource_1_bits_decodeResult_extend = laneRequestSourceWire_1_bits_decodeResult_extend;
  wire         validSource_1_bits_decodeResult_unOrderWrite = laneRequestSourceWire_1_bits_decodeResult_unOrderWrite;
  wire         validSource_1_bits_decodeResult_compress = laneRequestSourceWire_1_bits_decodeResult_compress;
  wire         validSource_1_bits_decodeResult_gather16 = laneRequestSourceWire_1_bits_decodeResult_gather16;
  wire         validSource_1_bits_decodeResult_gather = laneRequestSourceWire_1_bits_decodeResult_gather;
  wire         validSource_1_bits_decodeResult_slid = laneRequestSourceWire_1_bits_decodeResult_slid;
  wire         validSource_1_bits_decodeResult_targetRd = laneRequestSourceWire_1_bits_decodeResult_targetRd;
  wire         validSource_1_bits_decodeResult_widenReduce = laneRequestSourceWire_1_bits_decodeResult_widenReduce;
  wire         validSource_1_bits_decodeResult_red = laneRequestSourceWire_1_bits_decodeResult_red;
  wire         validSource_1_bits_decodeResult_nr = laneRequestSourceWire_1_bits_decodeResult_nr;
  wire         validSource_1_bits_decodeResult_itype = laneRequestSourceWire_1_bits_decodeResult_itype;
  wire         validSource_1_bits_decodeResult_unsigned1 = laneRequestSourceWire_1_bits_decodeResult_unsigned1;
  wire         validSource_1_bits_decodeResult_unsigned0 = laneRequestSourceWire_1_bits_decodeResult_unsigned0;
  wire         validSource_1_bits_decodeResult_other = laneRequestSourceWire_1_bits_decodeResult_other;
  wire         validSource_1_bits_decodeResult_multiCycle = laneRequestSourceWire_1_bits_decodeResult_multiCycle;
  wire         validSource_1_bits_decodeResult_divider = laneRequestSourceWire_1_bits_decodeResult_divider;
  wire         validSource_1_bits_decodeResult_multiplier = laneRequestSourceWire_1_bits_decodeResult_multiplier;
  wire         validSource_1_bits_decodeResult_shift = laneRequestSourceWire_1_bits_decodeResult_shift;
  wire         validSource_1_bits_decodeResult_adder = laneRequestSourceWire_1_bits_decodeResult_adder;
  wire         validSource_1_bits_decodeResult_logic = laneRequestSourceWire_1_bits_decodeResult_logic;
  wire         validSource_1_bits_loadStore = laneRequestSourceWire_1_bits_loadStore;
  wire         validSource_1_bits_issueInst = laneRequestSourceWire_1_bits_issueInst;
  wire         validSource_1_bits_store = laneRequestSourceWire_1_bits_store;
  wire         validSource_1_bits_special = laneRequestSourceWire_1_bits_special;
  wire         validSource_1_bits_lsWholeReg = laneRequestSourceWire_1_bits_lsWholeReg;
  wire [4:0]   validSource_1_bits_vs1 = laneRequestSourceWire_1_bits_vs1;
  wire [4:0]   validSource_1_bits_vs2 = laneRequestSourceWire_1_bits_vs2;
  wire [4:0]   validSource_1_bits_vd = laneRequestSourceWire_1_bits_vd;
  wire [1:0]   validSource_1_bits_loadStoreEEW = laneRequestSourceWire_1_bits_loadStoreEEW;
  wire         validSource_1_bits_mask = laneRequestSourceWire_1_bits_mask;
  wire [2:0]   validSource_1_bits_segment = laneRequestSourceWire_1_bits_segment;
  wire [31:0]  validSource_1_bits_readFromScalar = laneRequestSourceWire_1_bits_readFromScalar;
  wire [11:0]  validSource_1_bits_csrInterface_vl = laneRequestSourceWire_1_bits_csrInterface_vl;
  wire [11:0]  validSource_1_bits_csrInterface_vStart = laneRequestSourceWire_1_bits_csrInterface_vStart;
  wire [2:0]   validSource_1_bits_csrInterface_vlmul = laneRequestSourceWire_1_bits_csrInterface_vlmul;
  wire [1:0]   validSource_1_bits_csrInterface_vSew = laneRequestSourceWire_1_bits_csrInterface_vSew;
  wire [1:0]   validSource_1_bits_csrInterface_vxrm = laneRequestSourceWire_1_bits_csrInterface_vxrm;
  wire         validSource_1_bits_csrInterface_vta = laneRequestSourceWire_1_bits_csrInterface_vta;
  wire         validSource_1_bits_csrInterface_vma = laneRequestSourceWire_1_bits_csrInterface_vma;
  wire         tokenCheck_2;
  wire [2:0]   validSource_2_bits_instructionIndex = laneRequestSourceWire_2_bits_instructionIndex;
  wire         validSource_2_bits_decodeResult_specialSlot = laneRequestSourceWire_2_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_2_bits_decodeResult_topUop = laneRequestSourceWire_2_bits_decodeResult_topUop;
  wire         validSource_2_bits_decodeResult_popCount = laneRequestSourceWire_2_bits_decodeResult_popCount;
  wire         validSource_2_bits_decodeResult_ffo = laneRequestSourceWire_2_bits_decodeResult_ffo;
  wire         validSource_2_bits_decodeResult_average = laneRequestSourceWire_2_bits_decodeResult_average;
  wire         validSource_2_bits_decodeResult_reverse = laneRequestSourceWire_2_bits_decodeResult_reverse;
  wire         validSource_2_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_2_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_2_bits_decodeResult_scheduler = laneRequestSourceWire_2_bits_decodeResult_scheduler;
  wire         validSource_2_bits_decodeResult_sReadVD = laneRequestSourceWire_2_bits_decodeResult_sReadVD;
  wire         validSource_2_bits_decodeResult_vtype = laneRequestSourceWire_2_bits_decodeResult_vtype;
  wire         validSource_2_bits_decodeResult_sWrite = laneRequestSourceWire_2_bits_decodeResult_sWrite;
  wire         validSource_2_bits_decodeResult_crossRead = laneRequestSourceWire_2_bits_decodeResult_crossRead;
  wire         validSource_2_bits_decodeResult_crossWrite = laneRequestSourceWire_2_bits_decodeResult_crossWrite;
  wire         validSource_2_bits_decodeResult_maskUnit = laneRequestSourceWire_2_bits_decodeResult_maskUnit;
  wire         validSource_2_bits_decodeResult_special = laneRequestSourceWire_2_bits_decodeResult_special;
  wire         validSource_2_bits_decodeResult_saturate = laneRequestSourceWire_2_bits_decodeResult_saturate;
  wire         validSource_2_bits_decodeResult_vwmacc = laneRequestSourceWire_2_bits_decodeResult_vwmacc;
  wire         validSource_2_bits_decodeResult_readOnly = laneRequestSourceWire_2_bits_decodeResult_readOnly;
  wire         validSource_2_bits_decodeResult_maskSource = laneRequestSourceWire_2_bits_decodeResult_maskSource;
  wire         validSource_2_bits_decodeResult_maskDestination = laneRequestSourceWire_2_bits_decodeResult_maskDestination;
  wire         validSource_2_bits_decodeResult_maskLogic = laneRequestSourceWire_2_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_2_bits_decodeResult_uop = laneRequestSourceWire_2_bits_decodeResult_uop;
  wire         validSource_2_bits_decodeResult_iota = laneRequestSourceWire_2_bits_decodeResult_iota;
  wire         validSource_2_bits_decodeResult_mv = laneRequestSourceWire_2_bits_decodeResult_mv;
  wire         validSource_2_bits_decodeResult_extend = laneRequestSourceWire_2_bits_decodeResult_extend;
  wire         validSource_2_bits_decodeResult_unOrderWrite = laneRequestSourceWire_2_bits_decodeResult_unOrderWrite;
  wire         validSource_2_bits_decodeResult_compress = laneRequestSourceWire_2_bits_decodeResult_compress;
  wire         validSource_2_bits_decodeResult_gather16 = laneRequestSourceWire_2_bits_decodeResult_gather16;
  wire         validSource_2_bits_decodeResult_gather = laneRequestSourceWire_2_bits_decodeResult_gather;
  wire         validSource_2_bits_decodeResult_slid = laneRequestSourceWire_2_bits_decodeResult_slid;
  wire         validSource_2_bits_decodeResult_targetRd = laneRequestSourceWire_2_bits_decodeResult_targetRd;
  wire         validSource_2_bits_decodeResult_widenReduce = laneRequestSourceWire_2_bits_decodeResult_widenReduce;
  wire         validSource_2_bits_decodeResult_red = laneRequestSourceWire_2_bits_decodeResult_red;
  wire         validSource_2_bits_decodeResult_nr = laneRequestSourceWire_2_bits_decodeResult_nr;
  wire         validSource_2_bits_decodeResult_itype = laneRequestSourceWire_2_bits_decodeResult_itype;
  wire         validSource_2_bits_decodeResult_unsigned1 = laneRequestSourceWire_2_bits_decodeResult_unsigned1;
  wire         validSource_2_bits_decodeResult_unsigned0 = laneRequestSourceWire_2_bits_decodeResult_unsigned0;
  wire         validSource_2_bits_decodeResult_other = laneRequestSourceWire_2_bits_decodeResult_other;
  wire         validSource_2_bits_decodeResult_multiCycle = laneRequestSourceWire_2_bits_decodeResult_multiCycle;
  wire         validSource_2_bits_decodeResult_divider = laneRequestSourceWire_2_bits_decodeResult_divider;
  wire         validSource_2_bits_decodeResult_multiplier = laneRequestSourceWire_2_bits_decodeResult_multiplier;
  wire         validSource_2_bits_decodeResult_shift = laneRequestSourceWire_2_bits_decodeResult_shift;
  wire         validSource_2_bits_decodeResult_adder = laneRequestSourceWire_2_bits_decodeResult_adder;
  wire         validSource_2_bits_decodeResult_logic = laneRequestSourceWire_2_bits_decodeResult_logic;
  wire         validSource_2_bits_loadStore = laneRequestSourceWire_2_bits_loadStore;
  wire         validSource_2_bits_issueInst = laneRequestSourceWire_2_bits_issueInst;
  wire         validSource_2_bits_store = laneRequestSourceWire_2_bits_store;
  wire         validSource_2_bits_special = laneRequestSourceWire_2_bits_special;
  wire         validSource_2_bits_lsWholeReg = laneRequestSourceWire_2_bits_lsWholeReg;
  wire [4:0]   validSource_2_bits_vs1 = laneRequestSourceWire_2_bits_vs1;
  wire [4:0]   validSource_2_bits_vs2 = laneRequestSourceWire_2_bits_vs2;
  wire [4:0]   validSource_2_bits_vd = laneRequestSourceWire_2_bits_vd;
  wire [1:0]   validSource_2_bits_loadStoreEEW = laneRequestSourceWire_2_bits_loadStoreEEW;
  wire         validSource_2_bits_mask = laneRequestSourceWire_2_bits_mask;
  wire [2:0]   validSource_2_bits_segment = laneRequestSourceWire_2_bits_segment;
  wire [31:0]  validSource_2_bits_readFromScalar = laneRequestSourceWire_2_bits_readFromScalar;
  wire [11:0]  validSource_2_bits_csrInterface_vl = laneRequestSourceWire_2_bits_csrInterface_vl;
  wire [11:0]  validSource_2_bits_csrInterface_vStart = laneRequestSourceWire_2_bits_csrInterface_vStart;
  wire [2:0]   validSource_2_bits_csrInterface_vlmul = laneRequestSourceWire_2_bits_csrInterface_vlmul;
  wire [1:0]   validSource_2_bits_csrInterface_vSew = laneRequestSourceWire_2_bits_csrInterface_vSew;
  wire [1:0]   validSource_2_bits_csrInterface_vxrm = laneRequestSourceWire_2_bits_csrInterface_vxrm;
  wire         validSource_2_bits_csrInterface_vta = laneRequestSourceWire_2_bits_csrInterface_vta;
  wire         validSource_2_bits_csrInterface_vma = laneRequestSourceWire_2_bits_csrInterface_vma;
  wire         tokenCheck_3;
  wire [2:0]   validSource_3_bits_instructionIndex = laneRequestSourceWire_3_bits_instructionIndex;
  wire         validSource_3_bits_decodeResult_specialSlot = laneRequestSourceWire_3_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_3_bits_decodeResult_topUop = laneRequestSourceWire_3_bits_decodeResult_topUop;
  wire         validSource_3_bits_decodeResult_popCount = laneRequestSourceWire_3_bits_decodeResult_popCount;
  wire         validSource_3_bits_decodeResult_ffo = laneRequestSourceWire_3_bits_decodeResult_ffo;
  wire         validSource_3_bits_decodeResult_average = laneRequestSourceWire_3_bits_decodeResult_average;
  wire         validSource_3_bits_decodeResult_reverse = laneRequestSourceWire_3_bits_decodeResult_reverse;
  wire         validSource_3_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_3_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_3_bits_decodeResult_scheduler = laneRequestSourceWire_3_bits_decodeResult_scheduler;
  wire         validSource_3_bits_decodeResult_sReadVD = laneRequestSourceWire_3_bits_decodeResult_sReadVD;
  wire         validSource_3_bits_decodeResult_vtype = laneRequestSourceWire_3_bits_decodeResult_vtype;
  wire         validSource_3_bits_decodeResult_sWrite = laneRequestSourceWire_3_bits_decodeResult_sWrite;
  wire         validSource_3_bits_decodeResult_crossRead = laneRequestSourceWire_3_bits_decodeResult_crossRead;
  wire         validSource_3_bits_decodeResult_crossWrite = laneRequestSourceWire_3_bits_decodeResult_crossWrite;
  wire         validSource_3_bits_decodeResult_maskUnit = laneRequestSourceWire_3_bits_decodeResult_maskUnit;
  wire         validSource_3_bits_decodeResult_special = laneRequestSourceWire_3_bits_decodeResult_special;
  wire         validSource_3_bits_decodeResult_saturate = laneRequestSourceWire_3_bits_decodeResult_saturate;
  wire         validSource_3_bits_decodeResult_vwmacc = laneRequestSourceWire_3_bits_decodeResult_vwmacc;
  wire         validSource_3_bits_decodeResult_readOnly = laneRequestSourceWire_3_bits_decodeResult_readOnly;
  wire         validSource_3_bits_decodeResult_maskSource = laneRequestSourceWire_3_bits_decodeResult_maskSource;
  wire         validSource_3_bits_decodeResult_maskDestination = laneRequestSourceWire_3_bits_decodeResult_maskDestination;
  wire         validSource_3_bits_decodeResult_maskLogic = laneRequestSourceWire_3_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_3_bits_decodeResult_uop = laneRequestSourceWire_3_bits_decodeResult_uop;
  wire         validSource_3_bits_decodeResult_iota = laneRequestSourceWire_3_bits_decodeResult_iota;
  wire         validSource_3_bits_decodeResult_mv = laneRequestSourceWire_3_bits_decodeResult_mv;
  wire         validSource_3_bits_decodeResult_extend = laneRequestSourceWire_3_bits_decodeResult_extend;
  wire         validSource_3_bits_decodeResult_unOrderWrite = laneRequestSourceWire_3_bits_decodeResult_unOrderWrite;
  wire         validSource_3_bits_decodeResult_compress = laneRequestSourceWire_3_bits_decodeResult_compress;
  wire         validSource_3_bits_decodeResult_gather16 = laneRequestSourceWire_3_bits_decodeResult_gather16;
  wire         validSource_3_bits_decodeResult_gather = laneRequestSourceWire_3_bits_decodeResult_gather;
  wire         validSource_3_bits_decodeResult_slid = laneRequestSourceWire_3_bits_decodeResult_slid;
  wire         validSource_3_bits_decodeResult_targetRd = laneRequestSourceWire_3_bits_decodeResult_targetRd;
  wire         validSource_3_bits_decodeResult_widenReduce = laneRequestSourceWire_3_bits_decodeResult_widenReduce;
  wire         validSource_3_bits_decodeResult_red = laneRequestSourceWire_3_bits_decodeResult_red;
  wire         validSource_3_bits_decodeResult_nr = laneRequestSourceWire_3_bits_decodeResult_nr;
  wire         validSource_3_bits_decodeResult_itype = laneRequestSourceWire_3_bits_decodeResult_itype;
  wire         validSource_3_bits_decodeResult_unsigned1 = laneRequestSourceWire_3_bits_decodeResult_unsigned1;
  wire         validSource_3_bits_decodeResult_unsigned0 = laneRequestSourceWire_3_bits_decodeResult_unsigned0;
  wire         validSource_3_bits_decodeResult_other = laneRequestSourceWire_3_bits_decodeResult_other;
  wire         validSource_3_bits_decodeResult_multiCycle = laneRequestSourceWire_3_bits_decodeResult_multiCycle;
  wire         validSource_3_bits_decodeResult_divider = laneRequestSourceWire_3_bits_decodeResult_divider;
  wire         validSource_3_bits_decodeResult_multiplier = laneRequestSourceWire_3_bits_decodeResult_multiplier;
  wire         validSource_3_bits_decodeResult_shift = laneRequestSourceWire_3_bits_decodeResult_shift;
  wire         validSource_3_bits_decodeResult_adder = laneRequestSourceWire_3_bits_decodeResult_adder;
  wire         validSource_3_bits_decodeResult_logic = laneRequestSourceWire_3_bits_decodeResult_logic;
  wire         validSource_3_bits_loadStore = laneRequestSourceWire_3_bits_loadStore;
  wire         validSource_3_bits_issueInst = laneRequestSourceWire_3_bits_issueInst;
  wire         validSource_3_bits_store = laneRequestSourceWire_3_bits_store;
  wire         validSource_3_bits_special = laneRequestSourceWire_3_bits_special;
  wire         validSource_3_bits_lsWholeReg = laneRequestSourceWire_3_bits_lsWholeReg;
  wire [4:0]   validSource_3_bits_vs1 = laneRequestSourceWire_3_bits_vs1;
  wire [4:0]   validSource_3_bits_vs2 = laneRequestSourceWire_3_bits_vs2;
  wire [4:0]   validSource_3_bits_vd = laneRequestSourceWire_3_bits_vd;
  wire [1:0]   validSource_3_bits_loadStoreEEW = laneRequestSourceWire_3_bits_loadStoreEEW;
  wire         validSource_3_bits_mask = laneRequestSourceWire_3_bits_mask;
  wire [2:0]   validSource_3_bits_segment = laneRequestSourceWire_3_bits_segment;
  wire [31:0]  validSource_3_bits_readFromScalar = laneRequestSourceWire_3_bits_readFromScalar;
  wire [11:0]  validSource_3_bits_csrInterface_vl = laneRequestSourceWire_3_bits_csrInterface_vl;
  wire [11:0]  validSource_3_bits_csrInterface_vStart = laneRequestSourceWire_3_bits_csrInterface_vStart;
  wire [2:0]   validSource_3_bits_csrInterface_vlmul = laneRequestSourceWire_3_bits_csrInterface_vlmul;
  wire [1:0]   validSource_3_bits_csrInterface_vSew = laneRequestSourceWire_3_bits_csrInterface_vSew;
  wire [1:0]   validSource_3_bits_csrInterface_vxrm = laneRequestSourceWire_3_bits_csrInterface_vxrm;
  wire         validSource_3_bits_csrInterface_vta = laneRequestSourceWire_3_bits_csrInterface_vta;
  wire         validSource_3_bits_csrInterface_vma = laneRequestSourceWire_3_bits_csrInterface_vma;
  wire         tokenCheck_4;
  wire [2:0]   validSource_4_bits_instructionIndex = laneRequestSourceWire_4_bits_instructionIndex;
  wire         validSource_4_bits_decodeResult_specialSlot = laneRequestSourceWire_4_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_4_bits_decodeResult_topUop = laneRequestSourceWire_4_bits_decodeResult_topUop;
  wire         validSource_4_bits_decodeResult_popCount = laneRequestSourceWire_4_bits_decodeResult_popCount;
  wire         validSource_4_bits_decodeResult_ffo = laneRequestSourceWire_4_bits_decodeResult_ffo;
  wire         validSource_4_bits_decodeResult_average = laneRequestSourceWire_4_bits_decodeResult_average;
  wire         validSource_4_bits_decodeResult_reverse = laneRequestSourceWire_4_bits_decodeResult_reverse;
  wire         validSource_4_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_4_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_4_bits_decodeResult_scheduler = laneRequestSourceWire_4_bits_decodeResult_scheduler;
  wire         validSource_4_bits_decodeResult_sReadVD = laneRequestSourceWire_4_bits_decodeResult_sReadVD;
  wire         validSource_4_bits_decodeResult_vtype = laneRequestSourceWire_4_bits_decodeResult_vtype;
  wire         validSource_4_bits_decodeResult_sWrite = laneRequestSourceWire_4_bits_decodeResult_sWrite;
  wire         validSource_4_bits_decodeResult_crossRead = laneRequestSourceWire_4_bits_decodeResult_crossRead;
  wire         validSource_4_bits_decodeResult_crossWrite = laneRequestSourceWire_4_bits_decodeResult_crossWrite;
  wire         validSource_4_bits_decodeResult_maskUnit = laneRequestSourceWire_4_bits_decodeResult_maskUnit;
  wire         validSource_4_bits_decodeResult_special = laneRequestSourceWire_4_bits_decodeResult_special;
  wire         validSource_4_bits_decodeResult_saturate = laneRequestSourceWire_4_bits_decodeResult_saturate;
  wire         validSource_4_bits_decodeResult_vwmacc = laneRequestSourceWire_4_bits_decodeResult_vwmacc;
  wire         validSource_4_bits_decodeResult_readOnly = laneRequestSourceWire_4_bits_decodeResult_readOnly;
  wire         validSource_4_bits_decodeResult_maskSource = laneRequestSourceWire_4_bits_decodeResult_maskSource;
  wire         validSource_4_bits_decodeResult_maskDestination = laneRequestSourceWire_4_bits_decodeResult_maskDestination;
  wire         validSource_4_bits_decodeResult_maskLogic = laneRequestSourceWire_4_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_4_bits_decodeResult_uop = laneRequestSourceWire_4_bits_decodeResult_uop;
  wire         validSource_4_bits_decodeResult_iota = laneRequestSourceWire_4_bits_decodeResult_iota;
  wire         validSource_4_bits_decodeResult_mv = laneRequestSourceWire_4_bits_decodeResult_mv;
  wire         validSource_4_bits_decodeResult_extend = laneRequestSourceWire_4_bits_decodeResult_extend;
  wire         validSource_4_bits_decodeResult_unOrderWrite = laneRequestSourceWire_4_bits_decodeResult_unOrderWrite;
  wire         validSource_4_bits_decodeResult_compress = laneRequestSourceWire_4_bits_decodeResult_compress;
  wire         validSource_4_bits_decodeResult_gather16 = laneRequestSourceWire_4_bits_decodeResult_gather16;
  wire         validSource_4_bits_decodeResult_gather = laneRequestSourceWire_4_bits_decodeResult_gather;
  wire         validSource_4_bits_decodeResult_slid = laneRequestSourceWire_4_bits_decodeResult_slid;
  wire         validSource_4_bits_decodeResult_targetRd = laneRequestSourceWire_4_bits_decodeResult_targetRd;
  wire         validSource_4_bits_decodeResult_widenReduce = laneRequestSourceWire_4_bits_decodeResult_widenReduce;
  wire         validSource_4_bits_decodeResult_red = laneRequestSourceWire_4_bits_decodeResult_red;
  wire         validSource_4_bits_decodeResult_nr = laneRequestSourceWire_4_bits_decodeResult_nr;
  wire         validSource_4_bits_decodeResult_itype = laneRequestSourceWire_4_bits_decodeResult_itype;
  wire         validSource_4_bits_decodeResult_unsigned1 = laneRequestSourceWire_4_bits_decodeResult_unsigned1;
  wire         validSource_4_bits_decodeResult_unsigned0 = laneRequestSourceWire_4_bits_decodeResult_unsigned0;
  wire         validSource_4_bits_decodeResult_other = laneRequestSourceWire_4_bits_decodeResult_other;
  wire         validSource_4_bits_decodeResult_multiCycle = laneRequestSourceWire_4_bits_decodeResult_multiCycle;
  wire         validSource_4_bits_decodeResult_divider = laneRequestSourceWire_4_bits_decodeResult_divider;
  wire         validSource_4_bits_decodeResult_multiplier = laneRequestSourceWire_4_bits_decodeResult_multiplier;
  wire         validSource_4_bits_decodeResult_shift = laneRequestSourceWire_4_bits_decodeResult_shift;
  wire         validSource_4_bits_decodeResult_adder = laneRequestSourceWire_4_bits_decodeResult_adder;
  wire         validSource_4_bits_decodeResult_logic = laneRequestSourceWire_4_bits_decodeResult_logic;
  wire         validSource_4_bits_loadStore = laneRequestSourceWire_4_bits_loadStore;
  wire         validSource_4_bits_issueInst = laneRequestSourceWire_4_bits_issueInst;
  wire         validSource_4_bits_store = laneRequestSourceWire_4_bits_store;
  wire         validSource_4_bits_special = laneRequestSourceWire_4_bits_special;
  wire         validSource_4_bits_lsWholeReg = laneRequestSourceWire_4_bits_lsWholeReg;
  wire [4:0]   validSource_4_bits_vs1 = laneRequestSourceWire_4_bits_vs1;
  wire [4:0]   validSource_4_bits_vs2 = laneRequestSourceWire_4_bits_vs2;
  wire [4:0]   validSource_4_bits_vd = laneRequestSourceWire_4_bits_vd;
  wire [1:0]   validSource_4_bits_loadStoreEEW = laneRequestSourceWire_4_bits_loadStoreEEW;
  wire         validSource_4_bits_mask = laneRequestSourceWire_4_bits_mask;
  wire [2:0]   validSource_4_bits_segment = laneRequestSourceWire_4_bits_segment;
  wire [31:0]  validSource_4_bits_readFromScalar = laneRequestSourceWire_4_bits_readFromScalar;
  wire [11:0]  validSource_4_bits_csrInterface_vl = laneRequestSourceWire_4_bits_csrInterface_vl;
  wire [11:0]  validSource_4_bits_csrInterface_vStart = laneRequestSourceWire_4_bits_csrInterface_vStart;
  wire [2:0]   validSource_4_bits_csrInterface_vlmul = laneRequestSourceWire_4_bits_csrInterface_vlmul;
  wire [1:0]   validSource_4_bits_csrInterface_vSew = laneRequestSourceWire_4_bits_csrInterface_vSew;
  wire [1:0]   validSource_4_bits_csrInterface_vxrm = laneRequestSourceWire_4_bits_csrInterface_vxrm;
  wire         validSource_4_bits_csrInterface_vta = laneRequestSourceWire_4_bits_csrInterface_vta;
  wire         validSource_4_bits_csrInterface_vma = laneRequestSourceWire_4_bits_csrInterface_vma;
  wire         tokenCheck_5;
  wire [2:0]   validSource_5_bits_instructionIndex = laneRequestSourceWire_5_bits_instructionIndex;
  wire         validSource_5_bits_decodeResult_specialSlot = laneRequestSourceWire_5_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_5_bits_decodeResult_topUop = laneRequestSourceWire_5_bits_decodeResult_topUop;
  wire         validSource_5_bits_decodeResult_popCount = laneRequestSourceWire_5_bits_decodeResult_popCount;
  wire         validSource_5_bits_decodeResult_ffo = laneRequestSourceWire_5_bits_decodeResult_ffo;
  wire         validSource_5_bits_decodeResult_average = laneRequestSourceWire_5_bits_decodeResult_average;
  wire         validSource_5_bits_decodeResult_reverse = laneRequestSourceWire_5_bits_decodeResult_reverse;
  wire         validSource_5_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_5_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_5_bits_decodeResult_scheduler = laneRequestSourceWire_5_bits_decodeResult_scheduler;
  wire         validSource_5_bits_decodeResult_sReadVD = laneRequestSourceWire_5_bits_decodeResult_sReadVD;
  wire         validSource_5_bits_decodeResult_vtype = laneRequestSourceWire_5_bits_decodeResult_vtype;
  wire         validSource_5_bits_decodeResult_sWrite = laneRequestSourceWire_5_bits_decodeResult_sWrite;
  wire         validSource_5_bits_decodeResult_crossRead = laneRequestSourceWire_5_bits_decodeResult_crossRead;
  wire         validSource_5_bits_decodeResult_crossWrite = laneRequestSourceWire_5_bits_decodeResult_crossWrite;
  wire         validSource_5_bits_decodeResult_maskUnit = laneRequestSourceWire_5_bits_decodeResult_maskUnit;
  wire         validSource_5_bits_decodeResult_special = laneRequestSourceWire_5_bits_decodeResult_special;
  wire         validSource_5_bits_decodeResult_saturate = laneRequestSourceWire_5_bits_decodeResult_saturate;
  wire         validSource_5_bits_decodeResult_vwmacc = laneRequestSourceWire_5_bits_decodeResult_vwmacc;
  wire         validSource_5_bits_decodeResult_readOnly = laneRequestSourceWire_5_bits_decodeResult_readOnly;
  wire         validSource_5_bits_decodeResult_maskSource = laneRequestSourceWire_5_bits_decodeResult_maskSource;
  wire         validSource_5_bits_decodeResult_maskDestination = laneRequestSourceWire_5_bits_decodeResult_maskDestination;
  wire         validSource_5_bits_decodeResult_maskLogic = laneRequestSourceWire_5_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_5_bits_decodeResult_uop = laneRequestSourceWire_5_bits_decodeResult_uop;
  wire         validSource_5_bits_decodeResult_iota = laneRequestSourceWire_5_bits_decodeResult_iota;
  wire         validSource_5_bits_decodeResult_mv = laneRequestSourceWire_5_bits_decodeResult_mv;
  wire         validSource_5_bits_decodeResult_extend = laneRequestSourceWire_5_bits_decodeResult_extend;
  wire         validSource_5_bits_decodeResult_unOrderWrite = laneRequestSourceWire_5_bits_decodeResult_unOrderWrite;
  wire         validSource_5_bits_decodeResult_compress = laneRequestSourceWire_5_bits_decodeResult_compress;
  wire         validSource_5_bits_decodeResult_gather16 = laneRequestSourceWire_5_bits_decodeResult_gather16;
  wire         validSource_5_bits_decodeResult_gather = laneRequestSourceWire_5_bits_decodeResult_gather;
  wire         validSource_5_bits_decodeResult_slid = laneRequestSourceWire_5_bits_decodeResult_slid;
  wire         validSource_5_bits_decodeResult_targetRd = laneRequestSourceWire_5_bits_decodeResult_targetRd;
  wire         validSource_5_bits_decodeResult_widenReduce = laneRequestSourceWire_5_bits_decodeResult_widenReduce;
  wire         validSource_5_bits_decodeResult_red = laneRequestSourceWire_5_bits_decodeResult_red;
  wire         validSource_5_bits_decodeResult_nr = laneRequestSourceWire_5_bits_decodeResult_nr;
  wire         validSource_5_bits_decodeResult_itype = laneRequestSourceWire_5_bits_decodeResult_itype;
  wire         validSource_5_bits_decodeResult_unsigned1 = laneRequestSourceWire_5_bits_decodeResult_unsigned1;
  wire         validSource_5_bits_decodeResult_unsigned0 = laneRequestSourceWire_5_bits_decodeResult_unsigned0;
  wire         validSource_5_bits_decodeResult_other = laneRequestSourceWire_5_bits_decodeResult_other;
  wire         validSource_5_bits_decodeResult_multiCycle = laneRequestSourceWire_5_bits_decodeResult_multiCycle;
  wire         validSource_5_bits_decodeResult_divider = laneRequestSourceWire_5_bits_decodeResult_divider;
  wire         validSource_5_bits_decodeResult_multiplier = laneRequestSourceWire_5_bits_decodeResult_multiplier;
  wire         validSource_5_bits_decodeResult_shift = laneRequestSourceWire_5_bits_decodeResult_shift;
  wire         validSource_5_bits_decodeResult_adder = laneRequestSourceWire_5_bits_decodeResult_adder;
  wire         validSource_5_bits_decodeResult_logic = laneRequestSourceWire_5_bits_decodeResult_logic;
  wire         validSource_5_bits_loadStore = laneRequestSourceWire_5_bits_loadStore;
  wire         validSource_5_bits_issueInst = laneRequestSourceWire_5_bits_issueInst;
  wire         validSource_5_bits_store = laneRequestSourceWire_5_bits_store;
  wire         validSource_5_bits_special = laneRequestSourceWire_5_bits_special;
  wire         validSource_5_bits_lsWholeReg = laneRequestSourceWire_5_bits_lsWholeReg;
  wire [4:0]   validSource_5_bits_vs1 = laneRequestSourceWire_5_bits_vs1;
  wire [4:0]   validSource_5_bits_vs2 = laneRequestSourceWire_5_bits_vs2;
  wire [4:0]   validSource_5_bits_vd = laneRequestSourceWire_5_bits_vd;
  wire [1:0]   validSource_5_bits_loadStoreEEW = laneRequestSourceWire_5_bits_loadStoreEEW;
  wire         validSource_5_bits_mask = laneRequestSourceWire_5_bits_mask;
  wire [2:0]   validSource_5_bits_segment = laneRequestSourceWire_5_bits_segment;
  wire [31:0]  validSource_5_bits_readFromScalar = laneRequestSourceWire_5_bits_readFromScalar;
  wire [11:0]  validSource_5_bits_csrInterface_vl = laneRequestSourceWire_5_bits_csrInterface_vl;
  wire [11:0]  validSource_5_bits_csrInterface_vStart = laneRequestSourceWire_5_bits_csrInterface_vStart;
  wire [2:0]   validSource_5_bits_csrInterface_vlmul = laneRequestSourceWire_5_bits_csrInterface_vlmul;
  wire [1:0]   validSource_5_bits_csrInterface_vSew = laneRequestSourceWire_5_bits_csrInterface_vSew;
  wire [1:0]   validSource_5_bits_csrInterface_vxrm = laneRequestSourceWire_5_bits_csrInterface_vxrm;
  wire         validSource_5_bits_csrInterface_vta = laneRequestSourceWire_5_bits_csrInterface_vta;
  wire         validSource_5_bits_csrInterface_vma = laneRequestSourceWire_5_bits_csrInterface_vma;
  wire         tokenCheck_6;
  wire [2:0]   validSource_6_bits_instructionIndex = laneRequestSourceWire_6_bits_instructionIndex;
  wire         validSource_6_bits_decodeResult_specialSlot = laneRequestSourceWire_6_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_6_bits_decodeResult_topUop = laneRequestSourceWire_6_bits_decodeResult_topUop;
  wire         validSource_6_bits_decodeResult_popCount = laneRequestSourceWire_6_bits_decodeResult_popCount;
  wire         validSource_6_bits_decodeResult_ffo = laneRequestSourceWire_6_bits_decodeResult_ffo;
  wire         validSource_6_bits_decodeResult_average = laneRequestSourceWire_6_bits_decodeResult_average;
  wire         validSource_6_bits_decodeResult_reverse = laneRequestSourceWire_6_bits_decodeResult_reverse;
  wire         validSource_6_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_6_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_6_bits_decodeResult_scheduler = laneRequestSourceWire_6_bits_decodeResult_scheduler;
  wire         validSource_6_bits_decodeResult_sReadVD = laneRequestSourceWire_6_bits_decodeResult_sReadVD;
  wire         validSource_6_bits_decodeResult_vtype = laneRequestSourceWire_6_bits_decodeResult_vtype;
  wire         validSource_6_bits_decodeResult_sWrite = laneRequestSourceWire_6_bits_decodeResult_sWrite;
  wire         validSource_6_bits_decodeResult_crossRead = laneRequestSourceWire_6_bits_decodeResult_crossRead;
  wire         validSource_6_bits_decodeResult_crossWrite = laneRequestSourceWire_6_bits_decodeResult_crossWrite;
  wire         validSource_6_bits_decodeResult_maskUnit = laneRequestSourceWire_6_bits_decodeResult_maskUnit;
  wire         validSource_6_bits_decodeResult_special = laneRequestSourceWire_6_bits_decodeResult_special;
  wire         validSource_6_bits_decodeResult_saturate = laneRequestSourceWire_6_bits_decodeResult_saturate;
  wire         validSource_6_bits_decodeResult_vwmacc = laneRequestSourceWire_6_bits_decodeResult_vwmacc;
  wire         validSource_6_bits_decodeResult_readOnly = laneRequestSourceWire_6_bits_decodeResult_readOnly;
  wire         validSource_6_bits_decodeResult_maskSource = laneRequestSourceWire_6_bits_decodeResult_maskSource;
  wire         validSource_6_bits_decodeResult_maskDestination = laneRequestSourceWire_6_bits_decodeResult_maskDestination;
  wire         validSource_6_bits_decodeResult_maskLogic = laneRequestSourceWire_6_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_6_bits_decodeResult_uop = laneRequestSourceWire_6_bits_decodeResult_uop;
  wire         validSource_6_bits_decodeResult_iota = laneRequestSourceWire_6_bits_decodeResult_iota;
  wire         validSource_6_bits_decodeResult_mv = laneRequestSourceWire_6_bits_decodeResult_mv;
  wire         validSource_6_bits_decodeResult_extend = laneRequestSourceWire_6_bits_decodeResult_extend;
  wire         validSource_6_bits_decodeResult_unOrderWrite = laneRequestSourceWire_6_bits_decodeResult_unOrderWrite;
  wire         validSource_6_bits_decodeResult_compress = laneRequestSourceWire_6_bits_decodeResult_compress;
  wire         validSource_6_bits_decodeResult_gather16 = laneRequestSourceWire_6_bits_decodeResult_gather16;
  wire         validSource_6_bits_decodeResult_gather = laneRequestSourceWire_6_bits_decodeResult_gather;
  wire         validSource_6_bits_decodeResult_slid = laneRequestSourceWire_6_bits_decodeResult_slid;
  wire         validSource_6_bits_decodeResult_targetRd = laneRequestSourceWire_6_bits_decodeResult_targetRd;
  wire         validSource_6_bits_decodeResult_widenReduce = laneRequestSourceWire_6_bits_decodeResult_widenReduce;
  wire         validSource_6_bits_decodeResult_red = laneRequestSourceWire_6_bits_decodeResult_red;
  wire         validSource_6_bits_decodeResult_nr = laneRequestSourceWire_6_bits_decodeResult_nr;
  wire         validSource_6_bits_decodeResult_itype = laneRequestSourceWire_6_bits_decodeResult_itype;
  wire         validSource_6_bits_decodeResult_unsigned1 = laneRequestSourceWire_6_bits_decodeResult_unsigned1;
  wire         validSource_6_bits_decodeResult_unsigned0 = laneRequestSourceWire_6_bits_decodeResult_unsigned0;
  wire         validSource_6_bits_decodeResult_other = laneRequestSourceWire_6_bits_decodeResult_other;
  wire         validSource_6_bits_decodeResult_multiCycle = laneRequestSourceWire_6_bits_decodeResult_multiCycle;
  wire         validSource_6_bits_decodeResult_divider = laneRequestSourceWire_6_bits_decodeResult_divider;
  wire         validSource_6_bits_decodeResult_multiplier = laneRequestSourceWire_6_bits_decodeResult_multiplier;
  wire         validSource_6_bits_decodeResult_shift = laneRequestSourceWire_6_bits_decodeResult_shift;
  wire         validSource_6_bits_decodeResult_adder = laneRequestSourceWire_6_bits_decodeResult_adder;
  wire         validSource_6_bits_decodeResult_logic = laneRequestSourceWire_6_bits_decodeResult_logic;
  wire         validSource_6_bits_loadStore = laneRequestSourceWire_6_bits_loadStore;
  wire         validSource_6_bits_issueInst = laneRequestSourceWire_6_bits_issueInst;
  wire         validSource_6_bits_store = laneRequestSourceWire_6_bits_store;
  wire         validSource_6_bits_special = laneRequestSourceWire_6_bits_special;
  wire         validSource_6_bits_lsWholeReg = laneRequestSourceWire_6_bits_lsWholeReg;
  wire [4:0]   validSource_6_bits_vs1 = laneRequestSourceWire_6_bits_vs1;
  wire [4:0]   validSource_6_bits_vs2 = laneRequestSourceWire_6_bits_vs2;
  wire [4:0]   validSource_6_bits_vd = laneRequestSourceWire_6_bits_vd;
  wire [1:0]   validSource_6_bits_loadStoreEEW = laneRequestSourceWire_6_bits_loadStoreEEW;
  wire         validSource_6_bits_mask = laneRequestSourceWire_6_bits_mask;
  wire [2:0]   validSource_6_bits_segment = laneRequestSourceWire_6_bits_segment;
  wire [31:0]  validSource_6_bits_readFromScalar = laneRequestSourceWire_6_bits_readFromScalar;
  wire [11:0]  validSource_6_bits_csrInterface_vl = laneRequestSourceWire_6_bits_csrInterface_vl;
  wire [11:0]  validSource_6_bits_csrInterface_vStart = laneRequestSourceWire_6_bits_csrInterface_vStart;
  wire [2:0]   validSource_6_bits_csrInterface_vlmul = laneRequestSourceWire_6_bits_csrInterface_vlmul;
  wire [1:0]   validSource_6_bits_csrInterface_vSew = laneRequestSourceWire_6_bits_csrInterface_vSew;
  wire [1:0]   validSource_6_bits_csrInterface_vxrm = laneRequestSourceWire_6_bits_csrInterface_vxrm;
  wire         validSource_6_bits_csrInterface_vta = laneRequestSourceWire_6_bits_csrInterface_vta;
  wire         validSource_6_bits_csrInterface_vma = laneRequestSourceWire_6_bits_csrInterface_vma;
  wire         tokenCheck_7;
  wire [2:0]   validSource_7_bits_instructionIndex = laneRequestSourceWire_7_bits_instructionIndex;
  wire         validSource_7_bits_decodeResult_specialSlot = laneRequestSourceWire_7_bits_decodeResult_specialSlot;
  wire [4:0]   validSource_7_bits_decodeResult_topUop = laneRequestSourceWire_7_bits_decodeResult_topUop;
  wire         validSource_7_bits_decodeResult_popCount = laneRequestSourceWire_7_bits_decodeResult_popCount;
  wire         validSource_7_bits_decodeResult_ffo = laneRequestSourceWire_7_bits_decodeResult_ffo;
  wire         validSource_7_bits_decodeResult_average = laneRequestSourceWire_7_bits_decodeResult_average;
  wire         validSource_7_bits_decodeResult_reverse = laneRequestSourceWire_7_bits_decodeResult_reverse;
  wire         validSource_7_bits_decodeResult_dontNeedExecuteInLane = laneRequestSourceWire_7_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSource_7_bits_decodeResult_scheduler = laneRequestSourceWire_7_bits_decodeResult_scheduler;
  wire         validSource_7_bits_decodeResult_sReadVD = laneRequestSourceWire_7_bits_decodeResult_sReadVD;
  wire         validSource_7_bits_decodeResult_vtype = laneRequestSourceWire_7_bits_decodeResult_vtype;
  wire         validSource_7_bits_decodeResult_sWrite = laneRequestSourceWire_7_bits_decodeResult_sWrite;
  wire         validSource_7_bits_decodeResult_crossRead = laneRequestSourceWire_7_bits_decodeResult_crossRead;
  wire         validSource_7_bits_decodeResult_crossWrite = laneRequestSourceWire_7_bits_decodeResult_crossWrite;
  wire         validSource_7_bits_decodeResult_maskUnit = laneRequestSourceWire_7_bits_decodeResult_maskUnit;
  wire         validSource_7_bits_decodeResult_special = laneRequestSourceWire_7_bits_decodeResult_special;
  wire         validSource_7_bits_decodeResult_saturate = laneRequestSourceWire_7_bits_decodeResult_saturate;
  wire         validSource_7_bits_decodeResult_vwmacc = laneRequestSourceWire_7_bits_decodeResult_vwmacc;
  wire         validSource_7_bits_decodeResult_readOnly = laneRequestSourceWire_7_bits_decodeResult_readOnly;
  wire         validSource_7_bits_decodeResult_maskSource = laneRequestSourceWire_7_bits_decodeResult_maskSource;
  wire         validSource_7_bits_decodeResult_maskDestination = laneRequestSourceWire_7_bits_decodeResult_maskDestination;
  wire         validSource_7_bits_decodeResult_maskLogic = laneRequestSourceWire_7_bits_decodeResult_maskLogic;
  wire [3:0]   validSource_7_bits_decodeResult_uop = laneRequestSourceWire_7_bits_decodeResult_uop;
  wire         validSource_7_bits_decodeResult_iota = laneRequestSourceWire_7_bits_decodeResult_iota;
  wire         validSource_7_bits_decodeResult_mv = laneRequestSourceWire_7_bits_decodeResult_mv;
  wire         validSource_7_bits_decodeResult_extend = laneRequestSourceWire_7_bits_decodeResult_extend;
  wire         validSource_7_bits_decodeResult_unOrderWrite = laneRequestSourceWire_7_bits_decodeResult_unOrderWrite;
  wire         validSource_7_bits_decodeResult_compress = laneRequestSourceWire_7_bits_decodeResult_compress;
  wire         validSource_7_bits_decodeResult_gather16 = laneRequestSourceWire_7_bits_decodeResult_gather16;
  wire         validSource_7_bits_decodeResult_gather = laneRequestSourceWire_7_bits_decodeResult_gather;
  wire         validSource_7_bits_decodeResult_slid = laneRequestSourceWire_7_bits_decodeResult_slid;
  wire         validSource_7_bits_decodeResult_targetRd = laneRequestSourceWire_7_bits_decodeResult_targetRd;
  wire         validSource_7_bits_decodeResult_widenReduce = laneRequestSourceWire_7_bits_decodeResult_widenReduce;
  wire         validSource_7_bits_decodeResult_red = laneRequestSourceWire_7_bits_decodeResult_red;
  wire         validSource_7_bits_decodeResult_nr = laneRequestSourceWire_7_bits_decodeResult_nr;
  wire         validSource_7_bits_decodeResult_itype = laneRequestSourceWire_7_bits_decodeResult_itype;
  wire         validSource_7_bits_decodeResult_unsigned1 = laneRequestSourceWire_7_bits_decodeResult_unsigned1;
  wire         validSource_7_bits_decodeResult_unsigned0 = laneRequestSourceWire_7_bits_decodeResult_unsigned0;
  wire         validSource_7_bits_decodeResult_other = laneRequestSourceWire_7_bits_decodeResult_other;
  wire         validSource_7_bits_decodeResult_multiCycle = laneRequestSourceWire_7_bits_decodeResult_multiCycle;
  wire         validSource_7_bits_decodeResult_divider = laneRequestSourceWire_7_bits_decodeResult_divider;
  wire         validSource_7_bits_decodeResult_multiplier = laneRequestSourceWire_7_bits_decodeResult_multiplier;
  wire         validSource_7_bits_decodeResult_shift = laneRequestSourceWire_7_bits_decodeResult_shift;
  wire         validSource_7_bits_decodeResult_adder = laneRequestSourceWire_7_bits_decodeResult_adder;
  wire         validSource_7_bits_decodeResult_logic = laneRequestSourceWire_7_bits_decodeResult_logic;
  wire         validSource_7_bits_loadStore = laneRequestSourceWire_7_bits_loadStore;
  wire         validSource_7_bits_issueInst = laneRequestSourceWire_7_bits_issueInst;
  wire         validSource_7_bits_store = laneRequestSourceWire_7_bits_store;
  wire         validSource_7_bits_special = laneRequestSourceWire_7_bits_special;
  wire         validSource_7_bits_lsWholeReg = laneRequestSourceWire_7_bits_lsWholeReg;
  wire [4:0]   validSource_7_bits_vs1 = laneRequestSourceWire_7_bits_vs1;
  wire [4:0]   validSource_7_bits_vs2 = laneRequestSourceWire_7_bits_vs2;
  wire [4:0]   validSource_7_bits_vd = laneRequestSourceWire_7_bits_vd;
  wire [1:0]   validSource_7_bits_loadStoreEEW = laneRequestSourceWire_7_bits_loadStoreEEW;
  wire         validSource_7_bits_mask = laneRequestSourceWire_7_bits_mask;
  wire [2:0]   validSource_7_bits_segment = laneRequestSourceWire_7_bits_segment;
  wire [31:0]  validSource_7_bits_readFromScalar = laneRequestSourceWire_7_bits_readFromScalar;
  wire [11:0]  validSource_7_bits_csrInterface_vl = laneRequestSourceWire_7_bits_csrInterface_vl;
  wire [11:0]  validSource_7_bits_csrInterface_vStart = laneRequestSourceWire_7_bits_csrInterface_vStart;
  wire [2:0]   validSource_7_bits_csrInterface_vlmul = laneRequestSourceWire_7_bits_csrInterface_vlmul;
  wire [1:0]   validSource_7_bits_csrInterface_vSew = laneRequestSourceWire_7_bits_csrInterface_vSew;
  wire [1:0]   validSource_7_bits_csrInterface_vxrm = laneRequestSourceWire_7_bits_csrInterface_vxrm;
  wire         validSource_7_bits_csrInterface_vta = laneRequestSourceWire_7_bits_csrInterface_vta;
  wire         validSource_7_bits_csrInterface_vma = laneRequestSourceWire_7_bits_csrInterface_vma;
  wire         queue_deq_ready = laneRequestSinkWire_0_ready;
  wire         queue_deq_valid;
  wire [2:0]   queue_deq_bits_instructionIndex;
  wire         queue_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_deq_bits_decodeResult_topUop;
  wire         queue_deq_bits_decodeResult_popCount;
  wire         queue_deq_bits_decodeResult_ffo;
  wire         queue_deq_bits_decodeResult_average;
  wire         queue_deq_bits_decodeResult_reverse;
  wire         queue_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_deq_bits_decodeResult_scheduler;
  wire         queue_deq_bits_decodeResult_sReadVD;
  wire         queue_deq_bits_decodeResult_vtype;
  wire         queue_deq_bits_decodeResult_sWrite;
  wire         queue_deq_bits_decodeResult_crossRead;
  wire         queue_deq_bits_decodeResult_crossWrite;
  wire         queue_deq_bits_decodeResult_maskUnit;
  wire         queue_deq_bits_decodeResult_special;
  wire         queue_deq_bits_decodeResult_saturate;
  wire         queue_deq_bits_decodeResult_vwmacc;
  wire         queue_deq_bits_decodeResult_readOnly;
  wire         queue_deq_bits_decodeResult_maskSource;
  wire         queue_deq_bits_decodeResult_maskDestination;
  wire         queue_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_deq_bits_decodeResult_uop;
  wire         queue_deq_bits_decodeResult_iota;
  wire         queue_deq_bits_decodeResult_mv;
  wire         queue_deq_bits_decodeResult_extend;
  wire         queue_deq_bits_decodeResult_unOrderWrite;
  wire         queue_deq_bits_decodeResult_compress;
  wire         queue_deq_bits_decodeResult_gather16;
  wire         queue_deq_bits_decodeResult_gather;
  wire         queue_deq_bits_decodeResult_slid;
  wire         queue_deq_bits_decodeResult_targetRd;
  wire         queue_deq_bits_decodeResult_widenReduce;
  wire         queue_deq_bits_decodeResult_red;
  wire         queue_deq_bits_decodeResult_nr;
  wire         queue_deq_bits_decodeResult_itype;
  wire         queue_deq_bits_decodeResult_unsigned1;
  wire         queue_deq_bits_decodeResult_unsigned0;
  wire         queue_deq_bits_decodeResult_other;
  wire         queue_deq_bits_decodeResult_multiCycle;
  wire         queue_deq_bits_decodeResult_divider;
  wire         queue_deq_bits_decodeResult_multiplier;
  wire         queue_deq_bits_decodeResult_shift;
  wire         queue_deq_bits_decodeResult_adder;
  wire         queue_deq_bits_decodeResult_logic;
  wire         queue_deq_bits_loadStore;
  wire         queue_deq_bits_issueInst;
  wire         queue_deq_bits_store;
  wire         queue_deq_bits_special;
  wire         queue_deq_bits_lsWholeReg;
  wire [4:0]   queue_deq_bits_vs1;
  wire [4:0]   queue_deq_bits_vs2;
  wire [4:0]   queue_deq_bits_vd;
  wire [1:0]   queue_deq_bits_loadStoreEEW;
  wire         queue_deq_bits_mask;
  wire [2:0]   queue_deq_bits_segment;
  wire [31:0]  queue_deq_bits_readFromScalar;
  wire [11:0]  queue_deq_bits_csrInterface_vl;
  wire [11:0]  queue_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_deq_bits_csrInterface_vxrm;
  wire         queue_deq_bits_csrInterface_vta;
  wire         queue_deq_bits_csrInterface_vma;
  wire         queue_1_deq_ready = laneRequestSinkWire_1_ready;
  wire         queue_1_deq_valid;
  wire [2:0]   queue_1_deq_bits_instructionIndex;
  wire         queue_1_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_1_deq_bits_decodeResult_topUop;
  wire         queue_1_deq_bits_decodeResult_popCount;
  wire         queue_1_deq_bits_decodeResult_ffo;
  wire         queue_1_deq_bits_decodeResult_average;
  wire         queue_1_deq_bits_decodeResult_reverse;
  wire         queue_1_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_1_deq_bits_decodeResult_scheduler;
  wire         queue_1_deq_bits_decodeResult_sReadVD;
  wire         queue_1_deq_bits_decodeResult_vtype;
  wire         queue_1_deq_bits_decodeResult_sWrite;
  wire         queue_1_deq_bits_decodeResult_crossRead;
  wire         queue_1_deq_bits_decodeResult_crossWrite;
  wire         queue_1_deq_bits_decodeResult_maskUnit;
  wire         queue_1_deq_bits_decodeResult_special;
  wire         queue_1_deq_bits_decodeResult_saturate;
  wire         queue_1_deq_bits_decodeResult_vwmacc;
  wire         queue_1_deq_bits_decodeResult_readOnly;
  wire         queue_1_deq_bits_decodeResult_maskSource;
  wire         queue_1_deq_bits_decodeResult_maskDestination;
  wire         queue_1_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_1_deq_bits_decodeResult_uop;
  wire         queue_1_deq_bits_decodeResult_iota;
  wire         queue_1_deq_bits_decodeResult_mv;
  wire         queue_1_deq_bits_decodeResult_extend;
  wire         queue_1_deq_bits_decodeResult_unOrderWrite;
  wire         queue_1_deq_bits_decodeResult_compress;
  wire         queue_1_deq_bits_decodeResult_gather16;
  wire         queue_1_deq_bits_decodeResult_gather;
  wire         queue_1_deq_bits_decodeResult_slid;
  wire         queue_1_deq_bits_decodeResult_targetRd;
  wire         queue_1_deq_bits_decodeResult_widenReduce;
  wire         queue_1_deq_bits_decodeResult_red;
  wire         queue_1_deq_bits_decodeResult_nr;
  wire         queue_1_deq_bits_decodeResult_itype;
  wire         queue_1_deq_bits_decodeResult_unsigned1;
  wire         queue_1_deq_bits_decodeResult_unsigned0;
  wire         queue_1_deq_bits_decodeResult_other;
  wire         queue_1_deq_bits_decodeResult_multiCycle;
  wire         queue_1_deq_bits_decodeResult_divider;
  wire         queue_1_deq_bits_decodeResult_multiplier;
  wire         queue_1_deq_bits_decodeResult_shift;
  wire         queue_1_deq_bits_decodeResult_adder;
  wire         queue_1_deq_bits_decodeResult_logic;
  wire         queue_1_deq_bits_loadStore;
  wire         queue_1_deq_bits_issueInst;
  wire         queue_1_deq_bits_store;
  wire         queue_1_deq_bits_special;
  wire         queue_1_deq_bits_lsWholeReg;
  wire [4:0]   queue_1_deq_bits_vs1;
  wire [4:0]   queue_1_deq_bits_vs2;
  wire [4:0]   queue_1_deq_bits_vd;
  wire [1:0]   queue_1_deq_bits_loadStoreEEW;
  wire         queue_1_deq_bits_mask;
  wire [2:0]   queue_1_deq_bits_segment;
  wire [31:0]  queue_1_deq_bits_readFromScalar;
  wire [11:0]  queue_1_deq_bits_csrInterface_vl;
  wire [11:0]  queue_1_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_1_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_1_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_1_deq_bits_csrInterface_vxrm;
  wire         queue_1_deq_bits_csrInterface_vta;
  wire         queue_1_deq_bits_csrInterface_vma;
  wire         queue_2_deq_ready = laneRequestSinkWire_2_ready;
  wire         queue_2_deq_valid;
  wire [2:0]   queue_2_deq_bits_instructionIndex;
  wire         queue_2_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_2_deq_bits_decodeResult_topUop;
  wire         queue_2_deq_bits_decodeResult_popCount;
  wire         queue_2_deq_bits_decodeResult_ffo;
  wire         queue_2_deq_bits_decodeResult_average;
  wire         queue_2_deq_bits_decodeResult_reverse;
  wire         queue_2_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_2_deq_bits_decodeResult_scheduler;
  wire         queue_2_deq_bits_decodeResult_sReadVD;
  wire         queue_2_deq_bits_decodeResult_vtype;
  wire         queue_2_deq_bits_decodeResult_sWrite;
  wire         queue_2_deq_bits_decodeResult_crossRead;
  wire         queue_2_deq_bits_decodeResult_crossWrite;
  wire         queue_2_deq_bits_decodeResult_maskUnit;
  wire         queue_2_deq_bits_decodeResult_special;
  wire         queue_2_deq_bits_decodeResult_saturate;
  wire         queue_2_deq_bits_decodeResult_vwmacc;
  wire         queue_2_deq_bits_decodeResult_readOnly;
  wire         queue_2_deq_bits_decodeResult_maskSource;
  wire         queue_2_deq_bits_decodeResult_maskDestination;
  wire         queue_2_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_2_deq_bits_decodeResult_uop;
  wire         queue_2_deq_bits_decodeResult_iota;
  wire         queue_2_deq_bits_decodeResult_mv;
  wire         queue_2_deq_bits_decodeResult_extend;
  wire         queue_2_deq_bits_decodeResult_unOrderWrite;
  wire         queue_2_deq_bits_decodeResult_compress;
  wire         queue_2_deq_bits_decodeResult_gather16;
  wire         queue_2_deq_bits_decodeResult_gather;
  wire         queue_2_deq_bits_decodeResult_slid;
  wire         queue_2_deq_bits_decodeResult_targetRd;
  wire         queue_2_deq_bits_decodeResult_widenReduce;
  wire         queue_2_deq_bits_decodeResult_red;
  wire         queue_2_deq_bits_decodeResult_nr;
  wire         queue_2_deq_bits_decodeResult_itype;
  wire         queue_2_deq_bits_decodeResult_unsigned1;
  wire         queue_2_deq_bits_decodeResult_unsigned0;
  wire         queue_2_deq_bits_decodeResult_other;
  wire         queue_2_deq_bits_decodeResult_multiCycle;
  wire         queue_2_deq_bits_decodeResult_divider;
  wire         queue_2_deq_bits_decodeResult_multiplier;
  wire         queue_2_deq_bits_decodeResult_shift;
  wire         queue_2_deq_bits_decodeResult_adder;
  wire         queue_2_deq_bits_decodeResult_logic;
  wire         queue_2_deq_bits_loadStore;
  wire         queue_2_deq_bits_issueInst;
  wire         queue_2_deq_bits_store;
  wire         queue_2_deq_bits_special;
  wire         queue_2_deq_bits_lsWholeReg;
  wire [4:0]   queue_2_deq_bits_vs1;
  wire [4:0]   queue_2_deq_bits_vs2;
  wire [4:0]   queue_2_deq_bits_vd;
  wire [1:0]   queue_2_deq_bits_loadStoreEEW;
  wire         queue_2_deq_bits_mask;
  wire [2:0]   queue_2_deq_bits_segment;
  wire [31:0]  queue_2_deq_bits_readFromScalar;
  wire [11:0]  queue_2_deq_bits_csrInterface_vl;
  wire [11:0]  queue_2_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_2_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_2_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_2_deq_bits_csrInterface_vxrm;
  wire         queue_2_deq_bits_csrInterface_vta;
  wire         queue_2_deq_bits_csrInterface_vma;
  wire         queue_3_deq_ready = laneRequestSinkWire_3_ready;
  wire         queue_3_deq_valid;
  wire [2:0]   queue_3_deq_bits_instructionIndex;
  wire         queue_3_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_3_deq_bits_decodeResult_topUop;
  wire         queue_3_deq_bits_decodeResult_popCount;
  wire         queue_3_deq_bits_decodeResult_ffo;
  wire         queue_3_deq_bits_decodeResult_average;
  wire         queue_3_deq_bits_decodeResult_reverse;
  wire         queue_3_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_3_deq_bits_decodeResult_scheduler;
  wire         queue_3_deq_bits_decodeResult_sReadVD;
  wire         queue_3_deq_bits_decodeResult_vtype;
  wire         queue_3_deq_bits_decodeResult_sWrite;
  wire         queue_3_deq_bits_decodeResult_crossRead;
  wire         queue_3_deq_bits_decodeResult_crossWrite;
  wire         queue_3_deq_bits_decodeResult_maskUnit;
  wire         queue_3_deq_bits_decodeResult_special;
  wire         queue_3_deq_bits_decodeResult_saturate;
  wire         queue_3_deq_bits_decodeResult_vwmacc;
  wire         queue_3_deq_bits_decodeResult_readOnly;
  wire         queue_3_deq_bits_decodeResult_maskSource;
  wire         queue_3_deq_bits_decodeResult_maskDestination;
  wire         queue_3_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_3_deq_bits_decodeResult_uop;
  wire         queue_3_deq_bits_decodeResult_iota;
  wire         queue_3_deq_bits_decodeResult_mv;
  wire         queue_3_deq_bits_decodeResult_extend;
  wire         queue_3_deq_bits_decodeResult_unOrderWrite;
  wire         queue_3_deq_bits_decodeResult_compress;
  wire         queue_3_deq_bits_decodeResult_gather16;
  wire         queue_3_deq_bits_decodeResult_gather;
  wire         queue_3_deq_bits_decodeResult_slid;
  wire         queue_3_deq_bits_decodeResult_targetRd;
  wire         queue_3_deq_bits_decodeResult_widenReduce;
  wire         queue_3_deq_bits_decodeResult_red;
  wire         queue_3_deq_bits_decodeResult_nr;
  wire         queue_3_deq_bits_decodeResult_itype;
  wire         queue_3_deq_bits_decodeResult_unsigned1;
  wire         queue_3_deq_bits_decodeResult_unsigned0;
  wire         queue_3_deq_bits_decodeResult_other;
  wire         queue_3_deq_bits_decodeResult_multiCycle;
  wire         queue_3_deq_bits_decodeResult_divider;
  wire         queue_3_deq_bits_decodeResult_multiplier;
  wire         queue_3_deq_bits_decodeResult_shift;
  wire         queue_3_deq_bits_decodeResult_adder;
  wire         queue_3_deq_bits_decodeResult_logic;
  wire         queue_3_deq_bits_loadStore;
  wire         queue_3_deq_bits_issueInst;
  wire         queue_3_deq_bits_store;
  wire         queue_3_deq_bits_special;
  wire         queue_3_deq_bits_lsWholeReg;
  wire [4:0]   queue_3_deq_bits_vs1;
  wire [4:0]   queue_3_deq_bits_vs2;
  wire [4:0]   queue_3_deq_bits_vd;
  wire [1:0]   queue_3_deq_bits_loadStoreEEW;
  wire         queue_3_deq_bits_mask;
  wire [2:0]   queue_3_deq_bits_segment;
  wire [31:0]  queue_3_deq_bits_readFromScalar;
  wire [11:0]  queue_3_deq_bits_csrInterface_vl;
  wire [11:0]  queue_3_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_3_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_3_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_3_deq_bits_csrInterface_vxrm;
  wire         queue_3_deq_bits_csrInterface_vta;
  wire         queue_3_deq_bits_csrInterface_vma;
  wire         queue_4_deq_ready = laneRequestSinkWire_4_ready;
  wire         queue_4_deq_valid;
  wire [2:0]   queue_4_deq_bits_instructionIndex;
  wire         queue_4_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_4_deq_bits_decodeResult_topUop;
  wire         queue_4_deq_bits_decodeResult_popCount;
  wire         queue_4_deq_bits_decodeResult_ffo;
  wire         queue_4_deq_bits_decodeResult_average;
  wire         queue_4_deq_bits_decodeResult_reverse;
  wire         queue_4_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_4_deq_bits_decodeResult_scheduler;
  wire         queue_4_deq_bits_decodeResult_sReadVD;
  wire         queue_4_deq_bits_decodeResult_vtype;
  wire         queue_4_deq_bits_decodeResult_sWrite;
  wire         queue_4_deq_bits_decodeResult_crossRead;
  wire         queue_4_deq_bits_decodeResult_crossWrite;
  wire         queue_4_deq_bits_decodeResult_maskUnit;
  wire         queue_4_deq_bits_decodeResult_special;
  wire         queue_4_deq_bits_decodeResult_saturate;
  wire         queue_4_deq_bits_decodeResult_vwmacc;
  wire         queue_4_deq_bits_decodeResult_readOnly;
  wire         queue_4_deq_bits_decodeResult_maskSource;
  wire         queue_4_deq_bits_decodeResult_maskDestination;
  wire         queue_4_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_4_deq_bits_decodeResult_uop;
  wire         queue_4_deq_bits_decodeResult_iota;
  wire         queue_4_deq_bits_decodeResult_mv;
  wire         queue_4_deq_bits_decodeResult_extend;
  wire         queue_4_deq_bits_decodeResult_unOrderWrite;
  wire         queue_4_deq_bits_decodeResult_compress;
  wire         queue_4_deq_bits_decodeResult_gather16;
  wire         queue_4_deq_bits_decodeResult_gather;
  wire         queue_4_deq_bits_decodeResult_slid;
  wire         queue_4_deq_bits_decodeResult_targetRd;
  wire         queue_4_deq_bits_decodeResult_widenReduce;
  wire         queue_4_deq_bits_decodeResult_red;
  wire         queue_4_deq_bits_decodeResult_nr;
  wire         queue_4_deq_bits_decodeResult_itype;
  wire         queue_4_deq_bits_decodeResult_unsigned1;
  wire         queue_4_deq_bits_decodeResult_unsigned0;
  wire         queue_4_deq_bits_decodeResult_other;
  wire         queue_4_deq_bits_decodeResult_multiCycle;
  wire         queue_4_deq_bits_decodeResult_divider;
  wire         queue_4_deq_bits_decodeResult_multiplier;
  wire         queue_4_deq_bits_decodeResult_shift;
  wire         queue_4_deq_bits_decodeResult_adder;
  wire         queue_4_deq_bits_decodeResult_logic;
  wire         queue_4_deq_bits_loadStore;
  wire         queue_4_deq_bits_issueInst;
  wire         queue_4_deq_bits_store;
  wire         queue_4_deq_bits_special;
  wire         queue_4_deq_bits_lsWholeReg;
  wire [4:0]   queue_4_deq_bits_vs1;
  wire [4:0]   queue_4_deq_bits_vs2;
  wire [4:0]   queue_4_deq_bits_vd;
  wire [1:0]   queue_4_deq_bits_loadStoreEEW;
  wire         queue_4_deq_bits_mask;
  wire [2:0]   queue_4_deq_bits_segment;
  wire [31:0]  queue_4_deq_bits_readFromScalar;
  wire [11:0]  queue_4_deq_bits_csrInterface_vl;
  wire [11:0]  queue_4_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_4_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_4_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_4_deq_bits_csrInterface_vxrm;
  wire         queue_4_deq_bits_csrInterface_vta;
  wire         queue_4_deq_bits_csrInterface_vma;
  wire         queue_5_deq_ready = laneRequestSinkWire_5_ready;
  wire         queue_5_deq_valid;
  wire [2:0]   queue_5_deq_bits_instructionIndex;
  wire         queue_5_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_5_deq_bits_decodeResult_topUop;
  wire         queue_5_deq_bits_decodeResult_popCount;
  wire         queue_5_deq_bits_decodeResult_ffo;
  wire         queue_5_deq_bits_decodeResult_average;
  wire         queue_5_deq_bits_decodeResult_reverse;
  wire         queue_5_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_5_deq_bits_decodeResult_scheduler;
  wire         queue_5_deq_bits_decodeResult_sReadVD;
  wire         queue_5_deq_bits_decodeResult_vtype;
  wire         queue_5_deq_bits_decodeResult_sWrite;
  wire         queue_5_deq_bits_decodeResult_crossRead;
  wire         queue_5_deq_bits_decodeResult_crossWrite;
  wire         queue_5_deq_bits_decodeResult_maskUnit;
  wire         queue_5_deq_bits_decodeResult_special;
  wire         queue_5_deq_bits_decodeResult_saturate;
  wire         queue_5_deq_bits_decodeResult_vwmacc;
  wire         queue_5_deq_bits_decodeResult_readOnly;
  wire         queue_5_deq_bits_decodeResult_maskSource;
  wire         queue_5_deq_bits_decodeResult_maskDestination;
  wire         queue_5_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_5_deq_bits_decodeResult_uop;
  wire         queue_5_deq_bits_decodeResult_iota;
  wire         queue_5_deq_bits_decodeResult_mv;
  wire         queue_5_deq_bits_decodeResult_extend;
  wire         queue_5_deq_bits_decodeResult_unOrderWrite;
  wire         queue_5_deq_bits_decodeResult_compress;
  wire         queue_5_deq_bits_decodeResult_gather16;
  wire         queue_5_deq_bits_decodeResult_gather;
  wire         queue_5_deq_bits_decodeResult_slid;
  wire         queue_5_deq_bits_decodeResult_targetRd;
  wire         queue_5_deq_bits_decodeResult_widenReduce;
  wire         queue_5_deq_bits_decodeResult_red;
  wire         queue_5_deq_bits_decodeResult_nr;
  wire         queue_5_deq_bits_decodeResult_itype;
  wire         queue_5_deq_bits_decodeResult_unsigned1;
  wire         queue_5_deq_bits_decodeResult_unsigned0;
  wire         queue_5_deq_bits_decodeResult_other;
  wire         queue_5_deq_bits_decodeResult_multiCycle;
  wire         queue_5_deq_bits_decodeResult_divider;
  wire         queue_5_deq_bits_decodeResult_multiplier;
  wire         queue_5_deq_bits_decodeResult_shift;
  wire         queue_5_deq_bits_decodeResult_adder;
  wire         queue_5_deq_bits_decodeResult_logic;
  wire         queue_5_deq_bits_loadStore;
  wire         queue_5_deq_bits_issueInst;
  wire         queue_5_deq_bits_store;
  wire         queue_5_deq_bits_special;
  wire         queue_5_deq_bits_lsWholeReg;
  wire [4:0]   queue_5_deq_bits_vs1;
  wire [4:0]   queue_5_deq_bits_vs2;
  wire [4:0]   queue_5_deq_bits_vd;
  wire [1:0]   queue_5_deq_bits_loadStoreEEW;
  wire         queue_5_deq_bits_mask;
  wire [2:0]   queue_5_deq_bits_segment;
  wire [31:0]  queue_5_deq_bits_readFromScalar;
  wire [11:0]  queue_5_deq_bits_csrInterface_vl;
  wire [11:0]  queue_5_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_5_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_5_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_5_deq_bits_csrInterface_vxrm;
  wire         queue_5_deq_bits_csrInterface_vta;
  wire         queue_5_deq_bits_csrInterface_vma;
  wire         queue_6_deq_ready = laneRequestSinkWire_6_ready;
  wire         queue_6_deq_valid;
  wire [2:0]   queue_6_deq_bits_instructionIndex;
  wire         queue_6_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_6_deq_bits_decodeResult_topUop;
  wire         queue_6_deq_bits_decodeResult_popCount;
  wire         queue_6_deq_bits_decodeResult_ffo;
  wire         queue_6_deq_bits_decodeResult_average;
  wire         queue_6_deq_bits_decodeResult_reverse;
  wire         queue_6_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_6_deq_bits_decodeResult_scheduler;
  wire         queue_6_deq_bits_decodeResult_sReadVD;
  wire         queue_6_deq_bits_decodeResult_vtype;
  wire         queue_6_deq_bits_decodeResult_sWrite;
  wire         queue_6_deq_bits_decodeResult_crossRead;
  wire         queue_6_deq_bits_decodeResult_crossWrite;
  wire         queue_6_deq_bits_decodeResult_maskUnit;
  wire         queue_6_deq_bits_decodeResult_special;
  wire         queue_6_deq_bits_decodeResult_saturate;
  wire         queue_6_deq_bits_decodeResult_vwmacc;
  wire         queue_6_deq_bits_decodeResult_readOnly;
  wire         queue_6_deq_bits_decodeResult_maskSource;
  wire         queue_6_deq_bits_decodeResult_maskDestination;
  wire         queue_6_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_6_deq_bits_decodeResult_uop;
  wire         queue_6_deq_bits_decodeResult_iota;
  wire         queue_6_deq_bits_decodeResult_mv;
  wire         queue_6_deq_bits_decodeResult_extend;
  wire         queue_6_deq_bits_decodeResult_unOrderWrite;
  wire         queue_6_deq_bits_decodeResult_compress;
  wire         queue_6_deq_bits_decodeResult_gather16;
  wire         queue_6_deq_bits_decodeResult_gather;
  wire         queue_6_deq_bits_decodeResult_slid;
  wire         queue_6_deq_bits_decodeResult_targetRd;
  wire         queue_6_deq_bits_decodeResult_widenReduce;
  wire         queue_6_deq_bits_decodeResult_red;
  wire         queue_6_deq_bits_decodeResult_nr;
  wire         queue_6_deq_bits_decodeResult_itype;
  wire         queue_6_deq_bits_decodeResult_unsigned1;
  wire         queue_6_deq_bits_decodeResult_unsigned0;
  wire         queue_6_deq_bits_decodeResult_other;
  wire         queue_6_deq_bits_decodeResult_multiCycle;
  wire         queue_6_deq_bits_decodeResult_divider;
  wire         queue_6_deq_bits_decodeResult_multiplier;
  wire         queue_6_deq_bits_decodeResult_shift;
  wire         queue_6_deq_bits_decodeResult_adder;
  wire         queue_6_deq_bits_decodeResult_logic;
  wire         queue_6_deq_bits_loadStore;
  wire         queue_6_deq_bits_issueInst;
  wire         queue_6_deq_bits_store;
  wire         queue_6_deq_bits_special;
  wire         queue_6_deq_bits_lsWholeReg;
  wire [4:0]   queue_6_deq_bits_vs1;
  wire [4:0]   queue_6_deq_bits_vs2;
  wire [4:0]   queue_6_deq_bits_vd;
  wire [1:0]   queue_6_deq_bits_loadStoreEEW;
  wire         queue_6_deq_bits_mask;
  wire [2:0]   queue_6_deq_bits_segment;
  wire [31:0]  queue_6_deq_bits_readFromScalar;
  wire [11:0]  queue_6_deq_bits_csrInterface_vl;
  wire [11:0]  queue_6_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_6_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_6_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_6_deq_bits_csrInterface_vxrm;
  wire         queue_6_deq_bits_csrInterface_vta;
  wire         queue_6_deq_bits_csrInterface_vma;
  wire         queue_7_deq_ready = laneRequestSinkWire_7_ready;
  wire         queue_7_deq_valid;
  wire [2:0]   queue_7_deq_bits_instructionIndex;
  wire         queue_7_deq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_7_deq_bits_decodeResult_topUop;
  wire         queue_7_deq_bits_decodeResult_popCount;
  wire         queue_7_deq_bits_decodeResult_ffo;
  wire         queue_7_deq_bits_decodeResult_average;
  wire         queue_7_deq_bits_decodeResult_reverse;
  wire         queue_7_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_7_deq_bits_decodeResult_scheduler;
  wire         queue_7_deq_bits_decodeResult_sReadVD;
  wire         queue_7_deq_bits_decodeResult_vtype;
  wire         queue_7_deq_bits_decodeResult_sWrite;
  wire         queue_7_deq_bits_decodeResult_crossRead;
  wire         queue_7_deq_bits_decodeResult_crossWrite;
  wire         queue_7_deq_bits_decodeResult_maskUnit;
  wire         queue_7_deq_bits_decodeResult_special;
  wire         queue_7_deq_bits_decodeResult_saturate;
  wire         queue_7_deq_bits_decodeResult_vwmacc;
  wire         queue_7_deq_bits_decodeResult_readOnly;
  wire         queue_7_deq_bits_decodeResult_maskSource;
  wire         queue_7_deq_bits_decodeResult_maskDestination;
  wire         queue_7_deq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_7_deq_bits_decodeResult_uop;
  wire         queue_7_deq_bits_decodeResult_iota;
  wire         queue_7_deq_bits_decodeResult_mv;
  wire         queue_7_deq_bits_decodeResult_extend;
  wire         queue_7_deq_bits_decodeResult_unOrderWrite;
  wire         queue_7_deq_bits_decodeResult_compress;
  wire         queue_7_deq_bits_decodeResult_gather16;
  wire         queue_7_deq_bits_decodeResult_gather;
  wire         queue_7_deq_bits_decodeResult_slid;
  wire         queue_7_deq_bits_decodeResult_targetRd;
  wire         queue_7_deq_bits_decodeResult_widenReduce;
  wire         queue_7_deq_bits_decodeResult_red;
  wire         queue_7_deq_bits_decodeResult_nr;
  wire         queue_7_deq_bits_decodeResult_itype;
  wire         queue_7_deq_bits_decodeResult_unsigned1;
  wire         queue_7_deq_bits_decodeResult_unsigned0;
  wire         queue_7_deq_bits_decodeResult_other;
  wire         queue_7_deq_bits_decodeResult_multiCycle;
  wire         queue_7_deq_bits_decodeResult_divider;
  wire         queue_7_deq_bits_decodeResult_multiplier;
  wire         queue_7_deq_bits_decodeResult_shift;
  wire         queue_7_deq_bits_decodeResult_adder;
  wire         queue_7_deq_bits_decodeResult_logic;
  wire         queue_7_deq_bits_loadStore;
  wire         queue_7_deq_bits_issueInst;
  wire         queue_7_deq_bits_store;
  wire         queue_7_deq_bits_special;
  wire         queue_7_deq_bits_lsWholeReg;
  wire [4:0]   queue_7_deq_bits_vs1;
  wire [4:0]   queue_7_deq_bits_vs2;
  wire [4:0]   queue_7_deq_bits_vd;
  wire [1:0]   queue_7_deq_bits_loadStoreEEW;
  wire         queue_7_deq_bits_mask;
  wire [2:0]   queue_7_deq_bits_segment;
  wire [31:0]  queue_7_deq_bits_readFromScalar;
  wire [11:0]  queue_7_deq_bits_csrInterface_vl;
  wire [11:0]  queue_7_deq_bits_csrInterface_vStart;
  wire [2:0]   queue_7_deq_bits_csrInterface_vlmul;
  wire [1:0]   queue_7_deq_bits_csrInterface_vSew;
  wire [1:0]   queue_7_deq_bits_csrInterface_vxrm;
  wire         queue_7_deq_bits_csrInterface_vta;
  wire         queue_7_deq_bits_csrInterface_vma;
  wire         validSink_valid;
  wire [2:0]   validSink_bits_instructionIndex;
  wire         validSink_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_bits_decodeResult_topUop;
  wire         validSink_bits_decodeResult_popCount;
  wire         validSink_bits_decodeResult_ffo;
  wire         validSink_bits_decodeResult_average;
  wire         validSink_bits_decodeResult_reverse;
  wire         validSink_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_bits_decodeResult_scheduler;
  wire         validSink_bits_decodeResult_sReadVD;
  wire         validSink_bits_decodeResult_vtype;
  wire         validSink_bits_decodeResult_sWrite;
  wire         validSink_bits_decodeResult_crossRead;
  wire         validSink_bits_decodeResult_crossWrite;
  wire         validSink_bits_decodeResult_maskUnit;
  wire         validSink_bits_decodeResult_special;
  wire         validSink_bits_decodeResult_saturate;
  wire         validSink_bits_decodeResult_vwmacc;
  wire         validSink_bits_decodeResult_readOnly;
  wire         validSink_bits_decodeResult_maskSource;
  wire         validSink_bits_decodeResult_maskDestination;
  wire         validSink_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_bits_decodeResult_uop;
  wire         validSink_bits_decodeResult_iota;
  wire         validSink_bits_decodeResult_mv;
  wire         validSink_bits_decodeResult_extend;
  wire         validSink_bits_decodeResult_unOrderWrite;
  wire         validSink_bits_decodeResult_compress;
  wire         validSink_bits_decodeResult_gather16;
  wire         validSink_bits_decodeResult_gather;
  wire         validSink_bits_decodeResult_slid;
  wire         validSink_bits_decodeResult_targetRd;
  wire         validSink_bits_decodeResult_widenReduce;
  wire         validSink_bits_decodeResult_red;
  wire         validSink_bits_decodeResult_nr;
  wire         validSink_bits_decodeResult_itype;
  wire         validSink_bits_decodeResult_unsigned1;
  wire         validSink_bits_decodeResult_unsigned0;
  wire         validSink_bits_decodeResult_other;
  wire         validSink_bits_decodeResult_multiCycle;
  wire         validSink_bits_decodeResult_divider;
  wire         validSink_bits_decodeResult_multiplier;
  wire         validSink_bits_decodeResult_shift;
  wire         validSink_bits_decodeResult_adder;
  wire         validSink_bits_decodeResult_logic;
  wire         validSink_bits_loadStore;
  wire         validSink_bits_issueInst;
  wire         validSink_bits_store;
  wire         validSink_bits_special;
  wire         validSink_bits_lsWholeReg;
  wire [4:0]   validSink_bits_vs1;
  wire [4:0]   validSink_bits_vs2;
  wire [4:0]   validSink_bits_vd;
  wire [1:0]   validSink_bits_loadStoreEEW;
  wire         validSink_bits_mask;
  wire [2:0]   validSink_bits_segment;
  wire [31:0]  validSink_bits_readFromScalar;
  wire [11:0]  validSink_bits_csrInterface_vl;
  wire [11:0]  validSink_bits_csrInterface_vStart;
  wire [2:0]   validSink_bits_csrInterface_vlmul;
  wire [1:0]   validSink_bits_csrInterface_vSew;
  wire [1:0]   validSink_bits_csrInterface_vxrm;
  wire         validSink_bits_csrInterface_vta;
  wire         validSink_bits_csrInterface_vma;
  wire         laneRequestSinkWire_0_valid = queue_deq_valid;
  wire [2:0]   laneRequestSinkWire_0_bits_instructionIndex = queue_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_0_bits_decodeResult_specialSlot = queue_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_0_bits_decodeResult_topUop = queue_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_0_bits_decodeResult_popCount = queue_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_0_bits_decodeResult_ffo = queue_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_0_bits_decodeResult_average = queue_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_0_bits_decodeResult_reverse = queue_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_0_bits_decodeResult_dontNeedExecuteInLane = queue_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_0_bits_decodeResult_scheduler = queue_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_0_bits_decodeResult_sReadVD = queue_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_0_bits_decodeResult_vtype = queue_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_0_bits_decodeResult_sWrite = queue_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_0_bits_decodeResult_crossRead = queue_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_0_bits_decodeResult_crossWrite = queue_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_0_bits_decodeResult_maskUnit = queue_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_0_bits_decodeResult_special = queue_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_0_bits_decodeResult_saturate = queue_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_0_bits_decodeResult_vwmacc = queue_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_0_bits_decodeResult_readOnly = queue_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_0_bits_decodeResult_maskSource = queue_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_0_bits_decodeResult_maskDestination = queue_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_0_bits_decodeResult_maskLogic = queue_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_0_bits_decodeResult_uop = queue_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_0_bits_decodeResult_iota = queue_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_0_bits_decodeResult_mv = queue_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_0_bits_decodeResult_extend = queue_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_0_bits_decodeResult_unOrderWrite = queue_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_0_bits_decodeResult_compress = queue_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_0_bits_decodeResult_gather16 = queue_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_0_bits_decodeResult_gather = queue_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_0_bits_decodeResult_slid = queue_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_0_bits_decodeResult_targetRd = queue_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_0_bits_decodeResult_widenReduce = queue_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_0_bits_decodeResult_red = queue_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_0_bits_decodeResult_nr = queue_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_0_bits_decodeResult_itype = queue_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_0_bits_decodeResult_unsigned1 = queue_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_0_bits_decodeResult_unsigned0 = queue_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_0_bits_decodeResult_other = queue_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_0_bits_decodeResult_multiCycle = queue_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_0_bits_decodeResult_divider = queue_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_0_bits_decodeResult_multiplier = queue_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_0_bits_decodeResult_shift = queue_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_0_bits_decodeResult_adder = queue_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_0_bits_decodeResult_logic = queue_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_0_bits_loadStore = queue_deq_bits_loadStore;
  wire         laneRequestSinkWire_0_bits_issueInst = queue_deq_bits_issueInst;
  wire         laneRequestSinkWire_0_bits_store = queue_deq_bits_store;
  wire         laneRequestSinkWire_0_bits_special = queue_deq_bits_special;
  wire         laneRequestSinkWire_0_bits_lsWholeReg = queue_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_0_bits_vs1 = queue_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_0_bits_vs2 = queue_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_0_bits_vd = queue_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_0_bits_loadStoreEEW = queue_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_0_bits_mask = queue_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_0_bits_segment = queue_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_0_bits_readFromScalar = queue_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_0_bits_csrInterface_vl = queue_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_0_bits_csrInterface_vStart = queue_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_0_bits_csrInterface_vlmul = queue_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_0_bits_csrInterface_vSew = queue_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_0_bits_csrInterface_vxrm = queue_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_0_bits_csrInterface_vta = queue_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_0_bits_csrInterface_vma = queue_deq_bits_csrInterface_vma;
  wire [1:0]   queue_enq_bits_csrInterface_vxrm;
  wire         queue_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi = {queue_enq_bits_csrInterface_vxrm, queue_enq_bits_csrInterface_vta};
  wire         queue_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo = {queue_dataIn_lo_hi, queue_enq_bits_csrInterface_vma};
  wire [2:0]   queue_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo = {queue_enq_bits_csrInterface_vlmul, queue_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_enq_bits_csrInterface_vl;
  wire [11:0]  queue_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi = {queue_enq_bits_csrInterface_vl, queue_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi = {queue_dataIn_hi_hi, queue_dataIn_hi_lo};
  wire         queue_enq_bits_decodeResult_adder;
  wire         queue_enq_bits_decodeResult_logic;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo = {queue_enq_bits_decodeResult_adder, queue_enq_bits_decodeResult_logic};
  wire         queue_enq_bits_decodeResult_divider;
  wire         queue_enq_bits_decodeResult_multiplier;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi = {queue_enq_bits_decodeResult_divider, queue_enq_bits_decodeResult_multiplier};
  wire         queue_enq_bits_decodeResult_shift;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi = {queue_dataIn_lo_lo_lo_hi_hi, queue_enq_bits_decodeResult_shift};
  wire [4:0]   queue_dataIn_lo_lo_lo = {queue_dataIn_lo_lo_lo_hi, queue_dataIn_lo_lo_lo_lo};
  wire         queue_enq_bits_decodeResult_unsigned0;
  wire         queue_enq_bits_decodeResult_other;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi = {queue_enq_bits_decodeResult_unsigned0, queue_enq_bits_decodeResult_other};
  wire         queue_enq_bits_decodeResult_multiCycle;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo = {queue_dataIn_lo_lo_hi_lo_hi, queue_enq_bits_decodeResult_multiCycle};
  wire         queue_enq_bits_decodeResult_nr;
  wire         queue_enq_bits_decodeResult_itype;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi = {queue_enq_bits_decodeResult_nr, queue_enq_bits_decodeResult_itype};
  wire         queue_enq_bits_decodeResult_unsigned1;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi = {queue_dataIn_lo_lo_hi_hi_hi, queue_enq_bits_decodeResult_unsigned1};
  wire [5:0]   queue_dataIn_lo_lo_hi = {queue_dataIn_lo_lo_hi_hi, queue_dataIn_lo_lo_hi_lo};
  wire [10:0]  queue_dataIn_lo_lo = {queue_dataIn_lo_lo_hi, queue_dataIn_lo_lo_lo};
  wire         queue_enq_bits_decodeResult_widenReduce;
  wire         queue_enq_bits_decodeResult_red;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo = {queue_enq_bits_decodeResult_widenReduce, queue_enq_bits_decodeResult_red};
  wire         queue_enq_bits_decodeResult_gather;
  wire         queue_enq_bits_decodeResult_slid;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi = {queue_enq_bits_decodeResult_gather, queue_enq_bits_decodeResult_slid};
  wire         queue_enq_bits_decodeResult_targetRd;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi = {queue_dataIn_lo_hi_lo_hi_hi, queue_enq_bits_decodeResult_targetRd};
  wire [4:0]   queue_dataIn_lo_hi_lo = {queue_dataIn_lo_hi_lo_hi, queue_dataIn_lo_hi_lo_lo};
  wire         queue_enq_bits_decodeResult_unOrderWrite;
  wire         queue_enq_bits_decodeResult_compress;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi = {queue_enq_bits_decodeResult_unOrderWrite, queue_enq_bits_decodeResult_compress};
  wire         queue_enq_bits_decodeResult_gather16;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo = {queue_dataIn_lo_hi_hi_lo_hi, queue_enq_bits_decodeResult_gather16};
  wire         queue_enq_bits_decodeResult_iota;
  wire         queue_enq_bits_decodeResult_mv;
  wire [1:0]   queue_dataIn_lo_hi_hi_hi_hi = {queue_enq_bits_decodeResult_iota, queue_enq_bits_decodeResult_mv};
  wire         queue_enq_bits_decodeResult_extend;
  wire [2:0]   queue_dataIn_lo_hi_hi_hi = {queue_dataIn_lo_hi_hi_hi_hi, queue_enq_bits_decodeResult_extend};
  wire [5:0]   queue_dataIn_lo_hi_hi = {queue_dataIn_lo_hi_hi_hi, queue_dataIn_lo_hi_hi_lo};
  wire [10:0]  queue_dataIn_lo_hi_1 = {queue_dataIn_lo_hi_hi, queue_dataIn_lo_hi_lo};
  wire [21:0]  queue_dataIn_lo_1 = {queue_dataIn_lo_hi_1, queue_dataIn_lo_lo};
  wire         queue_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_hi_lo_lo_lo = {queue_enq_bits_decodeResult_maskLogic, queue_enq_bits_decodeResult_uop};
  wire         queue_enq_bits_decodeResult_readOnly;
  wire         queue_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi = {queue_enq_bits_decodeResult_readOnly, queue_enq_bits_decodeResult_maskSource};
  wire         queue_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi = {queue_dataIn_hi_lo_lo_hi_hi, queue_enq_bits_decodeResult_maskDestination};
  wire [7:0]   queue_dataIn_hi_lo_lo = {queue_dataIn_hi_lo_lo_hi, queue_dataIn_hi_lo_lo_lo};
  wire         queue_enq_bits_decodeResult_special;
  wire         queue_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi = {queue_enq_bits_decodeResult_special, queue_enq_bits_decodeResult_saturate};
  wire         queue_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo = {queue_dataIn_hi_lo_hi_lo_hi, queue_enq_bits_decodeResult_vwmacc};
  wire         queue_enq_bits_decodeResult_crossRead;
  wire         queue_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi = {queue_enq_bits_decodeResult_crossRead, queue_enq_bits_decodeResult_crossWrite};
  wire         queue_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi = {queue_dataIn_hi_lo_hi_hi_hi, queue_enq_bits_decodeResult_maskUnit};
  wire [5:0]   queue_dataIn_hi_lo_hi = {queue_dataIn_hi_lo_hi_hi, queue_dataIn_hi_lo_hi_lo};
  wire [13:0]  queue_dataIn_hi_lo_1 = {queue_dataIn_hi_lo_hi, queue_dataIn_hi_lo_lo};
  wire         queue_enq_bits_decodeResult_vtype;
  wire         queue_enq_bits_decodeResult_sWrite;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo = {queue_enq_bits_decodeResult_vtype, queue_enq_bits_decodeResult_sWrite};
  wire         queue_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_enq_bits_decodeResult_scheduler;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi = {queue_enq_bits_decodeResult_dontNeedExecuteInLane, queue_enq_bits_decodeResult_scheduler};
  wire         queue_enq_bits_decodeResult_sReadVD;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi = {queue_dataIn_hi_hi_lo_hi_hi, queue_enq_bits_decodeResult_sReadVD};
  wire [4:0]   queue_dataIn_hi_hi_lo = {queue_dataIn_hi_hi_lo_hi, queue_dataIn_hi_hi_lo_lo};
  wire         queue_enq_bits_decodeResult_ffo;
  wire         queue_enq_bits_decodeResult_average;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi = {queue_enq_bits_decodeResult_ffo, queue_enq_bits_decodeResult_average};
  wire         queue_enq_bits_decodeResult_reverse;
  wire [2:0]   queue_dataIn_hi_hi_hi_lo = {queue_dataIn_hi_hi_hi_lo_hi, queue_enq_bits_decodeResult_reverse};
  wire         queue_enq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_enq_bits_decodeResult_topUop;
  wire [5:0]   queue_dataIn_hi_hi_hi_hi_hi = {queue_enq_bits_decodeResult_specialSlot, queue_enq_bits_decodeResult_topUop};
  wire         queue_enq_bits_decodeResult_popCount;
  wire [6:0]   queue_dataIn_hi_hi_hi_hi = {queue_dataIn_hi_hi_hi_hi_hi, queue_enq_bits_decodeResult_popCount};
  wire [9:0]   queue_dataIn_hi_hi_hi = {queue_dataIn_hi_hi_hi_hi, queue_dataIn_hi_hi_hi_lo};
  wire [14:0]  queue_dataIn_hi_hi_1 = {queue_dataIn_hi_hi_hi, queue_dataIn_hi_hi_lo};
  wire [28:0]  queue_dataIn_hi_1 = {queue_dataIn_hi_hi_1, queue_dataIn_hi_lo_1};
  wire [2:0]   queue_enq_bits_segment;
  wire [31:0]  queue_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_1 = {queue_enq_bits_segment, queue_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_1 = {queue_dataIn_lo_lo_hi_1, queue_dataIn_hi, queue_dataIn_lo};
  wire [1:0]   queue_enq_bits_loadStoreEEW;
  wire         queue_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_1 = {queue_enq_bits_loadStoreEEW, queue_enq_bits_mask};
  wire [4:0]   queue_enq_bits_vs2;
  wire [4:0]   queue_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_1 = {queue_enq_bits_vs2, queue_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_2 = {queue_dataIn_lo_hi_hi_1, queue_dataIn_lo_hi_lo_1};
  wire [80:0]  queue_dataIn_lo_2 = {queue_dataIn_lo_hi_2, queue_dataIn_lo_lo_1};
  wire         queue_enq_bits_lsWholeReg;
  wire [4:0]   queue_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_1 = {queue_enq_bits_lsWholeReg, queue_enq_bits_vs1};
  wire         queue_enq_bits_store;
  wire         queue_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_1 = {queue_enq_bits_store, queue_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_2 = {queue_dataIn_hi_lo_hi_1, queue_dataIn_hi_lo_lo_1};
  wire         queue_enq_bits_loadStore;
  wire         queue_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_1 = {queue_enq_bits_loadStore, queue_enq_bits_issueInst};
  wire [2:0]   queue_enq_bits_instructionIndex;
  wire [53:0]  queue_dataIn_hi_hi_hi_1 = {queue_enq_bits_instructionIndex, queue_dataIn_hi_1, queue_dataIn_lo_1};
  wire [55:0]  queue_dataIn_hi_hi_2 = {queue_dataIn_hi_hi_hi_1, queue_dataIn_hi_hi_lo_1};
  wire [63:0]  queue_dataIn_hi_2 = {queue_dataIn_hi_hi_2, queue_dataIn_hi_lo_2};
  wire [144:0] queue_dataIn = {queue_dataIn_hi_2, queue_dataIn_lo_2};
  wire         queue_dataOut_csrInterface_vma = _queue_fifo_data_out[0];
  wire         queue_dataOut_csrInterface_vta = _queue_fifo_data_out[1];
  wire [1:0]   queue_dataOut_csrInterface_vxrm = _queue_fifo_data_out[3:2];
  wire [1:0]   queue_dataOut_csrInterface_vSew = _queue_fifo_data_out[5:4];
  wire [2:0]   queue_dataOut_csrInterface_vlmul = _queue_fifo_data_out[8:6];
  wire [11:0]  queue_dataOut_csrInterface_vStart = _queue_fifo_data_out[20:9];
  wire [11:0]  queue_dataOut_csrInterface_vl = _queue_fifo_data_out[32:21];
  wire [31:0]  queue_dataOut_readFromScalar = _queue_fifo_data_out[64:33];
  wire [2:0]   queue_dataOut_segment = _queue_fifo_data_out[67:65];
  wire         queue_dataOut_mask = _queue_fifo_data_out[68];
  wire [1:0]   queue_dataOut_loadStoreEEW = _queue_fifo_data_out[70:69];
  wire [4:0]   queue_dataOut_vd = _queue_fifo_data_out[75:71];
  wire [4:0]   queue_dataOut_vs2 = _queue_fifo_data_out[80:76];
  wire [4:0]   queue_dataOut_vs1 = _queue_fifo_data_out[85:81];
  wire         queue_dataOut_lsWholeReg = _queue_fifo_data_out[86];
  wire         queue_dataOut_special = _queue_fifo_data_out[87];
  wire         queue_dataOut_store = _queue_fifo_data_out[88];
  wire         queue_dataOut_issueInst = _queue_fifo_data_out[89];
  wire         queue_dataOut_loadStore = _queue_fifo_data_out[90];
  wire         queue_dataOut_decodeResult_logic = _queue_fifo_data_out[91];
  wire         queue_dataOut_decodeResult_adder = _queue_fifo_data_out[92];
  wire         queue_dataOut_decodeResult_shift = _queue_fifo_data_out[93];
  wire         queue_dataOut_decodeResult_multiplier = _queue_fifo_data_out[94];
  wire         queue_dataOut_decodeResult_divider = _queue_fifo_data_out[95];
  wire         queue_dataOut_decodeResult_multiCycle = _queue_fifo_data_out[96];
  wire         queue_dataOut_decodeResult_other = _queue_fifo_data_out[97];
  wire         queue_dataOut_decodeResult_unsigned0 = _queue_fifo_data_out[98];
  wire         queue_dataOut_decodeResult_unsigned1 = _queue_fifo_data_out[99];
  wire         queue_dataOut_decodeResult_itype = _queue_fifo_data_out[100];
  wire         queue_dataOut_decodeResult_nr = _queue_fifo_data_out[101];
  wire         queue_dataOut_decodeResult_red = _queue_fifo_data_out[102];
  wire         queue_dataOut_decodeResult_widenReduce = _queue_fifo_data_out[103];
  wire         queue_dataOut_decodeResult_targetRd = _queue_fifo_data_out[104];
  wire         queue_dataOut_decodeResult_slid = _queue_fifo_data_out[105];
  wire         queue_dataOut_decodeResult_gather = _queue_fifo_data_out[106];
  wire         queue_dataOut_decodeResult_gather16 = _queue_fifo_data_out[107];
  wire         queue_dataOut_decodeResult_compress = _queue_fifo_data_out[108];
  wire         queue_dataOut_decodeResult_unOrderWrite = _queue_fifo_data_out[109];
  wire         queue_dataOut_decodeResult_extend = _queue_fifo_data_out[110];
  wire         queue_dataOut_decodeResult_mv = _queue_fifo_data_out[111];
  wire         queue_dataOut_decodeResult_iota = _queue_fifo_data_out[112];
  wire [3:0]   queue_dataOut_decodeResult_uop = _queue_fifo_data_out[116:113];
  wire         queue_dataOut_decodeResult_maskLogic = _queue_fifo_data_out[117];
  wire         queue_dataOut_decodeResult_maskDestination = _queue_fifo_data_out[118];
  wire         queue_dataOut_decodeResult_maskSource = _queue_fifo_data_out[119];
  wire         queue_dataOut_decodeResult_readOnly = _queue_fifo_data_out[120];
  wire         queue_dataOut_decodeResult_vwmacc = _queue_fifo_data_out[121];
  wire         queue_dataOut_decodeResult_saturate = _queue_fifo_data_out[122];
  wire         queue_dataOut_decodeResult_special = _queue_fifo_data_out[123];
  wire         queue_dataOut_decodeResult_maskUnit = _queue_fifo_data_out[124];
  wire         queue_dataOut_decodeResult_crossWrite = _queue_fifo_data_out[125];
  wire         queue_dataOut_decodeResult_crossRead = _queue_fifo_data_out[126];
  wire         queue_dataOut_decodeResult_sWrite = _queue_fifo_data_out[127];
  wire         queue_dataOut_decodeResult_vtype = _queue_fifo_data_out[128];
  wire         queue_dataOut_decodeResult_sReadVD = _queue_fifo_data_out[129];
  wire         queue_dataOut_decodeResult_scheduler = _queue_fifo_data_out[130];
  wire         queue_dataOut_decodeResult_dontNeedExecuteInLane = _queue_fifo_data_out[131];
  wire         queue_dataOut_decodeResult_reverse = _queue_fifo_data_out[132];
  wire         queue_dataOut_decodeResult_average = _queue_fifo_data_out[133];
  wire         queue_dataOut_decodeResult_ffo = _queue_fifo_data_out[134];
  wire         queue_dataOut_decodeResult_popCount = _queue_fifo_data_out[135];
  wire [4:0]   queue_dataOut_decodeResult_topUop = _queue_fifo_data_out[140:136];
  wire         queue_dataOut_decodeResult_specialSlot = _queue_fifo_data_out[141];
  wire [2:0]   queue_dataOut_instructionIndex = _queue_fifo_data_out[144:142];
  wire         queue_enq_ready = ~_queue_fifo_full;
  wire         queue_enq_valid;
  assign queue_deq_valid = ~_queue_fifo_empty | queue_enq_valid;
  assign queue_deq_bits_instructionIndex = _queue_fifo_empty ? queue_enq_bits_instructionIndex : queue_dataOut_instructionIndex;
  assign queue_deq_bits_decodeResult_specialSlot = _queue_fifo_empty ? queue_enq_bits_decodeResult_specialSlot : queue_dataOut_decodeResult_specialSlot;
  assign queue_deq_bits_decodeResult_topUop = _queue_fifo_empty ? queue_enq_bits_decodeResult_topUop : queue_dataOut_decodeResult_topUop;
  assign queue_deq_bits_decodeResult_popCount = _queue_fifo_empty ? queue_enq_bits_decodeResult_popCount : queue_dataOut_decodeResult_popCount;
  assign queue_deq_bits_decodeResult_ffo = _queue_fifo_empty ? queue_enq_bits_decodeResult_ffo : queue_dataOut_decodeResult_ffo;
  assign queue_deq_bits_decodeResult_average = _queue_fifo_empty ? queue_enq_bits_decodeResult_average : queue_dataOut_decodeResult_average;
  assign queue_deq_bits_decodeResult_reverse = _queue_fifo_empty ? queue_enq_bits_decodeResult_reverse : queue_dataOut_decodeResult_reverse;
  assign queue_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_empty ? queue_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_decodeResult_dontNeedExecuteInLane;
  assign queue_deq_bits_decodeResult_scheduler = _queue_fifo_empty ? queue_enq_bits_decodeResult_scheduler : queue_dataOut_decodeResult_scheduler;
  assign queue_deq_bits_decodeResult_sReadVD = _queue_fifo_empty ? queue_enq_bits_decodeResult_sReadVD : queue_dataOut_decodeResult_sReadVD;
  assign queue_deq_bits_decodeResult_vtype = _queue_fifo_empty ? queue_enq_bits_decodeResult_vtype : queue_dataOut_decodeResult_vtype;
  assign queue_deq_bits_decodeResult_sWrite = _queue_fifo_empty ? queue_enq_bits_decodeResult_sWrite : queue_dataOut_decodeResult_sWrite;
  assign queue_deq_bits_decodeResult_crossRead = _queue_fifo_empty ? queue_enq_bits_decodeResult_crossRead : queue_dataOut_decodeResult_crossRead;
  assign queue_deq_bits_decodeResult_crossWrite = _queue_fifo_empty ? queue_enq_bits_decodeResult_crossWrite : queue_dataOut_decodeResult_crossWrite;
  assign queue_deq_bits_decodeResult_maskUnit = _queue_fifo_empty ? queue_enq_bits_decodeResult_maskUnit : queue_dataOut_decodeResult_maskUnit;
  assign queue_deq_bits_decodeResult_special = _queue_fifo_empty ? queue_enq_bits_decodeResult_special : queue_dataOut_decodeResult_special;
  assign queue_deq_bits_decodeResult_saturate = _queue_fifo_empty ? queue_enq_bits_decodeResult_saturate : queue_dataOut_decodeResult_saturate;
  assign queue_deq_bits_decodeResult_vwmacc = _queue_fifo_empty ? queue_enq_bits_decodeResult_vwmacc : queue_dataOut_decodeResult_vwmacc;
  assign queue_deq_bits_decodeResult_readOnly = _queue_fifo_empty ? queue_enq_bits_decodeResult_readOnly : queue_dataOut_decodeResult_readOnly;
  assign queue_deq_bits_decodeResult_maskSource = _queue_fifo_empty ? queue_enq_bits_decodeResult_maskSource : queue_dataOut_decodeResult_maskSource;
  assign queue_deq_bits_decodeResult_maskDestination = _queue_fifo_empty ? queue_enq_bits_decodeResult_maskDestination : queue_dataOut_decodeResult_maskDestination;
  assign queue_deq_bits_decodeResult_maskLogic = _queue_fifo_empty ? queue_enq_bits_decodeResult_maskLogic : queue_dataOut_decodeResult_maskLogic;
  assign queue_deq_bits_decodeResult_uop = _queue_fifo_empty ? queue_enq_bits_decodeResult_uop : queue_dataOut_decodeResult_uop;
  assign queue_deq_bits_decodeResult_iota = _queue_fifo_empty ? queue_enq_bits_decodeResult_iota : queue_dataOut_decodeResult_iota;
  assign queue_deq_bits_decodeResult_mv = _queue_fifo_empty ? queue_enq_bits_decodeResult_mv : queue_dataOut_decodeResult_mv;
  assign queue_deq_bits_decodeResult_extend = _queue_fifo_empty ? queue_enq_bits_decodeResult_extend : queue_dataOut_decodeResult_extend;
  assign queue_deq_bits_decodeResult_unOrderWrite = _queue_fifo_empty ? queue_enq_bits_decodeResult_unOrderWrite : queue_dataOut_decodeResult_unOrderWrite;
  assign queue_deq_bits_decodeResult_compress = _queue_fifo_empty ? queue_enq_bits_decodeResult_compress : queue_dataOut_decodeResult_compress;
  assign queue_deq_bits_decodeResult_gather16 = _queue_fifo_empty ? queue_enq_bits_decodeResult_gather16 : queue_dataOut_decodeResult_gather16;
  assign queue_deq_bits_decodeResult_gather = _queue_fifo_empty ? queue_enq_bits_decodeResult_gather : queue_dataOut_decodeResult_gather;
  assign queue_deq_bits_decodeResult_slid = _queue_fifo_empty ? queue_enq_bits_decodeResult_slid : queue_dataOut_decodeResult_slid;
  assign queue_deq_bits_decodeResult_targetRd = _queue_fifo_empty ? queue_enq_bits_decodeResult_targetRd : queue_dataOut_decodeResult_targetRd;
  assign queue_deq_bits_decodeResult_widenReduce = _queue_fifo_empty ? queue_enq_bits_decodeResult_widenReduce : queue_dataOut_decodeResult_widenReduce;
  assign queue_deq_bits_decodeResult_red = _queue_fifo_empty ? queue_enq_bits_decodeResult_red : queue_dataOut_decodeResult_red;
  assign queue_deq_bits_decodeResult_nr = _queue_fifo_empty ? queue_enq_bits_decodeResult_nr : queue_dataOut_decodeResult_nr;
  assign queue_deq_bits_decodeResult_itype = _queue_fifo_empty ? queue_enq_bits_decodeResult_itype : queue_dataOut_decodeResult_itype;
  assign queue_deq_bits_decodeResult_unsigned1 = _queue_fifo_empty ? queue_enq_bits_decodeResult_unsigned1 : queue_dataOut_decodeResult_unsigned1;
  assign queue_deq_bits_decodeResult_unsigned0 = _queue_fifo_empty ? queue_enq_bits_decodeResult_unsigned0 : queue_dataOut_decodeResult_unsigned0;
  assign queue_deq_bits_decodeResult_other = _queue_fifo_empty ? queue_enq_bits_decodeResult_other : queue_dataOut_decodeResult_other;
  assign queue_deq_bits_decodeResult_multiCycle = _queue_fifo_empty ? queue_enq_bits_decodeResult_multiCycle : queue_dataOut_decodeResult_multiCycle;
  assign queue_deq_bits_decodeResult_divider = _queue_fifo_empty ? queue_enq_bits_decodeResult_divider : queue_dataOut_decodeResult_divider;
  assign queue_deq_bits_decodeResult_multiplier = _queue_fifo_empty ? queue_enq_bits_decodeResult_multiplier : queue_dataOut_decodeResult_multiplier;
  assign queue_deq_bits_decodeResult_shift = _queue_fifo_empty ? queue_enq_bits_decodeResult_shift : queue_dataOut_decodeResult_shift;
  assign queue_deq_bits_decodeResult_adder = _queue_fifo_empty ? queue_enq_bits_decodeResult_adder : queue_dataOut_decodeResult_adder;
  assign queue_deq_bits_decodeResult_logic = _queue_fifo_empty ? queue_enq_bits_decodeResult_logic : queue_dataOut_decodeResult_logic;
  assign queue_deq_bits_loadStore = _queue_fifo_empty ? queue_enq_bits_loadStore : queue_dataOut_loadStore;
  assign queue_deq_bits_issueInst = _queue_fifo_empty ? queue_enq_bits_issueInst : queue_dataOut_issueInst;
  assign queue_deq_bits_store = _queue_fifo_empty ? queue_enq_bits_store : queue_dataOut_store;
  assign queue_deq_bits_special = _queue_fifo_empty ? queue_enq_bits_special : queue_dataOut_special;
  assign queue_deq_bits_lsWholeReg = _queue_fifo_empty ? queue_enq_bits_lsWholeReg : queue_dataOut_lsWholeReg;
  assign queue_deq_bits_vs1 = _queue_fifo_empty ? queue_enq_bits_vs1 : queue_dataOut_vs1;
  assign queue_deq_bits_vs2 = _queue_fifo_empty ? queue_enq_bits_vs2 : queue_dataOut_vs2;
  assign queue_deq_bits_vd = _queue_fifo_empty ? queue_enq_bits_vd : queue_dataOut_vd;
  assign queue_deq_bits_loadStoreEEW = _queue_fifo_empty ? queue_enq_bits_loadStoreEEW : queue_dataOut_loadStoreEEW;
  assign queue_deq_bits_mask = _queue_fifo_empty ? queue_enq_bits_mask : queue_dataOut_mask;
  assign queue_deq_bits_segment = _queue_fifo_empty ? queue_enq_bits_segment : queue_dataOut_segment;
  assign queue_deq_bits_readFromScalar = _queue_fifo_empty ? queue_enq_bits_readFromScalar : queue_dataOut_readFromScalar;
  assign queue_deq_bits_csrInterface_vl = _queue_fifo_empty ? queue_enq_bits_csrInterface_vl : queue_dataOut_csrInterface_vl;
  assign queue_deq_bits_csrInterface_vStart = _queue_fifo_empty ? queue_enq_bits_csrInterface_vStart : queue_dataOut_csrInterface_vStart;
  assign queue_deq_bits_csrInterface_vlmul = _queue_fifo_empty ? queue_enq_bits_csrInterface_vlmul : queue_dataOut_csrInterface_vlmul;
  assign queue_deq_bits_csrInterface_vSew = _queue_fifo_empty ? queue_enq_bits_csrInterface_vSew : queue_dataOut_csrInterface_vSew;
  assign queue_deq_bits_csrInterface_vxrm = _queue_fifo_empty ? queue_enq_bits_csrInterface_vxrm : queue_dataOut_csrInterface_vxrm;
  assign queue_deq_bits_csrInterface_vta = _queue_fifo_empty ? queue_enq_bits_csrInterface_vta : queue_dataOut_csrInterface_vta;
  assign queue_deq_bits_csrInterface_vma = _queue_fifo_empty ? queue_enq_bits_csrInterface_vma : queue_dataOut_csrInterface_vma;
  wire         laneVec_0_laneRequest_bits_issueInst = laneRequestSinkWire_0_ready & laneRequestSinkWire_0_valid;
  reg          releasePipe_pipe_v;
  wire         releasePipe_pipe_out_valid = releasePipe_pipe_v;
  wire         laneRequestSourceWire_0_ready;
  wire         validSource_valid = laneRequestSourceWire_0_ready & laneRequestSourceWire_0_valid;
  reg  [2:0]   tokenCheck_counter;
  wire [2:0]   tokenCheck_counterChange = validSource_valid ? 3'h1 : 3'h7;
  assign tokenCheck = ~(tokenCheck_counter[2]);
  assign laneRequestSourceWire_0_ready = tokenCheck;
  assign queue_enq_valid = validSink_valid;
  assign queue_enq_bits_instructionIndex = validSink_bits_instructionIndex;
  assign queue_enq_bits_decodeResult_specialSlot = validSink_bits_decodeResult_specialSlot;
  assign queue_enq_bits_decodeResult_topUop = validSink_bits_decodeResult_topUop;
  assign queue_enq_bits_decodeResult_popCount = validSink_bits_decodeResult_popCount;
  assign queue_enq_bits_decodeResult_ffo = validSink_bits_decodeResult_ffo;
  assign queue_enq_bits_decodeResult_average = validSink_bits_decodeResult_average;
  assign queue_enq_bits_decodeResult_reverse = validSink_bits_decodeResult_reverse;
  assign queue_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_enq_bits_decodeResult_scheduler = validSink_bits_decodeResult_scheduler;
  assign queue_enq_bits_decodeResult_sReadVD = validSink_bits_decodeResult_sReadVD;
  assign queue_enq_bits_decodeResult_vtype = validSink_bits_decodeResult_vtype;
  assign queue_enq_bits_decodeResult_sWrite = validSink_bits_decodeResult_sWrite;
  assign queue_enq_bits_decodeResult_crossRead = validSink_bits_decodeResult_crossRead;
  assign queue_enq_bits_decodeResult_crossWrite = validSink_bits_decodeResult_crossWrite;
  assign queue_enq_bits_decodeResult_maskUnit = validSink_bits_decodeResult_maskUnit;
  assign queue_enq_bits_decodeResult_special = validSink_bits_decodeResult_special;
  assign queue_enq_bits_decodeResult_saturate = validSink_bits_decodeResult_saturate;
  assign queue_enq_bits_decodeResult_vwmacc = validSink_bits_decodeResult_vwmacc;
  assign queue_enq_bits_decodeResult_readOnly = validSink_bits_decodeResult_readOnly;
  assign queue_enq_bits_decodeResult_maskSource = validSink_bits_decodeResult_maskSource;
  assign queue_enq_bits_decodeResult_maskDestination = validSink_bits_decodeResult_maskDestination;
  assign queue_enq_bits_decodeResult_maskLogic = validSink_bits_decodeResult_maskLogic;
  assign queue_enq_bits_decodeResult_uop = validSink_bits_decodeResult_uop;
  assign queue_enq_bits_decodeResult_iota = validSink_bits_decodeResult_iota;
  assign queue_enq_bits_decodeResult_mv = validSink_bits_decodeResult_mv;
  assign queue_enq_bits_decodeResult_extend = validSink_bits_decodeResult_extend;
  assign queue_enq_bits_decodeResult_unOrderWrite = validSink_bits_decodeResult_unOrderWrite;
  assign queue_enq_bits_decodeResult_compress = validSink_bits_decodeResult_compress;
  assign queue_enq_bits_decodeResult_gather16 = validSink_bits_decodeResult_gather16;
  assign queue_enq_bits_decodeResult_gather = validSink_bits_decodeResult_gather;
  assign queue_enq_bits_decodeResult_slid = validSink_bits_decodeResult_slid;
  assign queue_enq_bits_decodeResult_targetRd = validSink_bits_decodeResult_targetRd;
  assign queue_enq_bits_decodeResult_widenReduce = validSink_bits_decodeResult_widenReduce;
  assign queue_enq_bits_decodeResult_red = validSink_bits_decodeResult_red;
  assign queue_enq_bits_decodeResult_nr = validSink_bits_decodeResult_nr;
  assign queue_enq_bits_decodeResult_itype = validSink_bits_decodeResult_itype;
  assign queue_enq_bits_decodeResult_unsigned1 = validSink_bits_decodeResult_unsigned1;
  assign queue_enq_bits_decodeResult_unsigned0 = validSink_bits_decodeResult_unsigned0;
  assign queue_enq_bits_decodeResult_other = validSink_bits_decodeResult_other;
  assign queue_enq_bits_decodeResult_multiCycle = validSink_bits_decodeResult_multiCycle;
  assign queue_enq_bits_decodeResult_divider = validSink_bits_decodeResult_divider;
  assign queue_enq_bits_decodeResult_multiplier = validSink_bits_decodeResult_multiplier;
  assign queue_enq_bits_decodeResult_shift = validSink_bits_decodeResult_shift;
  assign queue_enq_bits_decodeResult_adder = validSink_bits_decodeResult_adder;
  assign queue_enq_bits_decodeResult_logic = validSink_bits_decodeResult_logic;
  assign queue_enq_bits_loadStore = validSink_bits_loadStore;
  assign queue_enq_bits_issueInst = validSink_bits_issueInst;
  assign queue_enq_bits_store = validSink_bits_store;
  assign queue_enq_bits_special = validSink_bits_special;
  assign queue_enq_bits_lsWholeReg = validSink_bits_lsWholeReg;
  assign queue_enq_bits_vs1 = validSink_bits_vs1;
  assign queue_enq_bits_vs2 = validSink_bits_vs2;
  assign queue_enq_bits_vd = validSink_bits_vd;
  assign queue_enq_bits_loadStoreEEW = validSink_bits_loadStoreEEW;
  assign queue_enq_bits_mask = validSink_bits_mask;
  assign queue_enq_bits_segment = validSink_bits_segment;
  assign queue_enq_bits_readFromScalar = validSink_bits_readFromScalar;
  assign queue_enq_bits_csrInterface_vl = validSink_bits_csrInterface_vl;
  assign queue_enq_bits_csrInterface_vStart = validSink_bits_csrInterface_vStart;
  assign queue_enq_bits_csrInterface_vlmul = validSink_bits_csrInterface_vlmul;
  assign queue_enq_bits_csrInterface_vSew = validSink_bits_csrInterface_vSew;
  assign queue_enq_bits_csrInterface_vxrm = validSink_bits_csrInterface_vxrm;
  assign queue_enq_bits_csrInterface_vta = validSink_bits_csrInterface_vta;
  assign queue_enq_bits_csrInterface_vma = validSink_bits_csrInterface_vma;
  reg          shifterReg_0_valid;
  assign validSink_valid = shifterReg_0_valid;
  reg  [2:0]   shifterReg_0_bits_instructionIndex;
  assign validSink_bits_instructionIndex = shifterReg_0_bits_instructionIndex;
  reg          shifterReg_0_bits_decodeResult_specialSlot;
  assign validSink_bits_decodeResult_specialSlot = shifterReg_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_0_bits_decodeResult_topUop;
  assign validSink_bits_decodeResult_topUop = shifterReg_0_bits_decodeResult_topUop;
  reg          shifterReg_0_bits_decodeResult_popCount;
  assign validSink_bits_decodeResult_popCount = shifterReg_0_bits_decodeResult_popCount;
  reg          shifterReg_0_bits_decodeResult_ffo;
  assign validSink_bits_decodeResult_ffo = shifterReg_0_bits_decodeResult_ffo;
  reg          shifterReg_0_bits_decodeResult_average;
  assign validSink_bits_decodeResult_average = shifterReg_0_bits_decodeResult_average;
  reg          shifterReg_0_bits_decodeResult_reverse;
  assign validSink_bits_decodeResult_reverse = shifterReg_0_bits_decodeResult_reverse;
  reg          shifterReg_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_bits_decodeResult_dontNeedExecuteInLane = shifterReg_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_0_bits_decodeResult_scheduler;
  assign validSink_bits_decodeResult_scheduler = shifterReg_0_bits_decodeResult_scheduler;
  reg          shifterReg_0_bits_decodeResult_sReadVD;
  assign validSink_bits_decodeResult_sReadVD = shifterReg_0_bits_decodeResult_sReadVD;
  reg          shifterReg_0_bits_decodeResult_vtype;
  assign validSink_bits_decodeResult_vtype = shifterReg_0_bits_decodeResult_vtype;
  reg          shifterReg_0_bits_decodeResult_sWrite;
  assign validSink_bits_decodeResult_sWrite = shifterReg_0_bits_decodeResult_sWrite;
  reg          shifterReg_0_bits_decodeResult_crossRead;
  assign validSink_bits_decodeResult_crossRead = shifterReg_0_bits_decodeResult_crossRead;
  reg          shifterReg_0_bits_decodeResult_crossWrite;
  assign validSink_bits_decodeResult_crossWrite = shifterReg_0_bits_decodeResult_crossWrite;
  reg          shifterReg_0_bits_decodeResult_maskUnit;
  assign validSink_bits_decodeResult_maskUnit = shifterReg_0_bits_decodeResult_maskUnit;
  reg          shifterReg_0_bits_decodeResult_special;
  assign validSink_bits_decodeResult_special = shifterReg_0_bits_decodeResult_special;
  reg          shifterReg_0_bits_decodeResult_saturate;
  assign validSink_bits_decodeResult_saturate = shifterReg_0_bits_decodeResult_saturate;
  reg          shifterReg_0_bits_decodeResult_vwmacc;
  assign validSink_bits_decodeResult_vwmacc = shifterReg_0_bits_decodeResult_vwmacc;
  reg          shifterReg_0_bits_decodeResult_readOnly;
  assign validSink_bits_decodeResult_readOnly = shifterReg_0_bits_decodeResult_readOnly;
  reg          shifterReg_0_bits_decodeResult_maskSource;
  assign validSink_bits_decodeResult_maskSource = shifterReg_0_bits_decodeResult_maskSource;
  reg          shifterReg_0_bits_decodeResult_maskDestination;
  assign validSink_bits_decodeResult_maskDestination = shifterReg_0_bits_decodeResult_maskDestination;
  reg          shifterReg_0_bits_decodeResult_maskLogic;
  assign validSink_bits_decodeResult_maskLogic = shifterReg_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_0_bits_decodeResult_uop;
  assign validSink_bits_decodeResult_uop = shifterReg_0_bits_decodeResult_uop;
  reg          shifterReg_0_bits_decodeResult_iota;
  assign validSink_bits_decodeResult_iota = shifterReg_0_bits_decodeResult_iota;
  reg          shifterReg_0_bits_decodeResult_mv;
  assign validSink_bits_decodeResult_mv = shifterReg_0_bits_decodeResult_mv;
  reg          shifterReg_0_bits_decodeResult_extend;
  assign validSink_bits_decodeResult_extend = shifterReg_0_bits_decodeResult_extend;
  reg          shifterReg_0_bits_decodeResult_unOrderWrite;
  assign validSink_bits_decodeResult_unOrderWrite = shifterReg_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_0_bits_decodeResult_compress;
  assign validSink_bits_decodeResult_compress = shifterReg_0_bits_decodeResult_compress;
  reg          shifterReg_0_bits_decodeResult_gather16;
  assign validSink_bits_decodeResult_gather16 = shifterReg_0_bits_decodeResult_gather16;
  reg          shifterReg_0_bits_decodeResult_gather;
  assign validSink_bits_decodeResult_gather = shifterReg_0_bits_decodeResult_gather;
  reg          shifterReg_0_bits_decodeResult_slid;
  assign validSink_bits_decodeResult_slid = shifterReg_0_bits_decodeResult_slid;
  reg          shifterReg_0_bits_decodeResult_targetRd;
  assign validSink_bits_decodeResult_targetRd = shifterReg_0_bits_decodeResult_targetRd;
  reg          shifterReg_0_bits_decodeResult_widenReduce;
  assign validSink_bits_decodeResult_widenReduce = shifterReg_0_bits_decodeResult_widenReduce;
  reg          shifterReg_0_bits_decodeResult_red;
  assign validSink_bits_decodeResult_red = shifterReg_0_bits_decodeResult_red;
  reg          shifterReg_0_bits_decodeResult_nr;
  assign validSink_bits_decodeResult_nr = shifterReg_0_bits_decodeResult_nr;
  reg          shifterReg_0_bits_decodeResult_itype;
  assign validSink_bits_decodeResult_itype = shifterReg_0_bits_decodeResult_itype;
  reg          shifterReg_0_bits_decodeResult_unsigned1;
  assign validSink_bits_decodeResult_unsigned1 = shifterReg_0_bits_decodeResult_unsigned1;
  reg          shifterReg_0_bits_decodeResult_unsigned0;
  assign validSink_bits_decodeResult_unsigned0 = shifterReg_0_bits_decodeResult_unsigned0;
  reg          shifterReg_0_bits_decodeResult_other;
  assign validSink_bits_decodeResult_other = shifterReg_0_bits_decodeResult_other;
  reg          shifterReg_0_bits_decodeResult_multiCycle;
  assign validSink_bits_decodeResult_multiCycle = shifterReg_0_bits_decodeResult_multiCycle;
  reg          shifterReg_0_bits_decodeResult_divider;
  assign validSink_bits_decodeResult_divider = shifterReg_0_bits_decodeResult_divider;
  reg          shifterReg_0_bits_decodeResult_multiplier;
  assign validSink_bits_decodeResult_multiplier = shifterReg_0_bits_decodeResult_multiplier;
  reg          shifterReg_0_bits_decodeResult_shift;
  assign validSink_bits_decodeResult_shift = shifterReg_0_bits_decodeResult_shift;
  reg          shifterReg_0_bits_decodeResult_adder;
  assign validSink_bits_decodeResult_adder = shifterReg_0_bits_decodeResult_adder;
  reg          shifterReg_0_bits_decodeResult_logic;
  assign validSink_bits_decodeResult_logic = shifterReg_0_bits_decodeResult_logic;
  reg          shifterReg_0_bits_loadStore;
  assign validSink_bits_loadStore = shifterReg_0_bits_loadStore;
  reg          shifterReg_0_bits_issueInst;
  assign validSink_bits_issueInst = shifterReg_0_bits_issueInst;
  reg          shifterReg_0_bits_store;
  assign validSink_bits_store = shifterReg_0_bits_store;
  reg          shifterReg_0_bits_special;
  assign validSink_bits_special = shifterReg_0_bits_special;
  reg          shifterReg_0_bits_lsWholeReg;
  assign validSink_bits_lsWholeReg = shifterReg_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_0_bits_vs1;
  assign validSink_bits_vs1 = shifterReg_0_bits_vs1;
  reg  [4:0]   shifterReg_0_bits_vs2;
  assign validSink_bits_vs2 = shifterReg_0_bits_vs2;
  reg  [4:0]   shifterReg_0_bits_vd;
  assign validSink_bits_vd = shifterReg_0_bits_vd;
  reg  [1:0]   shifterReg_0_bits_loadStoreEEW;
  assign validSink_bits_loadStoreEEW = shifterReg_0_bits_loadStoreEEW;
  reg          shifterReg_0_bits_mask;
  assign validSink_bits_mask = shifterReg_0_bits_mask;
  reg  [2:0]   shifterReg_0_bits_segment;
  assign validSink_bits_segment = shifterReg_0_bits_segment;
  reg  [31:0]  shifterReg_0_bits_readFromScalar;
  assign validSink_bits_readFromScalar = shifterReg_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_0_bits_csrInterface_vl;
  assign validSink_bits_csrInterface_vl = shifterReg_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_0_bits_csrInterface_vStart;
  assign validSink_bits_csrInterface_vStart = shifterReg_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_0_bits_csrInterface_vlmul;
  assign validSink_bits_csrInterface_vlmul = shifterReg_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_0_bits_csrInterface_vSew;
  assign validSink_bits_csrInterface_vSew = shifterReg_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_0_bits_csrInterface_vxrm;
  assign validSink_bits_csrInterface_vxrm = shifterReg_0_bits_csrInterface_vxrm;
  reg          shifterReg_0_bits_csrInterface_vta;
  assign validSink_bits_csrInterface_vta = shifterReg_0_bits_csrInterface_vta;
  reg          shifterReg_0_bits_csrInterface_vma;
  assign validSink_bits_csrInterface_vma = shifterReg_0_bits_csrInterface_vma;
  wire         shifterValid = shifterReg_0_valid | validSource_valid;
  wire         validSink_1_valid;
  wire [2:0]   validSink_1_bits_instructionIndex;
  wire         validSink_1_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_1_bits_decodeResult_topUop;
  wire         validSink_1_bits_decodeResult_popCount;
  wire         validSink_1_bits_decodeResult_ffo;
  wire         validSink_1_bits_decodeResult_average;
  wire         validSink_1_bits_decodeResult_reverse;
  wire         validSink_1_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_1_bits_decodeResult_scheduler;
  wire         validSink_1_bits_decodeResult_sReadVD;
  wire         validSink_1_bits_decodeResult_vtype;
  wire         validSink_1_bits_decodeResult_sWrite;
  wire         validSink_1_bits_decodeResult_crossRead;
  wire         validSink_1_bits_decodeResult_crossWrite;
  wire         validSink_1_bits_decodeResult_maskUnit;
  wire         validSink_1_bits_decodeResult_special;
  wire         validSink_1_bits_decodeResult_saturate;
  wire         validSink_1_bits_decodeResult_vwmacc;
  wire         validSink_1_bits_decodeResult_readOnly;
  wire         validSink_1_bits_decodeResult_maskSource;
  wire         validSink_1_bits_decodeResult_maskDestination;
  wire         validSink_1_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_1_bits_decodeResult_uop;
  wire         validSink_1_bits_decodeResult_iota;
  wire         validSink_1_bits_decodeResult_mv;
  wire         validSink_1_bits_decodeResult_extend;
  wire         validSink_1_bits_decodeResult_unOrderWrite;
  wire         validSink_1_bits_decodeResult_compress;
  wire         validSink_1_bits_decodeResult_gather16;
  wire         validSink_1_bits_decodeResult_gather;
  wire         validSink_1_bits_decodeResult_slid;
  wire         validSink_1_bits_decodeResult_targetRd;
  wire         validSink_1_bits_decodeResult_widenReduce;
  wire         validSink_1_bits_decodeResult_red;
  wire         validSink_1_bits_decodeResult_nr;
  wire         validSink_1_bits_decodeResult_itype;
  wire         validSink_1_bits_decodeResult_unsigned1;
  wire         validSink_1_bits_decodeResult_unsigned0;
  wire         validSink_1_bits_decodeResult_other;
  wire         validSink_1_bits_decodeResult_multiCycle;
  wire         validSink_1_bits_decodeResult_divider;
  wire         validSink_1_bits_decodeResult_multiplier;
  wire         validSink_1_bits_decodeResult_shift;
  wire         validSink_1_bits_decodeResult_adder;
  wire         validSink_1_bits_decodeResult_logic;
  wire         validSink_1_bits_loadStore;
  wire         validSink_1_bits_issueInst;
  wire         validSink_1_bits_store;
  wire         validSink_1_bits_special;
  wire         validSink_1_bits_lsWholeReg;
  wire [4:0]   validSink_1_bits_vs1;
  wire [4:0]   validSink_1_bits_vs2;
  wire [4:0]   validSink_1_bits_vd;
  wire [1:0]   validSink_1_bits_loadStoreEEW;
  wire         validSink_1_bits_mask;
  wire [2:0]   validSink_1_bits_segment;
  wire [31:0]  validSink_1_bits_readFromScalar;
  wire [11:0]  validSink_1_bits_csrInterface_vl;
  wire [11:0]  validSink_1_bits_csrInterface_vStart;
  wire [2:0]   validSink_1_bits_csrInterface_vlmul;
  wire [1:0]   validSink_1_bits_csrInterface_vSew;
  wire [1:0]   validSink_1_bits_csrInterface_vxrm;
  wire         validSink_1_bits_csrInterface_vta;
  wire         validSink_1_bits_csrInterface_vma;
  wire         laneRequestSinkWire_1_valid = queue_1_deq_valid;
  wire [2:0]   laneRequestSinkWire_1_bits_instructionIndex = queue_1_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_1_bits_decodeResult_specialSlot = queue_1_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_1_bits_decodeResult_topUop = queue_1_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_1_bits_decodeResult_popCount = queue_1_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_1_bits_decodeResult_ffo = queue_1_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_1_bits_decodeResult_average = queue_1_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_1_bits_decodeResult_reverse = queue_1_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_1_bits_decodeResult_dontNeedExecuteInLane = queue_1_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_1_bits_decodeResult_scheduler = queue_1_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_1_bits_decodeResult_sReadVD = queue_1_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_1_bits_decodeResult_vtype = queue_1_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_1_bits_decodeResult_sWrite = queue_1_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_1_bits_decodeResult_crossRead = queue_1_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_1_bits_decodeResult_crossWrite = queue_1_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_1_bits_decodeResult_maskUnit = queue_1_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_1_bits_decodeResult_special = queue_1_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_1_bits_decodeResult_saturate = queue_1_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_1_bits_decodeResult_vwmacc = queue_1_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_1_bits_decodeResult_readOnly = queue_1_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_1_bits_decodeResult_maskSource = queue_1_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_1_bits_decodeResult_maskDestination = queue_1_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_1_bits_decodeResult_maskLogic = queue_1_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_1_bits_decodeResult_uop = queue_1_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_1_bits_decodeResult_iota = queue_1_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_1_bits_decodeResult_mv = queue_1_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_1_bits_decodeResult_extend = queue_1_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_1_bits_decodeResult_unOrderWrite = queue_1_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_1_bits_decodeResult_compress = queue_1_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_1_bits_decodeResult_gather16 = queue_1_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_1_bits_decodeResult_gather = queue_1_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_1_bits_decodeResult_slid = queue_1_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_1_bits_decodeResult_targetRd = queue_1_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_1_bits_decodeResult_widenReduce = queue_1_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_1_bits_decodeResult_red = queue_1_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_1_bits_decodeResult_nr = queue_1_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_1_bits_decodeResult_itype = queue_1_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_1_bits_decodeResult_unsigned1 = queue_1_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_1_bits_decodeResult_unsigned0 = queue_1_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_1_bits_decodeResult_other = queue_1_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_1_bits_decodeResult_multiCycle = queue_1_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_1_bits_decodeResult_divider = queue_1_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_1_bits_decodeResult_multiplier = queue_1_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_1_bits_decodeResult_shift = queue_1_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_1_bits_decodeResult_adder = queue_1_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_1_bits_decodeResult_logic = queue_1_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_1_bits_loadStore = queue_1_deq_bits_loadStore;
  wire         laneRequestSinkWire_1_bits_issueInst = queue_1_deq_bits_issueInst;
  wire         laneRequestSinkWire_1_bits_store = queue_1_deq_bits_store;
  wire         laneRequestSinkWire_1_bits_special = queue_1_deq_bits_special;
  wire         laneRequestSinkWire_1_bits_lsWholeReg = queue_1_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_1_bits_vs1 = queue_1_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_1_bits_vs2 = queue_1_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_1_bits_vd = queue_1_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_1_bits_loadStoreEEW = queue_1_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_1_bits_mask = queue_1_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_1_bits_segment = queue_1_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_1_bits_readFromScalar = queue_1_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_1_bits_csrInterface_vl = queue_1_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_1_bits_csrInterface_vStart = queue_1_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_1_bits_csrInterface_vlmul = queue_1_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_1_bits_csrInterface_vSew = queue_1_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_1_bits_csrInterface_vxrm = queue_1_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_1_bits_csrInterface_vta = queue_1_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_1_bits_csrInterface_vma = queue_1_deq_bits_csrInterface_vma;
  wire [1:0]   queue_1_enq_bits_csrInterface_vxrm;
  wire         queue_1_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi_3 = {queue_1_enq_bits_csrInterface_vxrm, queue_1_enq_bits_csrInterface_vta};
  wire         queue_1_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo_3 = {queue_dataIn_lo_hi_3, queue_1_enq_bits_csrInterface_vma};
  wire [2:0]   queue_1_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_1_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo_3 = {queue_1_enq_bits_csrInterface_vlmul, queue_1_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_1_enq_bits_csrInterface_vl;
  wire [11:0]  queue_1_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi_3 = {queue_1_enq_bits_csrInterface_vl, queue_1_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi_3 = {queue_dataIn_hi_hi_3, queue_dataIn_hi_lo_3};
  wire         queue_1_enq_bits_decodeResult_adder;
  wire         queue_1_enq_bits_decodeResult_logic;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo_1 = {queue_1_enq_bits_decodeResult_adder, queue_1_enq_bits_decodeResult_logic};
  wire         queue_1_enq_bits_decodeResult_divider;
  wire         queue_1_enq_bits_decodeResult_multiplier;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi_1 = {queue_1_enq_bits_decodeResult_divider, queue_1_enq_bits_decodeResult_multiplier};
  wire         queue_1_enq_bits_decodeResult_shift;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi_1 = {queue_dataIn_lo_lo_lo_hi_hi_1, queue_1_enq_bits_decodeResult_shift};
  wire [4:0]   queue_dataIn_lo_lo_lo_1 = {queue_dataIn_lo_lo_lo_hi_1, queue_dataIn_lo_lo_lo_lo_1};
  wire         queue_1_enq_bits_decodeResult_unsigned0;
  wire         queue_1_enq_bits_decodeResult_other;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi_1 = {queue_1_enq_bits_decodeResult_unsigned0, queue_1_enq_bits_decodeResult_other};
  wire         queue_1_enq_bits_decodeResult_multiCycle;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo_1 = {queue_dataIn_lo_lo_hi_lo_hi_1, queue_1_enq_bits_decodeResult_multiCycle};
  wire         queue_1_enq_bits_decodeResult_nr;
  wire         queue_1_enq_bits_decodeResult_itype;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi_1 = {queue_1_enq_bits_decodeResult_nr, queue_1_enq_bits_decodeResult_itype};
  wire         queue_1_enq_bits_decodeResult_unsigned1;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi_1 = {queue_dataIn_lo_lo_hi_hi_hi_1, queue_1_enq_bits_decodeResult_unsigned1};
  wire [5:0]   queue_dataIn_lo_lo_hi_2 = {queue_dataIn_lo_lo_hi_hi_1, queue_dataIn_lo_lo_hi_lo_1};
  wire [10:0]  queue_dataIn_lo_lo_2 = {queue_dataIn_lo_lo_hi_2, queue_dataIn_lo_lo_lo_1};
  wire         queue_1_enq_bits_decodeResult_widenReduce;
  wire         queue_1_enq_bits_decodeResult_red;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo_1 = {queue_1_enq_bits_decodeResult_widenReduce, queue_1_enq_bits_decodeResult_red};
  wire         queue_1_enq_bits_decodeResult_gather;
  wire         queue_1_enq_bits_decodeResult_slid;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi_1 = {queue_1_enq_bits_decodeResult_gather, queue_1_enq_bits_decodeResult_slid};
  wire         queue_1_enq_bits_decodeResult_targetRd;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi_1 = {queue_dataIn_lo_hi_lo_hi_hi_1, queue_1_enq_bits_decodeResult_targetRd};
  wire [4:0]   queue_dataIn_lo_hi_lo_2 = {queue_dataIn_lo_hi_lo_hi_1, queue_dataIn_lo_hi_lo_lo_1};
  wire         queue_1_enq_bits_decodeResult_unOrderWrite;
  wire         queue_1_enq_bits_decodeResult_compress;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi_1 = {queue_1_enq_bits_decodeResult_unOrderWrite, queue_1_enq_bits_decodeResult_compress};
  wire         queue_1_enq_bits_decodeResult_gather16;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo_1 = {queue_dataIn_lo_hi_hi_lo_hi_1, queue_1_enq_bits_decodeResult_gather16};
  wire         queue_1_enq_bits_decodeResult_iota;
  wire         queue_1_enq_bits_decodeResult_mv;
  wire [1:0]   queue_dataIn_lo_hi_hi_hi_hi_1 = {queue_1_enq_bits_decodeResult_iota, queue_1_enq_bits_decodeResult_mv};
  wire         queue_1_enq_bits_decodeResult_extend;
  wire [2:0]   queue_dataIn_lo_hi_hi_hi_1 = {queue_dataIn_lo_hi_hi_hi_hi_1, queue_1_enq_bits_decodeResult_extend};
  wire [5:0]   queue_dataIn_lo_hi_hi_2 = {queue_dataIn_lo_hi_hi_hi_1, queue_dataIn_lo_hi_hi_lo_1};
  wire [10:0]  queue_dataIn_lo_hi_4 = {queue_dataIn_lo_hi_hi_2, queue_dataIn_lo_hi_lo_2};
  wire [21:0]  queue_dataIn_lo_4 = {queue_dataIn_lo_hi_4, queue_dataIn_lo_lo_2};
  wire         queue_1_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_1_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_hi_lo_lo_lo_1 = {queue_1_enq_bits_decodeResult_maskLogic, queue_1_enq_bits_decodeResult_uop};
  wire         queue_1_enq_bits_decodeResult_readOnly;
  wire         queue_1_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi_1 = {queue_1_enq_bits_decodeResult_readOnly, queue_1_enq_bits_decodeResult_maskSource};
  wire         queue_1_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi_1 = {queue_dataIn_hi_lo_lo_hi_hi_1, queue_1_enq_bits_decodeResult_maskDestination};
  wire [7:0]   queue_dataIn_hi_lo_lo_2 = {queue_dataIn_hi_lo_lo_hi_1, queue_dataIn_hi_lo_lo_lo_1};
  wire         queue_1_enq_bits_decodeResult_special;
  wire         queue_1_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi_1 = {queue_1_enq_bits_decodeResult_special, queue_1_enq_bits_decodeResult_saturate};
  wire         queue_1_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo_1 = {queue_dataIn_hi_lo_hi_lo_hi_1, queue_1_enq_bits_decodeResult_vwmacc};
  wire         queue_1_enq_bits_decodeResult_crossRead;
  wire         queue_1_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi_1 = {queue_1_enq_bits_decodeResult_crossRead, queue_1_enq_bits_decodeResult_crossWrite};
  wire         queue_1_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi_1 = {queue_dataIn_hi_lo_hi_hi_hi_1, queue_1_enq_bits_decodeResult_maskUnit};
  wire [5:0]   queue_dataIn_hi_lo_hi_2 = {queue_dataIn_hi_lo_hi_hi_1, queue_dataIn_hi_lo_hi_lo_1};
  wire [13:0]  queue_dataIn_hi_lo_4 = {queue_dataIn_hi_lo_hi_2, queue_dataIn_hi_lo_lo_2};
  wire         queue_1_enq_bits_decodeResult_vtype;
  wire         queue_1_enq_bits_decodeResult_sWrite;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo_1 = {queue_1_enq_bits_decodeResult_vtype, queue_1_enq_bits_decodeResult_sWrite};
  wire         queue_1_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_1_enq_bits_decodeResult_scheduler;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi_1 = {queue_1_enq_bits_decodeResult_dontNeedExecuteInLane, queue_1_enq_bits_decodeResult_scheduler};
  wire         queue_1_enq_bits_decodeResult_sReadVD;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi_1 = {queue_dataIn_hi_hi_lo_hi_hi_1, queue_1_enq_bits_decodeResult_sReadVD};
  wire [4:0]   queue_dataIn_hi_hi_lo_2 = {queue_dataIn_hi_hi_lo_hi_1, queue_dataIn_hi_hi_lo_lo_1};
  wire         queue_1_enq_bits_decodeResult_ffo;
  wire         queue_1_enq_bits_decodeResult_average;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi_1 = {queue_1_enq_bits_decodeResult_ffo, queue_1_enq_bits_decodeResult_average};
  wire         queue_1_enq_bits_decodeResult_reverse;
  wire [2:0]   queue_dataIn_hi_hi_hi_lo_1 = {queue_dataIn_hi_hi_hi_lo_hi_1, queue_1_enq_bits_decodeResult_reverse};
  wire         queue_1_enq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_1_enq_bits_decodeResult_topUop;
  wire [5:0]   queue_dataIn_hi_hi_hi_hi_hi_1 = {queue_1_enq_bits_decodeResult_specialSlot, queue_1_enq_bits_decodeResult_topUop};
  wire         queue_1_enq_bits_decodeResult_popCount;
  wire [6:0]   queue_dataIn_hi_hi_hi_hi_1 = {queue_dataIn_hi_hi_hi_hi_hi_1, queue_1_enq_bits_decodeResult_popCount};
  wire [9:0]   queue_dataIn_hi_hi_hi_2 = {queue_dataIn_hi_hi_hi_hi_1, queue_dataIn_hi_hi_hi_lo_1};
  wire [14:0]  queue_dataIn_hi_hi_4 = {queue_dataIn_hi_hi_hi_2, queue_dataIn_hi_hi_lo_2};
  wire [28:0]  queue_dataIn_hi_4 = {queue_dataIn_hi_hi_4, queue_dataIn_hi_lo_4};
  wire [2:0]   queue_1_enq_bits_segment;
  wire [31:0]  queue_1_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_3 = {queue_1_enq_bits_segment, queue_1_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_3 = {queue_dataIn_lo_lo_hi_3, queue_dataIn_hi_3, queue_dataIn_lo_3};
  wire [1:0]   queue_1_enq_bits_loadStoreEEW;
  wire         queue_1_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_3 = {queue_1_enq_bits_loadStoreEEW, queue_1_enq_bits_mask};
  wire [4:0]   queue_1_enq_bits_vs2;
  wire [4:0]   queue_1_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_3 = {queue_1_enq_bits_vs2, queue_1_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_5 = {queue_dataIn_lo_hi_hi_3, queue_dataIn_lo_hi_lo_3};
  wire [80:0]  queue_dataIn_lo_5 = {queue_dataIn_lo_hi_5, queue_dataIn_lo_lo_3};
  wire         queue_1_enq_bits_lsWholeReg;
  wire [4:0]   queue_1_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_3 = {queue_1_enq_bits_lsWholeReg, queue_1_enq_bits_vs1};
  wire         queue_1_enq_bits_store;
  wire         queue_1_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_3 = {queue_1_enq_bits_store, queue_1_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_5 = {queue_dataIn_hi_lo_hi_3, queue_dataIn_hi_lo_lo_3};
  wire         queue_1_enq_bits_loadStore;
  wire         queue_1_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_3 = {queue_1_enq_bits_loadStore, queue_1_enq_bits_issueInst};
  wire [2:0]   queue_1_enq_bits_instructionIndex;
  wire [53:0]  queue_dataIn_hi_hi_hi_3 = {queue_1_enq_bits_instructionIndex, queue_dataIn_hi_4, queue_dataIn_lo_4};
  wire [55:0]  queue_dataIn_hi_hi_5 = {queue_dataIn_hi_hi_hi_3, queue_dataIn_hi_hi_lo_3};
  wire [63:0]  queue_dataIn_hi_5 = {queue_dataIn_hi_hi_5, queue_dataIn_hi_lo_5};
  wire [144:0] queue_dataIn_1 = {queue_dataIn_hi_5, queue_dataIn_lo_5};
  wire         queue_dataOut_1_csrInterface_vma = _queue_fifo_1_data_out[0];
  wire         queue_dataOut_1_csrInterface_vta = _queue_fifo_1_data_out[1];
  wire [1:0]   queue_dataOut_1_csrInterface_vxrm = _queue_fifo_1_data_out[3:2];
  wire [1:0]   queue_dataOut_1_csrInterface_vSew = _queue_fifo_1_data_out[5:4];
  wire [2:0]   queue_dataOut_1_csrInterface_vlmul = _queue_fifo_1_data_out[8:6];
  wire [11:0]  queue_dataOut_1_csrInterface_vStart = _queue_fifo_1_data_out[20:9];
  wire [11:0]  queue_dataOut_1_csrInterface_vl = _queue_fifo_1_data_out[32:21];
  wire [31:0]  queue_dataOut_1_readFromScalar = _queue_fifo_1_data_out[64:33];
  wire [2:0]   queue_dataOut_1_segment = _queue_fifo_1_data_out[67:65];
  wire         queue_dataOut_1_mask = _queue_fifo_1_data_out[68];
  wire [1:0]   queue_dataOut_1_loadStoreEEW = _queue_fifo_1_data_out[70:69];
  wire [4:0]   queue_dataOut_1_vd = _queue_fifo_1_data_out[75:71];
  wire [4:0]   queue_dataOut_1_vs2 = _queue_fifo_1_data_out[80:76];
  wire [4:0]   queue_dataOut_1_vs1 = _queue_fifo_1_data_out[85:81];
  wire         queue_dataOut_1_lsWholeReg = _queue_fifo_1_data_out[86];
  wire         queue_dataOut_1_special = _queue_fifo_1_data_out[87];
  wire         queue_dataOut_1_store = _queue_fifo_1_data_out[88];
  wire         queue_dataOut_1_issueInst = _queue_fifo_1_data_out[89];
  wire         queue_dataOut_1_loadStore = _queue_fifo_1_data_out[90];
  wire         queue_dataOut_1_decodeResult_logic = _queue_fifo_1_data_out[91];
  wire         queue_dataOut_1_decodeResult_adder = _queue_fifo_1_data_out[92];
  wire         queue_dataOut_1_decodeResult_shift = _queue_fifo_1_data_out[93];
  wire         queue_dataOut_1_decodeResult_multiplier = _queue_fifo_1_data_out[94];
  wire         queue_dataOut_1_decodeResult_divider = _queue_fifo_1_data_out[95];
  wire         queue_dataOut_1_decodeResult_multiCycle = _queue_fifo_1_data_out[96];
  wire         queue_dataOut_1_decodeResult_other = _queue_fifo_1_data_out[97];
  wire         queue_dataOut_1_decodeResult_unsigned0 = _queue_fifo_1_data_out[98];
  wire         queue_dataOut_1_decodeResult_unsigned1 = _queue_fifo_1_data_out[99];
  wire         queue_dataOut_1_decodeResult_itype = _queue_fifo_1_data_out[100];
  wire         queue_dataOut_1_decodeResult_nr = _queue_fifo_1_data_out[101];
  wire         queue_dataOut_1_decodeResult_red = _queue_fifo_1_data_out[102];
  wire         queue_dataOut_1_decodeResult_widenReduce = _queue_fifo_1_data_out[103];
  wire         queue_dataOut_1_decodeResult_targetRd = _queue_fifo_1_data_out[104];
  wire         queue_dataOut_1_decodeResult_slid = _queue_fifo_1_data_out[105];
  wire         queue_dataOut_1_decodeResult_gather = _queue_fifo_1_data_out[106];
  wire         queue_dataOut_1_decodeResult_gather16 = _queue_fifo_1_data_out[107];
  wire         queue_dataOut_1_decodeResult_compress = _queue_fifo_1_data_out[108];
  wire         queue_dataOut_1_decodeResult_unOrderWrite = _queue_fifo_1_data_out[109];
  wire         queue_dataOut_1_decodeResult_extend = _queue_fifo_1_data_out[110];
  wire         queue_dataOut_1_decodeResult_mv = _queue_fifo_1_data_out[111];
  wire         queue_dataOut_1_decodeResult_iota = _queue_fifo_1_data_out[112];
  wire [3:0]   queue_dataOut_1_decodeResult_uop = _queue_fifo_1_data_out[116:113];
  wire         queue_dataOut_1_decodeResult_maskLogic = _queue_fifo_1_data_out[117];
  wire         queue_dataOut_1_decodeResult_maskDestination = _queue_fifo_1_data_out[118];
  wire         queue_dataOut_1_decodeResult_maskSource = _queue_fifo_1_data_out[119];
  wire         queue_dataOut_1_decodeResult_readOnly = _queue_fifo_1_data_out[120];
  wire         queue_dataOut_1_decodeResult_vwmacc = _queue_fifo_1_data_out[121];
  wire         queue_dataOut_1_decodeResult_saturate = _queue_fifo_1_data_out[122];
  wire         queue_dataOut_1_decodeResult_special = _queue_fifo_1_data_out[123];
  wire         queue_dataOut_1_decodeResult_maskUnit = _queue_fifo_1_data_out[124];
  wire         queue_dataOut_1_decodeResult_crossWrite = _queue_fifo_1_data_out[125];
  wire         queue_dataOut_1_decodeResult_crossRead = _queue_fifo_1_data_out[126];
  wire         queue_dataOut_1_decodeResult_sWrite = _queue_fifo_1_data_out[127];
  wire         queue_dataOut_1_decodeResult_vtype = _queue_fifo_1_data_out[128];
  wire         queue_dataOut_1_decodeResult_sReadVD = _queue_fifo_1_data_out[129];
  wire         queue_dataOut_1_decodeResult_scheduler = _queue_fifo_1_data_out[130];
  wire         queue_dataOut_1_decodeResult_dontNeedExecuteInLane = _queue_fifo_1_data_out[131];
  wire         queue_dataOut_1_decodeResult_reverse = _queue_fifo_1_data_out[132];
  wire         queue_dataOut_1_decodeResult_average = _queue_fifo_1_data_out[133];
  wire         queue_dataOut_1_decodeResult_ffo = _queue_fifo_1_data_out[134];
  wire         queue_dataOut_1_decodeResult_popCount = _queue_fifo_1_data_out[135];
  wire [4:0]   queue_dataOut_1_decodeResult_topUop = _queue_fifo_1_data_out[140:136];
  wire         queue_dataOut_1_decodeResult_specialSlot = _queue_fifo_1_data_out[141];
  wire [2:0]   queue_dataOut_1_instructionIndex = _queue_fifo_1_data_out[144:142];
  wire         queue_1_enq_ready = ~_queue_fifo_1_full;
  wire         queue_1_enq_valid;
  assign queue_1_deq_valid = ~_queue_fifo_1_empty | queue_1_enq_valid;
  assign queue_1_deq_bits_instructionIndex = _queue_fifo_1_empty ? queue_1_enq_bits_instructionIndex : queue_dataOut_1_instructionIndex;
  assign queue_1_deq_bits_decodeResult_specialSlot = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_specialSlot : queue_dataOut_1_decodeResult_specialSlot;
  assign queue_1_deq_bits_decodeResult_topUop = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_topUop : queue_dataOut_1_decodeResult_topUop;
  assign queue_1_deq_bits_decodeResult_popCount = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_popCount : queue_dataOut_1_decodeResult_popCount;
  assign queue_1_deq_bits_decodeResult_ffo = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_ffo : queue_dataOut_1_decodeResult_ffo;
  assign queue_1_deq_bits_decodeResult_average = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_average : queue_dataOut_1_decodeResult_average;
  assign queue_1_deq_bits_decodeResult_reverse = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_reverse : queue_dataOut_1_decodeResult_reverse;
  assign queue_1_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_1_decodeResult_dontNeedExecuteInLane;
  assign queue_1_deq_bits_decodeResult_scheduler = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_scheduler : queue_dataOut_1_decodeResult_scheduler;
  assign queue_1_deq_bits_decodeResult_sReadVD = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_sReadVD : queue_dataOut_1_decodeResult_sReadVD;
  assign queue_1_deq_bits_decodeResult_vtype = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_vtype : queue_dataOut_1_decodeResult_vtype;
  assign queue_1_deq_bits_decodeResult_sWrite = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_sWrite : queue_dataOut_1_decodeResult_sWrite;
  assign queue_1_deq_bits_decodeResult_crossRead = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_crossRead : queue_dataOut_1_decodeResult_crossRead;
  assign queue_1_deq_bits_decodeResult_crossWrite = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_crossWrite : queue_dataOut_1_decodeResult_crossWrite;
  assign queue_1_deq_bits_decodeResult_maskUnit = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_maskUnit : queue_dataOut_1_decodeResult_maskUnit;
  assign queue_1_deq_bits_decodeResult_special = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_special : queue_dataOut_1_decodeResult_special;
  assign queue_1_deq_bits_decodeResult_saturate = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_saturate : queue_dataOut_1_decodeResult_saturate;
  assign queue_1_deq_bits_decodeResult_vwmacc = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_vwmacc : queue_dataOut_1_decodeResult_vwmacc;
  assign queue_1_deq_bits_decodeResult_readOnly = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_readOnly : queue_dataOut_1_decodeResult_readOnly;
  assign queue_1_deq_bits_decodeResult_maskSource = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_maskSource : queue_dataOut_1_decodeResult_maskSource;
  assign queue_1_deq_bits_decodeResult_maskDestination = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_maskDestination : queue_dataOut_1_decodeResult_maskDestination;
  assign queue_1_deq_bits_decodeResult_maskLogic = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_maskLogic : queue_dataOut_1_decodeResult_maskLogic;
  assign queue_1_deq_bits_decodeResult_uop = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_uop : queue_dataOut_1_decodeResult_uop;
  assign queue_1_deq_bits_decodeResult_iota = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_iota : queue_dataOut_1_decodeResult_iota;
  assign queue_1_deq_bits_decodeResult_mv = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_mv : queue_dataOut_1_decodeResult_mv;
  assign queue_1_deq_bits_decodeResult_extend = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_extend : queue_dataOut_1_decodeResult_extend;
  assign queue_1_deq_bits_decodeResult_unOrderWrite = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_unOrderWrite : queue_dataOut_1_decodeResult_unOrderWrite;
  assign queue_1_deq_bits_decodeResult_compress = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_compress : queue_dataOut_1_decodeResult_compress;
  assign queue_1_deq_bits_decodeResult_gather16 = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_gather16 : queue_dataOut_1_decodeResult_gather16;
  assign queue_1_deq_bits_decodeResult_gather = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_gather : queue_dataOut_1_decodeResult_gather;
  assign queue_1_deq_bits_decodeResult_slid = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_slid : queue_dataOut_1_decodeResult_slid;
  assign queue_1_deq_bits_decodeResult_targetRd = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_targetRd : queue_dataOut_1_decodeResult_targetRd;
  assign queue_1_deq_bits_decodeResult_widenReduce = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_widenReduce : queue_dataOut_1_decodeResult_widenReduce;
  assign queue_1_deq_bits_decodeResult_red = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_red : queue_dataOut_1_decodeResult_red;
  assign queue_1_deq_bits_decodeResult_nr = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_nr : queue_dataOut_1_decodeResult_nr;
  assign queue_1_deq_bits_decodeResult_itype = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_itype : queue_dataOut_1_decodeResult_itype;
  assign queue_1_deq_bits_decodeResult_unsigned1 = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_unsigned1 : queue_dataOut_1_decodeResult_unsigned1;
  assign queue_1_deq_bits_decodeResult_unsigned0 = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_unsigned0 : queue_dataOut_1_decodeResult_unsigned0;
  assign queue_1_deq_bits_decodeResult_other = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_other : queue_dataOut_1_decodeResult_other;
  assign queue_1_deq_bits_decodeResult_multiCycle = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_multiCycle : queue_dataOut_1_decodeResult_multiCycle;
  assign queue_1_deq_bits_decodeResult_divider = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_divider : queue_dataOut_1_decodeResult_divider;
  assign queue_1_deq_bits_decodeResult_multiplier = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_multiplier : queue_dataOut_1_decodeResult_multiplier;
  assign queue_1_deq_bits_decodeResult_shift = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_shift : queue_dataOut_1_decodeResult_shift;
  assign queue_1_deq_bits_decodeResult_adder = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_adder : queue_dataOut_1_decodeResult_adder;
  assign queue_1_deq_bits_decodeResult_logic = _queue_fifo_1_empty ? queue_1_enq_bits_decodeResult_logic : queue_dataOut_1_decodeResult_logic;
  assign queue_1_deq_bits_loadStore = _queue_fifo_1_empty ? queue_1_enq_bits_loadStore : queue_dataOut_1_loadStore;
  assign queue_1_deq_bits_issueInst = _queue_fifo_1_empty ? queue_1_enq_bits_issueInst : queue_dataOut_1_issueInst;
  assign queue_1_deq_bits_store = _queue_fifo_1_empty ? queue_1_enq_bits_store : queue_dataOut_1_store;
  assign queue_1_deq_bits_special = _queue_fifo_1_empty ? queue_1_enq_bits_special : queue_dataOut_1_special;
  assign queue_1_deq_bits_lsWholeReg = _queue_fifo_1_empty ? queue_1_enq_bits_lsWholeReg : queue_dataOut_1_lsWholeReg;
  assign queue_1_deq_bits_vs1 = _queue_fifo_1_empty ? queue_1_enq_bits_vs1 : queue_dataOut_1_vs1;
  assign queue_1_deq_bits_vs2 = _queue_fifo_1_empty ? queue_1_enq_bits_vs2 : queue_dataOut_1_vs2;
  assign queue_1_deq_bits_vd = _queue_fifo_1_empty ? queue_1_enq_bits_vd : queue_dataOut_1_vd;
  assign queue_1_deq_bits_loadStoreEEW = _queue_fifo_1_empty ? queue_1_enq_bits_loadStoreEEW : queue_dataOut_1_loadStoreEEW;
  assign queue_1_deq_bits_mask = _queue_fifo_1_empty ? queue_1_enq_bits_mask : queue_dataOut_1_mask;
  assign queue_1_deq_bits_segment = _queue_fifo_1_empty ? queue_1_enq_bits_segment : queue_dataOut_1_segment;
  assign queue_1_deq_bits_readFromScalar = _queue_fifo_1_empty ? queue_1_enq_bits_readFromScalar : queue_dataOut_1_readFromScalar;
  assign queue_1_deq_bits_csrInterface_vl = _queue_fifo_1_empty ? queue_1_enq_bits_csrInterface_vl : queue_dataOut_1_csrInterface_vl;
  assign queue_1_deq_bits_csrInterface_vStart = _queue_fifo_1_empty ? queue_1_enq_bits_csrInterface_vStart : queue_dataOut_1_csrInterface_vStart;
  assign queue_1_deq_bits_csrInterface_vlmul = _queue_fifo_1_empty ? queue_1_enq_bits_csrInterface_vlmul : queue_dataOut_1_csrInterface_vlmul;
  assign queue_1_deq_bits_csrInterface_vSew = _queue_fifo_1_empty ? queue_1_enq_bits_csrInterface_vSew : queue_dataOut_1_csrInterface_vSew;
  assign queue_1_deq_bits_csrInterface_vxrm = _queue_fifo_1_empty ? queue_1_enq_bits_csrInterface_vxrm : queue_dataOut_1_csrInterface_vxrm;
  assign queue_1_deq_bits_csrInterface_vta = _queue_fifo_1_empty ? queue_1_enq_bits_csrInterface_vta : queue_dataOut_1_csrInterface_vta;
  assign queue_1_deq_bits_csrInterface_vma = _queue_fifo_1_empty ? queue_1_enq_bits_csrInterface_vma : queue_dataOut_1_csrInterface_vma;
  wire         laneVec_1_laneRequest_bits_issueInst = laneRequestSinkWire_1_ready & laneRequestSinkWire_1_valid;
  reg          releasePipe_pipe_v_1;
  wire         releasePipe_pipe_out_1_valid = releasePipe_pipe_v_1;
  wire         laneRequestSourceWire_1_ready;
  wire         validSource_1_valid = laneRequestSourceWire_1_ready & laneRequestSourceWire_1_valid;
  reg  [2:0]   tokenCheck_counter_1;
  wire [2:0]   tokenCheck_counterChange_1 = validSource_1_valid ? 3'h1 : 3'h7;
  assign tokenCheck_1 = ~(tokenCheck_counter_1[2]);
  assign laneRequestSourceWire_1_ready = tokenCheck_1;
  assign queue_1_enq_valid = validSink_1_valid;
  assign queue_1_enq_bits_instructionIndex = validSink_1_bits_instructionIndex;
  assign queue_1_enq_bits_decodeResult_specialSlot = validSink_1_bits_decodeResult_specialSlot;
  assign queue_1_enq_bits_decodeResult_topUop = validSink_1_bits_decodeResult_topUop;
  assign queue_1_enq_bits_decodeResult_popCount = validSink_1_bits_decodeResult_popCount;
  assign queue_1_enq_bits_decodeResult_ffo = validSink_1_bits_decodeResult_ffo;
  assign queue_1_enq_bits_decodeResult_average = validSink_1_bits_decodeResult_average;
  assign queue_1_enq_bits_decodeResult_reverse = validSink_1_bits_decodeResult_reverse;
  assign queue_1_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_1_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_1_enq_bits_decodeResult_scheduler = validSink_1_bits_decodeResult_scheduler;
  assign queue_1_enq_bits_decodeResult_sReadVD = validSink_1_bits_decodeResult_sReadVD;
  assign queue_1_enq_bits_decodeResult_vtype = validSink_1_bits_decodeResult_vtype;
  assign queue_1_enq_bits_decodeResult_sWrite = validSink_1_bits_decodeResult_sWrite;
  assign queue_1_enq_bits_decodeResult_crossRead = validSink_1_bits_decodeResult_crossRead;
  assign queue_1_enq_bits_decodeResult_crossWrite = validSink_1_bits_decodeResult_crossWrite;
  assign queue_1_enq_bits_decodeResult_maskUnit = validSink_1_bits_decodeResult_maskUnit;
  assign queue_1_enq_bits_decodeResult_special = validSink_1_bits_decodeResult_special;
  assign queue_1_enq_bits_decodeResult_saturate = validSink_1_bits_decodeResult_saturate;
  assign queue_1_enq_bits_decodeResult_vwmacc = validSink_1_bits_decodeResult_vwmacc;
  assign queue_1_enq_bits_decodeResult_readOnly = validSink_1_bits_decodeResult_readOnly;
  assign queue_1_enq_bits_decodeResult_maskSource = validSink_1_bits_decodeResult_maskSource;
  assign queue_1_enq_bits_decodeResult_maskDestination = validSink_1_bits_decodeResult_maskDestination;
  assign queue_1_enq_bits_decodeResult_maskLogic = validSink_1_bits_decodeResult_maskLogic;
  assign queue_1_enq_bits_decodeResult_uop = validSink_1_bits_decodeResult_uop;
  assign queue_1_enq_bits_decodeResult_iota = validSink_1_bits_decodeResult_iota;
  assign queue_1_enq_bits_decodeResult_mv = validSink_1_bits_decodeResult_mv;
  assign queue_1_enq_bits_decodeResult_extend = validSink_1_bits_decodeResult_extend;
  assign queue_1_enq_bits_decodeResult_unOrderWrite = validSink_1_bits_decodeResult_unOrderWrite;
  assign queue_1_enq_bits_decodeResult_compress = validSink_1_bits_decodeResult_compress;
  assign queue_1_enq_bits_decodeResult_gather16 = validSink_1_bits_decodeResult_gather16;
  assign queue_1_enq_bits_decodeResult_gather = validSink_1_bits_decodeResult_gather;
  assign queue_1_enq_bits_decodeResult_slid = validSink_1_bits_decodeResult_slid;
  assign queue_1_enq_bits_decodeResult_targetRd = validSink_1_bits_decodeResult_targetRd;
  assign queue_1_enq_bits_decodeResult_widenReduce = validSink_1_bits_decodeResult_widenReduce;
  assign queue_1_enq_bits_decodeResult_red = validSink_1_bits_decodeResult_red;
  assign queue_1_enq_bits_decodeResult_nr = validSink_1_bits_decodeResult_nr;
  assign queue_1_enq_bits_decodeResult_itype = validSink_1_bits_decodeResult_itype;
  assign queue_1_enq_bits_decodeResult_unsigned1 = validSink_1_bits_decodeResult_unsigned1;
  assign queue_1_enq_bits_decodeResult_unsigned0 = validSink_1_bits_decodeResult_unsigned0;
  assign queue_1_enq_bits_decodeResult_other = validSink_1_bits_decodeResult_other;
  assign queue_1_enq_bits_decodeResult_multiCycle = validSink_1_bits_decodeResult_multiCycle;
  assign queue_1_enq_bits_decodeResult_divider = validSink_1_bits_decodeResult_divider;
  assign queue_1_enq_bits_decodeResult_multiplier = validSink_1_bits_decodeResult_multiplier;
  assign queue_1_enq_bits_decodeResult_shift = validSink_1_bits_decodeResult_shift;
  assign queue_1_enq_bits_decodeResult_adder = validSink_1_bits_decodeResult_adder;
  assign queue_1_enq_bits_decodeResult_logic = validSink_1_bits_decodeResult_logic;
  assign queue_1_enq_bits_loadStore = validSink_1_bits_loadStore;
  assign queue_1_enq_bits_issueInst = validSink_1_bits_issueInst;
  assign queue_1_enq_bits_store = validSink_1_bits_store;
  assign queue_1_enq_bits_special = validSink_1_bits_special;
  assign queue_1_enq_bits_lsWholeReg = validSink_1_bits_lsWholeReg;
  assign queue_1_enq_bits_vs1 = validSink_1_bits_vs1;
  assign queue_1_enq_bits_vs2 = validSink_1_bits_vs2;
  assign queue_1_enq_bits_vd = validSink_1_bits_vd;
  assign queue_1_enq_bits_loadStoreEEW = validSink_1_bits_loadStoreEEW;
  assign queue_1_enq_bits_mask = validSink_1_bits_mask;
  assign queue_1_enq_bits_segment = validSink_1_bits_segment;
  assign queue_1_enq_bits_readFromScalar = validSink_1_bits_readFromScalar;
  assign queue_1_enq_bits_csrInterface_vl = validSink_1_bits_csrInterface_vl;
  assign queue_1_enq_bits_csrInterface_vStart = validSink_1_bits_csrInterface_vStart;
  assign queue_1_enq_bits_csrInterface_vlmul = validSink_1_bits_csrInterface_vlmul;
  assign queue_1_enq_bits_csrInterface_vSew = validSink_1_bits_csrInterface_vSew;
  assign queue_1_enq_bits_csrInterface_vxrm = validSink_1_bits_csrInterface_vxrm;
  assign queue_1_enq_bits_csrInterface_vta = validSink_1_bits_csrInterface_vta;
  assign queue_1_enq_bits_csrInterface_vma = validSink_1_bits_csrInterface_vma;
  reg          shifterReg_1_0_valid;
  assign validSink_1_valid = shifterReg_1_0_valid;
  reg  [2:0]   shifterReg_1_0_bits_instructionIndex;
  assign validSink_1_bits_instructionIndex = shifterReg_1_0_bits_instructionIndex;
  reg          shifterReg_1_0_bits_decodeResult_specialSlot;
  assign validSink_1_bits_decodeResult_specialSlot = shifterReg_1_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_1_0_bits_decodeResult_topUop;
  assign validSink_1_bits_decodeResult_topUop = shifterReg_1_0_bits_decodeResult_topUop;
  reg          shifterReg_1_0_bits_decodeResult_popCount;
  assign validSink_1_bits_decodeResult_popCount = shifterReg_1_0_bits_decodeResult_popCount;
  reg          shifterReg_1_0_bits_decodeResult_ffo;
  assign validSink_1_bits_decodeResult_ffo = shifterReg_1_0_bits_decodeResult_ffo;
  reg          shifterReg_1_0_bits_decodeResult_average;
  assign validSink_1_bits_decodeResult_average = shifterReg_1_0_bits_decodeResult_average;
  reg          shifterReg_1_0_bits_decodeResult_reverse;
  assign validSink_1_bits_decodeResult_reverse = shifterReg_1_0_bits_decodeResult_reverse;
  reg          shifterReg_1_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_1_bits_decodeResult_dontNeedExecuteInLane = shifterReg_1_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_1_0_bits_decodeResult_scheduler;
  assign validSink_1_bits_decodeResult_scheduler = shifterReg_1_0_bits_decodeResult_scheduler;
  reg          shifterReg_1_0_bits_decodeResult_sReadVD;
  assign validSink_1_bits_decodeResult_sReadVD = shifterReg_1_0_bits_decodeResult_sReadVD;
  reg          shifterReg_1_0_bits_decodeResult_vtype;
  assign validSink_1_bits_decodeResult_vtype = shifterReg_1_0_bits_decodeResult_vtype;
  reg          shifterReg_1_0_bits_decodeResult_sWrite;
  assign validSink_1_bits_decodeResult_sWrite = shifterReg_1_0_bits_decodeResult_sWrite;
  reg          shifterReg_1_0_bits_decodeResult_crossRead;
  assign validSink_1_bits_decodeResult_crossRead = shifterReg_1_0_bits_decodeResult_crossRead;
  reg          shifterReg_1_0_bits_decodeResult_crossWrite;
  assign validSink_1_bits_decodeResult_crossWrite = shifterReg_1_0_bits_decodeResult_crossWrite;
  reg          shifterReg_1_0_bits_decodeResult_maskUnit;
  assign validSink_1_bits_decodeResult_maskUnit = shifterReg_1_0_bits_decodeResult_maskUnit;
  reg          shifterReg_1_0_bits_decodeResult_special;
  assign validSink_1_bits_decodeResult_special = shifterReg_1_0_bits_decodeResult_special;
  reg          shifterReg_1_0_bits_decodeResult_saturate;
  assign validSink_1_bits_decodeResult_saturate = shifterReg_1_0_bits_decodeResult_saturate;
  reg          shifterReg_1_0_bits_decodeResult_vwmacc;
  assign validSink_1_bits_decodeResult_vwmacc = shifterReg_1_0_bits_decodeResult_vwmacc;
  reg          shifterReg_1_0_bits_decodeResult_readOnly;
  assign validSink_1_bits_decodeResult_readOnly = shifterReg_1_0_bits_decodeResult_readOnly;
  reg          shifterReg_1_0_bits_decodeResult_maskSource;
  assign validSink_1_bits_decodeResult_maskSource = shifterReg_1_0_bits_decodeResult_maskSource;
  reg          shifterReg_1_0_bits_decodeResult_maskDestination;
  assign validSink_1_bits_decodeResult_maskDestination = shifterReg_1_0_bits_decodeResult_maskDestination;
  reg          shifterReg_1_0_bits_decodeResult_maskLogic;
  assign validSink_1_bits_decodeResult_maskLogic = shifterReg_1_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_1_0_bits_decodeResult_uop;
  assign validSink_1_bits_decodeResult_uop = shifterReg_1_0_bits_decodeResult_uop;
  reg          shifterReg_1_0_bits_decodeResult_iota;
  assign validSink_1_bits_decodeResult_iota = shifterReg_1_0_bits_decodeResult_iota;
  reg          shifterReg_1_0_bits_decodeResult_mv;
  assign validSink_1_bits_decodeResult_mv = shifterReg_1_0_bits_decodeResult_mv;
  reg          shifterReg_1_0_bits_decodeResult_extend;
  assign validSink_1_bits_decodeResult_extend = shifterReg_1_0_bits_decodeResult_extend;
  reg          shifterReg_1_0_bits_decodeResult_unOrderWrite;
  assign validSink_1_bits_decodeResult_unOrderWrite = shifterReg_1_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_1_0_bits_decodeResult_compress;
  assign validSink_1_bits_decodeResult_compress = shifterReg_1_0_bits_decodeResult_compress;
  reg          shifterReg_1_0_bits_decodeResult_gather16;
  assign validSink_1_bits_decodeResult_gather16 = shifterReg_1_0_bits_decodeResult_gather16;
  reg          shifterReg_1_0_bits_decodeResult_gather;
  assign validSink_1_bits_decodeResult_gather = shifterReg_1_0_bits_decodeResult_gather;
  reg          shifterReg_1_0_bits_decodeResult_slid;
  assign validSink_1_bits_decodeResult_slid = shifterReg_1_0_bits_decodeResult_slid;
  reg          shifterReg_1_0_bits_decodeResult_targetRd;
  assign validSink_1_bits_decodeResult_targetRd = shifterReg_1_0_bits_decodeResult_targetRd;
  reg          shifterReg_1_0_bits_decodeResult_widenReduce;
  assign validSink_1_bits_decodeResult_widenReduce = shifterReg_1_0_bits_decodeResult_widenReduce;
  reg          shifterReg_1_0_bits_decodeResult_red;
  assign validSink_1_bits_decodeResult_red = shifterReg_1_0_bits_decodeResult_red;
  reg          shifterReg_1_0_bits_decodeResult_nr;
  assign validSink_1_bits_decodeResult_nr = shifterReg_1_0_bits_decodeResult_nr;
  reg          shifterReg_1_0_bits_decodeResult_itype;
  assign validSink_1_bits_decodeResult_itype = shifterReg_1_0_bits_decodeResult_itype;
  reg          shifterReg_1_0_bits_decodeResult_unsigned1;
  assign validSink_1_bits_decodeResult_unsigned1 = shifterReg_1_0_bits_decodeResult_unsigned1;
  reg          shifterReg_1_0_bits_decodeResult_unsigned0;
  assign validSink_1_bits_decodeResult_unsigned0 = shifterReg_1_0_bits_decodeResult_unsigned0;
  reg          shifterReg_1_0_bits_decodeResult_other;
  assign validSink_1_bits_decodeResult_other = shifterReg_1_0_bits_decodeResult_other;
  reg          shifterReg_1_0_bits_decodeResult_multiCycle;
  assign validSink_1_bits_decodeResult_multiCycle = shifterReg_1_0_bits_decodeResult_multiCycle;
  reg          shifterReg_1_0_bits_decodeResult_divider;
  assign validSink_1_bits_decodeResult_divider = shifterReg_1_0_bits_decodeResult_divider;
  reg          shifterReg_1_0_bits_decodeResult_multiplier;
  assign validSink_1_bits_decodeResult_multiplier = shifterReg_1_0_bits_decodeResult_multiplier;
  reg          shifterReg_1_0_bits_decodeResult_shift;
  assign validSink_1_bits_decodeResult_shift = shifterReg_1_0_bits_decodeResult_shift;
  reg          shifterReg_1_0_bits_decodeResult_adder;
  assign validSink_1_bits_decodeResult_adder = shifterReg_1_0_bits_decodeResult_adder;
  reg          shifterReg_1_0_bits_decodeResult_logic;
  assign validSink_1_bits_decodeResult_logic = shifterReg_1_0_bits_decodeResult_logic;
  reg          shifterReg_1_0_bits_loadStore;
  assign validSink_1_bits_loadStore = shifterReg_1_0_bits_loadStore;
  reg          shifterReg_1_0_bits_issueInst;
  assign validSink_1_bits_issueInst = shifterReg_1_0_bits_issueInst;
  reg          shifterReg_1_0_bits_store;
  assign validSink_1_bits_store = shifterReg_1_0_bits_store;
  reg          shifterReg_1_0_bits_special;
  assign validSink_1_bits_special = shifterReg_1_0_bits_special;
  reg          shifterReg_1_0_bits_lsWholeReg;
  assign validSink_1_bits_lsWholeReg = shifterReg_1_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_1_0_bits_vs1;
  assign validSink_1_bits_vs1 = shifterReg_1_0_bits_vs1;
  reg  [4:0]   shifterReg_1_0_bits_vs2;
  assign validSink_1_bits_vs2 = shifterReg_1_0_bits_vs2;
  reg  [4:0]   shifterReg_1_0_bits_vd;
  assign validSink_1_bits_vd = shifterReg_1_0_bits_vd;
  reg  [1:0]   shifterReg_1_0_bits_loadStoreEEW;
  assign validSink_1_bits_loadStoreEEW = shifterReg_1_0_bits_loadStoreEEW;
  reg          shifterReg_1_0_bits_mask;
  assign validSink_1_bits_mask = shifterReg_1_0_bits_mask;
  reg  [2:0]   shifterReg_1_0_bits_segment;
  assign validSink_1_bits_segment = shifterReg_1_0_bits_segment;
  reg  [31:0]  shifterReg_1_0_bits_readFromScalar;
  assign validSink_1_bits_readFromScalar = shifterReg_1_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_1_0_bits_csrInterface_vl;
  assign validSink_1_bits_csrInterface_vl = shifterReg_1_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_1_0_bits_csrInterface_vStart;
  assign validSink_1_bits_csrInterface_vStart = shifterReg_1_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_1_0_bits_csrInterface_vlmul;
  assign validSink_1_bits_csrInterface_vlmul = shifterReg_1_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_1_0_bits_csrInterface_vSew;
  assign validSink_1_bits_csrInterface_vSew = shifterReg_1_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_1_0_bits_csrInterface_vxrm;
  assign validSink_1_bits_csrInterface_vxrm = shifterReg_1_0_bits_csrInterface_vxrm;
  reg          shifterReg_1_0_bits_csrInterface_vta;
  assign validSink_1_bits_csrInterface_vta = shifterReg_1_0_bits_csrInterface_vta;
  reg          shifterReg_1_0_bits_csrInterface_vma;
  assign validSink_1_bits_csrInterface_vma = shifterReg_1_0_bits_csrInterface_vma;
  wire         shifterValid_1 = shifterReg_1_0_valid | validSource_1_valid;
  wire         validSink_2_valid;
  wire [2:0]   validSink_2_bits_instructionIndex;
  wire         validSink_2_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_2_bits_decodeResult_topUop;
  wire         validSink_2_bits_decodeResult_popCount;
  wire         validSink_2_bits_decodeResult_ffo;
  wire         validSink_2_bits_decodeResult_average;
  wire         validSink_2_bits_decodeResult_reverse;
  wire         validSink_2_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_2_bits_decodeResult_scheduler;
  wire         validSink_2_bits_decodeResult_sReadVD;
  wire         validSink_2_bits_decodeResult_vtype;
  wire         validSink_2_bits_decodeResult_sWrite;
  wire         validSink_2_bits_decodeResult_crossRead;
  wire         validSink_2_bits_decodeResult_crossWrite;
  wire         validSink_2_bits_decodeResult_maskUnit;
  wire         validSink_2_bits_decodeResult_special;
  wire         validSink_2_bits_decodeResult_saturate;
  wire         validSink_2_bits_decodeResult_vwmacc;
  wire         validSink_2_bits_decodeResult_readOnly;
  wire         validSink_2_bits_decodeResult_maskSource;
  wire         validSink_2_bits_decodeResult_maskDestination;
  wire         validSink_2_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_2_bits_decodeResult_uop;
  wire         validSink_2_bits_decodeResult_iota;
  wire         validSink_2_bits_decodeResult_mv;
  wire         validSink_2_bits_decodeResult_extend;
  wire         validSink_2_bits_decodeResult_unOrderWrite;
  wire         validSink_2_bits_decodeResult_compress;
  wire         validSink_2_bits_decodeResult_gather16;
  wire         validSink_2_bits_decodeResult_gather;
  wire         validSink_2_bits_decodeResult_slid;
  wire         validSink_2_bits_decodeResult_targetRd;
  wire         validSink_2_bits_decodeResult_widenReduce;
  wire         validSink_2_bits_decodeResult_red;
  wire         validSink_2_bits_decodeResult_nr;
  wire         validSink_2_bits_decodeResult_itype;
  wire         validSink_2_bits_decodeResult_unsigned1;
  wire         validSink_2_bits_decodeResult_unsigned0;
  wire         validSink_2_bits_decodeResult_other;
  wire         validSink_2_bits_decodeResult_multiCycle;
  wire         validSink_2_bits_decodeResult_divider;
  wire         validSink_2_bits_decodeResult_multiplier;
  wire         validSink_2_bits_decodeResult_shift;
  wire         validSink_2_bits_decodeResult_adder;
  wire         validSink_2_bits_decodeResult_logic;
  wire         validSink_2_bits_loadStore;
  wire         validSink_2_bits_issueInst;
  wire         validSink_2_bits_store;
  wire         validSink_2_bits_special;
  wire         validSink_2_bits_lsWholeReg;
  wire [4:0]   validSink_2_bits_vs1;
  wire [4:0]   validSink_2_bits_vs2;
  wire [4:0]   validSink_2_bits_vd;
  wire [1:0]   validSink_2_bits_loadStoreEEW;
  wire         validSink_2_bits_mask;
  wire [2:0]   validSink_2_bits_segment;
  wire [31:0]  validSink_2_bits_readFromScalar;
  wire [11:0]  validSink_2_bits_csrInterface_vl;
  wire [11:0]  validSink_2_bits_csrInterface_vStart;
  wire [2:0]   validSink_2_bits_csrInterface_vlmul;
  wire [1:0]   validSink_2_bits_csrInterface_vSew;
  wire [1:0]   validSink_2_bits_csrInterface_vxrm;
  wire         validSink_2_bits_csrInterface_vta;
  wire         validSink_2_bits_csrInterface_vma;
  wire         laneRequestSinkWire_2_valid = queue_2_deq_valid;
  wire [2:0]   laneRequestSinkWire_2_bits_instructionIndex = queue_2_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_2_bits_decodeResult_specialSlot = queue_2_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_2_bits_decodeResult_topUop = queue_2_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_2_bits_decodeResult_popCount = queue_2_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_2_bits_decodeResult_ffo = queue_2_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_2_bits_decodeResult_average = queue_2_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_2_bits_decodeResult_reverse = queue_2_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_2_bits_decodeResult_dontNeedExecuteInLane = queue_2_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_2_bits_decodeResult_scheduler = queue_2_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_2_bits_decodeResult_sReadVD = queue_2_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_2_bits_decodeResult_vtype = queue_2_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_2_bits_decodeResult_sWrite = queue_2_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_2_bits_decodeResult_crossRead = queue_2_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_2_bits_decodeResult_crossWrite = queue_2_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_2_bits_decodeResult_maskUnit = queue_2_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_2_bits_decodeResult_special = queue_2_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_2_bits_decodeResult_saturate = queue_2_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_2_bits_decodeResult_vwmacc = queue_2_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_2_bits_decodeResult_readOnly = queue_2_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_2_bits_decodeResult_maskSource = queue_2_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_2_bits_decodeResult_maskDestination = queue_2_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_2_bits_decodeResult_maskLogic = queue_2_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_2_bits_decodeResult_uop = queue_2_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_2_bits_decodeResult_iota = queue_2_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_2_bits_decodeResult_mv = queue_2_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_2_bits_decodeResult_extend = queue_2_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_2_bits_decodeResult_unOrderWrite = queue_2_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_2_bits_decodeResult_compress = queue_2_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_2_bits_decodeResult_gather16 = queue_2_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_2_bits_decodeResult_gather = queue_2_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_2_bits_decodeResult_slid = queue_2_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_2_bits_decodeResult_targetRd = queue_2_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_2_bits_decodeResult_widenReduce = queue_2_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_2_bits_decodeResult_red = queue_2_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_2_bits_decodeResult_nr = queue_2_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_2_bits_decodeResult_itype = queue_2_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_2_bits_decodeResult_unsigned1 = queue_2_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_2_bits_decodeResult_unsigned0 = queue_2_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_2_bits_decodeResult_other = queue_2_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_2_bits_decodeResult_multiCycle = queue_2_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_2_bits_decodeResult_divider = queue_2_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_2_bits_decodeResult_multiplier = queue_2_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_2_bits_decodeResult_shift = queue_2_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_2_bits_decodeResult_adder = queue_2_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_2_bits_decodeResult_logic = queue_2_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_2_bits_loadStore = queue_2_deq_bits_loadStore;
  wire         laneRequestSinkWire_2_bits_issueInst = queue_2_deq_bits_issueInst;
  wire         laneRequestSinkWire_2_bits_store = queue_2_deq_bits_store;
  wire         laneRequestSinkWire_2_bits_special = queue_2_deq_bits_special;
  wire         laneRequestSinkWire_2_bits_lsWholeReg = queue_2_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_2_bits_vs1 = queue_2_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_2_bits_vs2 = queue_2_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_2_bits_vd = queue_2_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_2_bits_loadStoreEEW = queue_2_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_2_bits_mask = queue_2_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_2_bits_segment = queue_2_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_2_bits_readFromScalar = queue_2_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_2_bits_csrInterface_vl = queue_2_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_2_bits_csrInterface_vStart = queue_2_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_2_bits_csrInterface_vlmul = queue_2_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_2_bits_csrInterface_vSew = queue_2_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_2_bits_csrInterface_vxrm = queue_2_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_2_bits_csrInterface_vta = queue_2_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_2_bits_csrInterface_vma = queue_2_deq_bits_csrInterface_vma;
  wire [1:0]   queue_2_enq_bits_csrInterface_vxrm;
  wire         queue_2_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi_6 = {queue_2_enq_bits_csrInterface_vxrm, queue_2_enq_bits_csrInterface_vta};
  wire         queue_2_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo_6 = {queue_dataIn_lo_hi_6, queue_2_enq_bits_csrInterface_vma};
  wire [2:0]   queue_2_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_2_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo_6 = {queue_2_enq_bits_csrInterface_vlmul, queue_2_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_2_enq_bits_csrInterface_vl;
  wire [11:0]  queue_2_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi_6 = {queue_2_enq_bits_csrInterface_vl, queue_2_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi_6 = {queue_dataIn_hi_hi_6, queue_dataIn_hi_lo_6};
  wire         queue_2_enq_bits_decodeResult_adder;
  wire         queue_2_enq_bits_decodeResult_logic;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo_2 = {queue_2_enq_bits_decodeResult_adder, queue_2_enq_bits_decodeResult_logic};
  wire         queue_2_enq_bits_decodeResult_divider;
  wire         queue_2_enq_bits_decodeResult_multiplier;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi_2 = {queue_2_enq_bits_decodeResult_divider, queue_2_enq_bits_decodeResult_multiplier};
  wire         queue_2_enq_bits_decodeResult_shift;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi_2 = {queue_dataIn_lo_lo_lo_hi_hi_2, queue_2_enq_bits_decodeResult_shift};
  wire [4:0]   queue_dataIn_lo_lo_lo_2 = {queue_dataIn_lo_lo_lo_hi_2, queue_dataIn_lo_lo_lo_lo_2};
  wire         queue_2_enq_bits_decodeResult_unsigned0;
  wire         queue_2_enq_bits_decodeResult_other;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi_2 = {queue_2_enq_bits_decodeResult_unsigned0, queue_2_enq_bits_decodeResult_other};
  wire         queue_2_enq_bits_decodeResult_multiCycle;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo_2 = {queue_dataIn_lo_lo_hi_lo_hi_2, queue_2_enq_bits_decodeResult_multiCycle};
  wire         queue_2_enq_bits_decodeResult_nr;
  wire         queue_2_enq_bits_decodeResult_itype;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi_2 = {queue_2_enq_bits_decodeResult_nr, queue_2_enq_bits_decodeResult_itype};
  wire         queue_2_enq_bits_decodeResult_unsigned1;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi_2 = {queue_dataIn_lo_lo_hi_hi_hi_2, queue_2_enq_bits_decodeResult_unsigned1};
  wire [5:0]   queue_dataIn_lo_lo_hi_4 = {queue_dataIn_lo_lo_hi_hi_2, queue_dataIn_lo_lo_hi_lo_2};
  wire [10:0]  queue_dataIn_lo_lo_4 = {queue_dataIn_lo_lo_hi_4, queue_dataIn_lo_lo_lo_2};
  wire         queue_2_enq_bits_decodeResult_widenReduce;
  wire         queue_2_enq_bits_decodeResult_red;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo_2 = {queue_2_enq_bits_decodeResult_widenReduce, queue_2_enq_bits_decodeResult_red};
  wire         queue_2_enq_bits_decodeResult_gather;
  wire         queue_2_enq_bits_decodeResult_slid;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi_2 = {queue_2_enq_bits_decodeResult_gather, queue_2_enq_bits_decodeResult_slid};
  wire         queue_2_enq_bits_decodeResult_targetRd;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi_2 = {queue_dataIn_lo_hi_lo_hi_hi_2, queue_2_enq_bits_decodeResult_targetRd};
  wire [4:0]   queue_dataIn_lo_hi_lo_4 = {queue_dataIn_lo_hi_lo_hi_2, queue_dataIn_lo_hi_lo_lo_2};
  wire         queue_2_enq_bits_decodeResult_unOrderWrite;
  wire         queue_2_enq_bits_decodeResult_compress;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi_2 = {queue_2_enq_bits_decodeResult_unOrderWrite, queue_2_enq_bits_decodeResult_compress};
  wire         queue_2_enq_bits_decodeResult_gather16;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo_2 = {queue_dataIn_lo_hi_hi_lo_hi_2, queue_2_enq_bits_decodeResult_gather16};
  wire         queue_2_enq_bits_decodeResult_iota;
  wire         queue_2_enq_bits_decodeResult_mv;
  wire [1:0]   queue_dataIn_lo_hi_hi_hi_hi_2 = {queue_2_enq_bits_decodeResult_iota, queue_2_enq_bits_decodeResult_mv};
  wire         queue_2_enq_bits_decodeResult_extend;
  wire [2:0]   queue_dataIn_lo_hi_hi_hi_2 = {queue_dataIn_lo_hi_hi_hi_hi_2, queue_2_enq_bits_decodeResult_extend};
  wire [5:0]   queue_dataIn_lo_hi_hi_4 = {queue_dataIn_lo_hi_hi_hi_2, queue_dataIn_lo_hi_hi_lo_2};
  wire [10:0]  queue_dataIn_lo_hi_7 = {queue_dataIn_lo_hi_hi_4, queue_dataIn_lo_hi_lo_4};
  wire [21:0]  queue_dataIn_lo_7 = {queue_dataIn_lo_hi_7, queue_dataIn_lo_lo_4};
  wire         queue_2_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_2_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_hi_lo_lo_lo_2 = {queue_2_enq_bits_decodeResult_maskLogic, queue_2_enq_bits_decodeResult_uop};
  wire         queue_2_enq_bits_decodeResult_readOnly;
  wire         queue_2_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi_2 = {queue_2_enq_bits_decodeResult_readOnly, queue_2_enq_bits_decodeResult_maskSource};
  wire         queue_2_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi_2 = {queue_dataIn_hi_lo_lo_hi_hi_2, queue_2_enq_bits_decodeResult_maskDestination};
  wire [7:0]   queue_dataIn_hi_lo_lo_4 = {queue_dataIn_hi_lo_lo_hi_2, queue_dataIn_hi_lo_lo_lo_2};
  wire         queue_2_enq_bits_decodeResult_special;
  wire         queue_2_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi_2 = {queue_2_enq_bits_decodeResult_special, queue_2_enq_bits_decodeResult_saturate};
  wire         queue_2_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo_2 = {queue_dataIn_hi_lo_hi_lo_hi_2, queue_2_enq_bits_decodeResult_vwmacc};
  wire         queue_2_enq_bits_decodeResult_crossRead;
  wire         queue_2_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi_2 = {queue_2_enq_bits_decodeResult_crossRead, queue_2_enq_bits_decodeResult_crossWrite};
  wire         queue_2_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi_2 = {queue_dataIn_hi_lo_hi_hi_hi_2, queue_2_enq_bits_decodeResult_maskUnit};
  wire [5:0]   queue_dataIn_hi_lo_hi_4 = {queue_dataIn_hi_lo_hi_hi_2, queue_dataIn_hi_lo_hi_lo_2};
  wire [13:0]  queue_dataIn_hi_lo_7 = {queue_dataIn_hi_lo_hi_4, queue_dataIn_hi_lo_lo_4};
  wire         queue_2_enq_bits_decodeResult_vtype;
  wire         queue_2_enq_bits_decodeResult_sWrite;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo_2 = {queue_2_enq_bits_decodeResult_vtype, queue_2_enq_bits_decodeResult_sWrite};
  wire         queue_2_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_2_enq_bits_decodeResult_scheduler;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi_2 = {queue_2_enq_bits_decodeResult_dontNeedExecuteInLane, queue_2_enq_bits_decodeResult_scheduler};
  wire         queue_2_enq_bits_decodeResult_sReadVD;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi_2 = {queue_dataIn_hi_hi_lo_hi_hi_2, queue_2_enq_bits_decodeResult_sReadVD};
  wire [4:0]   queue_dataIn_hi_hi_lo_4 = {queue_dataIn_hi_hi_lo_hi_2, queue_dataIn_hi_hi_lo_lo_2};
  wire         queue_2_enq_bits_decodeResult_ffo;
  wire         queue_2_enq_bits_decodeResult_average;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi_2 = {queue_2_enq_bits_decodeResult_ffo, queue_2_enq_bits_decodeResult_average};
  wire         queue_2_enq_bits_decodeResult_reverse;
  wire [2:0]   queue_dataIn_hi_hi_hi_lo_2 = {queue_dataIn_hi_hi_hi_lo_hi_2, queue_2_enq_bits_decodeResult_reverse};
  wire         queue_2_enq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_2_enq_bits_decodeResult_topUop;
  wire [5:0]   queue_dataIn_hi_hi_hi_hi_hi_2 = {queue_2_enq_bits_decodeResult_specialSlot, queue_2_enq_bits_decodeResult_topUop};
  wire         queue_2_enq_bits_decodeResult_popCount;
  wire [6:0]   queue_dataIn_hi_hi_hi_hi_2 = {queue_dataIn_hi_hi_hi_hi_hi_2, queue_2_enq_bits_decodeResult_popCount};
  wire [9:0]   queue_dataIn_hi_hi_hi_4 = {queue_dataIn_hi_hi_hi_hi_2, queue_dataIn_hi_hi_hi_lo_2};
  wire [14:0]  queue_dataIn_hi_hi_7 = {queue_dataIn_hi_hi_hi_4, queue_dataIn_hi_hi_lo_4};
  wire [28:0]  queue_dataIn_hi_7 = {queue_dataIn_hi_hi_7, queue_dataIn_hi_lo_7};
  wire [2:0]   queue_2_enq_bits_segment;
  wire [31:0]  queue_2_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_5 = {queue_2_enq_bits_segment, queue_2_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_5 = {queue_dataIn_lo_lo_hi_5, queue_dataIn_hi_6, queue_dataIn_lo_6};
  wire [1:0]   queue_2_enq_bits_loadStoreEEW;
  wire         queue_2_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_5 = {queue_2_enq_bits_loadStoreEEW, queue_2_enq_bits_mask};
  wire [4:0]   queue_2_enq_bits_vs2;
  wire [4:0]   queue_2_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_5 = {queue_2_enq_bits_vs2, queue_2_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_8 = {queue_dataIn_lo_hi_hi_5, queue_dataIn_lo_hi_lo_5};
  wire [80:0]  queue_dataIn_lo_8 = {queue_dataIn_lo_hi_8, queue_dataIn_lo_lo_5};
  wire         queue_2_enq_bits_lsWholeReg;
  wire [4:0]   queue_2_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_5 = {queue_2_enq_bits_lsWholeReg, queue_2_enq_bits_vs1};
  wire         queue_2_enq_bits_store;
  wire         queue_2_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_5 = {queue_2_enq_bits_store, queue_2_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_8 = {queue_dataIn_hi_lo_hi_5, queue_dataIn_hi_lo_lo_5};
  wire         queue_2_enq_bits_loadStore;
  wire         queue_2_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_5 = {queue_2_enq_bits_loadStore, queue_2_enq_bits_issueInst};
  wire [2:0]   queue_2_enq_bits_instructionIndex;
  wire [53:0]  queue_dataIn_hi_hi_hi_5 = {queue_2_enq_bits_instructionIndex, queue_dataIn_hi_7, queue_dataIn_lo_7};
  wire [55:0]  queue_dataIn_hi_hi_8 = {queue_dataIn_hi_hi_hi_5, queue_dataIn_hi_hi_lo_5};
  wire [63:0]  queue_dataIn_hi_8 = {queue_dataIn_hi_hi_8, queue_dataIn_hi_lo_8};
  wire [144:0] queue_dataIn_2 = {queue_dataIn_hi_8, queue_dataIn_lo_8};
  wire         queue_dataOut_2_csrInterface_vma = _queue_fifo_2_data_out[0];
  wire         queue_dataOut_2_csrInterface_vta = _queue_fifo_2_data_out[1];
  wire [1:0]   queue_dataOut_2_csrInterface_vxrm = _queue_fifo_2_data_out[3:2];
  wire [1:0]   queue_dataOut_2_csrInterface_vSew = _queue_fifo_2_data_out[5:4];
  wire [2:0]   queue_dataOut_2_csrInterface_vlmul = _queue_fifo_2_data_out[8:6];
  wire [11:0]  queue_dataOut_2_csrInterface_vStart = _queue_fifo_2_data_out[20:9];
  wire [11:0]  queue_dataOut_2_csrInterface_vl = _queue_fifo_2_data_out[32:21];
  wire [31:0]  queue_dataOut_2_readFromScalar = _queue_fifo_2_data_out[64:33];
  wire [2:0]   queue_dataOut_2_segment = _queue_fifo_2_data_out[67:65];
  wire         queue_dataOut_2_mask = _queue_fifo_2_data_out[68];
  wire [1:0]   queue_dataOut_2_loadStoreEEW = _queue_fifo_2_data_out[70:69];
  wire [4:0]   queue_dataOut_2_vd = _queue_fifo_2_data_out[75:71];
  wire [4:0]   queue_dataOut_2_vs2 = _queue_fifo_2_data_out[80:76];
  wire [4:0]   queue_dataOut_2_vs1 = _queue_fifo_2_data_out[85:81];
  wire         queue_dataOut_2_lsWholeReg = _queue_fifo_2_data_out[86];
  wire         queue_dataOut_2_special = _queue_fifo_2_data_out[87];
  wire         queue_dataOut_2_store = _queue_fifo_2_data_out[88];
  wire         queue_dataOut_2_issueInst = _queue_fifo_2_data_out[89];
  wire         queue_dataOut_2_loadStore = _queue_fifo_2_data_out[90];
  wire         queue_dataOut_2_decodeResult_logic = _queue_fifo_2_data_out[91];
  wire         queue_dataOut_2_decodeResult_adder = _queue_fifo_2_data_out[92];
  wire         queue_dataOut_2_decodeResult_shift = _queue_fifo_2_data_out[93];
  wire         queue_dataOut_2_decodeResult_multiplier = _queue_fifo_2_data_out[94];
  wire         queue_dataOut_2_decodeResult_divider = _queue_fifo_2_data_out[95];
  wire         queue_dataOut_2_decodeResult_multiCycle = _queue_fifo_2_data_out[96];
  wire         queue_dataOut_2_decodeResult_other = _queue_fifo_2_data_out[97];
  wire         queue_dataOut_2_decodeResult_unsigned0 = _queue_fifo_2_data_out[98];
  wire         queue_dataOut_2_decodeResult_unsigned1 = _queue_fifo_2_data_out[99];
  wire         queue_dataOut_2_decodeResult_itype = _queue_fifo_2_data_out[100];
  wire         queue_dataOut_2_decodeResult_nr = _queue_fifo_2_data_out[101];
  wire         queue_dataOut_2_decodeResult_red = _queue_fifo_2_data_out[102];
  wire         queue_dataOut_2_decodeResult_widenReduce = _queue_fifo_2_data_out[103];
  wire         queue_dataOut_2_decodeResult_targetRd = _queue_fifo_2_data_out[104];
  wire         queue_dataOut_2_decodeResult_slid = _queue_fifo_2_data_out[105];
  wire         queue_dataOut_2_decodeResult_gather = _queue_fifo_2_data_out[106];
  wire         queue_dataOut_2_decodeResult_gather16 = _queue_fifo_2_data_out[107];
  wire         queue_dataOut_2_decodeResult_compress = _queue_fifo_2_data_out[108];
  wire         queue_dataOut_2_decodeResult_unOrderWrite = _queue_fifo_2_data_out[109];
  wire         queue_dataOut_2_decodeResult_extend = _queue_fifo_2_data_out[110];
  wire         queue_dataOut_2_decodeResult_mv = _queue_fifo_2_data_out[111];
  wire         queue_dataOut_2_decodeResult_iota = _queue_fifo_2_data_out[112];
  wire [3:0]   queue_dataOut_2_decodeResult_uop = _queue_fifo_2_data_out[116:113];
  wire         queue_dataOut_2_decodeResult_maskLogic = _queue_fifo_2_data_out[117];
  wire         queue_dataOut_2_decodeResult_maskDestination = _queue_fifo_2_data_out[118];
  wire         queue_dataOut_2_decodeResult_maskSource = _queue_fifo_2_data_out[119];
  wire         queue_dataOut_2_decodeResult_readOnly = _queue_fifo_2_data_out[120];
  wire         queue_dataOut_2_decodeResult_vwmacc = _queue_fifo_2_data_out[121];
  wire         queue_dataOut_2_decodeResult_saturate = _queue_fifo_2_data_out[122];
  wire         queue_dataOut_2_decodeResult_special = _queue_fifo_2_data_out[123];
  wire         queue_dataOut_2_decodeResult_maskUnit = _queue_fifo_2_data_out[124];
  wire         queue_dataOut_2_decodeResult_crossWrite = _queue_fifo_2_data_out[125];
  wire         queue_dataOut_2_decodeResult_crossRead = _queue_fifo_2_data_out[126];
  wire         queue_dataOut_2_decodeResult_sWrite = _queue_fifo_2_data_out[127];
  wire         queue_dataOut_2_decodeResult_vtype = _queue_fifo_2_data_out[128];
  wire         queue_dataOut_2_decodeResult_sReadVD = _queue_fifo_2_data_out[129];
  wire         queue_dataOut_2_decodeResult_scheduler = _queue_fifo_2_data_out[130];
  wire         queue_dataOut_2_decodeResult_dontNeedExecuteInLane = _queue_fifo_2_data_out[131];
  wire         queue_dataOut_2_decodeResult_reverse = _queue_fifo_2_data_out[132];
  wire         queue_dataOut_2_decodeResult_average = _queue_fifo_2_data_out[133];
  wire         queue_dataOut_2_decodeResult_ffo = _queue_fifo_2_data_out[134];
  wire         queue_dataOut_2_decodeResult_popCount = _queue_fifo_2_data_out[135];
  wire [4:0]   queue_dataOut_2_decodeResult_topUop = _queue_fifo_2_data_out[140:136];
  wire         queue_dataOut_2_decodeResult_specialSlot = _queue_fifo_2_data_out[141];
  wire [2:0]   queue_dataOut_2_instructionIndex = _queue_fifo_2_data_out[144:142];
  wire         queue_2_enq_ready = ~_queue_fifo_2_full;
  wire         queue_2_enq_valid;
  assign queue_2_deq_valid = ~_queue_fifo_2_empty | queue_2_enq_valid;
  assign queue_2_deq_bits_instructionIndex = _queue_fifo_2_empty ? queue_2_enq_bits_instructionIndex : queue_dataOut_2_instructionIndex;
  assign queue_2_deq_bits_decodeResult_specialSlot = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_specialSlot : queue_dataOut_2_decodeResult_specialSlot;
  assign queue_2_deq_bits_decodeResult_topUop = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_topUop : queue_dataOut_2_decodeResult_topUop;
  assign queue_2_deq_bits_decodeResult_popCount = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_popCount : queue_dataOut_2_decodeResult_popCount;
  assign queue_2_deq_bits_decodeResult_ffo = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_ffo : queue_dataOut_2_decodeResult_ffo;
  assign queue_2_deq_bits_decodeResult_average = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_average : queue_dataOut_2_decodeResult_average;
  assign queue_2_deq_bits_decodeResult_reverse = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_reverse : queue_dataOut_2_decodeResult_reverse;
  assign queue_2_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_2_decodeResult_dontNeedExecuteInLane;
  assign queue_2_deq_bits_decodeResult_scheduler = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_scheduler : queue_dataOut_2_decodeResult_scheduler;
  assign queue_2_deq_bits_decodeResult_sReadVD = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_sReadVD : queue_dataOut_2_decodeResult_sReadVD;
  assign queue_2_deq_bits_decodeResult_vtype = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_vtype : queue_dataOut_2_decodeResult_vtype;
  assign queue_2_deq_bits_decodeResult_sWrite = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_sWrite : queue_dataOut_2_decodeResult_sWrite;
  assign queue_2_deq_bits_decodeResult_crossRead = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_crossRead : queue_dataOut_2_decodeResult_crossRead;
  assign queue_2_deq_bits_decodeResult_crossWrite = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_crossWrite : queue_dataOut_2_decodeResult_crossWrite;
  assign queue_2_deq_bits_decodeResult_maskUnit = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_maskUnit : queue_dataOut_2_decodeResult_maskUnit;
  assign queue_2_deq_bits_decodeResult_special = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_special : queue_dataOut_2_decodeResult_special;
  assign queue_2_deq_bits_decodeResult_saturate = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_saturate : queue_dataOut_2_decodeResult_saturate;
  assign queue_2_deq_bits_decodeResult_vwmacc = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_vwmacc : queue_dataOut_2_decodeResult_vwmacc;
  assign queue_2_deq_bits_decodeResult_readOnly = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_readOnly : queue_dataOut_2_decodeResult_readOnly;
  assign queue_2_deq_bits_decodeResult_maskSource = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_maskSource : queue_dataOut_2_decodeResult_maskSource;
  assign queue_2_deq_bits_decodeResult_maskDestination = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_maskDestination : queue_dataOut_2_decodeResult_maskDestination;
  assign queue_2_deq_bits_decodeResult_maskLogic = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_maskLogic : queue_dataOut_2_decodeResult_maskLogic;
  assign queue_2_deq_bits_decodeResult_uop = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_uop : queue_dataOut_2_decodeResult_uop;
  assign queue_2_deq_bits_decodeResult_iota = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_iota : queue_dataOut_2_decodeResult_iota;
  assign queue_2_deq_bits_decodeResult_mv = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_mv : queue_dataOut_2_decodeResult_mv;
  assign queue_2_deq_bits_decodeResult_extend = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_extend : queue_dataOut_2_decodeResult_extend;
  assign queue_2_deq_bits_decodeResult_unOrderWrite = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_unOrderWrite : queue_dataOut_2_decodeResult_unOrderWrite;
  assign queue_2_deq_bits_decodeResult_compress = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_compress : queue_dataOut_2_decodeResult_compress;
  assign queue_2_deq_bits_decodeResult_gather16 = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_gather16 : queue_dataOut_2_decodeResult_gather16;
  assign queue_2_deq_bits_decodeResult_gather = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_gather : queue_dataOut_2_decodeResult_gather;
  assign queue_2_deq_bits_decodeResult_slid = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_slid : queue_dataOut_2_decodeResult_slid;
  assign queue_2_deq_bits_decodeResult_targetRd = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_targetRd : queue_dataOut_2_decodeResult_targetRd;
  assign queue_2_deq_bits_decodeResult_widenReduce = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_widenReduce : queue_dataOut_2_decodeResult_widenReduce;
  assign queue_2_deq_bits_decodeResult_red = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_red : queue_dataOut_2_decodeResult_red;
  assign queue_2_deq_bits_decodeResult_nr = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_nr : queue_dataOut_2_decodeResult_nr;
  assign queue_2_deq_bits_decodeResult_itype = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_itype : queue_dataOut_2_decodeResult_itype;
  assign queue_2_deq_bits_decodeResult_unsigned1 = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_unsigned1 : queue_dataOut_2_decodeResult_unsigned1;
  assign queue_2_deq_bits_decodeResult_unsigned0 = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_unsigned0 : queue_dataOut_2_decodeResult_unsigned0;
  assign queue_2_deq_bits_decodeResult_other = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_other : queue_dataOut_2_decodeResult_other;
  assign queue_2_deq_bits_decodeResult_multiCycle = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_multiCycle : queue_dataOut_2_decodeResult_multiCycle;
  assign queue_2_deq_bits_decodeResult_divider = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_divider : queue_dataOut_2_decodeResult_divider;
  assign queue_2_deq_bits_decodeResult_multiplier = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_multiplier : queue_dataOut_2_decodeResult_multiplier;
  assign queue_2_deq_bits_decodeResult_shift = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_shift : queue_dataOut_2_decodeResult_shift;
  assign queue_2_deq_bits_decodeResult_adder = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_adder : queue_dataOut_2_decodeResult_adder;
  assign queue_2_deq_bits_decodeResult_logic = _queue_fifo_2_empty ? queue_2_enq_bits_decodeResult_logic : queue_dataOut_2_decodeResult_logic;
  assign queue_2_deq_bits_loadStore = _queue_fifo_2_empty ? queue_2_enq_bits_loadStore : queue_dataOut_2_loadStore;
  assign queue_2_deq_bits_issueInst = _queue_fifo_2_empty ? queue_2_enq_bits_issueInst : queue_dataOut_2_issueInst;
  assign queue_2_deq_bits_store = _queue_fifo_2_empty ? queue_2_enq_bits_store : queue_dataOut_2_store;
  assign queue_2_deq_bits_special = _queue_fifo_2_empty ? queue_2_enq_bits_special : queue_dataOut_2_special;
  assign queue_2_deq_bits_lsWholeReg = _queue_fifo_2_empty ? queue_2_enq_bits_lsWholeReg : queue_dataOut_2_lsWholeReg;
  assign queue_2_deq_bits_vs1 = _queue_fifo_2_empty ? queue_2_enq_bits_vs1 : queue_dataOut_2_vs1;
  assign queue_2_deq_bits_vs2 = _queue_fifo_2_empty ? queue_2_enq_bits_vs2 : queue_dataOut_2_vs2;
  assign queue_2_deq_bits_vd = _queue_fifo_2_empty ? queue_2_enq_bits_vd : queue_dataOut_2_vd;
  assign queue_2_deq_bits_loadStoreEEW = _queue_fifo_2_empty ? queue_2_enq_bits_loadStoreEEW : queue_dataOut_2_loadStoreEEW;
  assign queue_2_deq_bits_mask = _queue_fifo_2_empty ? queue_2_enq_bits_mask : queue_dataOut_2_mask;
  assign queue_2_deq_bits_segment = _queue_fifo_2_empty ? queue_2_enq_bits_segment : queue_dataOut_2_segment;
  assign queue_2_deq_bits_readFromScalar = _queue_fifo_2_empty ? queue_2_enq_bits_readFromScalar : queue_dataOut_2_readFromScalar;
  assign queue_2_deq_bits_csrInterface_vl = _queue_fifo_2_empty ? queue_2_enq_bits_csrInterface_vl : queue_dataOut_2_csrInterface_vl;
  assign queue_2_deq_bits_csrInterface_vStart = _queue_fifo_2_empty ? queue_2_enq_bits_csrInterface_vStart : queue_dataOut_2_csrInterface_vStart;
  assign queue_2_deq_bits_csrInterface_vlmul = _queue_fifo_2_empty ? queue_2_enq_bits_csrInterface_vlmul : queue_dataOut_2_csrInterface_vlmul;
  assign queue_2_deq_bits_csrInterface_vSew = _queue_fifo_2_empty ? queue_2_enq_bits_csrInterface_vSew : queue_dataOut_2_csrInterface_vSew;
  assign queue_2_deq_bits_csrInterface_vxrm = _queue_fifo_2_empty ? queue_2_enq_bits_csrInterface_vxrm : queue_dataOut_2_csrInterface_vxrm;
  assign queue_2_deq_bits_csrInterface_vta = _queue_fifo_2_empty ? queue_2_enq_bits_csrInterface_vta : queue_dataOut_2_csrInterface_vta;
  assign queue_2_deq_bits_csrInterface_vma = _queue_fifo_2_empty ? queue_2_enq_bits_csrInterface_vma : queue_dataOut_2_csrInterface_vma;
  wire         laneVec_2_laneRequest_bits_issueInst = laneRequestSinkWire_2_ready & laneRequestSinkWire_2_valid;
  reg          releasePipe_pipe_v_2;
  wire         releasePipe_pipe_out_2_valid = releasePipe_pipe_v_2;
  wire         laneRequestSourceWire_2_ready;
  wire         validSource_2_valid = laneRequestSourceWire_2_ready & laneRequestSourceWire_2_valid;
  reg  [2:0]   tokenCheck_counter_2;
  wire [2:0]   tokenCheck_counterChange_2 = validSource_2_valid ? 3'h1 : 3'h7;
  assign tokenCheck_2 = ~(tokenCheck_counter_2[2]);
  assign laneRequestSourceWire_2_ready = tokenCheck_2;
  assign queue_2_enq_valid = validSink_2_valid;
  assign queue_2_enq_bits_instructionIndex = validSink_2_bits_instructionIndex;
  assign queue_2_enq_bits_decodeResult_specialSlot = validSink_2_bits_decodeResult_specialSlot;
  assign queue_2_enq_bits_decodeResult_topUop = validSink_2_bits_decodeResult_topUop;
  assign queue_2_enq_bits_decodeResult_popCount = validSink_2_bits_decodeResult_popCount;
  assign queue_2_enq_bits_decodeResult_ffo = validSink_2_bits_decodeResult_ffo;
  assign queue_2_enq_bits_decodeResult_average = validSink_2_bits_decodeResult_average;
  assign queue_2_enq_bits_decodeResult_reverse = validSink_2_bits_decodeResult_reverse;
  assign queue_2_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_2_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_2_enq_bits_decodeResult_scheduler = validSink_2_bits_decodeResult_scheduler;
  assign queue_2_enq_bits_decodeResult_sReadVD = validSink_2_bits_decodeResult_sReadVD;
  assign queue_2_enq_bits_decodeResult_vtype = validSink_2_bits_decodeResult_vtype;
  assign queue_2_enq_bits_decodeResult_sWrite = validSink_2_bits_decodeResult_sWrite;
  assign queue_2_enq_bits_decodeResult_crossRead = validSink_2_bits_decodeResult_crossRead;
  assign queue_2_enq_bits_decodeResult_crossWrite = validSink_2_bits_decodeResult_crossWrite;
  assign queue_2_enq_bits_decodeResult_maskUnit = validSink_2_bits_decodeResult_maskUnit;
  assign queue_2_enq_bits_decodeResult_special = validSink_2_bits_decodeResult_special;
  assign queue_2_enq_bits_decodeResult_saturate = validSink_2_bits_decodeResult_saturate;
  assign queue_2_enq_bits_decodeResult_vwmacc = validSink_2_bits_decodeResult_vwmacc;
  assign queue_2_enq_bits_decodeResult_readOnly = validSink_2_bits_decodeResult_readOnly;
  assign queue_2_enq_bits_decodeResult_maskSource = validSink_2_bits_decodeResult_maskSource;
  assign queue_2_enq_bits_decodeResult_maskDestination = validSink_2_bits_decodeResult_maskDestination;
  assign queue_2_enq_bits_decodeResult_maskLogic = validSink_2_bits_decodeResult_maskLogic;
  assign queue_2_enq_bits_decodeResult_uop = validSink_2_bits_decodeResult_uop;
  assign queue_2_enq_bits_decodeResult_iota = validSink_2_bits_decodeResult_iota;
  assign queue_2_enq_bits_decodeResult_mv = validSink_2_bits_decodeResult_mv;
  assign queue_2_enq_bits_decodeResult_extend = validSink_2_bits_decodeResult_extend;
  assign queue_2_enq_bits_decodeResult_unOrderWrite = validSink_2_bits_decodeResult_unOrderWrite;
  assign queue_2_enq_bits_decodeResult_compress = validSink_2_bits_decodeResult_compress;
  assign queue_2_enq_bits_decodeResult_gather16 = validSink_2_bits_decodeResult_gather16;
  assign queue_2_enq_bits_decodeResult_gather = validSink_2_bits_decodeResult_gather;
  assign queue_2_enq_bits_decodeResult_slid = validSink_2_bits_decodeResult_slid;
  assign queue_2_enq_bits_decodeResult_targetRd = validSink_2_bits_decodeResult_targetRd;
  assign queue_2_enq_bits_decodeResult_widenReduce = validSink_2_bits_decodeResult_widenReduce;
  assign queue_2_enq_bits_decodeResult_red = validSink_2_bits_decodeResult_red;
  assign queue_2_enq_bits_decodeResult_nr = validSink_2_bits_decodeResult_nr;
  assign queue_2_enq_bits_decodeResult_itype = validSink_2_bits_decodeResult_itype;
  assign queue_2_enq_bits_decodeResult_unsigned1 = validSink_2_bits_decodeResult_unsigned1;
  assign queue_2_enq_bits_decodeResult_unsigned0 = validSink_2_bits_decodeResult_unsigned0;
  assign queue_2_enq_bits_decodeResult_other = validSink_2_bits_decodeResult_other;
  assign queue_2_enq_bits_decodeResult_multiCycle = validSink_2_bits_decodeResult_multiCycle;
  assign queue_2_enq_bits_decodeResult_divider = validSink_2_bits_decodeResult_divider;
  assign queue_2_enq_bits_decodeResult_multiplier = validSink_2_bits_decodeResult_multiplier;
  assign queue_2_enq_bits_decodeResult_shift = validSink_2_bits_decodeResult_shift;
  assign queue_2_enq_bits_decodeResult_adder = validSink_2_bits_decodeResult_adder;
  assign queue_2_enq_bits_decodeResult_logic = validSink_2_bits_decodeResult_logic;
  assign queue_2_enq_bits_loadStore = validSink_2_bits_loadStore;
  assign queue_2_enq_bits_issueInst = validSink_2_bits_issueInst;
  assign queue_2_enq_bits_store = validSink_2_bits_store;
  assign queue_2_enq_bits_special = validSink_2_bits_special;
  assign queue_2_enq_bits_lsWholeReg = validSink_2_bits_lsWholeReg;
  assign queue_2_enq_bits_vs1 = validSink_2_bits_vs1;
  assign queue_2_enq_bits_vs2 = validSink_2_bits_vs2;
  assign queue_2_enq_bits_vd = validSink_2_bits_vd;
  assign queue_2_enq_bits_loadStoreEEW = validSink_2_bits_loadStoreEEW;
  assign queue_2_enq_bits_mask = validSink_2_bits_mask;
  assign queue_2_enq_bits_segment = validSink_2_bits_segment;
  assign queue_2_enq_bits_readFromScalar = validSink_2_bits_readFromScalar;
  assign queue_2_enq_bits_csrInterface_vl = validSink_2_bits_csrInterface_vl;
  assign queue_2_enq_bits_csrInterface_vStart = validSink_2_bits_csrInterface_vStart;
  assign queue_2_enq_bits_csrInterface_vlmul = validSink_2_bits_csrInterface_vlmul;
  assign queue_2_enq_bits_csrInterface_vSew = validSink_2_bits_csrInterface_vSew;
  assign queue_2_enq_bits_csrInterface_vxrm = validSink_2_bits_csrInterface_vxrm;
  assign queue_2_enq_bits_csrInterface_vta = validSink_2_bits_csrInterface_vta;
  assign queue_2_enq_bits_csrInterface_vma = validSink_2_bits_csrInterface_vma;
  reg          shifterReg_2_0_valid;
  assign validSink_2_valid = shifterReg_2_0_valid;
  reg  [2:0]   shifterReg_2_0_bits_instructionIndex;
  assign validSink_2_bits_instructionIndex = shifterReg_2_0_bits_instructionIndex;
  reg          shifterReg_2_0_bits_decodeResult_specialSlot;
  assign validSink_2_bits_decodeResult_specialSlot = shifterReg_2_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_2_0_bits_decodeResult_topUop;
  assign validSink_2_bits_decodeResult_topUop = shifterReg_2_0_bits_decodeResult_topUop;
  reg          shifterReg_2_0_bits_decodeResult_popCount;
  assign validSink_2_bits_decodeResult_popCount = shifterReg_2_0_bits_decodeResult_popCount;
  reg          shifterReg_2_0_bits_decodeResult_ffo;
  assign validSink_2_bits_decodeResult_ffo = shifterReg_2_0_bits_decodeResult_ffo;
  reg          shifterReg_2_0_bits_decodeResult_average;
  assign validSink_2_bits_decodeResult_average = shifterReg_2_0_bits_decodeResult_average;
  reg          shifterReg_2_0_bits_decodeResult_reverse;
  assign validSink_2_bits_decodeResult_reverse = shifterReg_2_0_bits_decodeResult_reverse;
  reg          shifterReg_2_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_2_bits_decodeResult_dontNeedExecuteInLane = shifterReg_2_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_2_0_bits_decodeResult_scheduler;
  assign validSink_2_bits_decodeResult_scheduler = shifterReg_2_0_bits_decodeResult_scheduler;
  reg          shifterReg_2_0_bits_decodeResult_sReadVD;
  assign validSink_2_bits_decodeResult_sReadVD = shifterReg_2_0_bits_decodeResult_sReadVD;
  reg          shifterReg_2_0_bits_decodeResult_vtype;
  assign validSink_2_bits_decodeResult_vtype = shifterReg_2_0_bits_decodeResult_vtype;
  reg          shifterReg_2_0_bits_decodeResult_sWrite;
  assign validSink_2_bits_decodeResult_sWrite = shifterReg_2_0_bits_decodeResult_sWrite;
  reg          shifterReg_2_0_bits_decodeResult_crossRead;
  assign validSink_2_bits_decodeResult_crossRead = shifterReg_2_0_bits_decodeResult_crossRead;
  reg          shifterReg_2_0_bits_decodeResult_crossWrite;
  assign validSink_2_bits_decodeResult_crossWrite = shifterReg_2_0_bits_decodeResult_crossWrite;
  reg          shifterReg_2_0_bits_decodeResult_maskUnit;
  assign validSink_2_bits_decodeResult_maskUnit = shifterReg_2_0_bits_decodeResult_maskUnit;
  reg          shifterReg_2_0_bits_decodeResult_special;
  assign validSink_2_bits_decodeResult_special = shifterReg_2_0_bits_decodeResult_special;
  reg          shifterReg_2_0_bits_decodeResult_saturate;
  assign validSink_2_bits_decodeResult_saturate = shifterReg_2_0_bits_decodeResult_saturate;
  reg          shifterReg_2_0_bits_decodeResult_vwmacc;
  assign validSink_2_bits_decodeResult_vwmacc = shifterReg_2_0_bits_decodeResult_vwmacc;
  reg          shifterReg_2_0_bits_decodeResult_readOnly;
  assign validSink_2_bits_decodeResult_readOnly = shifterReg_2_0_bits_decodeResult_readOnly;
  reg          shifterReg_2_0_bits_decodeResult_maskSource;
  assign validSink_2_bits_decodeResult_maskSource = shifterReg_2_0_bits_decodeResult_maskSource;
  reg          shifterReg_2_0_bits_decodeResult_maskDestination;
  assign validSink_2_bits_decodeResult_maskDestination = shifterReg_2_0_bits_decodeResult_maskDestination;
  reg          shifterReg_2_0_bits_decodeResult_maskLogic;
  assign validSink_2_bits_decodeResult_maskLogic = shifterReg_2_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_2_0_bits_decodeResult_uop;
  assign validSink_2_bits_decodeResult_uop = shifterReg_2_0_bits_decodeResult_uop;
  reg          shifterReg_2_0_bits_decodeResult_iota;
  assign validSink_2_bits_decodeResult_iota = shifterReg_2_0_bits_decodeResult_iota;
  reg          shifterReg_2_0_bits_decodeResult_mv;
  assign validSink_2_bits_decodeResult_mv = shifterReg_2_0_bits_decodeResult_mv;
  reg          shifterReg_2_0_bits_decodeResult_extend;
  assign validSink_2_bits_decodeResult_extend = shifterReg_2_0_bits_decodeResult_extend;
  reg          shifterReg_2_0_bits_decodeResult_unOrderWrite;
  assign validSink_2_bits_decodeResult_unOrderWrite = shifterReg_2_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_2_0_bits_decodeResult_compress;
  assign validSink_2_bits_decodeResult_compress = shifterReg_2_0_bits_decodeResult_compress;
  reg          shifterReg_2_0_bits_decodeResult_gather16;
  assign validSink_2_bits_decodeResult_gather16 = shifterReg_2_0_bits_decodeResult_gather16;
  reg          shifterReg_2_0_bits_decodeResult_gather;
  assign validSink_2_bits_decodeResult_gather = shifterReg_2_0_bits_decodeResult_gather;
  reg          shifterReg_2_0_bits_decodeResult_slid;
  assign validSink_2_bits_decodeResult_slid = shifterReg_2_0_bits_decodeResult_slid;
  reg          shifterReg_2_0_bits_decodeResult_targetRd;
  assign validSink_2_bits_decodeResult_targetRd = shifterReg_2_0_bits_decodeResult_targetRd;
  reg          shifterReg_2_0_bits_decodeResult_widenReduce;
  assign validSink_2_bits_decodeResult_widenReduce = shifterReg_2_0_bits_decodeResult_widenReduce;
  reg          shifterReg_2_0_bits_decodeResult_red;
  assign validSink_2_bits_decodeResult_red = shifterReg_2_0_bits_decodeResult_red;
  reg          shifterReg_2_0_bits_decodeResult_nr;
  assign validSink_2_bits_decodeResult_nr = shifterReg_2_0_bits_decodeResult_nr;
  reg          shifterReg_2_0_bits_decodeResult_itype;
  assign validSink_2_bits_decodeResult_itype = shifterReg_2_0_bits_decodeResult_itype;
  reg          shifterReg_2_0_bits_decodeResult_unsigned1;
  assign validSink_2_bits_decodeResult_unsigned1 = shifterReg_2_0_bits_decodeResult_unsigned1;
  reg          shifterReg_2_0_bits_decodeResult_unsigned0;
  assign validSink_2_bits_decodeResult_unsigned0 = shifterReg_2_0_bits_decodeResult_unsigned0;
  reg          shifterReg_2_0_bits_decodeResult_other;
  assign validSink_2_bits_decodeResult_other = shifterReg_2_0_bits_decodeResult_other;
  reg          shifterReg_2_0_bits_decodeResult_multiCycle;
  assign validSink_2_bits_decodeResult_multiCycle = shifterReg_2_0_bits_decodeResult_multiCycle;
  reg          shifterReg_2_0_bits_decodeResult_divider;
  assign validSink_2_bits_decodeResult_divider = shifterReg_2_0_bits_decodeResult_divider;
  reg          shifterReg_2_0_bits_decodeResult_multiplier;
  assign validSink_2_bits_decodeResult_multiplier = shifterReg_2_0_bits_decodeResult_multiplier;
  reg          shifterReg_2_0_bits_decodeResult_shift;
  assign validSink_2_bits_decodeResult_shift = shifterReg_2_0_bits_decodeResult_shift;
  reg          shifterReg_2_0_bits_decodeResult_adder;
  assign validSink_2_bits_decodeResult_adder = shifterReg_2_0_bits_decodeResult_adder;
  reg          shifterReg_2_0_bits_decodeResult_logic;
  assign validSink_2_bits_decodeResult_logic = shifterReg_2_0_bits_decodeResult_logic;
  reg          shifterReg_2_0_bits_loadStore;
  assign validSink_2_bits_loadStore = shifterReg_2_0_bits_loadStore;
  reg          shifterReg_2_0_bits_issueInst;
  assign validSink_2_bits_issueInst = shifterReg_2_0_bits_issueInst;
  reg          shifterReg_2_0_bits_store;
  assign validSink_2_bits_store = shifterReg_2_0_bits_store;
  reg          shifterReg_2_0_bits_special;
  assign validSink_2_bits_special = shifterReg_2_0_bits_special;
  reg          shifterReg_2_0_bits_lsWholeReg;
  assign validSink_2_bits_lsWholeReg = shifterReg_2_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_2_0_bits_vs1;
  assign validSink_2_bits_vs1 = shifterReg_2_0_bits_vs1;
  reg  [4:0]   shifterReg_2_0_bits_vs2;
  assign validSink_2_bits_vs2 = shifterReg_2_0_bits_vs2;
  reg  [4:0]   shifterReg_2_0_bits_vd;
  assign validSink_2_bits_vd = shifterReg_2_0_bits_vd;
  reg  [1:0]   shifterReg_2_0_bits_loadStoreEEW;
  assign validSink_2_bits_loadStoreEEW = shifterReg_2_0_bits_loadStoreEEW;
  reg          shifterReg_2_0_bits_mask;
  assign validSink_2_bits_mask = shifterReg_2_0_bits_mask;
  reg  [2:0]   shifterReg_2_0_bits_segment;
  assign validSink_2_bits_segment = shifterReg_2_0_bits_segment;
  reg  [31:0]  shifterReg_2_0_bits_readFromScalar;
  assign validSink_2_bits_readFromScalar = shifterReg_2_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_2_0_bits_csrInterface_vl;
  assign validSink_2_bits_csrInterface_vl = shifterReg_2_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_2_0_bits_csrInterface_vStart;
  assign validSink_2_bits_csrInterface_vStart = shifterReg_2_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_2_0_bits_csrInterface_vlmul;
  assign validSink_2_bits_csrInterface_vlmul = shifterReg_2_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_2_0_bits_csrInterface_vSew;
  assign validSink_2_bits_csrInterface_vSew = shifterReg_2_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_2_0_bits_csrInterface_vxrm;
  assign validSink_2_bits_csrInterface_vxrm = shifterReg_2_0_bits_csrInterface_vxrm;
  reg          shifterReg_2_0_bits_csrInterface_vta;
  assign validSink_2_bits_csrInterface_vta = shifterReg_2_0_bits_csrInterface_vta;
  reg          shifterReg_2_0_bits_csrInterface_vma;
  assign validSink_2_bits_csrInterface_vma = shifterReg_2_0_bits_csrInterface_vma;
  wire         shifterValid_2 = shifterReg_2_0_valid | validSource_2_valid;
  wire         validSink_3_valid;
  wire [2:0]   validSink_3_bits_instructionIndex;
  wire         validSink_3_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_3_bits_decodeResult_topUop;
  wire         validSink_3_bits_decodeResult_popCount;
  wire         validSink_3_bits_decodeResult_ffo;
  wire         validSink_3_bits_decodeResult_average;
  wire         validSink_3_bits_decodeResult_reverse;
  wire         validSink_3_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_3_bits_decodeResult_scheduler;
  wire         validSink_3_bits_decodeResult_sReadVD;
  wire         validSink_3_bits_decodeResult_vtype;
  wire         validSink_3_bits_decodeResult_sWrite;
  wire         validSink_3_bits_decodeResult_crossRead;
  wire         validSink_3_bits_decodeResult_crossWrite;
  wire         validSink_3_bits_decodeResult_maskUnit;
  wire         validSink_3_bits_decodeResult_special;
  wire         validSink_3_bits_decodeResult_saturate;
  wire         validSink_3_bits_decodeResult_vwmacc;
  wire         validSink_3_bits_decodeResult_readOnly;
  wire         validSink_3_bits_decodeResult_maskSource;
  wire         validSink_3_bits_decodeResult_maskDestination;
  wire         validSink_3_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_3_bits_decodeResult_uop;
  wire         validSink_3_bits_decodeResult_iota;
  wire         validSink_3_bits_decodeResult_mv;
  wire         validSink_3_bits_decodeResult_extend;
  wire         validSink_3_bits_decodeResult_unOrderWrite;
  wire         validSink_3_bits_decodeResult_compress;
  wire         validSink_3_bits_decodeResult_gather16;
  wire         validSink_3_bits_decodeResult_gather;
  wire         validSink_3_bits_decodeResult_slid;
  wire         validSink_3_bits_decodeResult_targetRd;
  wire         validSink_3_bits_decodeResult_widenReduce;
  wire         validSink_3_bits_decodeResult_red;
  wire         validSink_3_bits_decodeResult_nr;
  wire         validSink_3_bits_decodeResult_itype;
  wire         validSink_3_bits_decodeResult_unsigned1;
  wire         validSink_3_bits_decodeResult_unsigned0;
  wire         validSink_3_bits_decodeResult_other;
  wire         validSink_3_bits_decodeResult_multiCycle;
  wire         validSink_3_bits_decodeResult_divider;
  wire         validSink_3_bits_decodeResult_multiplier;
  wire         validSink_3_bits_decodeResult_shift;
  wire         validSink_3_bits_decodeResult_adder;
  wire         validSink_3_bits_decodeResult_logic;
  wire         validSink_3_bits_loadStore;
  wire         validSink_3_bits_issueInst;
  wire         validSink_3_bits_store;
  wire         validSink_3_bits_special;
  wire         validSink_3_bits_lsWholeReg;
  wire [4:0]   validSink_3_bits_vs1;
  wire [4:0]   validSink_3_bits_vs2;
  wire [4:0]   validSink_3_bits_vd;
  wire [1:0]   validSink_3_bits_loadStoreEEW;
  wire         validSink_3_bits_mask;
  wire [2:0]   validSink_3_bits_segment;
  wire [31:0]  validSink_3_bits_readFromScalar;
  wire [11:0]  validSink_3_bits_csrInterface_vl;
  wire [11:0]  validSink_3_bits_csrInterface_vStart;
  wire [2:0]   validSink_3_bits_csrInterface_vlmul;
  wire [1:0]   validSink_3_bits_csrInterface_vSew;
  wire [1:0]   validSink_3_bits_csrInterface_vxrm;
  wire         validSink_3_bits_csrInterface_vta;
  wire         validSink_3_bits_csrInterface_vma;
  wire         laneRequestSinkWire_3_valid = queue_3_deq_valid;
  wire [2:0]   laneRequestSinkWire_3_bits_instructionIndex = queue_3_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_3_bits_decodeResult_specialSlot = queue_3_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_3_bits_decodeResult_topUop = queue_3_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_3_bits_decodeResult_popCount = queue_3_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_3_bits_decodeResult_ffo = queue_3_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_3_bits_decodeResult_average = queue_3_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_3_bits_decodeResult_reverse = queue_3_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_3_bits_decodeResult_dontNeedExecuteInLane = queue_3_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_3_bits_decodeResult_scheduler = queue_3_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_3_bits_decodeResult_sReadVD = queue_3_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_3_bits_decodeResult_vtype = queue_3_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_3_bits_decodeResult_sWrite = queue_3_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_3_bits_decodeResult_crossRead = queue_3_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_3_bits_decodeResult_crossWrite = queue_3_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_3_bits_decodeResult_maskUnit = queue_3_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_3_bits_decodeResult_special = queue_3_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_3_bits_decodeResult_saturate = queue_3_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_3_bits_decodeResult_vwmacc = queue_3_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_3_bits_decodeResult_readOnly = queue_3_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_3_bits_decodeResult_maskSource = queue_3_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_3_bits_decodeResult_maskDestination = queue_3_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_3_bits_decodeResult_maskLogic = queue_3_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_3_bits_decodeResult_uop = queue_3_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_3_bits_decodeResult_iota = queue_3_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_3_bits_decodeResult_mv = queue_3_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_3_bits_decodeResult_extend = queue_3_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_3_bits_decodeResult_unOrderWrite = queue_3_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_3_bits_decodeResult_compress = queue_3_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_3_bits_decodeResult_gather16 = queue_3_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_3_bits_decodeResult_gather = queue_3_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_3_bits_decodeResult_slid = queue_3_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_3_bits_decodeResult_targetRd = queue_3_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_3_bits_decodeResult_widenReduce = queue_3_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_3_bits_decodeResult_red = queue_3_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_3_bits_decodeResult_nr = queue_3_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_3_bits_decodeResult_itype = queue_3_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_3_bits_decodeResult_unsigned1 = queue_3_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_3_bits_decodeResult_unsigned0 = queue_3_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_3_bits_decodeResult_other = queue_3_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_3_bits_decodeResult_multiCycle = queue_3_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_3_bits_decodeResult_divider = queue_3_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_3_bits_decodeResult_multiplier = queue_3_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_3_bits_decodeResult_shift = queue_3_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_3_bits_decodeResult_adder = queue_3_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_3_bits_decodeResult_logic = queue_3_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_3_bits_loadStore = queue_3_deq_bits_loadStore;
  wire         laneRequestSinkWire_3_bits_issueInst = queue_3_deq_bits_issueInst;
  wire         laneRequestSinkWire_3_bits_store = queue_3_deq_bits_store;
  wire         laneRequestSinkWire_3_bits_special = queue_3_deq_bits_special;
  wire         laneRequestSinkWire_3_bits_lsWholeReg = queue_3_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_3_bits_vs1 = queue_3_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_3_bits_vs2 = queue_3_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_3_bits_vd = queue_3_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_3_bits_loadStoreEEW = queue_3_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_3_bits_mask = queue_3_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_3_bits_segment = queue_3_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_3_bits_readFromScalar = queue_3_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_3_bits_csrInterface_vl = queue_3_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_3_bits_csrInterface_vStart = queue_3_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_3_bits_csrInterface_vlmul = queue_3_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_3_bits_csrInterface_vSew = queue_3_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_3_bits_csrInterface_vxrm = queue_3_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_3_bits_csrInterface_vta = queue_3_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_3_bits_csrInterface_vma = queue_3_deq_bits_csrInterface_vma;
  wire [1:0]   queue_3_enq_bits_csrInterface_vxrm;
  wire         queue_3_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi_9 = {queue_3_enq_bits_csrInterface_vxrm, queue_3_enq_bits_csrInterface_vta};
  wire         queue_3_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo_9 = {queue_dataIn_lo_hi_9, queue_3_enq_bits_csrInterface_vma};
  wire [2:0]   queue_3_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_3_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo_9 = {queue_3_enq_bits_csrInterface_vlmul, queue_3_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_3_enq_bits_csrInterface_vl;
  wire [11:0]  queue_3_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi_9 = {queue_3_enq_bits_csrInterface_vl, queue_3_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi_9 = {queue_dataIn_hi_hi_9, queue_dataIn_hi_lo_9};
  wire         queue_3_enq_bits_decodeResult_adder;
  wire         queue_3_enq_bits_decodeResult_logic;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo_3 = {queue_3_enq_bits_decodeResult_adder, queue_3_enq_bits_decodeResult_logic};
  wire         queue_3_enq_bits_decodeResult_divider;
  wire         queue_3_enq_bits_decodeResult_multiplier;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi_3 = {queue_3_enq_bits_decodeResult_divider, queue_3_enq_bits_decodeResult_multiplier};
  wire         queue_3_enq_bits_decodeResult_shift;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi_3 = {queue_dataIn_lo_lo_lo_hi_hi_3, queue_3_enq_bits_decodeResult_shift};
  wire [4:0]   queue_dataIn_lo_lo_lo_3 = {queue_dataIn_lo_lo_lo_hi_3, queue_dataIn_lo_lo_lo_lo_3};
  wire         queue_3_enq_bits_decodeResult_unsigned0;
  wire         queue_3_enq_bits_decodeResult_other;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi_3 = {queue_3_enq_bits_decodeResult_unsigned0, queue_3_enq_bits_decodeResult_other};
  wire         queue_3_enq_bits_decodeResult_multiCycle;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo_3 = {queue_dataIn_lo_lo_hi_lo_hi_3, queue_3_enq_bits_decodeResult_multiCycle};
  wire         queue_3_enq_bits_decodeResult_nr;
  wire         queue_3_enq_bits_decodeResult_itype;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi_3 = {queue_3_enq_bits_decodeResult_nr, queue_3_enq_bits_decodeResult_itype};
  wire         queue_3_enq_bits_decodeResult_unsigned1;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi_3 = {queue_dataIn_lo_lo_hi_hi_hi_3, queue_3_enq_bits_decodeResult_unsigned1};
  wire [5:0]   queue_dataIn_lo_lo_hi_6 = {queue_dataIn_lo_lo_hi_hi_3, queue_dataIn_lo_lo_hi_lo_3};
  wire [10:0]  queue_dataIn_lo_lo_6 = {queue_dataIn_lo_lo_hi_6, queue_dataIn_lo_lo_lo_3};
  wire         queue_3_enq_bits_decodeResult_widenReduce;
  wire         queue_3_enq_bits_decodeResult_red;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo_3 = {queue_3_enq_bits_decodeResult_widenReduce, queue_3_enq_bits_decodeResult_red};
  wire         queue_3_enq_bits_decodeResult_gather;
  wire         queue_3_enq_bits_decodeResult_slid;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi_3 = {queue_3_enq_bits_decodeResult_gather, queue_3_enq_bits_decodeResult_slid};
  wire         queue_3_enq_bits_decodeResult_targetRd;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi_3 = {queue_dataIn_lo_hi_lo_hi_hi_3, queue_3_enq_bits_decodeResult_targetRd};
  wire [4:0]   queue_dataIn_lo_hi_lo_6 = {queue_dataIn_lo_hi_lo_hi_3, queue_dataIn_lo_hi_lo_lo_3};
  wire         queue_3_enq_bits_decodeResult_unOrderWrite;
  wire         queue_3_enq_bits_decodeResult_compress;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi_3 = {queue_3_enq_bits_decodeResult_unOrderWrite, queue_3_enq_bits_decodeResult_compress};
  wire         queue_3_enq_bits_decodeResult_gather16;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo_3 = {queue_dataIn_lo_hi_hi_lo_hi_3, queue_3_enq_bits_decodeResult_gather16};
  wire         queue_3_enq_bits_decodeResult_iota;
  wire         queue_3_enq_bits_decodeResult_mv;
  wire [1:0]   queue_dataIn_lo_hi_hi_hi_hi_3 = {queue_3_enq_bits_decodeResult_iota, queue_3_enq_bits_decodeResult_mv};
  wire         queue_3_enq_bits_decodeResult_extend;
  wire [2:0]   queue_dataIn_lo_hi_hi_hi_3 = {queue_dataIn_lo_hi_hi_hi_hi_3, queue_3_enq_bits_decodeResult_extend};
  wire [5:0]   queue_dataIn_lo_hi_hi_6 = {queue_dataIn_lo_hi_hi_hi_3, queue_dataIn_lo_hi_hi_lo_3};
  wire [10:0]  queue_dataIn_lo_hi_10 = {queue_dataIn_lo_hi_hi_6, queue_dataIn_lo_hi_lo_6};
  wire [21:0]  queue_dataIn_lo_10 = {queue_dataIn_lo_hi_10, queue_dataIn_lo_lo_6};
  wire         queue_3_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_3_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_hi_lo_lo_lo_3 = {queue_3_enq_bits_decodeResult_maskLogic, queue_3_enq_bits_decodeResult_uop};
  wire         queue_3_enq_bits_decodeResult_readOnly;
  wire         queue_3_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi_3 = {queue_3_enq_bits_decodeResult_readOnly, queue_3_enq_bits_decodeResult_maskSource};
  wire         queue_3_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi_3 = {queue_dataIn_hi_lo_lo_hi_hi_3, queue_3_enq_bits_decodeResult_maskDestination};
  wire [7:0]   queue_dataIn_hi_lo_lo_6 = {queue_dataIn_hi_lo_lo_hi_3, queue_dataIn_hi_lo_lo_lo_3};
  wire         queue_3_enq_bits_decodeResult_special;
  wire         queue_3_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi_3 = {queue_3_enq_bits_decodeResult_special, queue_3_enq_bits_decodeResult_saturate};
  wire         queue_3_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo_3 = {queue_dataIn_hi_lo_hi_lo_hi_3, queue_3_enq_bits_decodeResult_vwmacc};
  wire         queue_3_enq_bits_decodeResult_crossRead;
  wire         queue_3_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi_3 = {queue_3_enq_bits_decodeResult_crossRead, queue_3_enq_bits_decodeResult_crossWrite};
  wire         queue_3_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi_3 = {queue_dataIn_hi_lo_hi_hi_hi_3, queue_3_enq_bits_decodeResult_maskUnit};
  wire [5:0]   queue_dataIn_hi_lo_hi_6 = {queue_dataIn_hi_lo_hi_hi_3, queue_dataIn_hi_lo_hi_lo_3};
  wire [13:0]  queue_dataIn_hi_lo_10 = {queue_dataIn_hi_lo_hi_6, queue_dataIn_hi_lo_lo_6};
  wire         queue_3_enq_bits_decodeResult_vtype;
  wire         queue_3_enq_bits_decodeResult_sWrite;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo_3 = {queue_3_enq_bits_decodeResult_vtype, queue_3_enq_bits_decodeResult_sWrite};
  wire         queue_3_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_3_enq_bits_decodeResult_scheduler;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi_3 = {queue_3_enq_bits_decodeResult_dontNeedExecuteInLane, queue_3_enq_bits_decodeResult_scheduler};
  wire         queue_3_enq_bits_decodeResult_sReadVD;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi_3 = {queue_dataIn_hi_hi_lo_hi_hi_3, queue_3_enq_bits_decodeResult_sReadVD};
  wire [4:0]   queue_dataIn_hi_hi_lo_6 = {queue_dataIn_hi_hi_lo_hi_3, queue_dataIn_hi_hi_lo_lo_3};
  wire         queue_3_enq_bits_decodeResult_ffo;
  wire         queue_3_enq_bits_decodeResult_average;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi_3 = {queue_3_enq_bits_decodeResult_ffo, queue_3_enq_bits_decodeResult_average};
  wire         queue_3_enq_bits_decodeResult_reverse;
  wire [2:0]   queue_dataIn_hi_hi_hi_lo_3 = {queue_dataIn_hi_hi_hi_lo_hi_3, queue_3_enq_bits_decodeResult_reverse};
  wire         queue_3_enq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_3_enq_bits_decodeResult_topUop;
  wire [5:0]   queue_dataIn_hi_hi_hi_hi_hi_3 = {queue_3_enq_bits_decodeResult_specialSlot, queue_3_enq_bits_decodeResult_topUop};
  wire         queue_3_enq_bits_decodeResult_popCount;
  wire [6:0]   queue_dataIn_hi_hi_hi_hi_3 = {queue_dataIn_hi_hi_hi_hi_hi_3, queue_3_enq_bits_decodeResult_popCount};
  wire [9:0]   queue_dataIn_hi_hi_hi_6 = {queue_dataIn_hi_hi_hi_hi_3, queue_dataIn_hi_hi_hi_lo_3};
  wire [14:0]  queue_dataIn_hi_hi_10 = {queue_dataIn_hi_hi_hi_6, queue_dataIn_hi_hi_lo_6};
  wire [28:0]  queue_dataIn_hi_10 = {queue_dataIn_hi_hi_10, queue_dataIn_hi_lo_10};
  wire [2:0]   queue_3_enq_bits_segment;
  wire [31:0]  queue_3_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_7 = {queue_3_enq_bits_segment, queue_3_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_7 = {queue_dataIn_lo_lo_hi_7, queue_dataIn_hi_9, queue_dataIn_lo_9};
  wire [1:0]   queue_3_enq_bits_loadStoreEEW;
  wire         queue_3_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_7 = {queue_3_enq_bits_loadStoreEEW, queue_3_enq_bits_mask};
  wire [4:0]   queue_3_enq_bits_vs2;
  wire [4:0]   queue_3_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_7 = {queue_3_enq_bits_vs2, queue_3_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_11 = {queue_dataIn_lo_hi_hi_7, queue_dataIn_lo_hi_lo_7};
  wire [80:0]  queue_dataIn_lo_11 = {queue_dataIn_lo_hi_11, queue_dataIn_lo_lo_7};
  wire         queue_3_enq_bits_lsWholeReg;
  wire [4:0]   queue_3_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_7 = {queue_3_enq_bits_lsWholeReg, queue_3_enq_bits_vs1};
  wire         queue_3_enq_bits_store;
  wire         queue_3_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_7 = {queue_3_enq_bits_store, queue_3_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_11 = {queue_dataIn_hi_lo_hi_7, queue_dataIn_hi_lo_lo_7};
  wire         queue_3_enq_bits_loadStore;
  wire         queue_3_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_7 = {queue_3_enq_bits_loadStore, queue_3_enq_bits_issueInst};
  wire [2:0]   queue_3_enq_bits_instructionIndex;
  wire [53:0]  queue_dataIn_hi_hi_hi_7 = {queue_3_enq_bits_instructionIndex, queue_dataIn_hi_10, queue_dataIn_lo_10};
  wire [55:0]  queue_dataIn_hi_hi_11 = {queue_dataIn_hi_hi_hi_7, queue_dataIn_hi_hi_lo_7};
  wire [63:0]  queue_dataIn_hi_11 = {queue_dataIn_hi_hi_11, queue_dataIn_hi_lo_11};
  wire [144:0] queue_dataIn_3 = {queue_dataIn_hi_11, queue_dataIn_lo_11};
  wire         queue_dataOut_3_csrInterface_vma = _queue_fifo_3_data_out[0];
  wire         queue_dataOut_3_csrInterface_vta = _queue_fifo_3_data_out[1];
  wire [1:0]   queue_dataOut_3_csrInterface_vxrm = _queue_fifo_3_data_out[3:2];
  wire [1:0]   queue_dataOut_3_csrInterface_vSew = _queue_fifo_3_data_out[5:4];
  wire [2:0]   queue_dataOut_3_csrInterface_vlmul = _queue_fifo_3_data_out[8:6];
  wire [11:0]  queue_dataOut_3_csrInterface_vStart = _queue_fifo_3_data_out[20:9];
  wire [11:0]  queue_dataOut_3_csrInterface_vl = _queue_fifo_3_data_out[32:21];
  wire [31:0]  queue_dataOut_3_readFromScalar = _queue_fifo_3_data_out[64:33];
  wire [2:0]   queue_dataOut_3_segment = _queue_fifo_3_data_out[67:65];
  wire         queue_dataOut_3_mask = _queue_fifo_3_data_out[68];
  wire [1:0]   queue_dataOut_3_loadStoreEEW = _queue_fifo_3_data_out[70:69];
  wire [4:0]   queue_dataOut_3_vd = _queue_fifo_3_data_out[75:71];
  wire [4:0]   queue_dataOut_3_vs2 = _queue_fifo_3_data_out[80:76];
  wire [4:0]   queue_dataOut_3_vs1 = _queue_fifo_3_data_out[85:81];
  wire         queue_dataOut_3_lsWholeReg = _queue_fifo_3_data_out[86];
  wire         queue_dataOut_3_special = _queue_fifo_3_data_out[87];
  wire         queue_dataOut_3_store = _queue_fifo_3_data_out[88];
  wire         queue_dataOut_3_issueInst = _queue_fifo_3_data_out[89];
  wire         queue_dataOut_3_loadStore = _queue_fifo_3_data_out[90];
  wire         queue_dataOut_3_decodeResult_logic = _queue_fifo_3_data_out[91];
  wire         queue_dataOut_3_decodeResult_adder = _queue_fifo_3_data_out[92];
  wire         queue_dataOut_3_decodeResult_shift = _queue_fifo_3_data_out[93];
  wire         queue_dataOut_3_decodeResult_multiplier = _queue_fifo_3_data_out[94];
  wire         queue_dataOut_3_decodeResult_divider = _queue_fifo_3_data_out[95];
  wire         queue_dataOut_3_decodeResult_multiCycle = _queue_fifo_3_data_out[96];
  wire         queue_dataOut_3_decodeResult_other = _queue_fifo_3_data_out[97];
  wire         queue_dataOut_3_decodeResult_unsigned0 = _queue_fifo_3_data_out[98];
  wire         queue_dataOut_3_decodeResult_unsigned1 = _queue_fifo_3_data_out[99];
  wire         queue_dataOut_3_decodeResult_itype = _queue_fifo_3_data_out[100];
  wire         queue_dataOut_3_decodeResult_nr = _queue_fifo_3_data_out[101];
  wire         queue_dataOut_3_decodeResult_red = _queue_fifo_3_data_out[102];
  wire         queue_dataOut_3_decodeResult_widenReduce = _queue_fifo_3_data_out[103];
  wire         queue_dataOut_3_decodeResult_targetRd = _queue_fifo_3_data_out[104];
  wire         queue_dataOut_3_decodeResult_slid = _queue_fifo_3_data_out[105];
  wire         queue_dataOut_3_decodeResult_gather = _queue_fifo_3_data_out[106];
  wire         queue_dataOut_3_decodeResult_gather16 = _queue_fifo_3_data_out[107];
  wire         queue_dataOut_3_decodeResult_compress = _queue_fifo_3_data_out[108];
  wire         queue_dataOut_3_decodeResult_unOrderWrite = _queue_fifo_3_data_out[109];
  wire         queue_dataOut_3_decodeResult_extend = _queue_fifo_3_data_out[110];
  wire         queue_dataOut_3_decodeResult_mv = _queue_fifo_3_data_out[111];
  wire         queue_dataOut_3_decodeResult_iota = _queue_fifo_3_data_out[112];
  wire [3:0]   queue_dataOut_3_decodeResult_uop = _queue_fifo_3_data_out[116:113];
  wire         queue_dataOut_3_decodeResult_maskLogic = _queue_fifo_3_data_out[117];
  wire         queue_dataOut_3_decodeResult_maskDestination = _queue_fifo_3_data_out[118];
  wire         queue_dataOut_3_decodeResult_maskSource = _queue_fifo_3_data_out[119];
  wire         queue_dataOut_3_decodeResult_readOnly = _queue_fifo_3_data_out[120];
  wire         queue_dataOut_3_decodeResult_vwmacc = _queue_fifo_3_data_out[121];
  wire         queue_dataOut_3_decodeResult_saturate = _queue_fifo_3_data_out[122];
  wire         queue_dataOut_3_decodeResult_special = _queue_fifo_3_data_out[123];
  wire         queue_dataOut_3_decodeResult_maskUnit = _queue_fifo_3_data_out[124];
  wire         queue_dataOut_3_decodeResult_crossWrite = _queue_fifo_3_data_out[125];
  wire         queue_dataOut_3_decodeResult_crossRead = _queue_fifo_3_data_out[126];
  wire         queue_dataOut_3_decodeResult_sWrite = _queue_fifo_3_data_out[127];
  wire         queue_dataOut_3_decodeResult_vtype = _queue_fifo_3_data_out[128];
  wire         queue_dataOut_3_decodeResult_sReadVD = _queue_fifo_3_data_out[129];
  wire         queue_dataOut_3_decodeResult_scheduler = _queue_fifo_3_data_out[130];
  wire         queue_dataOut_3_decodeResult_dontNeedExecuteInLane = _queue_fifo_3_data_out[131];
  wire         queue_dataOut_3_decodeResult_reverse = _queue_fifo_3_data_out[132];
  wire         queue_dataOut_3_decodeResult_average = _queue_fifo_3_data_out[133];
  wire         queue_dataOut_3_decodeResult_ffo = _queue_fifo_3_data_out[134];
  wire         queue_dataOut_3_decodeResult_popCount = _queue_fifo_3_data_out[135];
  wire [4:0]   queue_dataOut_3_decodeResult_topUop = _queue_fifo_3_data_out[140:136];
  wire         queue_dataOut_3_decodeResult_specialSlot = _queue_fifo_3_data_out[141];
  wire [2:0]   queue_dataOut_3_instructionIndex = _queue_fifo_3_data_out[144:142];
  wire         queue_3_enq_ready = ~_queue_fifo_3_full;
  wire         queue_3_enq_valid;
  assign queue_3_deq_valid = ~_queue_fifo_3_empty | queue_3_enq_valid;
  assign queue_3_deq_bits_instructionIndex = _queue_fifo_3_empty ? queue_3_enq_bits_instructionIndex : queue_dataOut_3_instructionIndex;
  assign queue_3_deq_bits_decodeResult_specialSlot = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_specialSlot : queue_dataOut_3_decodeResult_specialSlot;
  assign queue_3_deq_bits_decodeResult_topUop = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_topUop : queue_dataOut_3_decodeResult_topUop;
  assign queue_3_deq_bits_decodeResult_popCount = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_popCount : queue_dataOut_3_decodeResult_popCount;
  assign queue_3_deq_bits_decodeResult_ffo = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_ffo : queue_dataOut_3_decodeResult_ffo;
  assign queue_3_deq_bits_decodeResult_average = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_average : queue_dataOut_3_decodeResult_average;
  assign queue_3_deq_bits_decodeResult_reverse = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_reverse : queue_dataOut_3_decodeResult_reverse;
  assign queue_3_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_3_decodeResult_dontNeedExecuteInLane;
  assign queue_3_deq_bits_decodeResult_scheduler = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_scheduler : queue_dataOut_3_decodeResult_scheduler;
  assign queue_3_deq_bits_decodeResult_sReadVD = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_sReadVD : queue_dataOut_3_decodeResult_sReadVD;
  assign queue_3_deq_bits_decodeResult_vtype = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_vtype : queue_dataOut_3_decodeResult_vtype;
  assign queue_3_deq_bits_decodeResult_sWrite = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_sWrite : queue_dataOut_3_decodeResult_sWrite;
  assign queue_3_deq_bits_decodeResult_crossRead = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_crossRead : queue_dataOut_3_decodeResult_crossRead;
  assign queue_3_deq_bits_decodeResult_crossWrite = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_crossWrite : queue_dataOut_3_decodeResult_crossWrite;
  assign queue_3_deq_bits_decodeResult_maskUnit = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_maskUnit : queue_dataOut_3_decodeResult_maskUnit;
  assign queue_3_deq_bits_decodeResult_special = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_special : queue_dataOut_3_decodeResult_special;
  assign queue_3_deq_bits_decodeResult_saturate = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_saturate : queue_dataOut_3_decodeResult_saturate;
  assign queue_3_deq_bits_decodeResult_vwmacc = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_vwmacc : queue_dataOut_3_decodeResult_vwmacc;
  assign queue_3_deq_bits_decodeResult_readOnly = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_readOnly : queue_dataOut_3_decodeResult_readOnly;
  assign queue_3_deq_bits_decodeResult_maskSource = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_maskSource : queue_dataOut_3_decodeResult_maskSource;
  assign queue_3_deq_bits_decodeResult_maskDestination = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_maskDestination : queue_dataOut_3_decodeResult_maskDestination;
  assign queue_3_deq_bits_decodeResult_maskLogic = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_maskLogic : queue_dataOut_3_decodeResult_maskLogic;
  assign queue_3_deq_bits_decodeResult_uop = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_uop : queue_dataOut_3_decodeResult_uop;
  assign queue_3_deq_bits_decodeResult_iota = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_iota : queue_dataOut_3_decodeResult_iota;
  assign queue_3_deq_bits_decodeResult_mv = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_mv : queue_dataOut_3_decodeResult_mv;
  assign queue_3_deq_bits_decodeResult_extend = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_extend : queue_dataOut_3_decodeResult_extend;
  assign queue_3_deq_bits_decodeResult_unOrderWrite = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_unOrderWrite : queue_dataOut_3_decodeResult_unOrderWrite;
  assign queue_3_deq_bits_decodeResult_compress = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_compress : queue_dataOut_3_decodeResult_compress;
  assign queue_3_deq_bits_decodeResult_gather16 = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_gather16 : queue_dataOut_3_decodeResult_gather16;
  assign queue_3_deq_bits_decodeResult_gather = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_gather : queue_dataOut_3_decodeResult_gather;
  assign queue_3_deq_bits_decodeResult_slid = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_slid : queue_dataOut_3_decodeResult_slid;
  assign queue_3_deq_bits_decodeResult_targetRd = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_targetRd : queue_dataOut_3_decodeResult_targetRd;
  assign queue_3_deq_bits_decodeResult_widenReduce = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_widenReduce : queue_dataOut_3_decodeResult_widenReduce;
  assign queue_3_deq_bits_decodeResult_red = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_red : queue_dataOut_3_decodeResult_red;
  assign queue_3_deq_bits_decodeResult_nr = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_nr : queue_dataOut_3_decodeResult_nr;
  assign queue_3_deq_bits_decodeResult_itype = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_itype : queue_dataOut_3_decodeResult_itype;
  assign queue_3_deq_bits_decodeResult_unsigned1 = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_unsigned1 : queue_dataOut_3_decodeResult_unsigned1;
  assign queue_3_deq_bits_decodeResult_unsigned0 = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_unsigned0 : queue_dataOut_3_decodeResult_unsigned0;
  assign queue_3_deq_bits_decodeResult_other = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_other : queue_dataOut_3_decodeResult_other;
  assign queue_3_deq_bits_decodeResult_multiCycle = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_multiCycle : queue_dataOut_3_decodeResult_multiCycle;
  assign queue_3_deq_bits_decodeResult_divider = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_divider : queue_dataOut_3_decodeResult_divider;
  assign queue_3_deq_bits_decodeResult_multiplier = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_multiplier : queue_dataOut_3_decodeResult_multiplier;
  assign queue_3_deq_bits_decodeResult_shift = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_shift : queue_dataOut_3_decodeResult_shift;
  assign queue_3_deq_bits_decodeResult_adder = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_adder : queue_dataOut_3_decodeResult_adder;
  assign queue_3_deq_bits_decodeResult_logic = _queue_fifo_3_empty ? queue_3_enq_bits_decodeResult_logic : queue_dataOut_3_decodeResult_logic;
  assign queue_3_deq_bits_loadStore = _queue_fifo_3_empty ? queue_3_enq_bits_loadStore : queue_dataOut_3_loadStore;
  assign queue_3_deq_bits_issueInst = _queue_fifo_3_empty ? queue_3_enq_bits_issueInst : queue_dataOut_3_issueInst;
  assign queue_3_deq_bits_store = _queue_fifo_3_empty ? queue_3_enq_bits_store : queue_dataOut_3_store;
  assign queue_3_deq_bits_special = _queue_fifo_3_empty ? queue_3_enq_bits_special : queue_dataOut_3_special;
  assign queue_3_deq_bits_lsWholeReg = _queue_fifo_3_empty ? queue_3_enq_bits_lsWholeReg : queue_dataOut_3_lsWholeReg;
  assign queue_3_deq_bits_vs1 = _queue_fifo_3_empty ? queue_3_enq_bits_vs1 : queue_dataOut_3_vs1;
  assign queue_3_deq_bits_vs2 = _queue_fifo_3_empty ? queue_3_enq_bits_vs2 : queue_dataOut_3_vs2;
  assign queue_3_deq_bits_vd = _queue_fifo_3_empty ? queue_3_enq_bits_vd : queue_dataOut_3_vd;
  assign queue_3_deq_bits_loadStoreEEW = _queue_fifo_3_empty ? queue_3_enq_bits_loadStoreEEW : queue_dataOut_3_loadStoreEEW;
  assign queue_3_deq_bits_mask = _queue_fifo_3_empty ? queue_3_enq_bits_mask : queue_dataOut_3_mask;
  assign queue_3_deq_bits_segment = _queue_fifo_3_empty ? queue_3_enq_bits_segment : queue_dataOut_3_segment;
  assign queue_3_deq_bits_readFromScalar = _queue_fifo_3_empty ? queue_3_enq_bits_readFromScalar : queue_dataOut_3_readFromScalar;
  assign queue_3_deq_bits_csrInterface_vl = _queue_fifo_3_empty ? queue_3_enq_bits_csrInterface_vl : queue_dataOut_3_csrInterface_vl;
  assign queue_3_deq_bits_csrInterface_vStart = _queue_fifo_3_empty ? queue_3_enq_bits_csrInterface_vStart : queue_dataOut_3_csrInterface_vStart;
  assign queue_3_deq_bits_csrInterface_vlmul = _queue_fifo_3_empty ? queue_3_enq_bits_csrInterface_vlmul : queue_dataOut_3_csrInterface_vlmul;
  assign queue_3_deq_bits_csrInterface_vSew = _queue_fifo_3_empty ? queue_3_enq_bits_csrInterface_vSew : queue_dataOut_3_csrInterface_vSew;
  assign queue_3_deq_bits_csrInterface_vxrm = _queue_fifo_3_empty ? queue_3_enq_bits_csrInterface_vxrm : queue_dataOut_3_csrInterface_vxrm;
  assign queue_3_deq_bits_csrInterface_vta = _queue_fifo_3_empty ? queue_3_enq_bits_csrInterface_vta : queue_dataOut_3_csrInterface_vta;
  assign queue_3_deq_bits_csrInterface_vma = _queue_fifo_3_empty ? queue_3_enq_bits_csrInterface_vma : queue_dataOut_3_csrInterface_vma;
  wire         laneVec_3_laneRequest_bits_issueInst = laneRequestSinkWire_3_ready & laneRequestSinkWire_3_valid;
  reg          releasePipe_pipe_v_3;
  wire         releasePipe_pipe_out_3_valid = releasePipe_pipe_v_3;
  wire         laneRequestSourceWire_3_ready;
  wire         validSource_3_valid = laneRequestSourceWire_3_ready & laneRequestSourceWire_3_valid;
  reg  [2:0]   tokenCheck_counter_3;
  wire [2:0]   tokenCheck_counterChange_3 = validSource_3_valid ? 3'h1 : 3'h7;
  assign tokenCheck_3 = ~(tokenCheck_counter_3[2]);
  assign laneRequestSourceWire_3_ready = tokenCheck_3;
  assign queue_3_enq_valid = validSink_3_valid;
  assign queue_3_enq_bits_instructionIndex = validSink_3_bits_instructionIndex;
  assign queue_3_enq_bits_decodeResult_specialSlot = validSink_3_bits_decodeResult_specialSlot;
  assign queue_3_enq_bits_decodeResult_topUop = validSink_3_bits_decodeResult_topUop;
  assign queue_3_enq_bits_decodeResult_popCount = validSink_3_bits_decodeResult_popCount;
  assign queue_3_enq_bits_decodeResult_ffo = validSink_3_bits_decodeResult_ffo;
  assign queue_3_enq_bits_decodeResult_average = validSink_3_bits_decodeResult_average;
  assign queue_3_enq_bits_decodeResult_reverse = validSink_3_bits_decodeResult_reverse;
  assign queue_3_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_3_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_3_enq_bits_decodeResult_scheduler = validSink_3_bits_decodeResult_scheduler;
  assign queue_3_enq_bits_decodeResult_sReadVD = validSink_3_bits_decodeResult_sReadVD;
  assign queue_3_enq_bits_decodeResult_vtype = validSink_3_bits_decodeResult_vtype;
  assign queue_3_enq_bits_decodeResult_sWrite = validSink_3_bits_decodeResult_sWrite;
  assign queue_3_enq_bits_decodeResult_crossRead = validSink_3_bits_decodeResult_crossRead;
  assign queue_3_enq_bits_decodeResult_crossWrite = validSink_3_bits_decodeResult_crossWrite;
  assign queue_3_enq_bits_decodeResult_maskUnit = validSink_3_bits_decodeResult_maskUnit;
  assign queue_3_enq_bits_decodeResult_special = validSink_3_bits_decodeResult_special;
  assign queue_3_enq_bits_decodeResult_saturate = validSink_3_bits_decodeResult_saturate;
  assign queue_3_enq_bits_decodeResult_vwmacc = validSink_3_bits_decodeResult_vwmacc;
  assign queue_3_enq_bits_decodeResult_readOnly = validSink_3_bits_decodeResult_readOnly;
  assign queue_3_enq_bits_decodeResult_maskSource = validSink_3_bits_decodeResult_maskSource;
  assign queue_3_enq_bits_decodeResult_maskDestination = validSink_3_bits_decodeResult_maskDestination;
  assign queue_3_enq_bits_decodeResult_maskLogic = validSink_3_bits_decodeResult_maskLogic;
  assign queue_3_enq_bits_decodeResult_uop = validSink_3_bits_decodeResult_uop;
  assign queue_3_enq_bits_decodeResult_iota = validSink_3_bits_decodeResult_iota;
  assign queue_3_enq_bits_decodeResult_mv = validSink_3_bits_decodeResult_mv;
  assign queue_3_enq_bits_decodeResult_extend = validSink_3_bits_decodeResult_extend;
  assign queue_3_enq_bits_decodeResult_unOrderWrite = validSink_3_bits_decodeResult_unOrderWrite;
  assign queue_3_enq_bits_decodeResult_compress = validSink_3_bits_decodeResult_compress;
  assign queue_3_enq_bits_decodeResult_gather16 = validSink_3_bits_decodeResult_gather16;
  assign queue_3_enq_bits_decodeResult_gather = validSink_3_bits_decodeResult_gather;
  assign queue_3_enq_bits_decodeResult_slid = validSink_3_bits_decodeResult_slid;
  assign queue_3_enq_bits_decodeResult_targetRd = validSink_3_bits_decodeResult_targetRd;
  assign queue_3_enq_bits_decodeResult_widenReduce = validSink_3_bits_decodeResult_widenReduce;
  assign queue_3_enq_bits_decodeResult_red = validSink_3_bits_decodeResult_red;
  assign queue_3_enq_bits_decodeResult_nr = validSink_3_bits_decodeResult_nr;
  assign queue_3_enq_bits_decodeResult_itype = validSink_3_bits_decodeResult_itype;
  assign queue_3_enq_bits_decodeResult_unsigned1 = validSink_3_bits_decodeResult_unsigned1;
  assign queue_3_enq_bits_decodeResult_unsigned0 = validSink_3_bits_decodeResult_unsigned0;
  assign queue_3_enq_bits_decodeResult_other = validSink_3_bits_decodeResult_other;
  assign queue_3_enq_bits_decodeResult_multiCycle = validSink_3_bits_decodeResult_multiCycle;
  assign queue_3_enq_bits_decodeResult_divider = validSink_3_bits_decodeResult_divider;
  assign queue_3_enq_bits_decodeResult_multiplier = validSink_3_bits_decodeResult_multiplier;
  assign queue_3_enq_bits_decodeResult_shift = validSink_3_bits_decodeResult_shift;
  assign queue_3_enq_bits_decodeResult_adder = validSink_3_bits_decodeResult_adder;
  assign queue_3_enq_bits_decodeResult_logic = validSink_3_bits_decodeResult_logic;
  assign queue_3_enq_bits_loadStore = validSink_3_bits_loadStore;
  assign queue_3_enq_bits_issueInst = validSink_3_bits_issueInst;
  assign queue_3_enq_bits_store = validSink_3_bits_store;
  assign queue_3_enq_bits_special = validSink_3_bits_special;
  assign queue_3_enq_bits_lsWholeReg = validSink_3_bits_lsWholeReg;
  assign queue_3_enq_bits_vs1 = validSink_3_bits_vs1;
  assign queue_3_enq_bits_vs2 = validSink_3_bits_vs2;
  assign queue_3_enq_bits_vd = validSink_3_bits_vd;
  assign queue_3_enq_bits_loadStoreEEW = validSink_3_bits_loadStoreEEW;
  assign queue_3_enq_bits_mask = validSink_3_bits_mask;
  assign queue_3_enq_bits_segment = validSink_3_bits_segment;
  assign queue_3_enq_bits_readFromScalar = validSink_3_bits_readFromScalar;
  assign queue_3_enq_bits_csrInterface_vl = validSink_3_bits_csrInterface_vl;
  assign queue_3_enq_bits_csrInterface_vStart = validSink_3_bits_csrInterface_vStart;
  assign queue_3_enq_bits_csrInterface_vlmul = validSink_3_bits_csrInterface_vlmul;
  assign queue_3_enq_bits_csrInterface_vSew = validSink_3_bits_csrInterface_vSew;
  assign queue_3_enq_bits_csrInterface_vxrm = validSink_3_bits_csrInterface_vxrm;
  assign queue_3_enq_bits_csrInterface_vta = validSink_3_bits_csrInterface_vta;
  assign queue_3_enq_bits_csrInterface_vma = validSink_3_bits_csrInterface_vma;
  reg          shifterReg_3_0_valid;
  assign validSink_3_valid = shifterReg_3_0_valid;
  reg  [2:0]   shifterReg_3_0_bits_instructionIndex;
  assign validSink_3_bits_instructionIndex = shifterReg_3_0_bits_instructionIndex;
  reg          shifterReg_3_0_bits_decodeResult_specialSlot;
  assign validSink_3_bits_decodeResult_specialSlot = shifterReg_3_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_3_0_bits_decodeResult_topUop;
  assign validSink_3_bits_decodeResult_topUop = shifterReg_3_0_bits_decodeResult_topUop;
  reg          shifterReg_3_0_bits_decodeResult_popCount;
  assign validSink_3_bits_decodeResult_popCount = shifterReg_3_0_bits_decodeResult_popCount;
  reg          shifterReg_3_0_bits_decodeResult_ffo;
  assign validSink_3_bits_decodeResult_ffo = shifterReg_3_0_bits_decodeResult_ffo;
  reg          shifterReg_3_0_bits_decodeResult_average;
  assign validSink_3_bits_decodeResult_average = shifterReg_3_0_bits_decodeResult_average;
  reg          shifterReg_3_0_bits_decodeResult_reverse;
  assign validSink_3_bits_decodeResult_reverse = shifterReg_3_0_bits_decodeResult_reverse;
  reg          shifterReg_3_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_3_bits_decodeResult_dontNeedExecuteInLane = shifterReg_3_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_3_0_bits_decodeResult_scheduler;
  assign validSink_3_bits_decodeResult_scheduler = shifterReg_3_0_bits_decodeResult_scheduler;
  reg          shifterReg_3_0_bits_decodeResult_sReadVD;
  assign validSink_3_bits_decodeResult_sReadVD = shifterReg_3_0_bits_decodeResult_sReadVD;
  reg          shifterReg_3_0_bits_decodeResult_vtype;
  assign validSink_3_bits_decodeResult_vtype = shifterReg_3_0_bits_decodeResult_vtype;
  reg          shifterReg_3_0_bits_decodeResult_sWrite;
  assign validSink_3_bits_decodeResult_sWrite = shifterReg_3_0_bits_decodeResult_sWrite;
  reg          shifterReg_3_0_bits_decodeResult_crossRead;
  assign validSink_3_bits_decodeResult_crossRead = shifterReg_3_0_bits_decodeResult_crossRead;
  reg          shifterReg_3_0_bits_decodeResult_crossWrite;
  assign validSink_3_bits_decodeResult_crossWrite = shifterReg_3_0_bits_decodeResult_crossWrite;
  reg          shifterReg_3_0_bits_decodeResult_maskUnit;
  assign validSink_3_bits_decodeResult_maskUnit = shifterReg_3_0_bits_decodeResult_maskUnit;
  reg          shifterReg_3_0_bits_decodeResult_special;
  assign validSink_3_bits_decodeResult_special = shifterReg_3_0_bits_decodeResult_special;
  reg          shifterReg_3_0_bits_decodeResult_saturate;
  assign validSink_3_bits_decodeResult_saturate = shifterReg_3_0_bits_decodeResult_saturate;
  reg          shifterReg_3_0_bits_decodeResult_vwmacc;
  assign validSink_3_bits_decodeResult_vwmacc = shifterReg_3_0_bits_decodeResult_vwmacc;
  reg          shifterReg_3_0_bits_decodeResult_readOnly;
  assign validSink_3_bits_decodeResult_readOnly = shifterReg_3_0_bits_decodeResult_readOnly;
  reg          shifterReg_3_0_bits_decodeResult_maskSource;
  assign validSink_3_bits_decodeResult_maskSource = shifterReg_3_0_bits_decodeResult_maskSource;
  reg          shifterReg_3_0_bits_decodeResult_maskDestination;
  assign validSink_3_bits_decodeResult_maskDestination = shifterReg_3_0_bits_decodeResult_maskDestination;
  reg          shifterReg_3_0_bits_decodeResult_maskLogic;
  assign validSink_3_bits_decodeResult_maskLogic = shifterReg_3_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_3_0_bits_decodeResult_uop;
  assign validSink_3_bits_decodeResult_uop = shifterReg_3_0_bits_decodeResult_uop;
  reg          shifterReg_3_0_bits_decodeResult_iota;
  assign validSink_3_bits_decodeResult_iota = shifterReg_3_0_bits_decodeResult_iota;
  reg          shifterReg_3_0_bits_decodeResult_mv;
  assign validSink_3_bits_decodeResult_mv = shifterReg_3_0_bits_decodeResult_mv;
  reg          shifterReg_3_0_bits_decodeResult_extend;
  assign validSink_3_bits_decodeResult_extend = shifterReg_3_0_bits_decodeResult_extend;
  reg          shifterReg_3_0_bits_decodeResult_unOrderWrite;
  assign validSink_3_bits_decodeResult_unOrderWrite = shifterReg_3_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_3_0_bits_decodeResult_compress;
  assign validSink_3_bits_decodeResult_compress = shifterReg_3_0_bits_decodeResult_compress;
  reg          shifterReg_3_0_bits_decodeResult_gather16;
  assign validSink_3_bits_decodeResult_gather16 = shifterReg_3_0_bits_decodeResult_gather16;
  reg          shifterReg_3_0_bits_decodeResult_gather;
  assign validSink_3_bits_decodeResult_gather = shifterReg_3_0_bits_decodeResult_gather;
  reg          shifterReg_3_0_bits_decodeResult_slid;
  assign validSink_3_bits_decodeResult_slid = shifterReg_3_0_bits_decodeResult_slid;
  reg          shifterReg_3_0_bits_decodeResult_targetRd;
  assign validSink_3_bits_decodeResult_targetRd = shifterReg_3_0_bits_decodeResult_targetRd;
  reg          shifterReg_3_0_bits_decodeResult_widenReduce;
  assign validSink_3_bits_decodeResult_widenReduce = shifterReg_3_0_bits_decodeResult_widenReduce;
  reg          shifterReg_3_0_bits_decodeResult_red;
  assign validSink_3_bits_decodeResult_red = shifterReg_3_0_bits_decodeResult_red;
  reg          shifterReg_3_0_bits_decodeResult_nr;
  assign validSink_3_bits_decodeResult_nr = shifterReg_3_0_bits_decodeResult_nr;
  reg          shifterReg_3_0_bits_decodeResult_itype;
  assign validSink_3_bits_decodeResult_itype = shifterReg_3_0_bits_decodeResult_itype;
  reg          shifterReg_3_0_bits_decodeResult_unsigned1;
  assign validSink_3_bits_decodeResult_unsigned1 = shifterReg_3_0_bits_decodeResult_unsigned1;
  reg          shifterReg_3_0_bits_decodeResult_unsigned0;
  assign validSink_3_bits_decodeResult_unsigned0 = shifterReg_3_0_bits_decodeResult_unsigned0;
  reg          shifterReg_3_0_bits_decodeResult_other;
  assign validSink_3_bits_decodeResult_other = shifterReg_3_0_bits_decodeResult_other;
  reg          shifterReg_3_0_bits_decodeResult_multiCycle;
  assign validSink_3_bits_decodeResult_multiCycle = shifterReg_3_0_bits_decodeResult_multiCycle;
  reg          shifterReg_3_0_bits_decodeResult_divider;
  assign validSink_3_bits_decodeResult_divider = shifterReg_3_0_bits_decodeResult_divider;
  reg          shifterReg_3_0_bits_decodeResult_multiplier;
  assign validSink_3_bits_decodeResult_multiplier = shifterReg_3_0_bits_decodeResult_multiplier;
  reg          shifterReg_3_0_bits_decodeResult_shift;
  assign validSink_3_bits_decodeResult_shift = shifterReg_3_0_bits_decodeResult_shift;
  reg          shifterReg_3_0_bits_decodeResult_adder;
  assign validSink_3_bits_decodeResult_adder = shifterReg_3_0_bits_decodeResult_adder;
  reg          shifterReg_3_0_bits_decodeResult_logic;
  assign validSink_3_bits_decodeResult_logic = shifterReg_3_0_bits_decodeResult_logic;
  reg          shifterReg_3_0_bits_loadStore;
  assign validSink_3_bits_loadStore = shifterReg_3_0_bits_loadStore;
  reg          shifterReg_3_0_bits_issueInst;
  assign validSink_3_bits_issueInst = shifterReg_3_0_bits_issueInst;
  reg          shifterReg_3_0_bits_store;
  assign validSink_3_bits_store = shifterReg_3_0_bits_store;
  reg          shifterReg_3_0_bits_special;
  assign validSink_3_bits_special = shifterReg_3_0_bits_special;
  reg          shifterReg_3_0_bits_lsWholeReg;
  assign validSink_3_bits_lsWholeReg = shifterReg_3_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_3_0_bits_vs1;
  assign validSink_3_bits_vs1 = shifterReg_3_0_bits_vs1;
  reg  [4:0]   shifterReg_3_0_bits_vs2;
  assign validSink_3_bits_vs2 = shifterReg_3_0_bits_vs2;
  reg  [4:0]   shifterReg_3_0_bits_vd;
  assign validSink_3_bits_vd = shifterReg_3_0_bits_vd;
  reg  [1:0]   shifterReg_3_0_bits_loadStoreEEW;
  assign validSink_3_bits_loadStoreEEW = shifterReg_3_0_bits_loadStoreEEW;
  reg          shifterReg_3_0_bits_mask;
  assign validSink_3_bits_mask = shifterReg_3_0_bits_mask;
  reg  [2:0]   shifterReg_3_0_bits_segment;
  assign validSink_3_bits_segment = shifterReg_3_0_bits_segment;
  reg  [31:0]  shifterReg_3_0_bits_readFromScalar;
  assign validSink_3_bits_readFromScalar = shifterReg_3_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_3_0_bits_csrInterface_vl;
  assign validSink_3_bits_csrInterface_vl = shifterReg_3_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_3_0_bits_csrInterface_vStart;
  assign validSink_3_bits_csrInterface_vStart = shifterReg_3_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_3_0_bits_csrInterface_vlmul;
  assign validSink_3_bits_csrInterface_vlmul = shifterReg_3_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_3_0_bits_csrInterface_vSew;
  assign validSink_3_bits_csrInterface_vSew = shifterReg_3_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_3_0_bits_csrInterface_vxrm;
  assign validSink_3_bits_csrInterface_vxrm = shifterReg_3_0_bits_csrInterface_vxrm;
  reg          shifterReg_3_0_bits_csrInterface_vta;
  assign validSink_3_bits_csrInterface_vta = shifterReg_3_0_bits_csrInterface_vta;
  reg          shifterReg_3_0_bits_csrInterface_vma;
  assign validSink_3_bits_csrInterface_vma = shifterReg_3_0_bits_csrInterface_vma;
  wire         shifterValid_3 = shifterReg_3_0_valid | validSource_3_valid;
  wire         validSink_4_valid;
  wire [2:0]   validSink_4_bits_instructionIndex;
  wire         validSink_4_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_4_bits_decodeResult_topUop;
  wire         validSink_4_bits_decodeResult_popCount;
  wire         validSink_4_bits_decodeResult_ffo;
  wire         validSink_4_bits_decodeResult_average;
  wire         validSink_4_bits_decodeResult_reverse;
  wire         validSink_4_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_4_bits_decodeResult_scheduler;
  wire         validSink_4_bits_decodeResult_sReadVD;
  wire         validSink_4_bits_decodeResult_vtype;
  wire         validSink_4_bits_decodeResult_sWrite;
  wire         validSink_4_bits_decodeResult_crossRead;
  wire         validSink_4_bits_decodeResult_crossWrite;
  wire         validSink_4_bits_decodeResult_maskUnit;
  wire         validSink_4_bits_decodeResult_special;
  wire         validSink_4_bits_decodeResult_saturate;
  wire         validSink_4_bits_decodeResult_vwmacc;
  wire         validSink_4_bits_decodeResult_readOnly;
  wire         validSink_4_bits_decodeResult_maskSource;
  wire         validSink_4_bits_decodeResult_maskDestination;
  wire         validSink_4_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_4_bits_decodeResult_uop;
  wire         validSink_4_bits_decodeResult_iota;
  wire         validSink_4_bits_decodeResult_mv;
  wire         validSink_4_bits_decodeResult_extend;
  wire         validSink_4_bits_decodeResult_unOrderWrite;
  wire         validSink_4_bits_decodeResult_compress;
  wire         validSink_4_bits_decodeResult_gather16;
  wire         validSink_4_bits_decodeResult_gather;
  wire         validSink_4_bits_decodeResult_slid;
  wire         validSink_4_bits_decodeResult_targetRd;
  wire         validSink_4_bits_decodeResult_widenReduce;
  wire         validSink_4_bits_decodeResult_red;
  wire         validSink_4_bits_decodeResult_nr;
  wire         validSink_4_bits_decodeResult_itype;
  wire         validSink_4_bits_decodeResult_unsigned1;
  wire         validSink_4_bits_decodeResult_unsigned0;
  wire         validSink_4_bits_decodeResult_other;
  wire         validSink_4_bits_decodeResult_multiCycle;
  wire         validSink_4_bits_decodeResult_divider;
  wire         validSink_4_bits_decodeResult_multiplier;
  wire         validSink_4_bits_decodeResult_shift;
  wire         validSink_4_bits_decodeResult_adder;
  wire         validSink_4_bits_decodeResult_logic;
  wire         validSink_4_bits_loadStore;
  wire         validSink_4_bits_issueInst;
  wire         validSink_4_bits_store;
  wire         validSink_4_bits_special;
  wire         validSink_4_bits_lsWholeReg;
  wire [4:0]   validSink_4_bits_vs1;
  wire [4:0]   validSink_4_bits_vs2;
  wire [4:0]   validSink_4_bits_vd;
  wire [1:0]   validSink_4_bits_loadStoreEEW;
  wire         validSink_4_bits_mask;
  wire [2:0]   validSink_4_bits_segment;
  wire [31:0]  validSink_4_bits_readFromScalar;
  wire [11:0]  validSink_4_bits_csrInterface_vl;
  wire [11:0]  validSink_4_bits_csrInterface_vStart;
  wire [2:0]   validSink_4_bits_csrInterface_vlmul;
  wire [1:0]   validSink_4_bits_csrInterface_vSew;
  wire [1:0]   validSink_4_bits_csrInterface_vxrm;
  wire         validSink_4_bits_csrInterface_vta;
  wire         validSink_4_bits_csrInterface_vma;
  wire         laneRequestSinkWire_4_valid = queue_4_deq_valid;
  wire [2:0]   laneRequestSinkWire_4_bits_instructionIndex = queue_4_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_4_bits_decodeResult_specialSlot = queue_4_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_4_bits_decodeResult_topUop = queue_4_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_4_bits_decodeResult_popCount = queue_4_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_4_bits_decodeResult_ffo = queue_4_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_4_bits_decodeResult_average = queue_4_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_4_bits_decodeResult_reverse = queue_4_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_4_bits_decodeResult_dontNeedExecuteInLane = queue_4_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_4_bits_decodeResult_scheduler = queue_4_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_4_bits_decodeResult_sReadVD = queue_4_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_4_bits_decodeResult_vtype = queue_4_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_4_bits_decodeResult_sWrite = queue_4_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_4_bits_decodeResult_crossRead = queue_4_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_4_bits_decodeResult_crossWrite = queue_4_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_4_bits_decodeResult_maskUnit = queue_4_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_4_bits_decodeResult_special = queue_4_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_4_bits_decodeResult_saturate = queue_4_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_4_bits_decodeResult_vwmacc = queue_4_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_4_bits_decodeResult_readOnly = queue_4_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_4_bits_decodeResult_maskSource = queue_4_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_4_bits_decodeResult_maskDestination = queue_4_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_4_bits_decodeResult_maskLogic = queue_4_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_4_bits_decodeResult_uop = queue_4_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_4_bits_decodeResult_iota = queue_4_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_4_bits_decodeResult_mv = queue_4_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_4_bits_decodeResult_extend = queue_4_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_4_bits_decodeResult_unOrderWrite = queue_4_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_4_bits_decodeResult_compress = queue_4_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_4_bits_decodeResult_gather16 = queue_4_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_4_bits_decodeResult_gather = queue_4_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_4_bits_decodeResult_slid = queue_4_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_4_bits_decodeResult_targetRd = queue_4_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_4_bits_decodeResult_widenReduce = queue_4_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_4_bits_decodeResult_red = queue_4_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_4_bits_decodeResult_nr = queue_4_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_4_bits_decodeResult_itype = queue_4_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_4_bits_decodeResult_unsigned1 = queue_4_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_4_bits_decodeResult_unsigned0 = queue_4_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_4_bits_decodeResult_other = queue_4_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_4_bits_decodeResult_multiCycle = queue_4_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_4_bits_decodeResult_divider = queue_4_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_4_bits_decodeResult_multiplier = queue_4_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_4_bits_decodeResult_shift = queue_4_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_4_bits_decodeResult_adder = queue_4_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_4_bits_decodeResult_logic = queue_4_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_4_bits_loadStore = queue_4_deq_bits_loadStore;
  wire         laneRequestSinkWire_4_bits_issueInst = queue_4_deq_bits_issueInst;
  wire         laneRequestSinkWire_4_bits_store = queue_4_deq_bits_store;
  wire         laneRequestSinkWire_4_bits_special = queue_4_deq_bits_special;
  wire         laneRequestSinkWire_4_bits_lsWholeReg = queue_4_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_4_bits_vs1 = queue_4_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_4_bits_vs2 = queue_4_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_4_bits_vd = queue_4_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_4_bits_loadStoreEEW = queue_4_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_4_bits_mask = queue_4_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_4_bits_segment = queue_4_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_4_bits_readFromScalar = queue_4_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_4_bits_csrInterface_vl = queue_4_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_4_bits_csrInterface_vStart = queue_4_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_4_bits_csrInterface_vlmul = queue_4_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_4_bits_csrInterface_vSew = queue_4_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_4_bits_csrInterface_vxrm = queue_4_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_4_bits_csrInterface_vta = queue_4_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_4_bits_csrInterface_vma = queue_4_deq_bits_csrInterface_vma;
  wire [1:0]   queue_4_enq_bits_csrInterface_vxrm;
  wire         queue_4_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi_12 = {queue_4_enq_bits_csrInterface_vxrm, queue_4_enq_bits_csrInterface_vta};
  wire         queue_4_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo_12 = {queue_dataIn_lo_hi_12, queue_4_enq_bits_csrInterface_vma};
  wire [2:0]   queue_4_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_4_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo_12 = {queue_4_enq_bits_csrInterface_vlmul, queue_4_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_4_enq_bits_csrInterface_vl;
  wire [11:0]  queue_4_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi_12 = {queue_4_enq_bits_csrInterface_vl, queue_4_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi_12 = {queue_dataIn_hi_hi_12, queue_dataIn_hi_lo_12};
  wire         queue_4_enq_bits_decodeResult_adder;
  wire         queue_4_enq_bits_decodeResult_logic;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo_4 = {queue_4_enq_bits_decodeResult_adder, queue_4_enq_bits_decodeResult_logic};
  wire         queue_4_enq_bits_decodeResult_divider;
  wire         queue_4_enq_bits_decodeResult_multiplier;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi_4 = {queue_4_enq_bits_decodeResult_divider, queue_4_enq_bits_decodeResult_multiplier};
  wire         queue_4_enq_bits_decodeResult_shift;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi_4 = {queue_dataIn_lo_lo_lo_hi_hi_4, queue_4_enq_bits_decodeResult_shift};
  wire [4:0]   queue_dataIn_lo_lo_lo_4 = {queue_dataIn_lo_lo_lo_hi_4, queue_dataIn_lo_lo_lo_lo_4};
  wire         queue_4_enq_bits_decodeResult_unsigned0;
  wire         queue_4_enq_bits_decodeResult_other;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi_4 = {queue_4_enq_bits_decodeResult_unsigned0, queue_4_enq_bits_decodeResult_other};
  wire         queue_4_enq_bits_decodeResult_multiCycle;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo_4 = {queue_dataIn_lo_lo_hi_lo_hi_4, queue_4_enq_bits_decodeResult_multiCycle};
  wire         queue_4_enq_bits_decodeResult_nr;
  wire         queue_4_enq_bits_decodeResult_itype;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi_4 = {queue_4_enq_bits_decodeResult_nr, queue_4_enq_bits_decodeResult_itype};
  wire         queue_4_enq_bits_decodeResult_unsigned1;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi_4 = {queue_dataIn_lo_lo_hi_hi_hi_4, queue_4_enq_bits_decodeResult_unsigned1};
  wire [5:0]   queue_dataIn_lo_lo_hi_8 = {queue_dataIn_lo_lo_hi_hi_4, queue_dataIn_lo_lo_hi_lo_4};
  wire [10:0]  queue_dataIn_lo_lo_8 = {queue_dataIn_lo_lo_hi_8, queue_dataIn_lo_lo_lo_4};
  wire         queue_4_enq_bits_decodeResult_widenReduce;
  wire         queue_4_enq_bits_decodeResult_red;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo_4 = {queue_4_enq_bits_decodeResult_widenReduce, queue_4_enq_bits_decodeResult_red};
  wire         queue_4_enq_bits_decodeResult_gather;
  wire         queue_4_enq_bits_decodeResult_slid;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi_4 = {queue_4_enq_bits_decodeResult_gather, queue_4_enq_bits_decodeResult_slid};
  wire         queue_4_enq_bits_decodeResult_targetRd;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi_4 = {queue_dataIn_lo_hi_lo_hi_hi_4, queue_4_enq_bits_decodeResult_targetRd};
  wire [4:0]   queue_dataIn_lo_hi_lo_8 = {queue_dataIn_lo_hi_lo_hi_4, queue_dataIn_lo_hi_lo_lo_4};
  wire         queue_4_enq_bits_decodeResult_unOrderWrite;
  wire         queue_4_enq_bits_decodeResult_compress;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi_4 = {queue_4_enq_bits_decodeResult_unOrderWrite, queue_4_enq_bits_decodeResult_compress};
  wire         queue_4_enq_bits_decodeResult_gather16;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo_4 = {queue_dataIn_lo_hi_hi_lo_hi_4, queue_4_enq_bits_decodeResult_gather16};
  wire         queue_4_enq_bits_decodeResult_iota;
  wire         queue_4_enq_bits_decodeResult_mv;
  wire [1:0]   queue_dataIn_lo_hi_hi_hi_hi_4 = {queue_4_enq_bits_decodeResult_iota, queue_4_enq_bits_decodeResult_mv};
  wire         queue_4_enq_bits_decodeResult_extend;
  wire [2:0]   queue_dataIn_lo_hi_hi_hi_4 = {queue_dataIn_lo_hi_hi_hi_hi_4, queue_4_enq_bits_decodeResult_extend};
  wire [5:0]   queue_dataIn_lo_hi_hi_8 = {queue_dataIn_lo_hi_hi_hi_4, queue_dataIn_lo_hi_hi_lo_4};
  wire [10:0]  queue_dataIn_lo_hi_13 = {queue_dataIn_lo_hi_hi_8, queue_dataIn_lo_hi_lo_8};
  wire [21:0]  queue_dataIn_lo_13 = {queue_dataIn_lo_hi_13, queue_dataIn_lo_lo_8};
  wire         queue_4_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_4_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_hi_lo_lo_lo_4 = {queue_4_enq_bits_decodeResult_maskLogic, queue_4_enq_bits_decodeResult_uop};
  wire         queue_4_enq_bits_decodeResult_readOnly;
  wire         queue_4_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi_4 = {queue_4_enq_bits_decodeResult_readOnly, queue_4_enq_bits_decodeResult_maskSource};
  wire         queue_4_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi_4 = {queue_dataIn_hi_lo_lo_hi_hi_4, queue_4_enq_bits_decodeResult_maskDestination};
  wire [7:0]   queue_dataIn_hi_lo_lo_8 = {queue_dataIn_hi_lo_lo_hi_4, queue_dataIn_hi_lo_lo_lo_4};
  wire         queue_4_enq_bits_decodeResult_special;
  wire         queue_4_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi_4 = {queue_4_enq_bits_decodeResult_special, queue_4_enq_bits_decodeResult_saturate};
  wire         queue_4_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo_4 = {queue_dataIn_hi_lo_hi_lo_hi_4, queue_4_enq_bits_decodeResult_vwmacc};
  wire         queue_4_enq_bits_decodeResult_crossRead;
  wire         queue_4_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi_4 = {queue_4_enq_bits_decodeResult_crossRead, queue_4_enq_bits_decodeResult_crossWrite};
  wire         queue_4_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi_4 = {queue_dataIn_hi_lo_hi_hi_hi_4, queue_4_enq_bits_decodeResult_maskUnit};
  wire [5:0]   queue_dataIn_hi_lo_hi_8 = {queue_dataIn_hi_lo_hi_hi_4, queue_dataIn_hi_lo_hi_lo_4};
  wire [13:0]  queue_dataIn_hi_lo_13 = {queue_dataIn_hi_lo_hi_8, queue_dataIn_hi_lo_lo_8};
  wire         queue_4_enq_bits_decodeResult_vtype;
  wire         queue_4_enq_bits_decodeResult_sWrite;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo_4 = {queue_4_enq_bits_decodeResult_vtype, queue_4_enq_bits_decodeResult_sWrite};
  wire         queue_4_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_4_enq_bits_decodeResult_scheduler;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi_4 = {queue_4_enq_bits_decodeResult_dontNeedExecuteInLane, queue_4_enq_bits_decodeResult_scheduler};
  wire         queue_4_enq_bits_decodeResult_sReadVD;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi_4 = {queue_dataIn_hi_hi_lo_hi_hi_4, queue_4_enq_bits_decodeResult_sReadVD};
  wire [4:0]   queue_dataIn_hi_hi_lo_8 = {queue_dataIn_hi_hi_lo_hi_4, queue_dataIn_hi_hi_lo_lo_4};
  wire         queue_4_enq_bits_decodeResult_ffo;
  wire         queue_4_enq_bits_decodeResult_average;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi_4 = {queue_4_enq_bits_decodeResult_ffo, queue_4_enq_bits_decodeResult_average};
  wire         queue_4_enq_bits_decodeResult_reverse;
  wire [2:0]   queue_dataIn_hi_hi_hi_lo_4 = {queue_dataIn_hi_hi_hi_lo_hi_4, queue_4_enq_bits_decodeResult_reverse};
  wire         queue_4_enq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_4_enq_bits_decodeResult_topUop;
  wire [5:0]   queue_dataIn_hi_hi_hi_hi_hi_4 = {queue_4_enq_bits_decodeResult_specialSlot, queue_4_enq_bits_decodeResult_topUop};
  wire         queue_4_enq_bits_decodeResult_popCount;
  wire [6:0]   queue_dataIn_hi_hi_hi_hi_4 = {queue_dataIn_hi_hi_hi_hi_hi_4, queue_4_enq_bits_decodeResult_popCount};
  wire [9:0]   queue_dataIn_hi_hi_hi_8 = {queue_dataIn_hi_hi_hi_hi_4, queue_dataIn_hi_hi_hi_lo_4};
  wire [14:0]  queue_dataIn_hi_hi_13 = {queue_dataIn_hi_hi_hi_8, queue_dataIn_hi_hi_lo_8};
  wire [28:0]  queue_dataIn_hi_13 = {queue_dataIn_hi_hi_13, queue_dataIn_hi_lo_13};
  wire [2:0]   queue_4_enq_bits_segment;
  wire [31:0]  queue_4_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_9 = {queue_4_enq_bits_segment, queue_4_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_9 = {queue_dataIn_lo_lo_hi_9, queue_dataIn_hi_12, queue_dataIn_lo_12};
  wire [1:0]   queue_4_enq_bits_loadStoreEEW;
  wire         queue_4_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_9 = {queue_4_enq_bits_loadStoreEEW, queue_4_enq_bits_mask};
  wire [4:0]   queue_4_enq_bits_vs2;
  wire [4:0]   queue_4_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_9 = {queue_4_enq_bits_vs2, queue_4_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_14 = {queue_dataIn_lo_hi_hi_9, queue_dataIn_lo_hi_lo_9};
  wire [80:0]  queue_dataIn_lo_14 = {queue_dataIn_lo_hi_14, queue_dataIn_lo_lo_9};
  wire         queue_4_enq_bits_lsWholeReg;
  wire [4:0]   queue_4_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_9 = {queue_4_enq_bits_lsWholeReg, queue_4_enq_bits_vs1};
  wire         queue_4_enq_bits_store;
  wire         queue_4_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_9 = {queue_4_enq_bits_store, queue_4_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_14 = {queue_dataIn_hi_lo_hi_9, queue_dataIn_hi_lo_lo_9};
  wire         queue_4_enq_bits_loadStore;
  wire         queue_4_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_9 = {queue_4_enq_bits_loadStore, queue_4_enq_bits_issueInst};
  wire [2:0]   queue_4_enq_bits_instructionIndex;
  wire [53:0]  queue_dataIn_hi_hi_hi_9 = {queue_4_enq_bits_instructionIndex, queue_dataIn_hi_13, queue_dataIn_lo_13};
  wire [55:0]  queue_dataIn_hi_hi_14 = {queue_dataIn_hi_hi_hi_9, queue_dataIn_hi_hi_lo_9};
  wire [63:0]  queue_dataIn_hi_14 = {queue_dataIn_hi_hi_14, queue_dataIn_hi_lo_14};
  wire [144:0] queue_dataIn_4 = {queue_dataIn_hi_14, queue_dataIn_lo_14};
  wire         queue_dataOut_4_csrInterface_vma = _queue_fifo_4_data_out[0];
  wire         queue_dataOut_4_csrInterface_vta = _queue_fifo_4_data_out[1];
  wire [1:0]   queue_dataOut_4_csrInterface_vxrm = _queue_fifo_4_data_out[3:2];
  wire [1:0]   queue_dataOut_4_csrInterface_vSew = _queue_fifo_4_data_out[5:4];
  wire [2:0]   queue_dataOut_4_csrInterface_vlmul = _queue_fifo_4_data_out[8:6];
  wire [11:0]  queue_dataOut_4_csrInterface_vStart = _queue_fifo_4_data_out[20:9];
  wire [11:0]  queue_dataOut_4_csrInterface_vl = _queue_fifo_4_data_out[32:21];
  wire [31:0]  queue_dataOut_4_readFromScalar = _queue_fifo_4_data_out[64:33];
  wire [2:0]   queue_dataOut_4_segment = _queue_fifo_4_data_out[67:65];
  wire         queue_dataOut_4_mask = _queue_fifo_4_data_out[68];
  wire [1:0]   queue_dataOut_4_loadStoreEEW = _queue_fifo_4_data_out[70:69];
  wire [4:0]   queue_dataOut_4_vd = _queue_fifo_4_data_out[75:71];
  wire [4:0]   queue_dataOut_4_vs2 = _queue_fifo_4_data_out[80:76];
  wire [4:0]   queue_dataOut_4_vs1 = _queue_fifo_4_data_out[85:81];
  wire         queue_dataOut_4_lsWholeReg = _queue_fifo_4_data_out[86];
  wire         queue_dataOut_4_special = _queue_fifo_4_data_out[87];
  wire         queue_dataOut_4_store = _queue_fifo_4_data_out[88];
  wire         queue_dataOut_4_issueInst = _queue_fifo_4_data_out[89];
  wire         queue_dataOut_4_loadStore = _queue_fifo_4_data_out[90];
  wire         queue_dataOut_4_decodeResult_logic = _queue_fifo_4_data_out[91];
  wire         queue_dataOut_4_decodeResult_adder = _queue_fifo_4_data_out[92];
  wire         queue_dataOut_4_decodeResult_shift = _queue_fifo_4_data_out[93];
  wire         queue_dataOut_4_decodeResult_multiplier = _queue_fifo_4_data_out[94];
  wire         queue_dataOut_4_decodeResult_divider = _queue_fifo_4_data_out[95];
  wire         queue_dataOut_4_decodeResult_multiCycle = _queue_fifo_4_data_out[96];
  wire         queue_dataOut_4_decodeResult_other = _queue_fifo_4_data_out[97];
  wire         queue_dataOut_4_decodeResult_unsigned0 = _queue_fifo_4_data_out[98];
  wire         queue_dataOut_4_decodeResult_unsigned1 = _queue_fifo_4_data_out[99];
  wire         queue_dataOut_4_decodeResult_itype = _queue_fifo_4_data_out[100];
  wire         queue_dataOut_4_decodeResult_nr = _queue_fifo_4_data_out[101];
  wire         queue_dataOut_4_decodeResult_red = _queue_fifo_4_data_out[102];
  wire         queue_dataOut_4_decodeResult_widenReduce = _queue_fifo_4_data_out[103];
  wire         queue_dataOut_4_decodeResult_targetRd = _queue_fifo_4_data_out[104];
  wire         queue_dataOut_4_decodeResult_slid = _queue_fifo_4_data_out[105];
  wire         queue_dataOut_4_decodeResult_gather = _queue_fifo_4_data_out[106];
  wire         queue_dataOut_4_decodeResult_gather16 = _queue_fifo_4_data_out[107];
  wire         queue_dataOut_4_decodeResult_compress = _queue_fifo_4_data_out[108];
  wire         queue_dataOut_4_decodeResult_unOrderWrite = _queue_fifo_4_data_out[109];
  wire         queue_dataOut_4_decodeResult_extend = _queue_fifo_4_data_out[110];
  wire         queue_dataOut_4_decodeResult_mv = _queue_fifo_4_data_out[111];
  wire         queue_dataOut_4_decodeResult_iota = _queue_fifo_4_data_out[112];
  wire [3:0]   queue_dataOut_4_decodeResult_uop = _queue_fifo_4_data_out[116:113];
  wire         queue_dataOut_4_decodeResult_maskLogic = _queue_fifo_4_data_out[117];
  wire         queue_dataOut_4_decodeResult_maskDestination = _queue_fifo_4_data_out[118];
  wire         queue_dataOut_4_decodeResult_maskSource = _queue_fifo_4_data_out[119];
  wire         queue_dataOut_4_decodeResult_readOnly = _queue_fifo_4_data_out[120];
  wire         queue_dataOut_4_decodeResult_vwmacc = _queue_fifo_4_data_out[121];
  wire         queue_dataOut_4_decodeResult_saturate = _queue_fifo_4_data_out[122];
  wire         queue_dataOut_4_decodeResult_special = _queue_fifo_4_data_out[123];
  wire         queue_dataOut_4_decodeResult_maskUnit = _queue_fifo_4_data_out[124];
  wire         queue_dataOut_4_decodeResult_crossWrite = _queue_fifo_4_data_out[125];
  wire         queue_dataOut_4_decodeResult_crossRead = _queue_fifo_4_data_out[126];
  wire         queue_dataOut_4_decodeResult_sWrite = _queue_fifo_4_data_out[127];
  wire         queue_dataOut_4_decodeResult_vtype = _queue_fifo_4_data_out[128];
  wire         queue_dataOut_4_decodeResult_sReadVD = _queue_fifo_4_data_out[129];
  wire         queue_dataOut_4_decodeResult_scheduler = _queue_fifo_4_data_out[130];
  wire         queue_dataOut_4_decodeResult_dontNeedExecuteInLane = _queue_fifo_4_data_out[131];
  wire         queue_dataOut_4_decodeResult_reverse = _queue_fifo_4_data_out[132];
  wire         queue_dataOut_4_decodeResult_average = _queue_fifo_4_data_out[133];
  wire         queue_dataOut_4_decodeResult_ffo = _queue_fifo_4_data_out[134];
  wire         queue_dataOut_4_decodeResult_popCount = _queue_fifo_4_data_out[135];
  wire [4:0]   queue_dataOut_4_decodeResult_topUop = _queue_fifo_4_data_out[140:136];
  wire         queue_dataOut_4_decodeResult_specialSlot = _queue_fifo_4_data_out[141];
  wire [2:0]   queue_dataOut_4_instructionIndex = _queue_fifo_4_data_out[144:142];
  wire         queue_4_enq_ready = ~_queue_fifo_4_full;
  wire         queue_4_enq_valid;
  assign queue_4_deq_valid = ~_queue_fifo_4_empty | queue_4_enq_valid;
  assign queue_4_deq_bits_instructionIndex = _queue_fifo_4_empty ? queue_4_enq_bits_instructionIndex : queue_dataOut_4_instructionIndex;
  assign queue_4_deq_bits_decodeResult_specialSlot = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_specialSlot : queue_dataOut_4_decodeResult_specialSlot;
  assign queue_4_deq_bits_decodeResult_topUop = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_topUop : queue_dataOut_4_decodeResult_topUop;
  assign queue_4_deq_bits_decodeResult_popCount = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_popCount : queue_dataOut_4_decodeResult_popCount;
  assign queue_4_deq_bits_decodeResult_ffo = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_ffo : queue_dataOut_4_decodeResult_ffo;
  assign queue_4_deq_bits_decodeResult_average = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_average : queue_dataOut_4_decodeResult_average;
  assign queue_4_deq_bits_decodeResult_reverse = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_reverse : queue_dataOut_4_decodeResult_reverse;
  assign queue_4_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_4_decodeResult_dontNeedExecuteInLane;
  assign queue_4_deq_bits_decodeResult_scheduler = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_scheduler : queue_dataOut_4_decodeResult_scheduler;
  assign queue_4_deq_bits_decodeResult_sReadVD = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_sReadVD : queue_dataOut_4_decodeResult_sReadVD;
  assign queue_4_deq_bits_decodeResult_vtype = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_vtype : queue_dataOut_4_decodeResult_vtype;
  assign queue_4_deq_bits_decodeResult_sWrite = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_sWrite : queue_dataOut_4_decodeResult_sWrite;
  assign queue_4_deq_bits_decodeResult_crossRead = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_crossRead : queue_dataOut_4_decodeResult_crossRead;
  assign queue_4_deq_bits_decodeResult_crossWrite = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_crossWrite : queue_dataOut_4_decodeResult_crossWrite;
  assign queue_4_deq_bits_decodeResult_maskUnit = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_maskUnit : queue_dataOut_4_decodeResult_maskUnit;
  assign queue_4_deq_bits_decodeResult_special = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_special : queue_dataOut_4_decodeResult_special;
  assign queue_4_deq_bits_decodeResult_saturate = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_saturate : queue_dataOut_4_decodeResult_saturate;
  assign queue_4_deq_bits_decodeResult_vwmacc = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_vwmacc : queue_dataOut_4_decodeResult_vwmacc;
  assign queue_4_deq_bits_decodeResult_readOnly = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_readOnly : queue_dataOut_4_decodeResult_readOnly;
  assign queue_4_deq_bits_decodeResult_maskSource = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_maskSource : queue_dataOut_4_decodeResult_maskSource;
  assign queue_4_deq_bits_decodeResult_maskDestination = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_maskDestination : queue_dataOut_4_decodeResult_maskDestination;
  assign queue_4_deq_bits_decodeResult_maskLogic = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_maskLogic : queue_dataOut_4_decodeResult_maskLogic;
  assign queue_4_deq_bits_decodeResult_uop = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_uop : queue_dataOut_4_decodeResult_uop;
  assign queue_4_deq_bits_decodeResult_iota = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_iota : queue_dataOut_4_decodeResult_iota;
  assign queue_4_deq_bits_decodeResult_mv = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_mv : queue_dataOut_4_decodeResult_mv;
  assign queue_4_deq_bits_decodeResult_extend = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_extend : queue_dataOut_4_decodeResult_extend;
  assign queue_4_deq_bits_decodeResult_unOrderWrite = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_unOrderWrite : queue_dataOut_4_decodeResult_unOrderWrite;
  assign queue_4_deq_bits_decodeResult_compress = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_compress : queue_dataOut_4_decodeResult_compress;
  assign queue_4_deq_bits_decodeResult_gather16 = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_gather16 : queue_dataOut_4_decodeResult_gather16;
  assign queue_4_deq_bits_decodeResult_gather = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_gather : queue_dataOut_4_decodeResult_gather;
  assign queue_4_deq_bits_decodeResult_slid = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_slid : queue_dataOut_4_decodeResult_slid;
  assign queue_4_deq_bits_decodeResult_targetRd = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_targetRd : queue_dataOut_4_decodeResult_targetRd;
  assign queue_4_deq_bits_decodeResult_widenReduce = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_widenReduce : queue_dataOut_4_decodeResult_widenReduce;
  assign queue_4_deq_bits_decodeResult_red = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_red : queue_dataOut_4_decodeResult_red;
  assign queue_4_deq_bits_decodeResult_nr = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_nr : queue_dataOut_4_decodeResult_nr;
  assign queue_4_deq_bits_decodeResult_itype = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_itype : queue_dataOut_4_decodeResult_itype;
  assign queue_4_deq_bits_decodeResult_unsigned1 = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_unsigned1 : queue_dataOut_4_decodeResult_unsigned1;
  assign queue_4_deq_bits_decodeResult_unsigned0 = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_unsigned0 : queue_dataOut_4_decodeResult_unsigned0;
  assign queue_4_deq_bits_decodeResult_other = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_other : queue_dataOut_4_decodeResult_other;
  assign queue_4_deq_bits_decodeResult_multiCycle = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_multiCycle : queue_dataOut_4_decodeResult_multiCycle;
  assign queue_4_deq_bits_decodeResult_divider = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_divider : queue_dataOut_4_decodeResult_divider;
  assign queue_4_deq_bits_decodeResult_multiplier = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_multiplier : queue_dataOut_4_decodeResult_multiplier;
  assign queue_4_deq_bits_decodeResult_shift = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_shift : queue_dataOut_4_decodeResult_shift;
  assign queue_4_deq_bits_decodeResult_adder = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_adder : queue_dataOut_4_decodeResult_adder;
  assign queue_4_deq_bits_decodeResult_logic = _queue_fifo_4_empty ? queue_4_enq_bits_decodeResult_logic : queue_dataOut_4_decodeResult_logic;
  assign queue_4_deq_bits_loadStore = _queue_fifo_4_empty ? queue_4_enq_bits_loadStore : queue_dataOut_4_loadStore;
  assign queue_4_deq_bits_issueInst = _queue_fifo_4_empty ? queue_4_enq_bits_issueInst : queue_dataOut_4_issueInst;
  assign queue_4_deq_bits_store = _queue_fifo_4_empty ? queue_4_enq_bits_store : queue_dataOut_4_store;
  assign queue_4_deq_bits_special = _queue_fifo_4_empty ? queue_4_enq_bits_special : queue_dataOut_4_special;
  assign queue_4_deq_bits_lsWholeReg = _queue_fifo_4_empty ? queue_4_enq_bits_lsWholeReg : queue_dataOut_4_lsWholeReg;
  assign queue_4_deq_bits_vs1 = _queue_fifo_4_empty ? queue_4_enq_bits_vs1 : queue_dataOut_4_vs1;
  assign queue_4_deq_bits_vs2 = _queue_fifo_4_empty ? queue_4_enq_bits_vs2 : queue_dataOut_4_vs2;
  assign queue_4_deq_bits_vd = _queue_fifo_4_empty ? queue_4_enq_bits_vd : queue_dataOut_4_vd;
  assign queue_4_deq_bits_loadStoreEEW = _queue_fifo_4_empty ? queue_4_enq_bits_loadStoreEEW : queue_dataOut_4_loadStoreEEW;
  assign queue_4_deq_bits_mask = _queue_fifo_4_empty ? queue_4_enq_bits_mask : queue_dataOut_4_mask;
  assign queue_4_deq_bits_segment = _queue_fifo_4_empty ? queue_4_enq_bits_segment : queue_dataOut_4_segment;
  assign queue_4_deq_bits_readFromScalar = _queue_fifo_4_empty ? queue_4_enq_bits_readFromScalar : queue_dataOut_4_readFromScalar;
  assign queue_4_deq_bits_csrInterface_vl = _queue_fifo_4_empty ? queue_4_enq_bits_csrInterface_vl : queue_dataOut_4_csrInterface_vl;
  assign queue_4_deq_bits_csrInterface_vStart = _queue_fifo_4_empty ? queue_4_enq_bits_csrInterface_vStart : queue_dataOut_4_csrInterface_vStart;
  assign queue_4_deq_bits_csrInterface_vlmul = _queue_fifo_4_empty ? queue_4_enq_bits_csrInterface_vlmul : queue_dataOut_4_csrInterface_vlmul;
  assign queue_4_deq_bits_csrInterface_vSew = _queue_fifo_4_empty ? queue_4_enq_bits_csrInterface_vSew : queue_dataOut_4_csrInterface_vSew;
  assign queue_4_deq_bits_csrInterface_vxrm = _queue_fifo_4_empty ? queue_4_enq_bits_csrInterface_vxrm : queue_dataOut_4_csrInterface_vxrm;
  assign queue_4_deq_bits_csrInterface_vta = _queue_fifo_4_empty ? queue_4_enq_bits_csrInterface_vta : queue_dataOut_4_csrInterface_vta;
  assign queue_4_deq_bits_csrInterface_vma = _queue_fifo_4_empty ? queue_4_enq_bits_csrInterface_vma : queue_dataOut_4_csrInterface_vma;
  wire         laneVec_4_laneRequest_bits_issueInst = laneRequestSinkWire_4_ready & laneRequestSinkWire_4_valid;
  reg          releasePipe_pipe_v_4;
  wire         releasePipe_pipe_out_4_valid = releasePipe_pipe_v_4;
  wire         laneRequestSourceWire_4_ready;
  wire         validSource_4_valid = laneRequestSourceWire_4_ready & laneRequestSourceWire_4_valid;
  reg  [2:0]   tokenCheck_counter_4;
  wire [2:0]   tokenCheck_counterChange_4 = validSource_4_valid ? 3'h1 : 3'h7;
  assign tokenCheck_4 = ~(tokenCheck_counter_4[2]);
  assign laneRequestSourceWire_4_ready = tokenCheck_4;
  assign queue_4_enq_valid = validSink_4_valid;
  assign queue_4_enq_bits_instructionIndex = validSink_4_bits_instructionIndex;
  assign queue_4_enq_bits_decodeResult_specialSlot = validSink_4_bits_decodeResult_specialSlot;
  assign queue_4_enq_bits_decodeResult_topUop = validSink_4_bits_decodeResult_topUop;
  assign queue_4_enq_bits_decodeResult_popCount = validSink_4_bits_decodeResult_popCount;
  assign queue_4_enq_bits_decodeResult_ffo = validSink_4_bits_decodeResult_ffo;
  assign queue_4_enq_bits_decodeResult_average = validSink_4_bits_decodeResult_average;
  assign queue_4_enq_bits_decodeResult_reverse = validSink_4_bits_decodeResult_reverse;
  assign queue_4_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_4_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_4_enq_bits_decodeResult_scheduler = validSink_4_bits_decodeResult_scheduler;
  assign queue_4_enq_bits_decodeResult_sReadVD = validSink_4_bits_decodeResult_sReadVD;
  assign queue_4_enq_bits_decodeResult_vtype = validSink_4_bits_decodeResult_vtype;
  assign queue_4_enq_bits_decodeResult_sWrite = validSink_4_bits_decodeResult_sWrite;
  assign queue_4_enq_bits_decodeResult_crossRead = validSink_4_bits_decodeResult_crossRead;
  assign queue_4_enq_bits_decodeResult_crossWrite = validSink_4_bits_decodeResult_crossWrite;
  assign queue_4_enq_bits_decodeResult_maskUnit = validSink_4_bits_decodeResult_maskUnit;
  assign queue_4_enq_bits_decodeResult_special = validSink_4_bits_decodeResult_special;
  assign queue_4_enq_bits_decodeResult_saturate = validSink_4_bits_decodeResult_saturate;
  assign queue_4_enq_bits_decodeResult_vwmacc = validSink_4_bits_decodeResult_vwmacc;
  assign queue_4_enq_bits_decodeResult_readOnly = validSink_4_bits_decodeResult_readOnly;
  assign queue_4_enq_bits_decodeResult_maskSource = validSink_4_bits_decodeResult_maskSource;
  assign queue_4_enq_bits_decodeResult_maskDestination = validSink_4_bits_decodeResult_maskDestination;
  assign queue_4_enq_bits_decodeResult_maskLogic = validSink_4_bits_decodeResult_maskLogic;
  assign queue_4_enq_bits_decodeResult_uop = validSink_4_bits_decodeResult_uop;
  assign queue_4_enq_bits_decodeResult_iota = validSink_4_bits_decodeResult_iota;
  assign queue_4_enq_bits_decodeResult_mv = validSink_4_bits_decodeResult_mv;
  assign queue_4_enq_bits_decodeResult_extend = validSink_4_bits_decodeResult_extend;
  assign queue_4_enq_bits_decodeResult_unOrderWrite = validSink_4_bits_decodeResult_unOrderWrite;
  assign queue_4_enq_bits_decodeResult_compress = validSink_4_bits_decodeResult_compress;
  assign queue_4_enq_bits_decodeResult_gather16 = validSink_4_bits_decodeResult_gather16;
  assign queue_4_enq_bits_decodeResult_gather = validSink_4_bits_decodeResult_gather;
  assign queue_4_enq_bits_decodeResult_slid = validSink_4_bits_decodeResult_slid;
  assign queue_4_enq_bits_decodeResult_targetRd = validSink_4_bits_decodeResult_targetRd;
  assign queue_4_enq_bits_decodeResult_widenReduce = validSink_4_bits_decodeResult_widenReduce;
  assign queue_4_enq_bits_decodeResult_red = validSink_4_bits_decodeResult_red;
  assign queue_4_enq_bits_decodeResult_nr = validSink_4_bits_decodeResult_nr;
  assign queue_4_enq_bits_decodeResult_itype = validSink_4_bits_decodeResult_itype;
  assign queue_4_enq_bits_decodeResult_unsigned1 = validSink_4_bits_decodeResult_unsigned1;
  assign queue_4_enq_bits_decodeResult_unsigned0 = validSink_4_bits_decodeResult_unsigned0;
  assign queue_4_enq_bits_decodeResult_other = validSink_4_bits_decodeResult_other;
  assign queue_4_enq_bits_decodeResult_multiCycle = validSink_4_bits_decodeResult_multiCycle;
  assign queue_4_enq_bits_decodeResult_divider = validSink_4_bits_decodeResult_divider;
  assign queue_4_enq_bits_decodeResult_multiplier = validSink_4_bits_decodeResult_multiplier;
  assign queue_4_enq_bits_decodeResult_shift = validSink_4_bits_decodeResult_shift;
  assign queue_4_enq_bits_decodeResult_adder = validSink_4_bits_decodeResult_adder;
  assign queue_4_enq_bits_decodeResult_logic = validSink_4_bits_decodeResult_logic;
  assign queue_4_enq_bits_loadStore = validSink_4_bits_loadStore;
  assign queue_4_enq_bits_issueInst = validSink_4_bits_issueInst;
  assign queue_4_enq_bits_store = validSink_4_bits_store;
  assign queue_4_enq_bits_special = validSink_4_bits_special;
  assign queue_4_enq_bits_lsWholeReg = validSink_4_bits_lsWholeReg;
  assign queue_4_enq_bits_vs1 = validSink_4_bits_vs1;
  assign queue_4_enq_bits_vs2 = validSink_4_bits_vs2;
  assign queue_4_enq_bits_vd = validSink_4_bits_vd;
  assign queue_4_enq_bits_loadStoreEEW = validSink_4_bits_loadStoreEEW;
  assign queue_4_enq_bits_mask = validSink_4_bits_mask;
  assign queue_4_enq_bits_segment = validSink_4_bits_segment;
  assign queue_4_enq_bits_readFromScalar = validSink_4_bits_readFromScalar;
  assign queue_4_enq_bits_csrInterface_vl = validSink_4_bits_csrInterface_vl;
  assign queue_4_enq_bits_csrInterface_vStart = validSink_4_bits_csrInterface_vStart;
  assign queue_4_enq_bits_csrInterface_vlmul = validSink_4_bits_csrInterface_vlmul;
  assign queue_4_enq_bits_csrInterface_vSew = validSink_4_bits_csrInterface_vSew;
  assign queue_4_enq_bits_csrInterface_vxrm = validSink_4_bits_csrInterface_vxrm;
  assign queue_4_enq_bits_csrInterface_vta = validSink_4_bits_csrInterface_vta;
  assign queue_4_enq_bits_csrInterface_vma = validSink_4_bits_csrInterface_vma;
  reg          shifterReg_4_0_valid;
  assign validSink_4_valid = shifterReg_4_0_valid;
  reg  [2:0]   shifterReg_4_0_bits_instructionIndex;
  assign validSink_4_bits_instructionIndex = shifterReg_4_0_bits_instructionIndex;
  reg          shifterReg_4_0_bits_decodeResult_specialSlot;
  assign validSink_4_bits_decodeResult_specialSlot = shifterReg_4_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_4_0_bits_decodeResult_topUop;
  assign validSink_4_bits_decodeResult_topUop = shifterReg_4_0_bits_decodeResult_topUop;
  reg          shifterReg_4_0_bits_decodeResult_popCount;
  assign validSink_4_bits_decodeResult_popCount = shifterReg_4_0_bits_decodeResult_popCount;
  reg          shifterReg_4_0_bits_decodeResult_ffo;
  assign validSink_4_bits_decodeResult_ffo = shifterReg_4_0_bits_decodeResult_ffo;
  reg          shifterReg_4_0_bits_decodeResult_average;
  assign validSink_4_bits_decodeResult_average = shifterReg_4_0_bits_decodeResult_average;
  reg          shifterReg_4_0_bits_decodeResult_reverse;
  assign validSink_4_bits_decodeResult_reverse = shifterReg_4_0_bits_decodeResult_reverse;
  reg          shifterReg_4_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_4_bits_decodeResult_dontNeedExecuteInLane = shifterReg_4_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_4_0_bits_decodeResult_scheduler;
  assign validSink_4_bits_decodeResult_scheduler = shifterReg_4_0_bits_decodeResult_scheduler;
  reg          shifterReg_4_0_bits_decodeResult_sReadVD;
  assign validSink_4_bits_decodeResult_sReadVD = shifterReg_4_0_bits_decodeResult_sReadVD;
  reg          shifterReg_4_0_bits_decodeResult_vtype;
  assign validSink_4_bits_decodeResult_vtype = shifterReg_4_0_bits_decodeResult_vtype;
  reg          shifterReg_4_0_bits_decodeResult_sWrite;
  assign validSink_4_bits_decodeResult_sWrite = shifterReg_4_0_bits_decodeResult_sWrite;
  reg          shifterReg_4_0_bits_decodeResult_crossRead;
  assign validSink_4_bits_decodeResult_crossRead = shifterReg_4_0_bits_decodeResult_crossRead;
  reg          shifterReg_4_0_bits_decodeResult_crossWrite;
  assign validSink_4_bits_decodeResult_crossWrite = shifterReg_4_0_bits_decodeResult_crossWrite;
  reg          shifterReg_4_0_bits_decodeResult_maskUnit;
  assign validSink_4_bits_decodeResult_maskUnit = shifterReg_4_0_bits_decodeResult_maskUnit;
  reg          shifterReg_4_0_bits_decodeResult_special;
  assign validSink_4_bits_decodeResult_special = shifterReg_4_0_bits_decodeResult_special;
  reg          shifterReg_4_0_bits_decodeResult_saturate;
  assign validSink_4_bits_decodeResult_saturate = shifterReg_4_0_bits_decodeResult_saturate;
  reg          shifterReg_4_0_bits_decodeResult_vwmacc;
  assign validSink_4_bits_decodeResult_vwmacc = shifterReg_4_0_bits_decodeResult_vwmacc;
  reg          shifterReg_4_0_bits_decodeResult_readOnly;
  assign validSink_4_bits_decodeResult_readOnly = shifterReg_4_0_bits_decodeResult_readOnly;
  reg          shifterReg_4_0_bits_decodeResult_maskSource;
  assign validSink_4_bits_decodeResult_maskSource = shifterReg_4_0_bits_decodeResult_maskSource;
  reg          shifterReg_4_0_bits_decodeResult_maskDestination;
  assign validSink_4_bits_decodeResult_maskDestination = shifterReg_4_0_bits_decodeResult_maskDestination;
  reg          shifterReg_4_0_bits_decodeResult_maskLogic;
  assign validSink_4_bits_decodeResult_maskLogic = shifterReg_4_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_4_0_bits_decodeResult_uop;
  assign validSink_4_bits_decodeResult_uop = shifterReg_4_0_bits_decodeResult_uop;
  reg          shifterReg_4_0_bits_decodeResult_iota;
  assign validSink_4_bits_decodeResult_iota = shifterReg_4_0_bits_decodeResult_iota;
  reg          shifterReg_4_0_bits_decodeResult_mv;
  assign validSink_4_bits_decodeResult_mv = shifterReg_4_0_bits_decodeResult_mv;
  reg          shifterReg_4_0_bits_decodeResult_extend;
  assign validSink_4_bits_decodeResult_extend = shifterReg_4_0_bits_decodeResult_extend;
  reg          shifterReg_4_0_bits_decodeResult_unOrderWrite;
  assign validSink_4_bits_decodeResult_unOrderWrite = shifterReg_4_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_4_0_bits_decodeResult_compress;
  assign validSink_4_bits_decodeResult_compress = shifterReg_4_0_bits_decodeResult_compress;
  reg          shifterReg_4_0_bits_decodeResult_gather16;
  assign validSink_4_bits_decodeResult_gather16 = shifterReg_4_0_bits_decodeResult_gather16;
  reg          shifterReg_4_0_bits_decodeResult_gather;
  assign validSink_4_bits_decodeResult_gather = shifterReg_4_0_bits_decodeResult_gather;
  reg          shifterReg_4_0_bits_decodeResult_slid;
  assign validSink_4_bits_decodeResult_slid = shifterReg_4_0_bits_decodeResult_slid;
  reg          shifterReg_4_0_bits_decodeResult_targetRd;
  assign validSink_4_bits_decodeResult_targetRd = shifterReg_4_0_bits_decodeResult_targetRd;
  reg          shifterReg_4_0_bits_decodeResult_widenReduce;
  assign validSink_4_bits_decodeResult_widenReduce = shifterReg_4_0_bits_decodeResult_widenReduce;
  reg          shifterReg_4_0_bits_decodeResult_red;
  assign validSink_4_bits_decodeResult_red = shifterReg_4_0_bits_decodeResult_red;
  reg          shifterReg_4_0_bits_decodeResult_nr;
  assign validSink_4_bits_decodeResult_nr = shifterReg_4_0_bits_decodeResult_nr;
  reg          shifterReg_4_0_bits_decodeResult_itype;
  assign validSink_4_bits_decodeResult_itype = shifterReg_4_0_bits_decodeResult_itype;
  reg          shifterReg_4_0_bits_decodeResult_unsigned1;
  assign validSink_4_bits_decodeResult_unsigned1 = shifterReg_4_0_bits_decodeResult_unsigned1;
  reg          shifterReg_4_0_bits_decodeResult_unsigned0;
  assign validSink_4_bits_decodeResult_unsigned0 = shifterReg_4_0_bits_decodeResult_unsigned0;
  reg          shifterReg_4_0_bits_decodeResult_other;
  assign validSink_4_bits_decodeResult_other = shifterReg_4_0_bits_decodeResult_other;
  reg          shifterReg_4_0_bits_decodeResult_multiCycle;
  assign validSink_4_bits_decodeResult_multiCycle = shifterReg_4_0_bits_decodeResult_multiCycle;
  reg          shifterReg_4_0_bits_decodeResult_divider;
  assign validSink_4_bits_decodeResult_divider = shifterReg_4_0_bits_decodeResult_divider;
  reg          shifterReg_4_0_bits_decodeResult_multiplier;
  assign validSink_4_bits_decodeResult_multiplier = shifterReg_4_0_bits_decodeResult_multiplier;
  reg          shifterReg_4_0_bits_decodeResult_shift;
  assign validSink_4_bits_decodeResult_shift = shifterReg_4_0_bits_decodeResult_shift;
  reg          shifterReg_4_0_bits_decodeResult_adder;
  assign validSink_4_bits_decodeResult_adder = shifterReg_4_0_bits_decodeResult_adder;
  reg          shifterReg_4_0_bits_decodeResult_logic;
  assign validSink_4_bits_decodeResult_logic = shifterReg_4_0_bits_decodeResult_logic;
  reg          shifterReg_4_0_bits_loadStore;
  assign validSink_4_bits_loadStore = shifterReg_4_0_bits_loadStore;
  reg          shifterReg_4_0_bits_issueInst;
  assign validSink_4_bits_issueInst = shifterReg_4_0_bits_issueInst;
  reg          shifterReg_4_0_bits_store;
  assign validSink_4_bits_store = shifterReg_4_0_bits_store;
  reg          shifterReg_4_0_bits_special;
  assign validSink_4_bits_special = shifterReg_4_0_bits_special;
  reg          shifterReg_4_0_bits_lsWholeReg;
  assign validSink_4_bits_lsWholeReg = shifterReg_4_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_4_0_bits_vs1;
  assign validSink_4_bits_vs1 = shifterReg_4_0_bits_vs1;
  reg  [4:0]   shifterReg_4_0_bits_vs2;
  assign validSink_4_bits_vs2 = shifterReg_4_0_bits_vs2;
  reg  [4:0]   shifterReg_4_0_bits_vd;
  assign validSink_4_bits_vd = shifterReg_4_0_bits_vd;
  reg  [1:0]   shifterReg_4_0_bits_loadStoreEEW;
  assign validSink_4_bits_loadStoreEEW = shifterReg_4_0_bits_loadStoreEEW;
  reg          shifterReg_4_0_bits_mask;
  assign validSink_4_bits_mask = shifterReg_4_0_bits_mask;
  reg  [2:0]   shifterReg_4_0_bits_segment;
  assign validSink_4_bits_segment = shifterReg_4_0_bits_segment;
  reg  [31:0]  shifterReg_4_0_bits_readFromScalar;
  assign validSink_4_bits_readFromScalar = shifterReg_4_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_4_0_bits_csrInterface_vl;
  assign validSink_4_bits_csrInterface_vl = shifterReg_4_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_4_0_bits_csrInterface_vStart;
  assign validSink_4_bits_csrInterface_vStart = shifterReg_4_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_4_0_bits_csrInterface_vlmul;
  assign validSink_4_bits_csrInterface_vlmul = shifterReg_4_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_4_0_bits_csrInterface_vSew;
  assign validSink_4_bits_csrInterface_vSew = shifterReg_4_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_4_0_bits_csrInterface_vxrm;
  assign validSink_4_bits_csrInterface_vxrm = shifterReg_4_0_bits_csrInterface_vxrm;
  reg          shifterReg_4_0_bits_csrInterface_vta;
  assign validSink_4_bits_csrInterface_vta = shifterReg_4_0_bits_csrInterface_vta;
  reg          shifterReg_4_0_bits_csrInterface_vma;
  assign validSink_4_bits_csrInterface_vma = shifterReg_4_0_bits_csrInterface_vma;
  wire         shifterValid_4 = shifterReg_4_0_valid | validSource_4_valid;
  wire         validSink_5_valid;
  wire [2:0]   validSink_5_bits_instructionIndex;
  wire         validSink_5_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_5_bits_decodeResult_topUop;
  wire         validSink_5_bits_decodeResult_popCount;
  wire         validSink_5_bits_decodeResult_ffo;
  wire         validSink_5_bits_decodeResult_average;
  wire         validSink_5_bits_decodeResult_reverse;
  wire         validSink_5_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_5_bits_decodeResult_scheduler;
  wire         validSink_5_bits_decodeResult_sReadVD;
  wire         validSink_5_bits_decodeResult_vtype;
  wire         validSink_5_bits_decodeResult_sWrite;
  wire         validSink_5_bits_decodeResult_crossRead;
  wire         validSink_5_bits_decodeResult_crossWrite;
  wire         validSink_5_bits_decodeResult_maskUnit;
  wire         validSink_5_bits_decodeResult_special;
  wire         validSink_5_bits_decodeResult_saturate;
  wire         validSink_5_bits_decodeResult_vwmacc;
  wire         validSink_5_bits_decodeResult_readOnly;
  wire         validSink_5_bits_decodeResult_maskSource;
  wire         validSink_5_bits_decodeResult_maskDestination;
  wire         validSink_5_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_5_bits_decodeResult_uop;
  wire         validSink_5_bits_decodeResult_iota;
  wire         validSink_5_bits_decodeResult_mv;
  wire         validSink_5_bits_decodeResult_extend;
  wire         validSink_5_bits_decodeResult_unOrderWrite;
  wire         validSink_5_bits_decodeResult_compress;
  wire         validSink_5_bits_decodeResult_gather16;
  wire         validSink_5_bits_decodeResult_gather;
  wire         validSink_5_bits_decodeResult_slid;
  wire         validSink_5_bits_decodeResult_targetRd;
  wire         validSink_5_bits_decodeResult_widenReduce;
  wire         validSink_5_bits_decodeResult_red;
  wire         validSink_5_bits_decodeResult_nr;
  wire         validSink_5_bits_decodeResult_itype;
  wire         validSink_5_bits_decodeResult_unsigned1;
  wire         validSink_5_bits_decodeResult_unsigned0;
  wire         validSink_5_bits_decodeResult_other;
  wire         validSink_5_bits_decodeResult_multiCycle;
  wire         validSink_5_bits_decodeResult_divider;
  wire         validSink_5_bits_decodeResult_multiplier;
  wire         validSink_5_bits_decodeResult_shift;
  wire         validSink_5_bits_decodeResult_adder;
  wire         validSink_5_bits_decodeResult_logic;
  wire         validSink_5_bits_loadStore;
  wire         validSink_5_bits_issueInst;
  wire         validSink_5_bits_store;
  wire         validSink_5_bits_special;
  wire         validSink_5_bits_lsWholeReg;
  wire [4:0]   validSink_5_bits_vs1;
  wire [4:0]   validSink_5_bits_vs2;
  wire [4:0]   validSink_5_bits_vd;
  wire [1:0]   validSink_5_bits_loadStoreEEW;
  wire         validSink_5_bits_mask;
  wire [2:0]   validSink_5_bits_segment;
  wire [31:0]  validSink_5_bits_readFromScalar;
  wire [11:0]  validSink_5_bits_csrInterface_vl;
  wire [11:0]  validSink_5_bits_csrInterface_vStart;
  wire [2:0]   validSink_5_bits_csrInterface_vlmul;
  wire [1:0]   validSink_5_bits_csrInterface_vSew;
  wire [1:0]   validSink_5_bits_csrInterface_vxrm;
  wire         validSink_5_bits_csrInterface_vta;
  wire         validSink_5_bits_csrInterface_vma;
  wire         laneRequestSinkWire_5_valid = queue_5_deq_valid;
  wire [2:0]   laneRequestSinkWire_5_bits_instructionIndex = queue_5_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_5_bits_decodeResult_specialSlot = queue_5_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_5_bits_decodeResult_topUop = queue_5_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_5_bits_decodeResult_popCount = queue_5_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_5_bits_decodeResult_ffo = queue_5_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_5_bits_decodeResult_average = queue_5_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_5_bits_decodeResult_reverse = queue_5_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_5_bits_decodeResult_dontNeedExecuteInLane = queue_5_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_5_bits_decodeResult_scheduler = queue_5_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_5_bits_decodeResult_sReadVD = queue_5_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_5_bits_decodeResult_vtype = queue_5_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_5_bits_decodeResult_sWrite = queue_5_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_5_bits_decodeResult_crossRead = queue_5_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_5_bits_decodeResult_crossWrite = queue_5_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_5_bits_decodeResult_maskUnit = queue_5_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_5_bits_decodeResult_special = queue_5_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_5_bits_decodeResult_saturate = queue_5_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_5_bits_decodeResult_vwmacc = queue_5_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_5_bits_decodeResult_readOnly = queue_5_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_5_bits_decodeResult_maskSource = queue_5_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_5_bits_decodeResult_maskDestination = queue_5_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_5_bits_decodeResult_maskLogic = queue_5_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_5_bits_decodeResult_uop = queue_5_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_5_bits_decodeResult_iota = queue_5_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_5_bits_decodeResult_mv = queue_5_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_5_bits_decodeResult_extend = queue_5_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_5_bits_decodeResult_unOrderWrite = queue_5_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_5_bits_decodeResult_compress = queue_5_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_5_bits_decodeResult_gather16 = queue_5_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_5_bits_decodeResult_gather = queue_5_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_5_bits_decodeResult_slid = queue_5_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_5_bits_decodeResult_targetRd = queue_5_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_5_bits_decodeResult_widenReduce = queue_5_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_5_bits_decodeResult_red = queue_5_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_5_bits_decodeResult_nr = queue_5_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_5_bits_decodeResult_itype = queue_5_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_5_bits_decodeResult_unsigned1 = queue_5_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_5_bits_decodeResult_unsigned0 = queue_5_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_5_bits_decodeResult_other = queue_5_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_5_bits_decodeResult_multiCycle = queue_5_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_5_bits_decodeResult_divider = queue_5_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_5_bits_decodeResult_multiplier = queue_5_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_5_bits_decodeResult_shift = queue_5_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_5_bits_decodeResult_adder = queue_5_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_5_bits_decodeResult_logic = queue_5_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_5_bits_loadStore = queue_5_deq_bits_loadStore;
  wire         laneRequestSinkWire_5_bits_issueInst = queue_5_deq_bits_issueInst;
  wire         laneRequestSinkWire_5_bits_store = queue_5_deq_bits_store;
  wire         laneRequestSinkWire_5_bits_special = queue_5_deq_bits_special;
  wire         laneRequestSinkWire_5_bits_lsWholeReg = queue_5_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_5_bits_vs1 = queue_5_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_5_bits_vs2 = queue_5_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_5_bits_vd = queue_5_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_5_bits_loadStoreEEW = queue_5_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_5_bits_mask = queue_5_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_5_bits_segment = queue_5_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_5_bits_readFromScalar = queue_5_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_5_bits_csrInterface_vl = queue_5_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_5_bits_csrInterface_vStart = queue_5_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_5_bits_csrInterface_vlmul = queue_5_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_5_bits_csrInterface_vSew = queue_5_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_5_bits_csrInterface_vxrm = queue_5_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_5_bits_csrInterface_vta = queue_5_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_5_bits_csrInterface_vma = queue_5_deq_bits_csrInterface_vma;
  wire [1:0]   queue_5_enq_bits_csrInterface_vxrm;
  wire         queue_5_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi_15 = {queue_5_enq_bits_csrInterface_vxrm, queue_5_enq_bits_csrInterface_vta};
  wire         queue_5_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo_15 = {queue_dataIn_lo_hi_15, queue_5_enq_bits_csrInterface_vma};
  wire [2:0]   queue_5_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_5_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo_15 = {queue_5_enq_bits_csrInterface_vlmul, queue_5_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_5_enq_bits_csrInterface_vl;
  wire [11:0]  queue_5_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi_15 = {queue_5_enq_bits_csrInterface_vl, queue_5_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi_15 = {queue_dataIn_hi_hi_15, queue_dataIn_hi_lo_15};
  wire         queue_5_enq_bits_decodeResult_adder;
  wire         queue_5_enq_bits_decodeResult_logic;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo_5 = {queue_5_enq_bits_decodeResult_adder, queue_5_enq_bits_decodeResult_logic};
  wire         queue_5_enq_bits_decodeResult_divider;
  wire         queue_5_enq_bits_decodeResult_multiplier;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi_5 = {queue_5_enq_bits_decodeResult_divider, queue_5_enq_bits_decodeResult_multiplier};
  wire         queue_5_enq_bits_decodeResult_shift;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi_5 = {queue_dataIn_lo_lo_lo_hi_hi_5, queue_5_enq_bits_decodeResult_shift};
  wire [4:0]   queue_dataIn_lo_lo_lo_5 = {queue_dataIn_lo_lo_lo_hi_5, queue_dataIn_lo_lo_lo_lo_5};
  wire         queue_5_enq_bits_decodeResult_unsigned0;
  wire         queue_5_enq_bits_decodeResult_other;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi_5 = {queue_5_enq_bits_decodeResult_unsigned0, queue_5_enq_bits_decodeResult_other};
  wire         queue_5_enq_bits_decodeResult_multiCycle;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo_5 = {queue_dataIn_lo_lo_hi_lo_hi_5, queue_5_enq_bits_decodeResult_multiCycle};
  wire         queue_5_enq_bits_decodeResult_nr;
  wire         queue_5_enq_bits_decodeResult_itype;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi_5 = {queue_5_enq_bits_decodeResult_nr, queue_5_enq_bits_decodeResult_itype};
  wire         queue_5_enq_bits_decodeResult_unsigned1;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi_5 = {queue_dataIn_lo_lo_hi_hi_hi_5, queue_5_enq_bits_decodeResult_unsigned1};
  wire [5:0]   queue_dataIn_lo_lo_hi_10 = {queue_dataIn_lo_lo_hi_hi_5, queue_dataIn_lo_lo_hi_lo_5};
  wire [10:0]  queue_dataIn_lo_lo_10 = {queue_dataIn_lo_lo_hi_10, queue_dataIn_lo_lo_lo_5};
  wire         queue_5_enq_bits_decodeResult_widenReduce;
  wire         queue_5_enq_bits_decodeResult_red;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo_5 = {queue_5_enq_bits_decodeResult_widenReduce, queue_5_enq_bits_decodeResult_red};
  wire         queue_5_enq_bits_decodeResult_gather;
  wire         queue_5_enq_bits_decodeResult_slid;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi_5 = {queue_5_enq_bits_decodeResult_gather, queue_5_enq_bits_decodeResult_slid};
  wire         queue_5_enq_bits_decodeResult_targetRd;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi_5 = {queue_dataIn_lo_hi_lo_hi_hi_5, queue_5_enq_bits_decodeResult_targetRd};
  wire [4:0]   queue_dataIn_lo_hi_lo_10 = {queue_dataIn_lo_hi_lo_hi_5, queue_dataIn_lo_hi_lo_lo_5};
  wire         queue_5_enq_bits_decodeResult_unOrderWrite;
  wire         queue_5_enq_bits_decodeResult_compress;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi_5 = {queue_5_enq_bits_decodeResult_unOrderWrite, queue_5_enq_bits_decodeResult_compress};
  wire         queue_5_enq_bits_decodeResult_gather16;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo_5 = {queue_dataIn_lo_hi_hi_lo_hi_5, queue_5_enq_bits_decodeResult_gather16};
  wire         queue_5_enq_bits_decodeResult_iota;
  wire         queue_5_enq_bits_decodeResult_mv;
  wire [1:0]   queue_dataIn_lo_hi_hi_hi_hi_5 = {queue_5_enq_bits_decodeResult_iota, queue_5_enq_bits_decodeResult_mv};
  wire         queue_5_enq_bits_decodeResult_extend;
  wire [2:0]   queue_dataIn_lo_hi_hi_hi_5 = {queue_dataIn_lo_hi_hi_hi_hi_5, queue_5_enq_bits_decodeResult_extend};
  wire [5:0]   queue_dataIn_lo_hi_hi_10 = {queue_dataIn_lo_hi_hi_hi_5, queue_dataIn_lo_hi_hi_lo_5};
  wire [10:0]  queue_dataIn_lo_hi_16 = {queue_dataIn_lo_hi_hi_10, queue_dataIn_lo_hi_lo_10};
  wire [21:0]  queue_dataIn_lo_16 = {queue_dataIn_lo_hi_16, queue_dataIn_lo_lo_10};
  wire         queue_5_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_5_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_hi_lo_lo_lo_5 = {queue_5_enq_bits_decodeResult_maskLogic, queue_5_enq_bits_decodeResult_uop};
  wire         queue_5_enq_bits_decodeResult_readOnly;
  wire         queue_5_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi_5 = {queue_5_enq_bits_decodeResult_readOnly, queue_5_enq_bits_decodeResult_maskSource};
  wire         queue_5_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi_5 = {queue_dataIn_hi_lo_lo_hi_hi_5, queue_5_enq_bits_decodeResult_maskDestination};
  wire [7:0]   queue_dataIn_hi_lo_lo_10 = {queue_dataIn_hi_lo_lo_hi_5, queue_dataIn_hi_lo_lo_lo_5};
  wire         queue_5_enq_bits_decodeResult_special;
  wire         queue_5_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi_5 = {queue_5_enq_bits_decodeResult_special, queue_5_enq_bits_decodeResult_saturate};
  wire         queue_5_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo_5 = {queue_dataIn_hi_lo_hi_lo_hi_5, queue_5_enq_bits_decodeResult_vwmacc};
  wire         queue_5_enq_bits_decodeResult_crossRead;
  wire         queue_5_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi_5 = {queue_5_enq_bits_decodeResult_crossRead, queue_5_enq_bits_decodeResult_crossWrite};
  wire         queue_5_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi_5 = {queue_dataIn_hi_lo_hi_hi_hi_5, queue_5_enq_bits_decodeResult_maskUnit};
  wire [5:0]   queue_dataIn_hi_lo_hi_10 = {queue_dataIn_hi_lo_hi_hi_5, queue_dataIn_hi_lo_hi_lo_5};
  wire [13:0]  queue_dataIn_hi_lo_16 = {queue_dataIn_hi_lo_hi_10, queue_dataIn_hi_lo_lo_10};
  wire         queue_5_enq_bits_decodeResult_vtype;
  wire         queue_5_enq_bits_decodeResult_sWrite;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo_5 = {queue_5_enq_bits_decodeResult_vtype, queue_5_enq_bits_decodeResult_sWrite};
  wire         queue_5_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_5_enq_bits_decodeResult_scheduler;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi_5 = {queue_5_enq_bits_decodeResult_dontNeedExecuteInLane, queue_5_enq_bits_decodeResult_scheduler};
  wire         queue_5_enq_bits_decodeResult_sReadVD;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi_5 = {queue_dataIn_hi_hi_lo_hi_hi_5, queue_5_enq_bits_decodeResult_sReadVD};
  wire [4:0]   queue_dataIn_hi_hi_lo_10 = {queue_dataIn_hi_hi_lo_hi_5, queue_dataIn_hi_hi_lo_lo_5};
  wire         queue_5_enq_bits_decodeResult_ffo;
  wire         queue_5_enq_bits_decodeResult_average;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi_5 = {queue_5_enq_bits_decodeResult_ffo, queue_5_enq_bits_decodeResult_average};
  wire         queue_5_enq_bits_decodeResult_reverse;
  wire [2:0]   queue_dataIn_hi_hi_hi_lo_5 = {queue_dataIn_hi_hi_hi_lo_hi_5, queue_5_enq_bits_decodeResult_reverse};
  wire         queue_5_enq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_5_enq_bits_decodeResult_topUop;
  wire [5:0]   queue_dataIn_hi_hi_hi_hi_hi_5 = {queue_5_enq_bits_decodeResult_specialSlot, queue_5_enq_bits_decodeResult_topUop};
  wire         queue_5_enq_bits_decodeResult_popCount;
  wire [6:0]   queue_dataIn_hi_hi_hi_hi_5 = {queue_dataIn_hi_hi_hi_hi_hi_5, queue_5_enq_bits_decodeResult_popCount};
  wire [9:0]   queue_dataIn_hi_hi_hi_10 = {queue_dataIn_hi_hi_hi_hi_5, queue_dataIn_hi_hi_hi_lo_5};
  wire [14:0]  queue_dataIn_hi_hi_16 = {queue_dataIn_hi_hi_hi_10, queue_dataIn_hi_hi_lo_10};
  wire [28:0]  queue_dataIn_hi_16 = {queue_dataIn_hi_hi_16, queue_dataIn_hi_lo_16};
  wire [2:0]   queue_5_enq_bits_segment;
  wire [31:0]  queue_5_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_11 = {queue_5_enq_bits_segment, queue_5_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_11 = {queue_dataIn_lo_lo_hi_11, queue_dataIn_hi_15, queue_dataIn_lo_15};
  wire [1:0]   queue_5_enq_bits_loadStoreEEW;
  wire         queue_5_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_11 = {queue_5_enq_bits_loadStoreEEW, queue_5_enq_bits_mask};
  wire [4:0]   queue_5_enq_bits_vs2;
  wire [4:0]   queue_5_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_11 = {queue_5_enq_bits_vs2, queue_5_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_17 = {queue_dataIn_lo_hi_hi_11, queue_dataIn_lo_hi_lo_11};
  wire [80:0]  queue_dataIn_lo_17 = {queue_dataIn_lo_hi_17, queue_dataIn_lo_lo_11};
  wire         queue_5_enq_bits_lsWholeReg;
  wire [4:0]   queue_5_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_11 = {queue_5_enq_bits_lsWholeReg, queue_5_enq_bits_vs1};
  wire         queue_5_enq_bits_store;
  wire         queue_5_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_11 = {queue_5_enq_bits_store, queue_5_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_17 = {queue_dataIn_hi_lo_hi_11, queue_dataIn_hi_lo_lo_11};
  wire         queue_5_enq_bits_loadStore;
  wire         queue_5_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_11 = {queue_5_enq_bits_loadStore, queue_5_enq_bits_issueInst};
  wire [2:0]   queue_5_enq_bits_instructionIndex;
  wire [53:0]  queue_dataIn_hi_hi_hi_11 = {queue_5_enq_bits_instructionIndex, queue_dataIn_hi_16, queue_dataIn_lo_16};
  wire [55:0]  queue_dataIn_hi_hi_17 = {queue_dataIn_hi_hi_hi_11, queue_dataIn_hi_hi_lo_11};
  wire [63:0]  queue_dataIn_hi_17 = {queue_dataIn_hi_hi_17, queue_dataIn_hi_lo_17};
  wire [144:0] queue_dataIn_5 = {queue_dataIn_hi_17, queue_dataIn_lo_17};
  wire         queue_dataOut_5_csrInterface_vma = _queue_fifo_5_data_out[0];
  wire         queue_dataOut_5_csrInterface_vta = _queue_fifo_5_data_out[1];
  wire [1:0]   queue_dataOut_5_csrInterface_vxrm = _queue_fifo_5_data_out[3:2];
  wire [1:0]   queue_dataOut_5_csrInterface_vSew = _queue_fifo_5_data_out[5:4];
  wire [2:0]   queue_dataOut_5_csrInterface_vlmul = _queue_fifo_5_data_out[8:6];
  wire [11:0]  queue_dataOut_5_csrInterface_vStart = _queue_fifo_5_data_out[20:9];
  wire [11:0]  queue_dataOut_5_csrInterface_vl = _queue_fifo_5_data_out[32:21];
  wire [31:0]  queue_dataOut_5_readFromScalar = _queue_fifo_5_data_out[64:33];
  wire [2:0]   queue_dataOut_5_segment = _queue_fifo_5_data_out[67:65];
  wire         queue_dataOut_5_mask = _queue_fifo_5_data_out[68];
  wire [1:0]   queue_dataOut_5_loadStoreEEW = _queue_fifo_5_data_out[70:69];
  wire [4:0]   queue_dataOut_5_vd = _queue_fifo_5_data_out[75:71];
  wire [4:0]   queue_dataOut_5_vs2 = _queue_fifo_5_data_out[80:76];
  wire [4:0]   queue_dataOut_5_vs1 = _queue_fifo_5_data_out[85:81];
  wire         queue_dataOut_5_lsWholeReg = _queue_fifo_5_data_out[86];
  wire         queue_dataOut_5_special = _queue_fifo_5_data_out[87];
  wire         queue_dataOut_5_store = _queue_fifo_5_data_out[88];
  wire         queue_dataOut_5_issueInst = _queue_fifo_5_data_out[89];
  wire         queue_dataOut_5_loadStore = _queue_fifo_5_data_out[90];
  wire         queue_dataOut_5_decodeResult_logic = _queue_fifo_5_data_out[91];
  wire         queue_dataOut_5_decodeResult_adder = _queue_fifo_5_data_out[92];
  wire         queue_dataOut_5_decodeResult_shift = _queue_fifo_5_data_out[93];
  wire         queue_dataOut_5_decodeResult_multiplier = _queue_fifo_5_data_out[94];
  wire         queue_dataOut_5_decodeResult_divider = _queue_fifo_5_data_out[95];
  wire         queue_dataOut_5_decodeResult_multiCycle = _queue_fifo_5_data_out[96];
  wire         queue_dataOut_5_decodeResult_other = _queue_fifo_5_data_out[97];
  wire         queue_dataOut_5_decodeResult_unsigned0 = _queue_fifo_5_data_out[98];
  wire         queue_dataOut_5_decodeResult_unsigned1 = _queue_fifo_5_data_out[99];
  wire         queue_dataOut_5_decodeResult_itype = _queue_fifo_5_data_out[100];
  wire         queue_dataOut_5_decodeResult_nr = _queue_fifo_5_data_out[101];
  wire         queue_dataOut_5_decodeResult_red = _queue_fifo_5_data_out[102];
  wire         queue_dataOut_5_decodeResult_widenReduce = _queue_fifo_5_data_out[103];
  wire         queue_dataOut_5_decodeResult_targetRd = _queue_fifo_5_data_out[104];
  wire         queue_dataOut_5_decodeResult_slid = _queue_fifo_5_data_out[105];
  wire         queue_dataOut_5_decodeResult_gather = _queue_fifo_5_data_out[106];
  wire         queue_dataOut_5_decodeResult_gather16 = _queue_fifo_5_data_out[107];
  wire         queue_dataOut_5_decodeResult_compress = _queue_fifo_5_data_out[108];
  wire         queue_dataOut_5_decodeResult_unOrderWrite = _queue_fifo_5_data_out[109];
  wire         queue_dataOut_5_decodeResult_extend = _queue_fifo_5_data_out[110];
  wire         queue_dataOut_5_decodeResult_mv = _queue_fifo_5_data_out[111];
  wire         queue_dataOut_5_decodeResult_iota = _queue_fifo_5_data_out[112];
  wire [3:0]   queue_dataOut_5_decodeResult_uop = _queue_fifo_5_data_out[116:113];
  wire         queue_dataOut_5_decodeResult_maskLogic = _queue_fifo_5_data_out[117];
  wire         queue_dataOut_5_decodeResult_maskDestination = _queue_fifo_5_data_out[118];
  wire         queue_dataOut_5_decodeResult_maskSource = _queue_fifo_5_data_out[119];
  wire         queue_dataOut_5_decodeResult_readOnly = _queue_fifo_5_data_out[120];
  wire         queue_dataOut_5_decodeResult_vwmacc = _queue_fifo_5_data_out[121];
  wire         queue_dataOut_5_decodeResult_saturate = _queue_fifo_5_data_out[122];
  wire         queue_dataOut_5_decodeResult_special = _queue_fifo_5_data_out[123];
  wire         queue_dataOut_5_decodeResult_maskUnit = _queue_fifo_5_data_out[124];
  wire         queue_dataOut_5_decodeResult_crossWrite = _queue_fifo_5_data_out[125];
  wire         queue_dataOut_5_decodeResult_crossRead = _queue_fifo_5_data_out[126];
  wire         queue_dataOut_5_decodeResult_sWrite = _queue_fifo_5_data_out[127];
  wire         queue_dataOut_5_decodeResult_vtype = _queue_fifo_5_data_out[128];
  wire         queue_dataOut_5_decodeResult_sReadVD = _queue_fifo_5_data_out[129];
  wire         queue_dataOut_5_decodeResult_scheduler = _queue_fifo_5_data_out[130];
  wire         queue_dataOut_5_decodeResult_dontNeedExecuteInLane = _queue_fifo_5_data_out[131];
  wire         queue_dataOut_5_decodeResult_reverse = _queue_fifo_5_data_out[132];
  wire         queue_dataOut_5_decodeResult_average = _queue_fifo_5_data_out[133];
  wire         queue_dataOut_5_decodeResult_ffo = _queue_fifo_5_data_out[134];
  wire         queue_dataOut_5_decodeResult_popCount = _queue_fifo_5_data_out[135];
  wire [4:0]   queue_dataOut_5_decodeResult_topUop = _queue_fifo_5_data_out[140:136];
  wire         queue_dataOut_5_decodeResult_specialSlot = _queue_fifo_5_data_out[141];
  wire [2:0]   queue_dataOut_5_instructionIndex = _queue_fifo_5_data_out[144:142];
  wire         queue_5_enq_ready = ~_queue_fifo_5_full;
  wire         queue_5_enq_valid;
  assign queue_5_deq_valid = ~_queue_fifo_5_empty | queue_5_enq_valid;
  assign queue_5_deq_bits_instructionIndex = _queue_fifo_5_empty ? queue_5_enq_bits_instructionIndex : queue_dataOut_5_instructionIndex;
  assign queue_5_deq_bits_decodeResult_specialSlot = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_specialSlot : queue_dataOut_5_decodeResult_specialSlot;
  assign queue_5_deq_bits_decodeResult_topUop = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_topUop : queue_dataOut_5_decodeResult_topUop;
  assign queue_5_deq_bits_decodeResult_popCount = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_popCount : queue_dataOut_5_decodeResult_popCount;
  assign queue_5_deq_bits_decodeResult_ffo = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_ffo : queue_dataOut_5_decodeResult_ffo;
  assign queue_5_deq_bits_decodeResult_average = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_average : queue_dataOut_5_decodeResult_average;
  assign queue_5_deq_bits_decodeResult_reverse = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_reverse : queue_dataOut_5_decodeResult_reverse;
  assign queue_5_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_5_decodeResult_dontNeedExecuteInLane;
  assign queue_5_deq_bits_decodeResult_scheduler = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_scheduler : queue_dataOut_5_decodeResult_scheduler;
  assign queue_5_deq_bits_decodeResult_sReadVD = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_sReadVD : queue_dataOut_5_decodeResult_sReadVD;
  assign queue_5_deq_bits_decodeResult_vtype = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_vtype : queue_dataOut_5_decodeResult_vtype;
  assign queue_5_deq_bits_decodeResult_sWrite = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_sWrite : queue_dataOut_5_decodeResult_sWrite;
  assign queue_5_deq_bits_decodeResult_crossRead = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_crossRead : queue_dataOut_5_decodeResult_crossRead;
  assign queue_5_deq_bits_decodeResult_crossWrite = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_crossWrite : queue_dataOut_5_decodeResult_crossWrite;
  assign queue_5_deq_bits_decodeResult_maskUnit = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_maskUnit : queue_dataOut_5_decodeResult_maskUnit;
  assign queue_5_deq_bits_decodeResult_special = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_special : queue_dataOut_5_decodeResult_special;
  assign queue_5_deq_bits_decodeResult_saturate = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_saturate : queue_dataOut_5_decodeResult_saturate;
  assign queue_5_deq_bits_decodeResult_vwmacc = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_vwmacc : queue_dataOut_5_decodeResult_vwmacc;
  assign queue_5_deq_bits_decodeResult_readOnly = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_readOnly : queue_dataOut_5_decodeResult_readOnly;
  assign queue_5_deq_bits_decodeResult_maskSource = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_maskSource : queue_dataOut_5_decodeResult_maskSource;
  assign queue_5_deq_bits_decodeResult_maskDestination = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_maskDestination : queue_dataOut_5_decodeResult_maskDestination;
  assign queue_5_deq_bits_decodeResult_maskLogic = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_maskLogic : queue_dataOut_5_decodeResult_maskLogic;
  assign queue_5_deq_bits_decodeResult_uop = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_uop : queue_dataOut_5_decodeResult_uop;
  assign queue_5_deq_bits_decodeResult_iota = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_iota : queue_dataOut_5_decodeResult_iota;
  assign queue_5_deq_bits_decodeResult_mv = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_mv : queue_dataOut_5_decodeResult_mv;
  assign queue_5_deq_bits_decodeResult_extend = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_extend : queue_dataOut_5_decodeResult_extend;
  assign queue_5_deq_bits_decodeResult_unOrderWrite = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_unOrderWrite : queue_dataOut_5_decodeResult_unOrderWrite;
  assign queue_5_deq_bits_decodeResult_compress = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_compress : queue_dataOut_5_decodeResult_compress;
  assign queue_5_deq_bits_decodeResult_gather16 = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_gather16 : queue_dataOut_5_decodeResult_gather16;
  assign queue_5_deq_bits_decodeResult_gather = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_gather : queue_dataOut_5_decodeResult_gather;
  assign queue_5_deq_bits_decodeResult_slid = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_slid : queue_dataOut_5_decodeResult_slid;
  assign queue_5_deq_bits_decodeResult_targetRd = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_targetRd : queue_dataOut_5_decodeResult_targetRd;
  assign queue_5_deq_bits_decodeResult_widenReduce = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_widenReduce : queue_dataOut_5_decodeResult_widenReduce;
  assign queue_5_deq_bits_decodeResult_red = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_red : queue_dataOut_5_decodeResult_red;
  assign queue_5_deq_bits_decodeResult_nr = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_nr : queue_dataOut_5_decodeResult_nr;
  assign queue_5_deq_bits_decodeResult_itype = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_itype : queue_dataOut_5_decodeResult_itype;
  assign queue_5_deq_bits_decodeResult_unsigned1 = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_unsigned1 : queue_dataOut_5_decodeResult_unsigned1;
  assign queue_5_deq_bits_decodeResult_unsigned0 = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_unsigned0 : queue_dataOut_5_decodeResult_unsigned0;
  assign queue_5_deq_bits_decodeResult_other = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_other : queue_dataOut_5_decodeResult_other;
  assign queue_5_deq_bits_decodeResult_multiCycle = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_multiCycle : queue_dataOut_5_decodeResult_multiCycle;
  assign queue_5_deq_bits_decodeResult_divider = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_divider : queue_dataOut_5_decodeResult_divider;
  assign queue_5_deq_bits_decodeResult_multiplier = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_multiplier : queue_dataOut_5_decodeResult_multiplier;
  assign queue_5_deq_bits_decodeResult_shift = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_shift : queue_dataOut_5_decodeResult_shift;
  assign queue_5_deq_bits_decodeResult_adder = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_adder : queue_dataOut_5_decodeResult_adder;
  assign queue_5_deq_bits_decodeResult_logic = _queue_fifo_5_empty ? queue_5_enq_bits_decodeResult_logic : queue_dataOut_5_decodeResult_logic;
  assign queue_5_deq_bits_loadStore = _queue_fifo_5_empty ? queue_5_enq_bits_loadStore : queue_dataOut_5_loadStore;
  assign queue_5_deq_bits_issueInst = _queue_fifo_5_empty ? queue_5_enq_bits_issueInst : queue_dataOut_5_issueInst;
  assign queue_5_deq_bits_store = _queue_fifo_5_empty ? queue_5_enq_bits_store : queue_dataOut_5_store;
  assign queue_5_deq_bits_special = _queue_fifo_5_empty ? queue_5_enq_bits_special : queue_dataOut_5_special;
  assign queue_5_deq_bits_lsWholeReg = _queue_fifo_5_empty ? queue_5_enq_bits_lsWholeReg : queue_dataOut_5_lsWholeReg;
  assign queue_5_deq_bits_vs1 = _queue_fifo_5_empty ? queue_5_enq_bits_vs1 : queue_dataOut_5_vs1;
  assign queue_5_deq_bits_vs2 = _queue_fifo_5_empty ? queue_5_enq_bits_vs2 : queue_dataOut_5_vs2;
  assign queue_5_deq_bits_vd = _queue_fifo_5_empty ? queue_5_enq_bits_vd : queue_dataOut_5_vd;
  assign queue_5_deq_bits_loadStoreEEW = _queue_fifo_5_empty ? queue_5_enq_bits_loadStoreEEW : queue_dataOut_5_loadStoreEEW;
  assign queue_5_deq_bits_mask = _queue_fifo_5_empty ? queue_5_enq_bits_mask : queue_dataOut_5_mask;
  assign queue_5_deq_bits_segment = _queue_fifo_5_empty ? queue_5_enq_bits_segment : queue_dataOut_5_segment;
  assign queue_5_deq_bits_readFromScalar = _queue_fifo_5_empty ? queue_5_enq_bits_readFromScalar : queue_dataOut_5_readFromScalar;
  assign queue_5_deq_bits_csrInterface_vl = _queue_fifo_5_empty ? queue_5_enq_bits_csrInterface_vl : queue_dataOut_5_csrInterface_vl;
  assign queue_5_deq_bits_csrInterface_vStart = _queue_fifo_5_empty ? queue_5_enq_bits_csrInterface_vStart : queue_dataOut_5_csrInterface_vStart;
  assign queue_5_deq_bits_csrInterface_vlmul = _queue_fifo_5_empty ? queue_5_enq_bits_csrInterface_vlmul : queue_dataOut_5_csrInterface_vlmul;
  assign queue_5_deq_bits_csrInterface_vSew = _queue_fifo_5_empty ? queue_5_enq_bits_csrInterface_vSew : queue_dataOut_5_csrInterface_vSew;
  assign queue_5_deq_bits_csrInterface_vxrm = _queue_fifo_5_empty ? queue_5_enq_bits_csrInterface_vxrm : queue_dataOut_5_csrInterface_vxrm;
  assign queue_5_deq_bits_csrInterface_vta = _queue_fifo_5_empty ? queue_5_enq_bits_csrInterface_vta : queue_dataOut_5_csrInterface_vta;
  assign queue_5_deq_bits_csrInterface_vma = _queue_fifo_5_empty ? queue_5_enq_bits_csrInterface_vma : queue_dataOut_5_csrInterface_vma;
  wire         laneVec_5_laneRequest_bits_issueInst = laneRequestSinkWire_5_ready & laneRequestSinkWire_5_valid;
  reg          releasePipe_pipe_v_5;
  wire         releasePipe_pipe_out_5_valid = releasePipe_pipe_v_5;
  wire         laneRequestSourceWire_5_ready;
  wire         validSource_5_valid = laneRequestSourceWire_5_ready & laneRequestSourceWire_5_valid;
  reg  [2:0]   tokenCheck_counter_5;
  wire [2:0]   tokenCheck_counterChange_5 = validSource_5_valid ? 3'h1 : 3'h7;
  assign tokenCheck_5 = ~(tokenCheck_counter_5[2]);
  assign laneRequestSourceWire_5_ready = tokenCheck_5;
  assign queue_5_enq_valid = validSink_5_valid;
  assign queue_5_enq_bits_instructionIndex = validSink_5_bits_instructionIndex;
  assign queue_5_enq_bits_decodeResult_specialSlot = validSink_5_bits_decodeResult_specialSlot;
  assign queue_5_enq_bits_decodeResult_topUop = validSink_5_bits_decodeResult_topUop;
  assign queue_5_enq_bits_decodeResult_popCount = validSink_5_bits_decodeResult_popCount;
  assign queue_5_enq_bits_decodeResult_ffo = validSink_5_bits_decodeResult_ffo;
  assign queue_5_enq_bits_decodeResult_average = validSink_5_bits_decodeResult_average;
  assign queue_5_enq_bits_decodeResult_reverse = validSink_5_bits_decodeResult_reverse;
  assign queue_5_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_5_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_5_enq_bits_decodeResult_scheduler = validSink_5_bits_decodeResult_scheduler;
  assign queue_5_enq_bits_decodeResult_sReadVD = validSink_5_bits_decodeResult_sReadVD;
  assign queue_5_enq_bits_decodeResult_vtype = validSink_5_bits_decodeResult_vtype;
  assign queue_5_enq_bits_decodeResult_sWrite = validSink_5_bits_decodeResult_sWrite;
  assign queue_5_enq_bits_decodeResult_crossRead = validSink_5_bits_decodeResult_crossRead;
  assign queue_5_enq_bits_decodeResult_crossWrite = validSink_5_bits_decodeResult_crossWrite;
  assign queue_5_enq_bits_decodeResult_maskUnit = validSink_5_bits_decodeResult_maskUnit;
  assign queue_5_enq_bits_decodeResult_special = validSink_5_bits_decodeResult_special;
  assign queue_5_enq_bits_decodeResult_saturate = validSink_5_bits_decodeResult_saturate;
  assign queue_5_enq_bits_decodeResult_vwmacc = validSink_5_bits_decodeResult_vwmacc;
  assign queue_5_enq_bits_decodeResult_readOnly = validSink_5_bits_decodeResult_readOnly;
  assign queue_5_enq_bits_decodeResult_maskSource = validSink_5_bits_decodeResult_maskSource;
  assign queue_5_enq_bits_decodeResult_maskDestination = validSink_5_bits_decodeResult_maskDestination;
  assign queue_5_enq_bits_decodeResult_maskLogic = validSink_5_bits_decodeResult_maskLogic;
  assign queue_5_enq_bits_decodeResult_uop = validSink_5_bits_decodeResult_uop;
  assign queue_5_enq_bits_decodeResult_iota = validSink_5_bits_decodeResult_iota;
  assign queue_5_enq_bits_decodeResult_mv = validSink_5_bits_decodeResult_mv;
  assign queue_5_enq_bits_decodeResult_extend = validSink_5_bits_decodeResult_extend;
  assign queue_5_enq_bits_decodeResult_unOrderWrite = validSink_5_bits_decodeResult_unOrderWrite;
  assign queue_5_enq_bits_decodeResult_compress = validSink_5_bits_decodeResult_compress;
  assign queue_5_enq_bits_decodeResult_gather16 = validSink_5_bits_decodeResult_gather16;
  assign queue_5_enq_bits_decodeResult_gather = validSink_5_bits_decodeResult_gather;
  assign queue_5_enq_bits_decodeResult_slid = validSink_5_bits_decodeResult_slid;
  assign queue_5_enq_bits_decodeResult_targetRd = validSink_5_bits_decodeResult_targetRd;
  assign queue_5_enq_bits_decodeResult_widenReduce = validSink_5_bits_decodeResult_widenReduce;
  assign queue_5_enq_bits_decodeResult_red = validSink_5_bits_decodeResult_red;
  assign queue_5_enq_bits_decodeResult_nr = validSink_5_bits_decodeResult_nr;
  assign queue_5_enq_bits_decodeResult_itype = validSink_5_bits_decodeResult_itype;
  assign queue_5_enq_bits_decodeResult_unsigned1 = validSink_5_bits_decodeResult_unsigned1;
  assign queue_5_enq_bits_decodeResult_unsigned0 = validSink_5_bits_decodeResult_unsigned0;
  assign queue_5_enq_bits_decodeResult_other = validSink_5_bits_decodeResult_other;
  assign queue_5_enq_bits_decodeResult_multiCycle = validSink_5_bits_decodeResult_multiCycle;
  assign queue_5_enq_bits_decodeResult_divider = validSink_5_bits_decodeResult_divider;
  assign queue_5_enq_bits_decodeResult_multiplier = validSink_5_bits_decodeResult_multiplier;
  assign queue_5_enq_bits_decodeResult_shift = validSink_5_bits_decodeResult_shift;
  assign queue_5_enq_bits_decodeResult_adder = validSink_5_bits_decodeResult_adder;
  assign queue_5_enq_bits_decodeResult_logic = validSink_5_bits_decodeResult_logic;
  assign queue_5_enq_bits_loadStore = validSink_5_bits_loadStore;
  assign queue_5_enq_bits_issueInst = validSink_5_bits_issueInst;
  assign queue_5_enq_bits_store = validSink_5_bits_store;
  assign queue_5_enq_bits_special = validSink_5_bits_special;
  assign queue_5_enq_bits_lsWholeReg = validSink_5_bits_lsWholeReg;
  assign queue_5_enq_bits_vs1 = validSink_5_bits_vs1;
  assign queue_5_enq_bits_vs2 = validSink_5_bits_vs2;
  assign queue_5_enq_bits_vd = validSink_5_bits_vd;
  assign queue_5_enq_bits_loadStoreEEW = validSink_5_bits_loadStoreEEW;
  assign queue_5_enq_bits_mask = validSink_5_bits_mask;
  assign queue_5_enq_bits_segment = validSink_5_bits_segment;
  assign queue_5_enq_bits_readFromScalar = validSink_5_bits_readFromScalar;
  assign queue_5_enq_bits_csrInterface_vl = validSink_5_bits_csrInterface_vl;
  assign queue_5_enq_bits_csrInterface_vStart = validSink_5_bits_csrInterface_vStart;
  assign queue_5_enq_bits_csrInterface_vlmul = validSink_5_bits_csrInterface_vlmul;
  assign queue_5_enq_bits_csrInterface_vSew = validSink_5_bits_csrInterface_vSew;
  assign queue_5_enq_bits_csrInterface_vxrm = validSink_5_bits_csrInterface_vxrm;
  assign queue_5_enq_bits_csrInterface_vta = validSink_5_bits_csrInterface_vta;
  assign queue_5_enq_bits_csrInterface_vma = validSink_5_bits_csrInterface_vma;
  reg          shifterReg_5_0_valid;
  assign validSink_5_valid = shifterReg_5_0_valid;
  reg  [2:0]   shifterReg_5_0_bits_instructionIndex;
  assign validSink_5_bits_instructionIndex = shifterReg_5_0_bits_instructionIndex;
  reg          shifterReg_5_0_bits_decodeResult_specialSlot;
  assign validSink_5_bits_decodeResult_specialSlot = shifterReg_5_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_5_0_bits_decodeResult_topUop;
  assign validSink_5_bits_decodeResult_topUop = shifterReg_5_0_bits_decodeResult_topUop;
  reg          shifterReg_5_0_bits_decodeResult_popCount;
  assign validSink_5_bits_decodeResult_popCount = shifterReg_5_0_bits_decodeResult_popCount;
  reg          shifterReg_5_0_bits_decodeResult_ffo;
  assign validSink_5_bits_decodeResult_ffo = shifterReg_5_0_bits_decodeResult_ffo;
  reg          shifterReg_5_0_bits_decodeResult_average;
  assign validSink_5_bits_decodeResult_average = shifterReg_5_0_bits_decodeResult_average;
  reg          shifterReg_5_0_bits_decodeResult_reverse;
  assign validSink_5_bits_decodeResult_reverse = shifterReg_5_0_bits_decodeResult_reverse;
  reg          shifterReg_5_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_5_bits_decodeResult_dontNeedExecuteInLane = shifterReg_5_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_5_0_bits_decodeResult_scheduler;
  assign validSink_5_bits_decodeResult_scheduler = shifterReg_5_0_bits_decodeResult_scheduler;
  reg          shifterReg_5_0_bits_decodeResult_sReadVD;
  assign validSink_5_bits_decodeResult_sReadVD = shifterReg_5_0_bits_decodeResult_sReadVD;
  reg          shifterReg_5_0_bits_decodeResult_vtype;
  assign validSink_5_bits_decodeResult_vtype = shifterReg_5_0_bits_decodeResult_vtype;
  reg          shifterReg_5_0_bits_decodeResult_sWrite;
  assign validSink_5_bits_decodeResult_sWrite = shifterReg_5_0_bits_decodeResult_sWrite;
  reg          shifterReg_5_0_bits_decodeResult_crossRead;
  assign validSink_5_bits_decodeResult_crossRead = shifterReg_5_0_bits_decodeResult_crossRead;
  reg          shifterReg_5_0_bits_decodeResult_crossWrite;
  assign validSink_5_bits_decodeResult_crossWrite = shifterReg_5_0_bits_decodeResult_crossWrite;
  reg          shifterReg_5_0_bits_decodeResult_maskUnit;
  assign validSink_5_bits_decodeResult_maskUnit = shifterReg_5_0_bits_decodeResult_maskUnit;
  reg          shifterReg_5_0_bits_decodeResult_special;
  assign validSink_5_bits_decodeResult_special = shifterReg_5_0_bits_decodeResult_special;
  reg          shifterReg_5_0_bits_decodeResult_saturate;
  assign validSink_5_bits_decodeResult_saturate = shifterReg_5_0_bits_decodeResult_saturate;
  reg          shifterReg_5_0_bits_decodeResult_vwmacc;
  assign validSink_5_bits_decodeResult_vwmacc = shifterReg_5_0_bits_decodeResult_vwmacc;
  reg          shifterReg_5_0_bits_decodeResult_readOnly;
  assign validSink_5_bits_decodeResult_readOnly = shifterReg_5_0_bits_decodeResult_readOnly;
  reg          shifterReg_5_0_bits_decodeResult_maskSource;
  assign validSink_5_bits_decodeResult_maskSource = shifterReg_5_0_bits_decodeResult_maskSource;
  reg          shifterReg_5_0_bits_decodeResult_maskDestination;
  assign validSink_5_bits_decodeResult_maskDestination = shifterReg_5_0_bits_decodeResult_maskDestination;
  reg          shifterReg_5_0_bits_decodeResult_maskLogic;
  assign validSink_5_bits_decodeResult_maskLogic = shifterReg_5_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_5_0_bits_decodeResult_uop;
  assign validSink_5_bits_decodeResult_uop = shifterReg_5_0_bits_decodeResult_uop;
  reg          shifterReg_5_0_bits_decodeResult_iota;
  assign validSink_5_bits_decodeResult_iota = shifterReg_5_0_bits_decodeResult_iota;
  reg          shifterReg_5_0_bits_decodeResult_mv;
  assign validSink_5_bits_decodeResult_mv = shifterReg_5_0_bits_decodeResult_mv;
  reg          shifterReg_5_0_bits_decodeResult_extend;
  assign validSink_5_bits_decodeResult_extend = shifterReg_5_0_bits_decodeResult_extend;
  reg          shifterReg_5_0_bits_decodeResult_unOrderWrite;
  assign validSink_5_bits_decodeResult_unOrderWrite = shifterReg_5_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_5_0_bits_decodeResult_compress;
  assign validSink_5_bits_decodeResult_compress = shifterReg_5_0_bits_decodeResult_compress;
  reg          shifterReg_5_0_bits_decodeResult_gather16;
  assign validSink_5_bits_decodeResult_gather16 = shifterReg_5_0_bits_decodeResult_gather16;
  reg          shifterReg_5_0_bits_decodeResult_gather;
  assign validSink_5_bits_decodeResult_gather = shifterReg_5_0_bits_decodeResult_gather;
  reg          shifterReg_5_0_bits_decodeResult_slid;
  assign validSink_5_bits_decodeResult_slid = shifterReg_5_0_bits_decodeResult_slid;
  reg          shifterReg_5_0_bits_decodeResult_targetRd;
  assign validSink_5_bits_decodeResult_targetRd = shifterReg_5_0_bits_decodeResult_targetRd;
  reg          shifterReg_5_0_bits_decodeResult_widenReduce;
  assign validSink_5_bits_decodeResult_widenReduce = shifterReg_5_0_bits_decodeResult_widenReduce;
  reg          shifterReg_5_0_bits_decodeResult_red;
  assign validSink_5_bits_decodeResult_red = shifterReg_5_0_bits_decodeResult_red;
  reg          shifterReg_5_0_bits_decodeResult_nr;
  assign validSink_5_bits_decodeResult_nr = shifterReg_5_0_bits_decodeResult_nr;
  reg          shifterReg_5_0_bits_decodeResult_itype;
  assign validSink_5_bits_decodeResult_itype = shifterReg_5_0_bits_decodeResult_itype;
  reg          shifterReg_5_0_bits_decodeResult_unsigned1;
  assign validSink_5_bits_decodeResult_unsigned1 = shifterReg_5_0_bits_decodeResult_unsigned1;
  reg          shifterReg_5_0_bits_decodeResult_unsigned0;
  assign validSink_5_bits_decodeResult_unsigned0 = shifterReg_5_0_bits_decodeResult_unsigned0;
  reg          shifterReg_5_0_bits_decodeResult_other;
  assign validSink_5_bits_decodeResult_other = shifterReg_5_0_bits_decodeResult_other;
  reg          shifterReg_5_0_bits_decodeResult_multiCycle;
  assign validSink_5_bits_decodeResult_multiCycle = shifterReg_5_0_bits_decodeResult_multiCycle;
  reg          shifterReg_5_0_bits_decodeResult_divider;
  assign validSink_5_bits_decodeResult_divider = shifterReg_5_0_bits_decodeResult_divider;
  reg          shifterReg_5_0_bits_decodeResult_multiplier;
  assign validSink_5_bits_decodeResult_multiplier = shifterReg_5_0_bits_decodeResult_multiplier;
  reg          shifterReg_5_0_bits_decodeResult_shift;
  assign validSink_5_bits_decodeResult_shift = shifterReg_5_0_bits_decodeResult_shift;
  reg          shifterReg_5_0_bits_decodeResult_adder;
  assign validSink_5_bits_decodeResult_adder = shifterReg_5_0_bits_decodeResult_adder;
  reg          shifterReg_5_0_bits_decodeResult_logic;
  assign validSink_5_bits_decodeResult_logic = shifterReg_5_0_bits_decodeResult_logic;
  reg          shifterReg_5_0_bits_loadStore;
  assign validSink_5_bits_loadStore = shifterReg_5_0_bits_loadStore;
  reg          shifterReg_5_0_bits_issueInst;
  assign validSink_5_bits_issueInst = shifterReg_5_0_bits_issueInst;
  reg          shifterReg_5_0_bits_store;
  assign validSink_5_bits_store = shifterReg_5_0_bits_store;
  reg          shifterReg_5_0_bits_special;
  assign validSink_5_bits_special = shifterReg_5_0_bits_special;
  reg          shifterReg_5_0_bits_lsWholeReg;
  assign validSink_5_bits_lsWholeReg = shifterReg_5_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_5_0_bits_vs1;
  assign validSink_5_bits_vs1 = shifterReg_5_0_bits_vs1;
  reg  [4:0]   shifterReg_5_0_bits_vs2;
  assign validSink_5_bits_vs2 = shifterReg_5_0_bits_vs2;
  reg  [4:0]   shifterReg_5_0_bits_vd;
  assign validSink_5_bits_vd = shifterReg_5_0_bits_vd;
  reg  [1:0]   shifterReg_5_0_bits_loadStoreEEW;
  assign validSink_5_bits_loadStoreEEW = shifterReg_5_0_bits_loadStoreEEW;
  reg          shifterReg_5_0_bits_mask;
  assign validSink_5_bits_mask = shifterReg_5_0_bits_mask;
  reg  [2:0]   shifterReg_5_0_bits_segment;
  assign validSink_5_bits_segment = shifterReg_5_0_bits_segment;
  reg  [31:0]  shifterReg_5_0_bits_readFromScalar;
  assign validSink_5_bits_readFromScalar = shifterReg_5_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_5_0_bits_csrInterface_vl;
  assign validSink_5_bits_csrInterface_vl = shifterReg_5_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_5_0_bits_csrInterface_vStart;
  assign validSink_5_bits_csrInterface_vStart = shifterReg_5_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_5_0_bits_csrInterface_vlmul;
  assign validSink_5_bits_csrInterface_vlmul = shifterReg_5_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_5_0_bits_csrInterface_vSew;
  assign validSink_5_bits_csrInterface_vSew = shifterReg_5_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_5_0_bits_csrInterface_vxrm;
  assign validSink_5_bits_csrInterface_vxrm = shifterReg_5_0_bits_csrInterface_vxrm;
  reg          shifterReg_5_0_bits_csrInterface_vta;
  assign validSink_5_bits_csrInterface_vta = shifterReg_5_0_bits_csrInterface_vta;
  reg          shifterReg_5_0_bits_csrInterface_vma;
  assign validSink_5_bits_csrInterface_vma = shifterReg_5_0_bits_csrInterface_vma;
  wire         shifterValid_5 = shifterReg_5_0_valid | validSource_5_valid;
  wire         validSink_6_valid;
  wire [2:0]   validSink_6_bits_instructionIndex;
  wire         validSink_6_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_6_bits_decodeResult_topUop;
  wire         validSink_6_bits_decodeResult_popCount;
  wire         validSink_6_bits_decodeResult_ffo;
  wire         validSink_6_bits_decodeResult_average;
  wire         validSink_6_bits_decodeResult_reverse;
  wire         validSink_6_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_6_bits_decodeResult_scheduler;
  wire         validSink_6_bits_decodeResult_sReadVD;
  wire         validSink_6_bits_decodeResult_vtype;
  wire         validSink_6_bits_decodeResult_sWrite;
  wire         validSink_6_bits_decodeResult_crossRead;
  wire         validSink_6_bits_decodeResult_crossWrite;
  wire         validSink_6_bits_decodeResult_maskUnit;
  wire         validSink_6_bits_decodeResult_special;
  wire         validSink_6_bits_decodeResult_saturate;
  wire         validSink_6_bits_decodeResult_vwmacc;
  wire         validSink_6_bits_decodeResult_readOnly;
  wire         validSink_6_bits_decodeResult_maskSource;
  wire         validSink_6_bits_decodeResult_maskDestination;
  wire         validSink_6_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_6_bits_decodeResult_uop;
  wire         validSink_6_bits_decodeResult_iota;
  wire         validSink_6_bits_decodeResult_mv;
  wire         validSink_6_bits_decodeResult_extend;
  wire         validSink_6_bits_decodeResult_unOrderWrite;
  wire         validSink_6_bits_decodeResult_compress;
  wire         validSink_6_bits_decodeResult_gather16;
  wire         validSink_6_bits_decodeResult_gather;
  wire         validSink_6_bits_decodeResult_slid;
  wire         validSink_6_bits_decodeResult_targetRd;
  wire         validSink_6_bits_decodeResult_widenReduce;
  wire         validSink_6_bits_decodeResult_red;
  wire         validSink_6_bits_decodeResult_nr;
  wire         validSink_6_bits_decodeResult_itype;
  wire         validSink_6_bits_decodeResult_unsigned1;
  wire         validSink_6_bits_decodeResult_unsigned0;
  wire         validSink_6_bits_decodeResult_other;
  wire         validSink_6_bits_decodeResult_multiCycle;
  wire         validSink_6_bits_decodeResult_divider;
  wire         validSink_6_bits_decodeResult_multiplier;
  wire         validSink_6_bits_decodeResult_shift;
  wire         validSink_6_bits_decodeResult_adder;
  wire         validSink_6_bits_decodeResult_logic;
  wire         validSink_6_bits_loadStore;
  wire         validSink_6_bits_issueInst;
  wire         validSink_6_bits_store;
  wire         validSink_6_bits_special;
  wire         validSink_6_bits_lsWholeReg;
  wire [4:0]   validSink_6_bits_vs1;
  wire [4:0]   validSink_6_bits_vs2;
  wire [4:0]   validSink_6_bits_vd;
  wire [1:0]   validSink_6_bits_loadStoreEEW;
  wire         validSink_6_bits_mask;
  wire [2:0]   validSink_6_bits_segment;
  wire [31:0]  validSink_6_bits_readFromScalar;
  wire [11:0]  validSink_6_bits_csrInterface_vl;
  wire [11:0]  validSink_6_bits_csrInterface_vStart;
  wire [2:0]   validSink_6_bits_csrInterface_vlmul;
  wire [1:0]   validSink_6_bits_csrInterface_vSew;
  wire [1:0]   validSink_6_bits_csrInterface_vxrm;
  wire         validSink_6_bits_csrInterface_vta;
  wire         validSink_6_bits_csrInterface_vma;
  wire         laneRequestSinkWire_6_valid = queue_6_deq_valid;
  wire [2:0]   laneRequestSinkWire_6_bits_instructionIndex = queue_6_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_6_bits_decodeResult_specialSlot = queue_6_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_6_bits_decodeResult_topUop = queue_6_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_6_bits_decodeResult_popCount = queue_6_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_6_bits_decodeResult_ffo = queue_6_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_6_bits_decodeResult_average = queue_6_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_6_bits_decodeResult_reverse = queue_6_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_6_bits_decodeResult_dontNeedExecuteInLane = queue_6_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_6_bits_decodeResult_scheduler = queue_6_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_6_bits_decodeResult_sReadVD = queue_6_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_6_bits_decodeResult_vtype = queue_6_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_6_bits_decodeResult_sWrite = queue_6_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_6_bits_decodeResult_crossRead = queue_6_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_6_bits_decodeResult_crossWrite = queue_6_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_6_bits_decodeResult_maskUnit = queue_6_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_6_bits_decodeResult_special = queue_6_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_6_bits_decodeResult_saturate = queue_6_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_6_bits_decodeResult_vwmacc = queue_6_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_6_bits_decodeResult_readOnly = queue_6_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_6_bits_decodeResult_maskSource = queue_6_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_6_bits_decodeResult_maskDestination = queue_6_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_6_bits_decodeResult_maskLogic = queue_6_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_6_bits_decodeResult_uop = queue_6_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_6_bits_decodeResult_iota = queue_6_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_6_bits_decodeResult_mv = queue_6_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_6_bits_decodeResult_extend = queue_6_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_6_bits_decodeResult_unOrderWrite = queue_6_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_6_bits_decodeResult_compress = queue_6_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_6_bits_decodeResult_gather16 = queue_6_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_6_bits_decodeResult_gather = queue_6_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_6_bits_decodeResult_slid = queue_6_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_6_bits_decodeResult_targetRd = queue_6_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_6_bits_decodeResult_widenReduce = queue_6_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_6_bits_decodeResult_red = queue_6_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_6_bits_decodeResult_nr = queue_6_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_6_bits_decodeResult_itype = queue_6_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_6_bits_decodeResult_unsigned1 = queue_6_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_6_bits_decodeResult_unsigned0 = queue_6_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_6_bits_decodeResult_other = queue_6_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_6_bits_decodeResult_multiCycle = queue_6_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_6_bits_decodeResult_divider = queue_6_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_6_bits_decodeResult_multiplier = queue_6_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_6_bits_decodeResult_shift = queue_6_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_6_bits_decodeResult_adder = queue_6_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_6_bits_decodeResult_logic = queue_6_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_6_bits_loadStore = queue_6_deq_bits_loadStore;
  wire         laneRequestSinkWire_6_bits_issueInst = queue_6_deq_bits_issueInst;
  wire         laneRequestSinkWire_6_bits_store = queue_6_deq_bits_store;
  wire         laneRequestSinkWire_6_bits_special = queue_6_deq_bits_special;
  wire         laneRequestSinkWire_6_bits_lsWholeReg = queue_6_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_6_bits_vs1 = queue_6_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_6_bits_vs2 = queue_6_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_6_bits_vd = queue_6_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_6_bits_loadStoreEEW = queue_6_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_6_bits_mask = queue_6_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_6_bits_segment = queue_6_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_6_bits_readFromScalar = queue_6_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_6_bits_csrInterface_vl = queue_6_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_6_bits_csrInterface_vStart = queue_6_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_6_bits_csrInterface_vlmul = queue_6_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_6_bits_csrInterface_vSew = queue_6_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_6_bits_csrInterface_vxrm = queue_6_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_6_bits_csrInterface_vta = queue_6_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_6_bits_csrInterface_vma = queue_6_deq_bits_csrInterface_vma;
  wire [1:0]   queue_6_enq_bits_csrInterface_vxrm;
  wire         queue_6_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi_18 = {queue_6_enq_bits_csrInterface_vxrm, queue_6_enq_bits_csrInterface_vta};
  wire         queue_6_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo_18 = {queue_dataIn_lo_hi_18, queue_6_enq_bits_csrInterface_vma};
  wire [2:0]   queue_6_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_6_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo_18 = {queue_6_enq_bits_csrInterface_vlmul, queue_6_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_6_enq_bits_csrInterface_vl;
  wire [11:0]  queue_6_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi_18 = {queue_6_enq_bits_csrInterface_vl, queue_6_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi_18 = {queue_dataIn_hi_hi_18, queue_dataIn_hi_lo_18};
  wire         queue_6_enq_bits_decodeResult_adder;
  wire         queue_6_enq_bits_decodeResult_logic;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo_6 = {queue_6_enq_bits_decodeResult_adder, queue_6_enq_bits_decodeResult_logic};
  wire         queue_6_enq_bits_decodeResult_divider;
  wire         queue_6_enq_bits_decodeResult_multiplier;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi_6 = {queue_6_enq_bits_decodeResult_divider, queue_6_enq_bits_decodeResult_multiplier};
  wire         queue_6_enq_bits_decodeResult_shift;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi_6 = {queue_dataIn_lo_lo_lo_hi_hi_6, queue_6_enq_bits_decodeResult_shift};
  wire [4:0]   queue_dataIn_lo_lo_lo_6 = {queue_dataIn_lo_lo_lo_hi_6, queue_dataIn_lo_lo_lo_lo_6};
  wire         queue_6_enq_bits_decodeResult_unsigned0;
  wire         queue_6_enq_bits_decodeResult_other;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi_6 = {queue_6_enq_bits_decodeResult_unsigned0, queue_6_enq_bits_decodeResult_other};
  wire         queue_6_enq_bits_decodeResult_multiCycle;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo_6 = {queue_dataIn_lo_lo_hi_lo_hi_6, queue_6_enq_bits_decodeResult_multiCycle};
  wire         queue_6_enq_bits_decodeResult_nr;
  wire         queue_6_enq_bits_decodeResult_itype;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi_6 = {queue_6_enq_bits_decodeResult_nr, queue_6_enq_bits_decodeResult_itype};
  wire         queue_6_enq_bits_decodeResult_unsigned1;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi_6 = {queue_dataIn_lo_lo_hi_hi_hi_6, queue_6_enq_bits_decodeResult_unsigned1};
  wire [5:0]   queue_dataIn_lo_lo_hi_12 = {queue_dataIn_lo_lo_hi_hi_6, queue_dataIn_lo_lo_hi_lo_6};
  wire [10:0]  queue_dataIn_lo_lo_12 = {queue_dataIn_lo_lo_hi_12, queue_dataIn_lo_lo_lo_6};
  wire         queue_6_enq_bits_decodeResult_widenReduce;
  wire         queue_6_enq_bits_decodeResult_red;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo_6 = {queue_6_enq_bits_decodeResult_widenReduce, queue_6_enq_bits_decodeResult_red};
  wire         queue_6_enq_bits_decodeResult_gather;
  wire         queue_6_enq_bits_decodeResult_slid;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi_6 = {queue_6_enq_bits_decodeResult_gather, queue_6_enq_bits_decodeResult_slid};
  wire         queue_6_enq_bits_decodeResult_targetRd;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi_6 = {queue_dataIn_lo_hi_lo_hi_hi_6, queue_6_enq_bits_decodeResult_targetRd};
  wire [4:0]   queue_dataIn_lo_hi_lo_12 = {queue_dataIn_lo_hi_lo_hi_6, queue_dataIn_lo_hi_lo_lo_6};
  wire         queue_6_enq_bits_decodeResult_unOrderWrite;
  wire         queue_6_enq_bits_decodeResult_compress;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi_6 = {queue_6_enq_bits_decodeResult_unOrderWrite, queue_6_enq_bits_decodeResult_compress};
  wire         queue_6_enq_bits_decodeResult_gather16;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo_6 = {queue_dataIn_lo_hi_hi_lo_hi_6, queue_6_enq_bits_decodeResult_gather16};
  wire         queue_6_enq_bits_decodeResult_iota;
  wire         queue_6_enq_bits_decodeResult_mv;
  wire [1:0]   queue_dataIn_lo_hi_hi_hi_hi_6 = {queue_6_enq_bits_decodeResult_iota, queue_6_enq_bits_decodeResult_mv};
  wire         queue_6_enq_bits_decodeResult_extend;
  wire [2:0]   queue_dataIn_lo_hi_hi_hi_6 = {queue_dataIn_lo_hi_hi_hi_hi_6, queue_6_enq_bits_decodeResult_extend};
  wire [5:0]   queue_dataIn_lo_hi_hi_12 = {queue_dataIn_lo_hi_hi_hi_6, queue_dataIn_lo_hi_hi_lo_6};
  wire [10:0]  queue_dataIn_lo_hi_19 = {queue_dataIn_lo_hi_hi_12, queue_dataIn_lo_hi_lo_12};
  wire [21:0]  queue_dataIn_lo_19 = {queue_dataIn_lo_hi_19, queue_dataIn_lo_lo_12};
  wire         queue_6_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_6_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_hi_lo_lo_lo_6 = {queue_6_enq_bits_decodeResult_maskLogic, queue_6_enq_bits_decodeResult_uop};
  wire         queue_6_enq_bits_decodeResult_readOnly;
  wire         queue_6_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi_6 = {queue_6_enq_bits_decodeResult_readOnly, queue_6_enq_bits_decodeResult_maskSource};
  wire         queue_6_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi_6 = {queue_dataIn_hi_lo_lo_hi_hi_6, queue_6_enq_bits_decodeResult_maskDestination};
  wire [7:0]   queue_dataIn_hi_lo_lo_12 = {queue_dataIn_hi_lo_lo_hi_6, queue_dataIn_hi_lo_lo_lo_6};
  wire         queue_6_enq_bits_decodeResult_special;
  wire         queue_6_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi_6 = {queue_6_enq_bits_decodeResult_special, queue_6_enq_bits_decodeResult_saturate};
  wire         queue_6_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo_6 = {queue_dataIn_hi_lo_hi_lo_hi_6, queue_6_enq_bits_decodeResult_vwmacc};
  wire         queue_6_enq_bits_decodeResult_crossRead;
  wire         queue_6_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi_6 = {queue_6_enq_bits_decodeResult_crossRead, queue_6_enq_bits_decodeResult_crossWrite};
  wire         queue_6_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi_6 = {queue_dataIn_hi_lo_hi_hi_hi_6, queue_6_enq_bits_decodeResult_maskUnit};
  wire [5:0]   queue_dataIn_hi_lo_hi_12 = {queue_dataIn_hi_lo_hi_hi_6, queue_dataIn_hi_lo_hi_lo_6};
  wire [13:0]  queue_dataIn_hi_lo_19 = {queue_dataIn_hi_lo_hi_12, queue_dataIn_hi_lo_lo_12};
  wire         queue_6_enq_bits_decodeResult_vtype;
  wire         queue_6_enq_bits_decodeResult_sWrite;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo_6 = {queue_6_enq_bits_decodeResult_vtype, queue_6_enq_bits_decodeResult_sWrite};
  wire         queue_6_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_6_enq_bits_decodeResult_scheduler;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi_6 = {queue_6_enq_bits_decodeResult_dontNeedExecuteInLane, queue_6_enq_bits_decodeResult_scheduler};
  wire         queue_6_enq_bits_decodeResult_sReadVD;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi_6 = {queue_dataIn_hi_hi_lo_hi_hi_6, queue_6_enq_bits_decodeResult_sReadVD};
  wire [4:0]   queue_dataIn_hi_hi_lo_12 = {queue_dataIn_hi_hi_lo_hi_6, queue_dataIn_hi_hi_lo_lo_6};
  wire         queue_6_enq_bits_decodeResult_ffo;
  wire         queue_6_enq_bits_decodeResult_average;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi_6 = {queue_6_enq_bits_decodeResult_ffo, queue_6_enq_bits_decodeResult_average};
  wire         queue_6_enq_bits_decodeResult_reverse;
  wire [2:0]   queue_dataIn_hi_hi_hi_lo_6 = {queue_dataIn_hi_hi_hi_lo_hi_6, queue_6_enq_bits_decodeResult_reverse};
  wire         queue_6_enq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_6_enq_bits_decodeResult_topUop;
  wire [5:0]   queue_dataIn_hi_hi_hi_hi_hi_6 = {queue_6_enq_bits_decodeResult_specialSlot, queue_6_enq_bits_decodeResult_topUop};
  wire         queue_6_enq_bits_decodeResult_popCount;
  wire [6:0]   queue_dataIn_hi_hi_hi_hi_6 = {queue_dataIn_hi_hi_hi_hi_hi_6, queue_6_enq_bits_decodeResult_popCount};
  wire [9:0]   queue_dataIn_hi_hi_hi_12 = {queue_dataIn_hi_hi_hi_hi_6, queue_dataIn_hi_hi_hi_lo_6};
  wire [14:0]  queue_dataIn_hi_hi_19 = {queue_dataIn_hi_hi_hi_12, queue_dataIn_hi_hi_lo_12};
  wire [28:0]  queue_dataIn_hi_19 = {queue_dataIn_hi_hi_19, queue_dataIn_hi_lo_19};
  wire [2:0]   queue_6_enq_bits_segment;
  wire [31:0]  queue_6_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_13 = {queue_6_enq_bits_segment, queue_6_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_13 = {queue_dataIn_lo_lo_hi_13, queue_dataIn_hi_18, queue_dataIn_lo_18};
  wire [1:0]   queue_6_enq_bits_loadStoreEEW;
  wire         queue_6_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_13 = {queue_6_enq_bits_loadStoreEEW, queue_6_enq_bits_mask};
  wire [4:0]   queue_6_enq_bits_vs2;
  wire [4:0]   queue_6_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_13 = {queue_6_enq_bits_vs2, queue_6_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_20 = {queue_dataIn_lo_hi_hi_13, queue_dataIn_lo_hi_lo_13};
  wire [80:0]  queue_dataIn_lo_20 = {queue_dataIn_lo_hi_20, queue_dataIn_lo_lo_13};
  wire         queue_6_enq_bits_lsWholeReg;
  wire [4:0]   queue_6_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_13 = {queue_6_enq_bits_lsWholeReg, queue_6_enq_bits_vs1};
  wire         queue_6_enq_bits_store;
  wire         queue_6_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_13 = {queue_6_enq_bits_store, queue_6_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_20 = {queue_dataIn_hi_lo_hi_13, queue_dataIn_hi_lo_lo_13};
  wire         queue_6_enq_bits_loadStore;
  wire         queue_6_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_13 = {queue_6_enq_bits_loadStore, queue_6_enq_bits_issueInst};
  wire [2:0]   queue_6_enq_bits_instructionIndex;
  wire [53:0]  queue_dataIn_hi_hi_hi_13 = {queue_6_enq_bits_instructionIndex, queue_dataIn_hi_19, queue_dataIn_lo_19};
  wire [55:0]  queue_dataIn_hi_hi_20 = {queue_dataIn_hi_hi_hi_13, queue_dataIn_hi_hi_lo_13};
  wire [63:0]  queue_dataIn_hi_20 = {queue_dataIn_hi_hi_20, queue_dataIn_hi_lo_20};
  wire [144:0] queue_dataIn_6 = {queue_dataIn_hi_20, queue_dataIn_lo_20};
  wire         queue_dataOut_6_csrInterface_vma = _queue_fifo_6_data_out[0];
  wire         queue_dataOut_6_csrInterface_vta = _queue_fifo_6_data_out[1];
  wire [1:0]   queue_dataOut_6_csrInterface_vxrm = _queue_fifo_6_data_out[3:2];
  wire [1:0]   queue_dataOut_6_csrInterface_vSew = _queue_fifo_6_data_out[5:4];
  wire [2:0]   queue_dataOut_6_csrInterface_vlmul = _queue_fifo_6_data_out[8:6];
  wire [11:0]  queue_dataOut_6_csrInterface_vStart = _queue_fifo_6_data_out[20:9];
  wire [11:0]  queue_dataOut_6_csrInterface_vl = _queue_fifo_6_data_out[32:21];
  wire [31:0]  queue_dataOut_6_readFromScalar = _queue_fifo_6_data_out[64:33];
  wire [2:0]   queue_dataOut_6_segment = _queue_fifo_6_data_out[67:65];
  wire         queue_dataOut_6_mask = _queue_fifo_6_data_out[68];
  wire [1:0]   queue_dataOut_6_loadStoreEEW = _queue_fifo_6_data_out[70:69];
  wire [4:0]   queue_dataOut_6_vd = _queue_fifo_6_data_out[75:71];
  wire [4:0]   queue_dataOut_6_vs2 = _queue_fifo_6_data_out[80:76];
  wire [4:0]   queue_dataOut_6_vs1 = _queue_fifo_6_data_out[85:81];
  wire         queue_dataOut_6_lsWholeReg = _queue_fifo_6_data_out[86];
  wire         queue_dataOut_6_special = _queue_fifo_6_data_out[87];
  wire         queue_dataOut_6_store = _queue_fifo_6_data_out[88];
  wire         queue_dataOut_6_issueInst = _queue_fifo_6_data_out[89];
  wire         queue_dataOut_6_loadStore = _queue_fifo_6_data_out[90];
  wire         queue_dataOut_6_decodeResult_logic = _queue_fifo_6_data_out[91];
  wire         queue_dataOut_6_decodeResult_adder = _queue_fifo_6_data_out[92];
  wire         queue_dataOut_6_decodeResult_shift = _queue_fifo_6_data_out[93];
  wire         queue_dataOut_6_decodeResult_multiplier = _queue_fifo_6_data_out[94];
  wire         queue_dataOut_6_decodeResult_divider = _queue_fifo_6_data_out[95];
  wire         queue_dataOut_6_decodeResult_multiCycle = _queue_fifo_6_data_out[96];
  wire         queue_dataOut_6_decodeResult_other = _queue_fifo_6_data_out[97];
  wire         queue_dataOut_6_decodeResult_unsigned0 = _queue_fifo_6_data_out[98];
  wire         queue_dataOut_6_decodeResult_unsigned1 = _queue_fifo_6_data_out[99];
  wire         queue_dataOut_6_decodeResult_itype = _queue_fifo_6_data_out[100];
  wire         queue_dataOut_6_decodeResult_nr = _queue_fifo_6_data_out[101];
  wire         queue_dataOut_6_decodeResult_red = _queue_fifo_6_data_out[102];
  wire         queue_dataOut_6_decodeResult_widenReduce = _queue_fifo_6_data_out[103];
  wire         queue_dataOut_6_decodeResult_targetRd = _queue_fifo_6_data_out[104];
  wire         queue_dataOut_6_decodeResult_slid = _queue_fifo_6_data_out[105];
  wire         queue_dataOut_6_decodeResult_gather = _queue_fifo_6_data_out[106];
  wire         queue_dataOut_6_decodeResult_gather16 = _queue_fifo_6_data_out[107];
  wire         queue_dataOut_6_decodeResult_compress = _queue_fifo_6_data_out[108];
  wire         queue_dataOut_6_decodeResult_unOrderWrite = _queue_fifo_6_data_out[109];
  wire         queue_dataOut_6_decodeResult_extend = _queue_fifo_6_data_out[110];
  wire         queue_dataOut_6_decodeResult_mv = _queue_fifo_6_data_out[111];
  wire         queue_dataOut_6_decodeResult_iota = _queue_fifo_6_data_out[112];
  wire [3:0]   queue_dataOut_6_decodeResult_uop = _queue_fifo_6_data_out[116:113];
  wire         queue_dataOut_6_decodeResult_maskLogic = _queue_fifo_6_data_out[117];
  wire         queue_dataOut_6_decodeResult_maskDestination = _queue_fifo_6_data_out[118];
  wire         queue_dataOut_6_decodeResult_maskSource = _queue_fifo_6_data_out[119];
  wire         queue_dataOut_6_decodeResult_readOnly = _queue_fifo_6_data_out[120];
  wire         queue_dataOut_6_decodeResult_vwmacc = _queue_fifo_6_data_out[121];
  wire         queue_dataOut_6_decodeResult_saturate = _queue_fifo_6_data_out[122];
  wire         queue_dataOut_6_decodeResult_special = _queue_fifo_6_data_out[123];
  wire         queue_dataOut_6_decodeResult_maskUnit = _queue_fifo_6_data_out[124];
  wire         queue_dataOut_6_decodeResult_crossWrite = _queue_fifo_6_data_out[125];
  wire         queue_dataOut_6_decodeResult_crossRead = _queue_fifo_6_data_out[126];
  wire         queue_dataOut_6_decodeResult_sWrite = _queue_fifo_6_data_out[127];
  wire         queue_dataOut_6_decodeResult_vtype = _queue_fifo_6_data_out[128];
  wire         queue_dataOut_6_decodeResult_sReadVD = _queue_fifo_6_data_out[129];
  wire         queue_dataOut_6_decodeResult_scheduler = _queue_fifo_6_data_out[130];
  wire         queue_dataOut_6_decodeResult_dontNeedExecuteInLane = _queue_fifo_6_data_out[131];
  wire         queue_dataOut_6_decodeResult_reverse = _queue_fifo_6_data_out[132];
  wire         queue_dataOut_6_decodeResult_average = _queue_fifo_6_data_out[133];
  wire         queue_dataOut_6_decodeResult_ffo = _queue_fifo_6_data_out[134];
  wire         queue_dataOut_6_decodeResult_popCount = _queue_fifo_6_data_out[135];
  wire [4:0]   queue_dataOut_6_decodeResult_topUop = _queue_fifo_6_data_out[140:136];
  wire         queue_dataOut_6_decodeResult_specialSlot = _queue_fifo_6_data_out[141];
  wire [2:0]   queue_dataOut_6_instructionIndex = _queue_fifo_6_data_out[144:142];
  wire         queue_6_enq_ready = ~_queue_fifo_6_full;
  wire         queue_6_enq_valid;
  assign queue_6_deq_valid = ~_queue_fifo_6_empty | queue_6_enq_valid;
  assign queue_6_deq_bits_instructionIndex = _queue_fifo_6_empty ? queue_6_enq_bits_instructionIndex : queue_dataOut_6_instructionIndex;
  assign queue_6_deq_bits_decodeResult_specialSlot = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_specialSlot : queue_dataOut_6_decodeResult_specialSlot;
  assign queue_6_deq_bits_decodeResult_topUop = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_topUop : queue_dataOut_6_decodeResult_topUop;
  assign queue_6_deq_bits_decodeResult_popCount = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_popCount : queue_dataOut_6_decodeResult_popCount;
  assign queue_6_deq_bits_decodeResult_ffo = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_ffo : queue_dataOut_6_decodeResult_ffo;
  assign queue_6_deq_bits_decodeResult_average = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_average : queue_dataOut_6_decodeResult_average;
  assign queue_6_deq_bits_decodeResult_reverse = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_reverse : queue_dataOut_6_decodeResult_reverse;
  assign queue_6_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_6_decodeResult_dontNeedExecuteInLane;
  assign queue_6_deq_bits_decodeResult_scheduler = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_scheduler : queue_dataOut_6_decodeResult_scheduler;
  assign queue_6_deq_bits_decodeResult_sReadVD = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_sReadVD : queue_dataOut_6_decodeResult_sReadVD;
  assign queue_6_deq_bits_decodeResult_vtype = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_vtype : queue_dataOut_6_decodeResult_vtype;
  assign queue_6_deq_bits_decodeResult_sWrite = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_sWrite : queue_dataOut_6_decodeResult_sWrite;
  assign queue_6_deq_bits_decodeResult_crossRead = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_crossRead : queue_dataOut_6_decodeResult_crossRead;
  assign queue_6_deq_bits_decodeResult_crossWrite = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_crossWrite : queue_dataOut_6_decodeResult_crossWrite;
  assign queue_6_deq_bits_decodeResult_maskUnit = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_maskUnit : queue_dataOut_6_decodeResult_maskUnit;
  assign queue_6_deq_bits_decodeResult_special = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_special : queue_dataOut_6_decodeResult_special;
  assign queue_6_deq_bits_decodeResult_saturate = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_saturate : queue_dataOut_6_decodeResult_saturate;
  assign queue_6_deq_bits_decodeResult_vwmacc = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_vwmacc : queue_dataOut_6_decodeResult_vwmacc;
  assign queue_6_deq_bits_decodeResult_readOnly = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_readOnly : queue_dataOut_6_decodeResult_readOnly;
  assign queue_6_deq_bits_decodeResult_maskSource = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_maskSource : queue_dataOut_6_decodeResult_maskSource;
  assign queue_6_deq_bits_decodeResult_maskDestination = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_maskDestination : queue_dataOut_6_decodeResult_maskDestination;
  assign queue_6_deq_bits_decodeResult_maskLogic = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_maskLogic : queue_dataOut_6_decodeResult_maskLogic;
  assign queue_6_deq_bits_decodeResult_uop = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_uop : queue_dataOut_6_decodeResult_uop;
  assign queue_6_deq_bits_decodeResult_iota = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_iota : queue_dataOut_6_decodeResult_iota;
  assign queue_6_deq_bits_decodeResult_mv = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_mv : queue_dataOut_6_decodeResult_mv;
  assign queue_6_deq_bits_decodeResult_extend = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_extend : queue_dataOut_6_decodeResult_extend;
  assign queue_6_deq_bits_decodeResult_unOrderWrite = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_unOrderWrite : queue_dataOut_6_decodeResult_unOrderWrite;
  assign queue_6_deq_bits_decodeResult_compress = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_compress : queue_dataOut_6_decodeResult_compress;
  assign queue_6_deq_bits_decodeResult_gather16 = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_gather16 : queue_dataOut_6_decodeResult_gather16;
  assign queue_6_deq_bits_decodeResult_gather = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_gather : queue_dataOut_6_decodeResult_gather;
  assign queue_6_deq_bits_decodeResult_slid = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_slid : queue_dataOut_6_decodeResult_slid;
  assign queue_6_deq_bits_decodeResult_targetRd = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_targetRd : queue_dataOut_6_decodeResult_targetRd;
  assign queue_6_deq_bits_decodeResult_widenReduce = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_widenReduce : queue_dataOut_6_decodeResult_widenReduce;
  assign queue_6_deq_bits_decodeResult_red = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_red : queue_dataOut_6_decodeResult_red;
  assign queue_6_deq_bits_decodeResult_nr = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_nr : queue_dataOut_6_decodeResult_nr;
  assign queue_6_deq_bits_decodeResult_itype = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_itype : queue_dataOut_6_decodeResult_itype;
  assign queue_6_deq_bits_decodeResult_unsigned1 = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_unsigned1 : queue_dataOut_6_decodeResult_unsigned1;
  assign queue_6_deq_bits_decodeResult_unsigned0 = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_unsigned0 : queue_dataOut_6_decodeResult_unsigned0;
  assign queue_6_deq_bits_decodeResult_other = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_other : queue_dataOut_6_decodeResult_other;
  assign queue_6_deq_bits_decodeResult_multiCycle = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_multiCycle : queue_dataOut_6_decodeResult_multiCycle;
  assign queue_6_deq_bits_decodeResult_divider = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_divider : queue_dataOut_6_decodeResult_divider;
  assign queue_6_deq_bits_decodeResult_multiplier = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_multiplier : queue_dataOut_6_decodeResult_multiplier;
  assign queue_6_deq_bits_decodeResult_shift = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_shift : queue_dataOut_6_decodeResult_shift;
  assign queue_6_deq_bits_decodeResult_adder = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_adder : queue_dataOut_6_decodeResult_adder;
  assign queue_6_deq_bits_decodeResult_logic = _queue_fifo_6_empty ? queue_6_enq_bits_decodeResult_logic : queue_dataOut_6_decodeResult_logic;
  assign queue_6_deq_bits_loadStore = _queue_fifo_6_empty ? queue_6_enq_bits_loadStore : queue_dataOut_6_loadStore;
  assign queue_6_deq_bits_issueInst = _queue_fifo_6_empty ? queue_6_enq_bits_issueInst : queue_dataOut_6_issueInst;
  assign queue_6_deq_bits_store = _queue_fifo_6_empty ? queue_6_enq_bits_store : queue_dataOut_6_store;
  assign queue_6_deq_bits_special = _queue_fifo_6_empty ? queue_6_enq_bits_special : queue_dataOut_6_special;
  assign queue_6_deq_bits_lsWholeReg = _queue_fifo_6_empty ? queue_6_enq_bits_lsWholeReg : queue_dataOut_6_lsWholeReg;
  assign queue_6_deq_bits_vs1 = _queue_fifo_6_empty ? queue_6_enq_bits_vs1 : queue_dataOut_6_vs1;
  assign queue_6_deq_bits_vs2 = _queue_fifo_6_empty ? queue_6_enq_bits_vs2 : queue_dataOut_6_vs2;
  assign queue_6_deq_bits_vd = _queue_fifo_6_empty ? queue_6_enq_bits_vd : queue_dataOut_6_vd;
  assign queue_6_deq_bits_loadStoreEEW = _queue_fifo_6_empty ? queue_6_enq_bits_loadStoreEEW : queue_dataOut_6_loadStoreEEW;
  assign queue_6_deq_bits_mask = _queue_fifo_6_empty ? queue_6_enq_bits_mask : queue_dataOut_6_mask;
  assign queue_6_deq_bits_segment = _queue_fifo_6_empty ? queue_6_enq_bits_segment : queue_dataOut_6_segment;
  assign queue_6_deq_bits_readFromScalar = _queue_fifo_6_empty ? queue_6_enq_bits_readFromScalar : queue_dataOut_6_readFromScalar;
  assign queue_6_deq_bits_csrInterface_vl = _queue_fifo_6_empty ? queue_6_enq_bits_csrInterface_vl : queue_dataOut_6_csrInterface_vl;
  assign queue_6_deq_bits_csrInterface_vStart = _queue_fifo_6_empty ? queue_6_enq_bits_csrInterface_vStart : queue_dataOut_6_csrInterface_vStart;
  assign queue_6_deq_bits_csrInterface_vlmul = _queue_fifo_6_empty ? queue_6_enq_bits_csrInterface_vlmul : queue_dataOut_6_csrInterface_vlmul;
  assign queue_6_deq_bits_csrInterface_vSew = _queue_fifo_6_empty ? queue_6_enq_bits_csrInterface_vSew : queue_dataOut_6_csrInterface_vSew;
  assign queue_6_deq_bits_csrInterface_vxrm = _queue_fifo_6_empty ? queue_6_enq_bits_csrInterface_vxrm : queue_dataOut_6_csrInterface_vxrm;
  assign queue_6_deq_bits_csrInterface_vta = _queue_fifo_6_empty ? queue_6_enq_bits_csrInterface_vta : queue_dataOut_6_csrInterface_vta;
  assign queue_6_deq_bits_csrInterface_vma = _queue_fifo_6_empty ? queue_6_enq_bits_csrInterface_vma : queue_dataOut_6_csrInterface_vma;
  wire         laneVec_6_laneRequest_bits_issueInst = laneRequestSinkWire_6_ready & laneRequestSinkWire_6_valid;
  reg          releasePipe_pipe_v_6;
  wire         releasePipe_pipe_out_6_valid = releasePipe_pipe_v_6;
  wire         laneRequestSourceWire_6_ready;
  wire         validSource_6_valid = laneRequestSourceWire_6_ready & laneRequestSourceWire_6_valid;
  reg  [2:0]   tokenCheck_counter_6;
  wire [2:0]   tokenCheck_counterChange_6 = validSource_6_valid ? 3'h1 : 3'h7;
  assign tokenCheck_6 = ~(tokenCheck_counter_6[2]);
  assign laneRequestSourceWire_6_ready = tokenCheck_6;
  assign queue_6_enq_valid = validSink_6_valid;
  assign queue_6_enq_bits_instructionIndex = validSink_6_bits_instructionIndex;
  assign queue_6_enq_bits_decodeResult_specialSlot = validSink_6_bits_decodeResult_specialSlot;
  assign queue_6_enq_bits_decodeResult_topUop = validSink_6_bits_decodeResult_topUop;
  assign queue_6_enq_bits_decodeResult_popCount = validSink_6_bits_decodeResult_popCount;
  assign queue_6_enq_bits_decodeResult_ffo = validSink_6_bits_decodeResult_ffo;
  assign queue_6_enq_bits_decodeResult_average = validSink_6_bits_decodeResult_average;
  assign queue_6_enq_bits_decodeResult_reverse = validSink_6_bits_decodeResult_reverse;
  assign queue_6_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_6_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_6_enq_bits_decodeResult_scheduler = validSink_6_bits_decodeResult_scheduler;
  assign queue_6_enq_bits_decodeResult_sReadVD = validSink_6_bits_decodeResult_sReadVD;
  assign queue_6_enq_bits_decodeResult_vtype = validSink_6_bits_decodeResult_vtype;
  assign queue_6_enq_bits_decodeResult_sWrite = validSink_6_bits_decodeResult_sWrite;
  assign queue_6_enq_bits_decodeResult_crossRead = validSink_6_bits_decodeResult_crossRead;
  assign queue_6_enq_bits_decodeResult_crossWrite = validSink_6_bits_decodeResult_crossWrite;
  assign queue_6_enq_bits_decodeResult_maskUnit = validSink_6_bits_decodeResult_maskUnit;
  assign queue_6_enq_bits_decodeResult_special = validSink_6_bits_decodeResult_special;
  assign queue_6_enq_bits_decodeResult_saturate = validSink_6_bits_decodeResult_saturate;
  assign queue_6_enq_bits_decodeResult_vwmacc = validSink_6_bits_decodeResult_vwmacc;
  assign queue_6_enq_bits_decodeResult_readOnly = validSink_6_bits_decodeResult_readOnly;
  assign queue_6_enq_bits_decodeResult_maskSource = validSink_6_bits_decodeResult_maskSource;
  assign queue_6_enq_bits_decodeResult_maskDestination = validSink_6_bits_decodeResult_maskDestination;
  assign queue_6_enq_bits_decodeResult_maskLogic = validSink_6_bits_decodeResult_maskLogic;
  assign queue_6_enq_bits_decodeResult_uop = validSink_6_bits_decodeResult_uop;
  assign queue_6_enq_bits_decodeResult_iota = validSink_6_bits_decodeResult_iota;
  assign queue_6_enq_bits_decodeResult_mv = validSink_6_bits_decodeResult_mv;
  assign queue_6_enq_bits_decodeResult_extend = validSink_6_bits_decodeResult_extend;
  assign queue_6_enq_bits_decodeResult_unOrderWrite = validSink_6_bits_decodeResult_unOrderWrite;
  assign queue_6_enq_bits_decodeResult_compress = validSink_6_bits_decodeResult_compress;
  assign queue_6_enq_bits_decodeResult_gather16 = validSink_6_bits_decodeResult_gather16;
  assign queue_6_enq_bits_decodeResult_gather = validSink_6_bits_decodeResult_gather;
  assign queue_6_enq_bits_decodeResult_slid = validSink_6_bits_decodeResult_slid;
  assign queue_6_enq_bits_decodeResult_targetRd = validSink_6_bits_decodeResult_targetRd;
  assign queue_6_enq_bits_decodeResult_widenReduce = validSink_6_bits_decodeResult_widenReduce;
  assign queue_6_enq_bits_decodeResult_red = validSink_6_bits_decodeResult_red;
  assign queue_6_enq_bits_decodeResult_nr = validSink_6_bits_decodeResult_nr;
  assign queue_6_enq_bits_decodeResult_itype = validSink_6_bits_decodeResult_itype;
  assign queue_6_enq_bits_decodeResult_unsigned1 = validSink_6_bits_decodeResult_unsigned1;
  assign queue_6_enq_bits_decodeResult_unsigned0 = validSink_6_bits_decodeResult_unsigned0;
  assign queue_6_enq_bits_decodeResult_other = validSink_6_bits_decodeResult_other;
  assign queue_6_enq_bits_decodeResult_multiCycle = validSink_6_bits_decodeResult_multiCycle;
  assign queue_6_enq_bits_decodeResult_divider = validSink_6_bits_decodeResult_divider;
  assign queue_6_enq_bits_decodeResult_multiplier = validSink_6_bits_decodeResult_multiplier;
  assign queue_6_enq_bits_decodeResult_shift = validSink_6_bits_decodeResult_shift;
  assign queue_6_enq_bits_decodeResult_adder = validSink_6_bits_decodeResult_adder;
  assign queue_6_enq_bits_decodeResult_logic = validSink_6_bits_decodeResult_logic;
  assign queue_6_enq_bits_loadStore = validSink_6_bits_loadStore;
  assign queue_6_enq_bits_issueInst = validSink_6_bits_issueInst;
  assign queue_6_enq_bits_store = validSink_6_bits_store;
  assign queue_6_enq_bits_special = validSink_6_bits_special;
  assign queue_6_enq_bits_lsWholeReg = validSink_6_bits_lsWholeReg;
  assign queue_6_enq_bits_vs1 = validSink_6_bits_vs1;
  assign queue_6_enq_bits_vs2 = validSink_6_bits_vs2;
  assign queue_6_enq_bits_vd = validSink_6_bits_vd;
  assign queue_6_enq_bits_loadStoreEEW = validSink_6_bits_loadStoreEEW;
  assign queue_6_enq_bits_mask = validSink_6_bits_mask;
  assign queue_6_enq_bits_segment = validSink_6_bits_segment;
  assign queue_6_enq_bits_readFromScalar = validSink_6_bits_readFromScalar;
  assign queue_6_enq_bits_csrInterface_vl = validSink_6_bits_csrInterface_vl;
  assign queue_6_enq_bits_csrInterface_vStart = validSink_6_bits_csrInterface_vStart;
  assign queue_6_enq_bits_csrInterface_vlmul = validSink_6_bits_csrInterface_vlmul;
  assign queue_6_enq_bits_csrInterface_vSew = validSink_6_bits_csrInterface_vSew;
  assign queue_6_enq_bits_csrInterface_vxrm = validSink_6_bits_csrInterface_vxrm;
  assign queue_6_enq_bits_csrInterface_vta = validSink_6_bits_csrInterface_vta;
  assign queue_6_enq_bits_csrInterface_vma = validSink_6_bits_csrInterface_vma;
  reg          shifterReg_6_0_valid;
  assign validSink_6_valid = shifterReg_6_0_valid;
  reg  [2:0]   shifterReg_6_0_bits_instructionIndex;
  assign validSink_6_bits_instructionIndex = shifterReg_6_0_bits_instructionIndex;
  reg          shifterReg_6_0_bits_decodeResult_specialSlot;
  assign validSink_6_bits_decodeResult_specialSlot = shifterReg_6_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_6_0_bits_decodeResult_topUop;
  assign validSink_6_bits_decodeResult_topUop = shifterReg_6_0_bits_decodeResult_topUop;
  reg          shifterReg_6_0_bits_decodeResult_popCount;
  assign validSink_6_bits_decodeResult_popCount = shifterReg_6_0_bits_decodeResult_popCount;
  reg          shifterReg_6_0_bits_decodeResult_ffo;
  assign validSink_6_bits_decodeResult_ffo = shifterReg_6_0_bits_decodeResult_ffo;
  reg          shifterReg_6_0_bits_decodeResult_average;
  assign validSink_6_bits_decodeResult_average = shifterReg_6_0_bits_decodeResult_average;
  reg          shifterReg_6_0_bits_decodeResult_reverse;
  assign validSink_6_bits_decodeResult_reverse = shifterReg_6_0_bits_decodeResult_reverse;
  reg          shifterReg_6_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_6_bits_decodeResult_dontNeedExecuteInLane = shifterReg_6_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_6_0_bits_decodeResult_scheduler;
  assign validSink_6_bits_decodeResult_scheduler = shifterReg_6_0_bits_decodeResult_scheduler;
  reg          shifterReg_6_0_bits_decodeResult_sReadVD;
  assign validSink_6_bits_decodeResult_sReadVD = shifterReg_6_0_bits_decodeResult_sReadVD;
  reg          shifterReg_6_0_bits_decodeResult_vtype;
  assign validSink_6_bits_decodeResult_vtype = shifterReg_6_0_bits_decodeResult_vtype;
  reg          shifterReg_6_0_bits_decodeResult_sWrite;
  assign validSink_6_bits_decodeResult_sWrite = shifterReg_6_0_bits_decodeResult_sWrite;
  reg          shifterReg_6_0_bits_decodeResult_crossRead;
  assign validSink_6_bits_decodeResult_crossRead = shifterReg_6_0_bits_decodeResult_crossRead;
  reg          shifterReg_6_0_bits_decodeResult_crossWrite;
  assign validSink_6_bits_decodeResult_crossWrite = shifterReg_6_0_bits_decodeResult_crossWrite;
  reg          shifterReg_6_0_bits_decodeResult_maskUnit;
  assign validSink_6_bits_decodeResult_maskUnit = shifterReg_6_0_bits_decodeResult_maskUnit;
  reg          shifterReg_6_0_bits_decodeResult_special;
  assign validSink_6_bits_decodeResult_special = shifterReg_6_0_bits_decodeResult_special;
  reg          shifterReg_6_0_bits_decodeResult_saturate;
  assign validSink_6_bits_decodeResult_saturate = shifterReg_6_0_bits_decodeResult_saturate;
  reg          shifterReg_6_0_bits_decodeResult_vwmacc;
  assign validSink_6_bits_decodeResult_vwmacc = shifterReg_6_0_bits_decodeResult_vwmacc;
  reg          shifterReg_6_0_bits_decodeResult_readOnly;
  assign validSink_6_bits_decodeResult_readOnly = shifterReg_6_0_bits_decodeResult_readOnly;
  reg          shifterReg_6_0_bits_decodeResult_maskSource;
  assign validSink_6_bits_decodeResult_maskSource = shifterReg_6_0_bits_decodeResult_maskSource;
  reg          shifterReg_6_0_bits_decodeResult_maskDestination;
  assign validSink_6_bits_decodeResult_maskDestination = shifterReg_6_0_bits_decodeResult_maskDestination;
  reg          shifterReg_6_0_bits_decodeResult_maskLogic;
  assign validSink_6_bits_decodeResult_maskLogic = shifterReg_6_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_6_0_bits_decodeResult_uop;
  assign validSink_6_bits_decodeResult_uop = shifterReg_6_0_bits_decodeResult_uop;
  reg          shifterReg_6_0_bits_decodeResult_iota;
  assign validSink_6_bits_decodeResult_iota = shifterReg_6_0_bits_decodeResult_iota;
  reg          shifterReg_6_0_bits_decodeResult_mv;
  assign validSink_6_bits_decodeResult_mv = shifterReg_6_0_bits_decodeResult_mv;
  reg          shifterReg_6_0_bits_decodeResult_extend;
  assign validSink_6_bits_decodeResult_extend = shifterReg_6_0_bits_decodeResult_extend;
  reg          shifterReg_6_0_bits_decodeResult_unOrderWrite;
  assign validSink_6_bits_decodeResult_unOrderWrite = shifterReg_6_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_6_0_bits_decodeResult_compress;
  assign validSink_6_bits_decodeResult_compress = shifterReg_6_0_bits_decodeResult_compress;
  reg          shifterReg_6_0_bits_decodeResult_gather16;
  assign validSink_6_bits_decodeResult_gather16 = shifterReg_6_0_bits_decodeResult_gather16;
  reg          shifterReg_6_0_bits_decodeResult_gather;
  assign validSink_6_bits_decodeResult_gather = shifterReg_6_0_bits_decodeResult_gather;
  reg          shifterReg_6_0_bits_decodeResult_slid;
  assign validSink_6_bits_decodeResult_slid = shifterReg_6_0_bits_decodeResult_slid;
  reg          shifterReg_6_0_bits_decodeResult_targetRd;
  assign validSink_6_bits_decodeResult_targetRd = shifterReg_6_0_bits_decodeResult_targetRd;
  reg          shifterReg_6_0_bits_decodeResult_widenReduce;
  assign validSink_6_bits_decodeResult_widenReduce = shifterReg_6_0_bits_decodeResult_widenReduce;
  reg          shifterReg_6_0_bits_decodeResult_red;
  assign validSink_6_bits_decodeResult_red = shifterReg_6_0_bits_decodeResult_red;
  reg          shifterReg_6_0_bits_decodeResult_nr;
  assign validSink_6_bits_decodeResult_nr = shifterReg_6_0_bits_decodeResult_nr;
  reg          shifterReg_6_0_bits_decodeResult_itype;
  assign validSink_6_bits_decodeResult_itype = shifterReg_6_0_bits_decodeResult_itype;
  reg          shifterReg_6_0_bits_decodeResult_unsigned1;
  assign validSink_6_bits_decodeResult_unsigned1 = shifterReg_6_0_bits_decodeResult_unsigned1;
  reg          shifterReg_6_0_bits_decodeResult_unsigned0;
  assign validSink_6_bits_decodeResult_unsigned0 = shifterReg_6_0_bits_decodeResult_unsigned0;
  reg          shifterReg_6_0_bits_decodeResult_other;
  assign validSink_6_bits_decodeResult_other = shifterReg_6_0_bits_decodeResult_other;
  reg          shifterReg_6_0_bits_decodeResult_multiCycle;
  assign validSink_6_bits_decodeResult_multiCycle = shifterReg_6_0_bits_decodeResult_multiCycle;
  reg          shifterReg_6_0_bits_decodeResult_divider;
  assign validSink_6_bits_decodeResult_divider = shifterReg_6_0_bits_decodeResult_divider;
  reg          shifterReg_6_0_bits_decodeResult_multiplier;
  assign validSink_6_bits_decodeResult_multiplier = shifterReg_6_0_bits_decodeResult_multiplier;
  reg          shifterReg_6_0_bits_decodeResult_shift;
  assign validSink_6_bits_decodeResult_shift = shifterReg_6_0_bits_decodeResult_shift;
  reg          shifterReg_6_0_bits_decodeResult_adder;
  assign validSink_6_bits_decodeResult_adder = shifterReg_6_0_bits_decodeResult_adder;
  reg          shifterReg_6_0_bits_decodeResult_logic;
  assign validSink_6_bits_decodeResult_logic = shifterReg_6_0_bits_decodeResult_logic;
  reg          shifterReg_6_0_bits_loadStore;
  assign validSink_6_bits_loadStore = shifterReg_6_0_bits_loadStore;
  reg          shifterReg_6_0_bits_issueInst;
  assign validSink_6_bits_issueInst = shifterReg_6_0_bits_issueInst;
  reg          shifterReg_6_0_bits_store;
  assign validSink_6_bits_store = shifterReg_6_0_bits_store;
  reg          shifterReg_6_0_bits_special;
  assign validSink_6_bits_special = shifterReg_6_0_bits_special;
  reg          shifterReg_6_0_bits_lsWholeReg;
  assign validSink_6_bits_lsWholeReg = shifterReg_6_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_6_0_bits_vs1;
  assign validSink_6_bits_vs1 = shifterReg_6_0_bits_vs1;
  reg  [4:0]   shifterReg_6_0_bits_vs2;
  assign validSink_6_bits_vs2 = shifterReg_6_0_bits_vs2;
  reg  [4:0]   shifterReg_6_0_bits_vd;
  assign validSink_6_bits_vd = shifterReg_6_0_bits_vd;
  reg  [1:0]   shifterReg_6_0_bits_loadStoreEEW;
  assign validSink_6_bits_loadStoreEEW = shifterReg_6_0_bits_loadStoreEEW;
  reg          shifterReg_6_0_bits_mask;
  assign validSink_6_bits_mask = shifterReg_6_0_bits_mask;
  reg  [2:0]   shifterReg_6_0_bits_segment;
  assign validSink_6_bits_segment = shifterReg_6_0_bits_segment;
  reg  [31:0]  shifterReg_6_0_bits_readFromScalar;
  assign validSink_6_bits_readFromScalar = shifterReg_6_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_6_0_bits_csrInterface_vl;
  assign validSink_6_bits_csrInterface_vl = shifterReg_6_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_6_0_bits_csrInterface_vStart;
  assign validSink_6_bits_csrInterface_vStart = shifterReg_6_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_6_0_bits_csrInterface_vlmul;
  assign validSink_6_bits_csrInterface_vlmul = shifterReg_6_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_6_0_bits_csrInterface_vSew;
  assign validSink_6_bits_csrInterface_vSew = shifterReg_6_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_6_0_bits_csrInterface_vxrm;
  assign validSink_6_bits_csrInterface_vxrm = shifterReg_6_0_bits_csrInterface_vxrm;
  reg          shifterReg_6_0_bits_csrInterface_vta;
  assign validSink_6_bits_csrInterface_vta = shifterReg_6_0_bits_csrInterface_vta;
  reg          shifterReg_6_0_bits_csrInterface_vma;
  assign validSink_6_bits_csrInterface_vma = shifterReg_6_0_bits_csrInterface_vma;
  wire         shifterValid_6 = shifterReg_6_0_valid | validSource_6_valid;
  wire         validSink_7_valid;
  wire [2:0]   validSink_7_bits_instructionIndex;
  wire         validSink_7_bits_decodeResult_specialSlot;
  wire [4:0]   validSink_7_bits_decodeResult_topUop;
  wire         validSink_7_bits_decodeResult_popCount;
  wire         validSink_7_bits_decodeResult_ffo;
  wire         validSink_7_bits_decodeResult_average;
  wire         validSink_7_bits_decodeResult_reverse;
  wire         validSink_7_bits_decodeResult_dontNeedExecuteInLane;
  wire         validSink_7_bits_decodeResult_scheduler;
  wire         validSink_7_bits_decodeResult_sReadVD;
  wire         validSink_7_bits_decodeResult_vtype;
  wire         validSink_7_bits_decodeResult_sWrite;
  wire         validSink_7_bits_decodeResult_crossRead;
  wire         validSink_7_bits_decodeResult_crossWrite;
  wire         validSink_7_bits_decodeResult_maskUnit;
  wire         validSink_7_bits_decodeResult_special;
  wire         validSink_7_bits_decodeResult_saturate;
  wire         validSink_7_bits_decodeResult_vwmacc;
  wire         validSink_7_bits_decodeResult_readOnly;
  wire         validSink_7_bits_decodeResult_maskSource;
  wire         validSink_7_bits_decodeResult_maskDestination;
  wire         validSink_7_bits_decodeResult_maskLogic;
  wire [3:0]   validSink_7_bits_decodeResult_uop;
  wire         validSink_7_bits_decodeResult_iota;
  wire         validSink_7_bits_decodeResult_mv;
  wire         validSink_7_bits_decodeResult_extend;
  wire         validSink_7_bits_decodeResult_unOrderWrite;
  wire         validSink_7_bits_decodeResult_compress;
  wire         validSink_7_bits_decodeResult_gather16;
  wire         validSink_7_bits_decodeResult_gather;
  wire         validSink_7_bits_decodeResult_slid;
  wire         validSink_7_bits_decodeResult_targetRd;
  wire         validSink_7_bits_decodeResult_widenReduce;
  wire         validSink_7_bits_decodeResult_red;
  wire         validSink_7_bits_decodeResult_nr;
  wire         validSink_7_bits_decodeResult_itype;
  wire         validSink_7_bits_decodeResult_unsigned1;
  wire         validSink_7_bits_decodeResult_unsigned0;
  wire         validSink_7_bits_decodeResult_other;
  wire         validSink_7_bits_decodeResult_multiCycle;
  wire         validSink_7_bits_decodeResult_divider;
  wire         validSink_7_bits_decodeResult_multiplier;
  wire         validSink_7_bits_decodeResult_shift;
  wire         validSink_7_bits_decodeResult_adder;
  wire         validSink_7_bits_decodeResult_logic;
  wire         validSink_7_bits_loadStore;
  wire         validSink_7_bits_issueInst;
  wire         validSink_7_bits_store;
  wire         validSink_7_bits_special;
  wire         validSink_7_bits_lsWholeReg;
  wire [4:0]   validSink_7_bits_vs1;
  wire [4:0]   validSink_7_bits_vs2;
  wire [4:0]   validSink_7_bits_vd;
  wire [1:0]   validSink_7_bits_loadStoreEEW;
  wire         validSink_7_bits_mask;
  wire [2:0]   validSink_7_bits_segment;
  wire [31:0]  validSink_7_bits_readFromScalar;
  wire [11:0]  validSink_7_bits_csrInterface_vl;
  wire [11:0]  validSink_7_bits_csrInterface_vStart;
  wire [2:0]   validSink_7_bits_csrInterface_vlmul;
  wire [1:0]   validSink_7_bits_csrInterface_vSew;
  wire [1:0]   validSink_7_bits_csrInterface_vxrm;
  wire         validSink_7_bits_csrInterface_vta;
  wire         validSink_7_bits_csrInterface_vma;
  wire         laneRequestSinkWire_7_valid = queue_7_deq_valid;
  wire [2:0]   laneRequestSinkWire_7_bits_instructionIndex = queue_7_deq_bits_instructionIndex;
  wire         laneRequestSinkWire_7_bits_decodeResult_specialSlot = queue_7_deq_bits_decodeResult_specialSlot;
  wire [4:0]   laneRequestSinkWire_7_bits_decodeResult_topUop = queue_7_deq_bits_decodeResult_topUop;
  wire         laneRequestSinkWire_7_bits_decodeResult_popCount = queue_7_deq_bits_decodeResult_popCount;
  wire         laneRequestSinkWire_7_bits_decodeResult_ffo = queue_7_deq_bits_decodeResult_ffo;
  wire         laneRequestSinkWire_7_bits_decodeResult_average = queue_7_deq_bits_decodeResult_average;
  wire         laneRequestSinkWire_7_bits_decodeResult_reverse = queue_7_deq_bits_decodeResult_reverse;
  wire         laneRequestSinkWire_7_bits_decodeResult_dontNeedExecuteInLane = queue_7_deq_bits_decodeResult_dontNeedExecuteInLane;
  wire         laneRequestSinkWire_7_bits_decodeResult_scheduler = queue_7_deq_bits_decodeResult_scheduler;
  wire         laneRequestSinkWire_7_bits_decodeResult_sReadVD = queue_7_deq_bits_decodeResult_sReadVD;
  wire         laneRequestSinkWire_7_bits_decodeResult_vtype = queue_7_deq_bits_decodeResult_vtype;
  wire         laneRequestSinkWire_7_bits_decodeResult_sWrite = queue_7_deq_bits_decodeResult_sWrite;
  wire         laneRequestSinkWire_7_bits_decodeResult_crossRead = queue_7_deq_bits_decodeResult_crossRead;
  wire         laneRequestSinkWire_7_bits_decodeResult_crossWrite = queue_7_deq_bits_decodeResult_crossWrite;
  wire         laneRequestSinkWire_7_bits_decodeResult_maskUnit = queue_7_deq_bits_decodeResult_maskUnit;
  wire         laneRequestSinkWire_7_bits_decodeResult_special = queue_7_deq_bits_decodeResult_special;
  wire         laneRequestSinkWire_7_bits_decodeResult_saturate = queue_7_deq_bits_decodeResult_saturate;
  wire         laneRequestSinkWire_7_bits_decodeResult_vwmacc = queue_7_deq_bits_decodeResult_vwmacc;
  wire         laneRequestSinkWire_7_bits_decodeResult_readOnly = queue_7_deq_bits_decodeResult_readOnly;
  wire         laneRequestSinkWire_7_bits_decodeResult_maskSource = queue_7_deq_bits_decodeResult_maskSource;
  wire         laneRequestSinkWire_7_bits_decodeResult_maskDestination = queue_7_deq_bits_decodeResult_maskDestination;
  wire         laneRequestSinkWire_7_bits_decodeResult_maskLogic = queue_7_deq_bits_decodeResult_maskLogic;
  wire [3:0]   laneRequestSinkWire_7_bits_decodeResult_uop = queue_7_deq_bits_decodeResult_uop;
  wire         laneRequestSinkWire_7_bits_decodeResult_iota = queue_7_deq_bits_decodeResult_iota;
  wire         laneRequestSinkWire_7_bits_decodeResult_mv = queue_7_deq_bits_decodeResult_mv;
  wire         laneRequestSinkWire_7_bits_decodeResult_extend = queue_7_deq_bits_decodeResult_extend;
  wire         laneRequestSinkWire_7_bits_decodeResult_unOrderWrite = queue_7_deq_bits_decodeResult_unOrderWrite;
  wire         laneRequestSinkWire_7_bits_decodeResult_compress = queue_7_deq_bits_decodeResult_compress;
  wire         laneRequestSinkWire_7_bits_decodeResult_gather16 = queue_7_deq_bits_decodeResult_gather16;
  wire         laneRequestSinkWire_7_bits_decodeResult_gather = queue_7_deq_bits_decodeResult_gather;
  wire         laneRequestSinkWire_7_bits_decodeResult_slid = queue_7_deq_bits_decodeResult_slid;
  wire         laneRequestSinkWire_7_bits_decodeResult_targetRd = queue_7_deq_bits_decodeResult_targetRd;
  wire         laneRequestSinkWire_7_bits_decodeResult_widenReduce = queue_7_deq_bits_decodeResult_widenReduce;
  wire         laneRequestSinkWire_7_bits_decodeResult_red = queue_7_deq_bits_decodeResult_red;
  wire         laneRequestSinkWire_7_bits_decodeResult_nr = queue_7_deq_bits_decodeResult_nr;
  wire         laneRequestSinkWire_7_bits_decodeResult_itype = queue_7_deq_bits_decodeResult_itype;
  wire         laneRequestSinkWire_7_bits_decodeResult_unsigned1 = queue_7_deq_bits_decodeResult_unsigned1;
  wire         laneRequestSinkWire_7_bits_decodeResult_unsigned0 = queue_7_deq_bits_decodeResult_unsigned0;
  wire         laneRequestSinkWire_7_bits_decodeResult_other = queue_7_deq_bits_decodeResult_other;
  wire         laneRequestSinkWire_7_bits_decodeResult_multiCycle = queue_7_deq_bits_decodeResult_multiCycle;
  wire         laneRequestSinkWire_7_bits_decodeResult_divider = queue_7_deq_bits_decodeResult_divider;
  wire         laneRequestSinkWire_7_bits_decodeResult_multiplier = queue_7_deq_bits_decodeResult_multiplier;
  wire         laneRequestSinkWire_7_bits_decodeResult_shift = queue_7_deq_bits_decodeResult_shift;
  wire         laneRequestSinkWire_7_bits_decodeResult_adder = queue_7_deq_bits_decodeResult_adder;
  wire         laneRequestSinkWire_7_bits_decodeResult_logic = queue_7_deq_bits_decodeResult_logic;
  wire         laneRequestSinkWire_7_bits_loadStore = queue_7_deq_bits_loadStore;
  wire         laneRequestSinkWire_7_bits_issueInst = queue_7_deq_bits_issueInst;
  wire         laneRequestSinkWire_7_bits_store = queue_7_deq_bits_store;
  wire         laneRequestSinkWire_7_bits_special = queue_7_deq_bits_special;
  wire         laneRequestSinkWire_7_bits_lsWholeReg = queue_7_deq_bits_lsWholeReg;
  wire [4:0]   laneRequestSinkWire_7_bits_vs1 = queue_7_deq_bits_vs1;
  wire [4:0]   laneRequestSinkWire_7_bits_vs2 = queue_7_deq_bits_vs2;
  wire [4:0]   laneRequestSinkWire_7_bits_vd = queue_7_deq_bits_vd;
  wire [1:0]   laneRequestSinkWire_7_bits_loadStoreEEW = queue_7_deq_bits_loadStoreEEW;
  wire         laneRequestSinkWire_7_bits_mask = queue_7_deq_bits_mask;
  wire [2:0]   laneRequestSinkWire_7_bits_segment = queue_7_deq_bits_segment;
  wire [31:0]  laneRequestSinkWire_7_bits_readFromScalar = queue_7_deq_bits_readFromScalar;
  wire [11:0]  laneRequestSinkWire_7_bits_csrInterface_vl = queue_7_deq_bits_csrInterface_vl;
  wire [11:0]  laneRequestSinkWire_7_bits_csrInterface_vStart = queue_7_deq_bits_csrInterface_vStart;
  wire [2:0]   laneRequestSinkWire_7_bits_csrInterface_vlmul = queue_7_deq_bits_csrInterface_vlmul;
  wire [1:0]   laneRequestSinkWire_7_bits_csrInterface_vSew = queue_7_deq_bits_csrInterface_vSew;
  wire [1:0]   laneRequestSinkWire_7_bits_csrInterface_vxrm = queue_7_deq_bits_csrInterface_vxrm;
  wire         laneRequestSinkWire_7_bits_csrInterface_vta = queue_7_deq_bits_csrInterface_vta;
  wire         laneRequestSinkWire_7_bits_csrInterface_vma = queue_7_deq_bits_csrInterface_vma;
  wire [1:0]   queue_7_enq_bits_csrInterface_vxrm;
  wire         queue_7_enq_bits_csrInterface_vta;
  wire [2:0]   queue_dataIn_lo_hi_21 = {queue_7_enq_bits_csrInterface_vxrm, queue_7_enq_bits_csrInterface_vta};
  wire         queue_7_enq_bits_csrInterface_vma;
  wire [3:0]   queue_dataIn_lo_21 = {queue_dataIn_lo_hi_21, queue_7_enq_bits_csrInterface_vma};
  wire [2:0]   queue_7_enq_bits_csrInterface_vlmul;
  wire [1:0]   queue_7_enq_bits_csrInterface_vSew;
  wire [4:0]   queue_dataIn_hi_lo_21 = {queue_7_enq_bits_csrInterface_vlmul, queue_7_enq_bits_csrInterface_vSew};
  wire [11:0]  queue_7_enq_bits_csrInterface_vl;
  wire [11:0]  queue_7_enq_bits_csrInterface_vStart;
  wire [23:0]  queue_dataIn_hi_hi_21 = {queue_7_enq_bits_csrInterface_vl, queue_7_enq_bits_csrInterface_vStart};
  wire [28:0]  queue_dataIn_hi_21 = {queue_dataIn_hi_hi_21, queue_dataIn_hi_lo_21};
  wire         queue_7_enq_bits_decodeResult_adder;
  wire         queue_7_enq_bits_decodeResult_logic;
  wire [1:0]   queue_dataIn_lo_lo_lo_lo_7 = {queue_7_enq_bits_decodeResult_adder, queue_7_enq_bits_decodeResult_logic};
  wire         queue_7_enq_bits_decodeResult_divider;
  wire         queue_7_enq_bits_decodeResult_multiplier;
  wire [1:0]   queue_dataIn_lo_lo_lo_hi_hi_7 = {queue_7_enq_bits_decodeResult_divider, queue_7_enq_bits_decodeResult_multiplier};
  wire         queue_7_enq_bits_decodeResult_shift;
  wire [2:0]   queue_dataIn_lo_lo_lo_hi_7 = {queue_dataIn_lo_lo_lo_hi_hi_7, queue_7_enq_bits_decodeResult_shift};
  wire [4:0]   queue_dataIn_lo_lo_lo_7 = {queue_dataIn_lo_lo_lo_hi_7, queue_dataIn_lo_lo_lo_lo_7};
  wire         queue_7_enq_bits_decodeResult_unsigned0;
  wire         queue_7_enq_bits_decodeResult_other;
  wire [1:0]   queue_dataIn_lo_lo_hi_lo_hi_7 = {queue_7_enq_bits_decodeResult_unsigned0, queue_7_enq_bits_decodeResult_other};
  wire         queue_7_enq_bits_decodeResult_multiCycle;
  wire [2:0]   queue_dataIn_lo_lo_hi_lo_7 = {queue_dataIn_lo_lo_hi_lo_hi_7, queue_7_enq_bits_decodeResult_multiCycle};
  wire         queue_7_enq_bits_decodeResult_nr;
  wire         queue_7_enq_bits_decodeResult_itype;
  wire [1:0]   queue_dataIn_lo_lo_hi_hi_hi_7 = {queue_7_enq_bits_decodeResult_nr, queue_7_enq_bits_decodeResult_itype};
  wire         queue_7_enq_bits_decodeResult_unsigned1;
  wire [2:0]   queue_dataIn_lo_lo_hi_hi_7 = {queue_dataIn_lo_lo_hi_hi_hi_7, queue_7_enq_bits_decodeResult_unsigned1};
  wire [5:0]   queue_dataIn_lo_lo_hi_14 = {queue_dataIn_lo_lo_hi_hi_7, queue_dataIn_lo_lo_hi_lo_7};
  wire [10:0]  queue_dataIn_lo_lo_14 = {queue_dataIn_lo_lo_hi_14, queue_dataIn_lo_lo_lo_7};
  wire         queue_7_enq_bits_decodeResult_widenReduce;
  wire         queue_7_enq_bits_decodeResult_red;
  wire [1:0]   queue_dataIn_lo_hi_lo_lo_7 = {queue_7_enq_bits_decodeResult_widenReduce, queue_7_enq_bits_decodeResult_red};
  wire         queue_7_enq_bits_decodeResult_gather;
  wire         queue_7_enq_bits_decodeResult_slid;
  wire [1:0]   queue_dataIn_lo_hi_lo_hi_hi_7 = {queue_7_enq_bits_decodeResult_gather, queue_7_enq_bits_decodeResult_slid};
  wire         queue_7_enq_bits_decodeResult_targetRd;
  wire [2:0]   queue_dataIn_lo_hi_lo_hi_7 = {queue_dataIn_lo_hi_lo_hi_hi_7, queue_7_enq_bits_decodeResult_targetRd};
  wire [4:0]   queue_dataIn_lo_hi_lo_14 = {queue_dataIn_lo_hi_lo_hi_7, queue_dataIn_lo_hi_lo_lo_7};
  wire         queue_7_enq_bits_decodeResult_unOrderWrite;
  wire         queue_7_enq_bits_decodeResult_compress;
  wire [1:0]   queue_dataIn_lo_hi_hi_lo_hi_7 = {queue_7_enq_bits_decodeResult_unOrderWrite, queue_7_enq_bits_decodeResult_compress};
  wire         queue_7_enq_bits_decodeResult_gather16;
  wire [2:0]   queue_dataIn_lo_hi_hi_lo_7 = {queue_dataIn_lo_hi_hi_lo_hi_7, queue_7_enq_bits_decodeResult_gather16};
  wire         queue_7_enq_bits_decodeResult_iota;
  wire         queue_7_enq_bits_decodeResult_mv;
  wire [1:0]   queue_dataIn_lo_hi_hi_hi_hi_7 = {queue_7_enq_bits_decodeResult_iota, queue_7_enq_bits_decodeResult_mv};
  wire         queue_7_enq_bits_decodeResult_extend;
  wire [2:0]   queue_dataIn_lo_hi_hi_hi_7 = {queue_dataIn_lo_hi_hi_hi_hi_7, queue_7_enq_bits_decodeResult_extend};
  wire [5:0]   queue_dataIn_lo_hi_hi_14 = {queue_dataIn_lo_hi_hi_hi_7, queue_dataIn_lo_hi_hi_lo_7};
  wire [10:0]  queue_dataIn_lo_hi_22 = {queue_dataIn_lo_hi_hi_14, queue_dataIn_lo_hi_lo_14};
  wire [21:0]  queue_dataIn_lo_22 = {queue_dataIn_lo_hi_22, queue_dataIn_lo_lo_14};
  wire         queue_7_enq_bits_decodeResult_maskLogic;
  wire [3:0]   queue_7_enq_bits_decodeResult_uop;
  wire [4:0]   queue_dataIn_hi_lo_lo_lo_7 = {queue_7_enq_bits_decodeResult_maskLogic, queue_7_enq_bits_decodeResult_uop};
  wire         queue_7_enq_bits_decodeResult_readOnly;
  wire         queue_7_enq_bits_decodeResult_maskSource;
  wire [1:0]   queue_dataIn_hi_lo_lo_hi_hi_7 = {queue_7_enq_bits_decodeResult_readOnly, queue_7_enq_bits_decodeResult_maskSource};
  wire         queue_7_enq_bits_decodeResult_maskDestination;
  wire [2:0]   queue_dataIn_hi_lo_lo_hi_7 = {queue_dataIn_hi_lo_lo_hi_hi_7, queue_7_enq_bits_decodeResult_maskDestination};
  wire [7:0]   queue_dataIn_hi_lo_lo_14 = {queue_dataIn_hi_lo_lo_hi_7, queue_dataIn_hi_lo_lo_lo_7};
  wire         queue_7_enq_bits_decodeResult_special;
  wire         queue_7_enq_bits_decodeResult_saturate;
  wire [1:0]   queue_dataIn_hi_lo_hi_lo_hi_7 = {queue_7_enq_bits_decodeResult_special, queue_7_enq_bits_decodeResult_saturate};
  wire         queue_7_enq_bits_decodeResult_vwmacc;
  wire [2:0]   queue_dataIn_hi_lo_hi_lo_7 = {queue_dataIn_hi_lo_hi_lo_hi_7, queue_7_enq_bits_decodeResult_vwmacc};
  wire         queue_7_enq_bits_decodeResult_crossRead;
  wire         queue_7_enq_bits_decodeResult_crossWrite;
  wire [1:0]   queue_dataIn_hi_lo_hi_hi_hi_7 = {queue_7_enq_bits_decodeResult_crossRead, queue_7_enq_bits_decodeResult_crossWrite};
  wire         queue_7_enq_bits_decodeResult_maskUnit;
  wire [2:0]   queue_dataIn_hi_lo_hi_hi_7 = {queue_dataIn_hi_lo_hi_hi_hi_7, queue_7_enq_bits_decodeResult_maskUnit};
  wire [5:0]   queue_dataIn_hi_lo_hi_14 = {queue_dataIn_hi_lo_hi_hi_7, queue_dataIn_hi_lo_hi_lo_7};
  wire [13:0]  queue_dataIn_hi_lo_22 = {queue_dataIn_hi_lo_hi_14, queue_dataIn_hi_lo_lo_14};
  wire         queue_7_enq_bits_decodeResult_vtype;
  wire         queue_7_enq_bits_decodeResult_sWrite;
  wire [1:0]   queue_dataIn_hi_hi_lo_lo_7 = {queue_7_enq_bits_decodeResult_vtype, queue_7_enq_bits_decodeResult_sWrite};
  wire         queue_7_enq_bits_decodeResult_dontNeedExecuteInLane;
  wire         queue_7_enq_bits_decodeResult_scheduler;
  wire [1:0]   queue_dataIn_hi_hi_lo_hi_hi_7 = {queue_7_enq_bits_decodeResult_dontNeedExecuteInLane, queue_7_enq_bits_decodeResult_scheduler};
  wire         queue_7_enq_bits_decodeResult_sReadVD;
  wire [2:0]   queue_dataIn_hi_hi_lo_hi_7 = {queue_dataIn_hi_hi_lo_hi_hi_7, queue_7_enq_bits_decodeResult_sReadVD};
  wire [4:0]   queue_dataIn_hi_hi_lo_14 = {queue_dataIn_hi_hi_lo_hi_7, queue_dataIn_hi_hi_lo_lo_7};
  wire         queue_7_enq_bits_decodeResult_ffo;
  wire         queue_7_enq_bits_decodeResult_average;
  wire [1:0]   queue_dataIn_hi_hi_hi_lo_hi_7 = {queue_7_enq_bits_decodeResult_ffo, queue_7_enq_bits_decodeResult_average};
  wire         queue_7_enq_bits_decodeResult_reverse;
  wire [2:0]   queue_dataIn_hi_hi_hi_lo_7 = {queue_dataIn_hi_hi_hi_lo_hi_7, queue_7_enq_bits_decodeResult_reverse};
  wire         queue_7_enq_bits_decodeResult_specialSlot;
  wire [4:0]   queue_7_enq_bits_decodeResult_topUop;
  wire [5:0]   queue_dataIn_hi_hi_hi_hi_hi_7 = {queue_7_enq_bits_decodeResult_specialSlot, queue_7_enq_bits_decodeResult_topUop};
  wire         queue_7_enq_bits_decodeResult_popCount;
  wire [6:0]   queue_dataIn_hi_hi_hi_hi_7 = {queue_dataIn_hi_hi_hi_hi_hi_7, queue_7_enq_bits_decodeResult_popCount};
  wire [9:0]   queue_dataIn_hi_hi_hi_14 = {queue_dataIn_hi_hi_hi_hi_7, queue_dataIn_hi_hi_hi_lo_7};
  wire [14:0]  queue_dataIn_hi_hi_22 = {queue_dataIn_hi_hi_hi_14, queue_dataIn_hi_hi_lo_14};
  wire [28:0]  queue_dataIn_hi_22 = {queue_dataIn_hi_hi_22, queue_dataIn_hi_lo_22};
  wire [2:0]   queue_7_enq_bits_segment;
  wire [31:0]  queue_7_enq_bits_readFromScalar;
  wire [34:0]  queue_dataIn_lo_lo_hi_15 = {queue_7_enq_bits_segment, queue_7_enq_bits_readFromScalar};
  wire [67:0]  queue_dataIn_lo_lo_15 = {queue_dataIn_lo_lo_hi_15, queue_dataIn_hi_21, queue_dataIn_lo_21};
  wire [1:0]   queue_7_enq_bits_loadStoreEEW;
  wire         queue_7_enq_bits_mask;
  wire [2:0]   queue_dataIn_lo_hi_lo_15 = {queue_7_enq_bits_loadStoreEEW, queue_7_enq_bits_mask};
  wire [4:0]   queue_7_enq_bits_vs2;
  wire [4:0]   queue_7_enq_bits_vd;
  wire [9:0]   queue_dataIn_lo_hi_hi_15 = {queue_7_enq_bits_vs2, queue_7_enq_bits_vd};
  wire [12:0]  queue_dataIn_lo_hi_23 = {queue_dataIn_lo_hi_hi_15, queue_dataIn_lo_hi_lo_15};
  wire [80:0]  queue_dataIn_lo_23 = {queue_dataIn_lo_hi_23, queue_dataIn_lo_lo_15};
  wire         queue_7_enq_bits_lsWholeReg;
  wire [4:0]   queue_7_enq_bits_vs1;
  wire [5:0]   queue_dataIn_hi_lo_lo_15 = {queue_7_enq_bits_lsWholeReg, queue_7_enq_bits_vs1};
  wire         queue_7_enq_bits_store;
  wire         queue_7_enq_bits_special;
  wire [1:0]   queue_dataIn_hi_lo_hi_15 = {queue_7_enq_bits_store, queue_7_enq_bits_special};
  wire [7:0]   queue_dataIn_hi_lo_23 = {queue_dataIn_hi_lo_hi_15, queue_dataIn_hi_lo_lo_15};
  wire         queue_7_enq_bits_loadStore;
  wire         queue_7_enq_bits_issueInst;
  wire [1:0]   queue_dataIn_hi_hi_lo_15 = {queue_7_enq_bits_loadStore, queue_7_enq_bits_issueInst};
  wire [2:0]   queue_7_enq_bits_instructionIndex;
  wire [53:0]  queue_dataIn_hi_hi_hi_15 = {queue_7_enq_bits_instructionIndex, queue_dataIn_hi_22, queue_dataIn_lo_22};
  wire [55:0]  queue_dataIn_hi_hi_23 = {queue_dataIn_hi_hi_hi_15, queue_dataIn_hi_hi_lo_15};
  wire [63:0]  queue_dataIn_hi_23 = {queue_dataIn_hi_hi_23, queue_dataIn_hi_lo_23};
  wire [144:0] queue_dataIn_7 = {queue_dataIn_hi_23, queue_dataIn_lo_23};
  wire         queue_dataOut_7_csrInterface_vma = _queue_fifo_7_data_out[0];
  wire         queue_dataOut_7_csrInterface_vta = _queue_fifo_7_data_out[1];
  wire [1:0]   queue_dataOut_7_csrInterface_vxrm = _queue_fifo_7_data_out[3:2];
  wire [1:0]   queue_dataOut_7_csrInterface_vSew = _queue_fifo_7_data_out[5:4];
  wire [2:0]   queue_dataOut_7_csrInterface_vlmul = _queue_fifo_7_data_out[8:6];
  wire [11:0]  queue_dataOut_7_csrInterface_vStart = _queue_fifo_7_data_out[20:9];
  wire [11:0]  queue_dataOut_7_csrInterface_vl = _queue_fifo_7_data_out[32:21];
  wire [31:0]  queue_dataOut_7_readFromScalar = _queue_fifo_7_data_out[64:33];
  wire [2:0]   queue_dataOut_7_segment = _queue_fifo_7_data_out[67:65];
  wire         queue_dataOut_7_mask = _queue_fifo_7_data_out[68];
  wire [1:0]   queue_dataOut_7_loadStoreEEW = _queue_fifo_7_data_out[70:69];
  wire [4:0]   queue_dataOut_7_vd = _queue_fifo_7_data_out[75:71];
  wire [4:0]   queue_dataOut_7_vs2 = _queue_fifo_7_data_out[80:76];
  wire [4:0]   queue_dataOut_7_vs1 = _queue_fifo_7_data_out[85:81];
  wire         queue_dataOut_7_lsWholeReg = _queue_fifo_7_data_out[86];
  wire         queue_dataOut_7_special = _queue_fifo_7_data_out[87];
  wire         queue_dataOut_7_store = _queue_fifo_7_data_out[88];
  wire         queue_dataOut_7_issueInst = _queue_fifo_7_data_out[89];
  wire         queue_dataOut_7_loadStore = _queue_fifo_7_data_out[90];
  wire         queue_dataOut_7_decodeResult_logic = _queue_fifo_7_data_out[91];
  wire         queue_dataOut_7_decodeResult_adder = _queue_fifo_7_data_out[92];
  wire         queue_dataOut_7_decodeResult_shift = _queue_fifo_7_data_out[93];
  wire         queue_dataOut_7_decodeResult_multiplier = _queue_fifo_7_data_out[94];
  wire         queue_dataOut_7_decodeResult_divider = _queue_fifo_7_data_out[95];
  wire         queue_dataOut_7_decodeResult_multiCycle = _queue_fifo_7_data_out[96];
  wire         queue_dataOut_7_decodeResult_other = _queue_fifo_7_data_out[97];
  wire         queue_dataOut_7_decodeResult_unsigned0 = _queue_fifo_7_data_out[98];
  wire         queue_dataOut_7_decodeResult_unsigned1 = _queue_fifo_7_data_out[99];
  wire         queue_dataOut_7_decodeResult_itype = _queue_fifo_7_data_out[100];
  wire         queue_dataOut_7_decodeResult_nr = _queue_fifo_7_data_out[101];
  wire         queue_dataOut_7_decodeResult_red = _queue_fifo_7_data_out[102];
  wire         queue_dataOut_7_decodeResult_widenReduce = _queue_fifo_7_data_out[103];
  wire         queue_dataOut_7_decodeResult_targetRd = _queue_fifo_7_data_out[104];
  wire         queue_dataOut_7_decodeResult_slid = _queue_fifo_7_data_out[105];
  wire         queue_dataOut_7_decodeResult_gather = _queue_fifo_7_data_out[106];
  wire         queue_dataOut_7_decodeResult_gather16 = _queue_fifo_7_data_out[107];
  wire         queue_dataOut_7_decodeResult_compress = _queue_fifo_7_data_out[108];
  wire         queue_dataOut_7_decodeResult_unOrderWrite = _queue_fifo_7_data_out[109];
  wire         queue_dataOut_7_decodeResult_extend = _queue_fifo_7_data_out[110];
  wire         queue_dataOut_7_decodeResult_mv = _queue_fifo_7_data_out[111];
  wire         queue_dataOut_7_decodeResult_iota = _queue_fifo_7_data_out[112];
  wire [3:0]   queue_dataOut_7_decodeResult_uop = _queue_fifo_7_data_out[116:113];
  wire         queue_dataOut_7_decodeResult_maskLogic = _queue_fifo_7_data_out[117];
  wire         queue_dataOut_7_decodeResult_maskDestination = _queue_fifo_7_data_out[118];
  wire         queue_dataOut_7_decodeResult_maskSource = _queue_fifo_7_data_out[119];
  wire         queue_dataOut_7_decodeResult_readOnly = _queue_fifo_7_data_out[120];
  wire         queue_dataOut_7_decodeResult_vwmacc = _queue_fifo_7_data_out[121];
  wire         queue_dataOut_7_decodeResult_saturate = _queue_fifo_7_data_out[122];
  wire         queue_dataOut_7_decodeResult_special = _queue_fifo_7_data_out[123];
  wire         queue_dataOut_7_decodeResult_maskUnit = _queue_fifo_7_data_out[124];
  wire         queue_dataOut_7_decodeResult_crossWrite = _queue_fifo_7_data_out[125];
  wire         queue_dataOut_7_decodeResult_crossRead = _queue_fifo_7_data_out[126];
  wire         queue_dataOut_7_decodeResult_sWrite = _queue_fifo_7_data_out[127];
  wire         queue_dataOut_7_decodeResult_vtype = _queue_fifo_7_data_out[128];
  wire         queue_dataOut_7_decodeResult_sReadVD = _queue_fifo_7_data_out[129];
  wire         queue_dataOut_7_decodeResult_scheduler = _queue_fifo_7_data_out[130];
  wire         queue_dataOut_7_decodeResult_dontNeedExecuteInLane = _queue_fifo_7_data_out[131];
  wire         queue_dataOut_7_decodeResult_reverse = _queue_fifo_7_data_out[132];
  wire         queue_dataOut_7_decodeResult_average = _queue_fifo_7_data_out[133];
  wire         queue_dataOut_7_decodeResult_ffo = _queue_fifo_7_data_out[134];
  wire         queue_dataOut_7_decodeResult_popCount = _queue_fifo_7_data_out[135];
  wire [4:0]   queue_dataOut_7_decodeResult_topUop = _queue_fifo_7_data_out[140:136];
  wire         queue_dataOut_7_decodeResult_specialSlot = _queue_fifo_7_data_out[141];
  wire [2:0]   queue_dataOut_7_instructionIndex = _queue_fifo_7_data_out[144:142];
  wire         queue_7_enq_ready = ~_queue_fifo_7_full;
  wire         queue_7_enq_valid;
  assign queue_7_deq_valid = ~_queue_fifo_7_empty | queue_7_enq_valid;
  assign queue_7_deq_bits_instructionIndex = _queue_fifo_7_empty ? queue_7_enq_bits_instructionIndex : queue_dataOut_7_instructionIndex;
  assign queue_7_deq_bits_decodeResult_specialSlot = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_specialSlot : queue_dataOut_7_decodeResult_specialSlot;
  assign queue_7_deq_bits_decodeResult_topUop = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_topUop : queue_dataOut_7_decodeResult_topUop;
  assign queue_7_deq_bits_decodeResult_popCount = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_popCount : queue_dataOut_7_decodeResult_popCount;
  assign queue_7_deq_bits_decodeResult_ffo = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_ffo : queue_dataOut_7_decodeResult_ffo;
  assign queue_7_deq_bits_decodeResult_average = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_average : queue_dataOut_7_decodeResult_average;
  assign queue_7_deq_bits_decodeResult_reverse = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_reverse : queue_dataOut_7_decodeResult_reverse;
  assign queue_7_deq_bits_decodeResult_dontNeedExecuteInLane = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_dontNeedExecuteInLane : queue_dataOut_7_decodeResult_dontNeedExecuteInLane;
  assign queue_7_deq_bits_decodeResult_scheduler = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_scheduler : queue_dataOut_7_decodeResult_scheduler;
  assign queue_7_deq_bits_decodeResult_sReadVD = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_sReadVD : queue_dataOut_7_decodeResult_sReadVD;
  assign queue_7_deq_bits_decodeResult_vtype = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_vtype : queue_dataOut_7_decodeResult_vtype;
  assign queue_7_deq_bits_decodeResult_sWrite = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_sWrite : queue_dataOut_7_decodeResult_sWrite;
  assign queue_7_deq_bits_decodeResult_crossRead = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_crossRead : queue_dataOut_7_decodeResult_crossRead;
  assign queue_7_deq_bits_decodeResult_crossWrite = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_crossWrite : queue_dataOut_7_decodeResult_crossWrite;
  assign queue_7_deq_bits_decodeResult_maskUnit = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_maskUnit : queue_dataOut_7_decodeResult_maskUnit;
  assign queue_7_deq_bits_decodeResult_special = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_special : queue_dataOut_7_decodeResult_special;
  assign queue_7_deq_bits_decodeResult_saturate = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_saturate : queue_dataOut_7_decodeResult_saturate;
  assign queue_7_deq_bits_decodeResult_vwmacc = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_vwmacc : queue_dataOut_7_decodeResult_vwmacc;
  assign queue_7_deq_bits_decodeResult_readOnly = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_readOnly : queue_dataOut_7_decodeResult_readOnly;
  assign queue_7_deq_bits_decodeResult_maskSource = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_maskSource : queue_dataOut_7_decodeResult_maskSource;
  assign queue_7_deq_bits_decodeResult_maskDestination = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_maskDestination : queue_dataOut_7_decodeResult_maskDestination;
  assign queue_7_deq_bits_decodeResult_maskLogic = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_maskLogic : queue_dataOut_7_decodeResult_maskLogic;
  assign queue_7_deq_bits_decodeResult_uop = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_uop : queue_dataOut_7_decodeResult_uop;
  assign queue_7_deq_bits_decodeResult_iota = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_iota : queue_dataOut_7_decodeResult_iota;
  assign queue_7_deq_bits_decodeResult_mv = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_mv : queue_dataOut_7_decodeResult_mv;
  assign queue_7_deq_bits_decodeResult_extend = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_extend : queue_dataOut_7_decodeResult_extend;
  assign queue_7_deq_bits_decodeResult_unOrderWrite = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_unOrderWrite : queue_dataOut_7_decodeResult_unOrderWrite;
  assign queue_7_deq_bits_decodeResult_compress = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_compress : queue_dataOut_7_decodeResult_compress;
  assign queue_7_deq_bits_decodeResult_gather16 = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_gather16 : queue_dataOut_7_decodeResult_gather16;
  assign queue_7_deq_bits_decodeResult_gather = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_gather : queue_dataOut_7_decodeResult_gather;
  assign queue_7_deq_bits_decodeResult_slid = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_slid : queue_dataOut_7_decodeResult_slid;
  assign queue_7_deq_bits_decodeResult_targetRd = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_targetRd : queue_dataOut_7_decodeResult_targetRd;
  assign queue_7_deq_bits_decodeResult_widenReduce = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_widenReduce : queue_dataOut_7_decodeResult_widenReduce;
  assign queue_7_deq_bits_decodeResult_red = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_red : queue_dataOut_7_decodeResult_red;
  assign queue_7_deq_bits_decodeResult_nr = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_nr : queue_dataOut_7_decodeResult_nr;
  assign queue_7_deq_bits_decodeResult_itype = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_itype : queue_dataOut_7_decodeResult_itype;
  assign queue_7_deq_bits_decodeResult_unsigned1 = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_unsigned1 : queue_dataOut_7_decodeResult_unsigned1;
  assign queue_7_deq_bits_decodeResult_unsigned0 = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_unsigned0 : queue_dataOut_7_decodeResult_unsigned0;
  assign queue_7_deq_bits_decodeResult_other = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_other : queue_dataOut_7_decodeResult_other;
  assign queue_7_deq_bits_decodeResult_multiCycle = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_multiCycle : queue_dataOut_7_decodeResult_multiCycle;
  assign queue_7_deq_bits_decodeResult_divider = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_divider : queue_dataOut_7_decodeResult_divider;
  assign queue_7_deq_bits_decodeResult_multiplier = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_multiplier : queue_dataOut_7_decodeResult_multiplier;
  assign queue_7_deq_bits_decodeResult_shift = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_shift : queue_dataOut_7_decodeResult_shift;
  assign queue_7_deq_bits_decodeResult_adder = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_adder : queue_dataOut_7_decodeResult_adder;
  assign queue_7_deq_bits_decodeResult_logic = _queue_fifo_7_empty ? queue_7_enq_bits_decodeResult_logic : queue_dataOut_7_decodeResult_logic;
  assign queue_7_deq_bits_loadStore = _queue_fifo_7_empty ? queue_7_enq_bits_loadStore : queue_dataOut_7_loadStore;
  assign queue_7_deq_bits_issueInst = _queue_fifo_7_empty ? queue_7_enq_bits_issueInst : queue_dataOut_7_issueInst;
  assign queue_7_deq_bits_store = _queue_fifo_7_empty ? queue_7_enq_bits_store : queue_dataOut_7_store;
  assign queue_7_deq_bits_special = _queue_fifo_7_empty ? queue_7_enq_bits_special : queue_dataOut_7_special;
  assign queue_7_deq_bits_lsWholeReg = _queue_fifo_7_empty ? queue_7_enq_bits_lsWholeReg : queue_dataOut_7_lsWholeReg;
  assign queue_7_deq_bits_vs1 = _queue_fifo_7_empty ? queue_7_enq_bits_vs1 : queue_dataOut_7_vs1;
  assign queue_7_deq_bits_vs2 = _queue_fifo_7_empty ? queue_7_enq_bits_vs2 : queue_dataOut_7_vs2;
  assign queue_7_deq_bits_vd = _queue_fifo_7_empty ? queue_7_enq_bits_vd : queue_dataOut_7_vd;
  assign queue_7_deq_bits_loadStoreEEW = _queue_fifo_7_empty ? queue_7_enq_bits_loadStoreEEW : queue_dataOut_7_loadStoreEEW;
  assign queue_7_deq_bits_mask = _queue_fifo_7_empty ? queue_7_enq_bits_mask : queue_dataOut_7_mask;
  assign queue_7_deq_bits_segment = _queue_fifo_7_empty ? queue_7_enq_bits_segment : queue_dataOut_7_segment;
  assign queue_7_deq_bits_readFromScalar = _queue_fifo_7_empty ? queue_7_enq_bits_readFromScalar : queue_dataOut_7_readFromScalar;
  assign queue_7_deq_bits_csrInterface_vl = _queue_fifo_7_empty ? queue_7_enq_bits_csrInterface_vl : queue_dataOut_7_csrInterface_vl;
  assign queue_7_deq_bits_csrInterface_vStart = _queue_fifo_7_empty ? queue_7_enq_bits_csrInterface_vStart : queue_dataOut_7_csrInterface_vStart;
  assign queue_7_deq_bits_csrInterface_vlmul = _queue_fifo_7_empty ? queue_7_enq_bits_csrInterface_vlmul : queue_dataOut_7_csrInterface_vlmul;
  assign queue_7_deq_bits_csrInterface_vSew = _queue_fifo_7_empty ? queue_7_enq_bits_csrInterface_vSew : queue_dataOut_7_csrInterface_vSew;
  assign queue_7_deq_bits_csrInterface_vxrm = _queue_fifo_7_empty ? queue_7_enq_bits_csrInterface_vxrm : queue_dataOut_7_csrInterface_vxrm;
  assign queue_7_deq_bits_csrInterface_vta = _queue_fifo_7_empty ? queue_7_enq_bits_csrInterface_vta : queue_dataOut_7_csrInterface_vta;
  assign queue_7_deq_bits_csrInterface_vma = _queue_fifo_7_empty ? queue_7_enq_bits_csrInterface_vma : queue_dataOut_7_csrInterface_vma;
  wire         laneVec_7_laneRequest_bits_issueInst = laneRequestSinkWire_7_ready & laneRequestSinkWire_7_valid;
  reg          releasePipe_pipe_v_7;
  wire         releasePipe_pipe_out_7_valid = releasePipe_pipe_v_7;
  wire         laneRequestSourceWire_7_ready;
  wire         validSource_7_valid = laneRequestSourceWire_7_ready & laneRequestSourceWire_7_valid;
  reg  [2:0]   tokenCheck_counter_7;
  wire [2:0]   tokenCheck_counterChange_7 = validSource_7_valid ? 3'h1 : 3'h7;
  assign tokenCheck_7 = ~(tokenCheck_counter_7[2]);
  assign laneRequestSourceWire_7_ready = tokenCheck_7;
  assign queue_7_enq_valid = validSink_7_valid;
  assign queue_7_enq_bits_instructionIndex = validSink_7_bits_instructionIndex;
  assign queue_7_enq_bits_decodeResult_specialSlot = validSink_7_bits_decodeResult_specialSlot;
  assign queue_7_enq_bits_decodeResult_topUop = validSink_7_bits_decodeResult_topUop;
  assign queue_7_enq_bits_decodeResult_popCount = validSink_7_bits_decodeResult_popCount;
  assign queue_7_enq_bits_decodeResult_ffo = validSink_7_bits_decodeResult_ffo;
  assign queue_7_enq_bits_decodeResult_average = validSink_7_bits_decodeResult_average;
  assign queue_7_enq_bits_decodeResult_reverse = validSink_7_bits_decodeResult_reverse;
  assign queue_7_enq_bits_decodeResult_dontNeedExecuteInLane = validSink_7_bits_decodeResult_dontNeedExecuteInLane;
  assign queue_7_enq_bits_decodeResult_scheduler = validSink_7_bits_decodeResult_scheduler;
  assign queue_7_enq_bits_decodeResult_sReadVD = validSink_7_bits_decodeResult_sReadVD;
  assign queue_7_enq_bits_decodeResult_vtype = validSink_7_bits_decodeResult_vtype;
  assign queue_7_enq_bits_decodeResult_sWrite = validSink_7_bits_decodeResult_sWrite;
  assign queue_7_enq_bits_decodeResult_crossRead = validSink_7_bits_decodeResult_crossRead;
  assign queue_7_enq_bits_decodeResult_crossWrite = validSink_7_bits_decodeResult_crossWrite;
  assign queue_7_enq_bits_decodeResult_maskUnit = validSink_7_bits_decodeResult_maskUnit;
  assign queue_7_enq_bits_decodeResult_special = validSink_7_bits_decodeResult_special;
  assign queue_7_enq_bits_decodeResult_saturate = validSink_7_bits_decodeResult_saturate;
  assign queue_7_enq_bits_decodeResult_vwmacc = validSink_7_bits_decodeResult_vwmacc;
  assign queue_7_enq_bits_decodeResult_readOnly = validSink_7_bits_decodeResult_readOnly;
  assign queue_7_enq_bits_decodeResult_maskSource = validSink_7_bits_decodeResult_maskSource;
  assign queue_7_enq_bits_decodeResult_maskDestination = validSink_7_bits_decodeResult_maskDestination;
  assign queue_7_enq_bits_decodeResult_maskLogic = validSink_7_bits_decodeResult_maskLogic;
  assign queue_7_enq_bits_decodeResult_uop = validSink_7_bits_decodeResult_uop;
  assign queue_7_enq_bits_decodeResult_iota = validSink_7_bits_decodeResult_iota;
  assign queue_7_enq_bits_decodeResult_mv = validSink_7_bits_decodeResult_mv;
  assign queue_7_enq_bits_decodeResult_extend = validSink_7_bits_decodeResult_extend;
  assign queue_7_enq_bits_decodeResult_unOrderWrite = validSink_7_bits_decodeResult_unOrderWrite;
  assign queue_7_enq_bits_decodeResult_compress = validSink_7_bits_decodeResult_compress;
  assign queue_7_enq_bits_decodeResult_gather16 = validSink_7_bits_decodeResult_gather16;
  assign queue_7_enq_bits_decodeResult_gather = validSink_7_bits_decodeResult_gather;
  assign queue_7_enq_bits_decodeResult_slid = validSink_7_bits_decodeResult_slid;
  assign queue_7_enq_bits_decodeResult_targetRd = validSink_7_bits_decodeResult_targetRd;
  assign queue_7_enq_bits_decodeResult_widenReduce = validSink_7_bits_decodeResult_widenReduce;
  assign queue_7_enq_bits_decodeResult_red = validSink_7_bits_decodeResult_red;
  assign queue_7_enq_bits_decodeResult_nr = validSink_7_bits_decodeResult_nr;
  assign queue_7_enq_bits_decodeResult_itype = validSink_7_bits_decodeResult_itype;
  assign queue_7_enq_bits_decodeResult_unsigned1 = validSink_7_bits_decodeResult_unsigned1;
  assign queue_7_enq_bits_decodeResult_unsigned0 = validSink_7_bits_decodeResult_unsigned0;
  assign queue_7_enq_bits_decodeResult_other = validSink_7_bits_decodeResult_other;
  assign queue_7_enq_bits_decodeResult_multiCycle = validSink_7_bits_decodeResult_multiCycle;
  assign queue_7_enq_bits_decodeResult_divider = validSink_7_bits_decodeResult_divider;
  assign queue_7_enq_bits_decodeResult_multiplier = validSink_7_bits_decodeResult_multiplier;
  assign queue_7_enq_bits_decodeResult_shift = validSink_7_bits_decodeResult_shift;
  assign queue_7_enq_bits_decodeResult_adder = validSink_7_bits_decodeResult_adder;
  assign queue_7_enq_bits_decodeResult_logic = validSink_7_bits_decodeResult_logic;
  assign queue_7_enq_bits_loadStore = validSink_7_bits_loadStore;
  assign queue_7_enq_bits_issueInst = validSink_7_bits_issueInst;
  assign queue_7_enq_bits_store = validSink_7_bits_store;
  assign queue_7_enq_bits_special = validSink_7_bits_special;
  assign queue_7_enq_bits_lsWholeReg = validSink_7_bits_lsWholeReg;
  assign queue_7_enq_bits_vs1 = validSink_7_bits_vs1;
  assign queue_7_enq_bits_vs2 = validSink_7_bits_vs2;
  assign queue_7_enq_bits_vd = validSink_7_bits_vd;
  assign queue_7_enq_bits_loadStoreEEW = validSink_7_bits_loadStoreEEW;
  assign queue_7_enq_bits_mask = validSink_7_bits_mask;
  assign queue_7_enq_bits_segment = validSink_7_bits_segment;
  assign queue_7_enq_bits_readFromScalar = validSink_7_bits_readFromScalar;
  assign queue_7_enq_bits_csrInterface_vl = validSink_7_bits_csrInterface_vl;
  assign queue_7_enq_bits_csrInterface_vStart = validSink_7_bits_csrInterface_vStart;
  assign queue_7_enq_bits_csrInterface_vlmul = validSink_7_bits_csrInterface_vlmul;
  assign queue_7_enq_bits_csrInterface_vSew = validSink_7_bits_csrInterface_vSew;
  assign queue_7_enq_bits_csrInterface_vxrm = validSink_7_bits_csrInterface_vxrm;
  assign queue_7_enq_bits_csrInterface_vta = validSink_7_bits_csrInterface_vta;
  assign queue_7_enq_bits_csrInterface_vma = validSink_7_bits_csrInterface_vma;
  reg          shifterReg_7_0_valid;
  assign validSink_7_valid = shifterReg_7_0_valid;
  reg  [2:0]   shifterReg_7_0_bits_instructionIndex;
  assign validSink_7_bits_instructionIndex = shifterReg_7_0_bits_instructionIndex;
  reg          shifterReg_7_0_bits_decodeResult_specialSlot;
  assign validSink_7_bits_decodeResult_specialSlot = shifterReg_7_0_bits_decodeResult_specialSlot;
  reg  [4:0]   shifterReg_7_0_bits_decodeResult_topUop;
  assign validSink_7_bits_decodeResult_topUop = shifterReg_7_0_bits_decodeResult_topUop;
  reg          shifterReg_7_0_bits_decodeResult_popCount;
  assign validSink_7_bits_decodeResult_popCount = shifterReg_7_0_bits_decodeResult_popCount;
  reg          shifterReg_7_0_bits_decodeResult_ffo;
  assign validSink_7_bits_decodeResult_ffo = shifterReg_7_0_bits_decodeResult_ffo;
  reg          shifterReg_7_0_bits_decodeResult_average;
  assign validSink_7_bits_decodeResult_average = shifterReg_7_0_bits_decodeResult_average;
  reg          shifterReg_7_0_bits_decodeResult_reverse;
  assign validSink_7_bits_decodeResult_reverse = shifterReg_7_0_bits_decodeResult_reverse;
  reg          shifterReg_7_0_bits_decodeResult_dontNeedExecuteInLane;
  assign validSink_7_bits_decodeResult_dontNeedExecuteInLane = shifterReg_7_0_bits_decodeResult_dontNeedExecuteInLane;
  reg          shifterReg_7_0_bits_decodeResult_scheduler;
  assign validSink_7_bits_decodeResult_scheduler = shifterReg_7_0_bits_decodeResult_scheduler;
  reg          shifterReg_7_0_bits_decodeResult_sReadVD;
  assign validSink_7_bits_decodeResult_sReadVD = shifterReg_7_0_bits_decodeResult_sReadVD;
  reg          shifterReg_7_0_bits_decodeResult_vtype;
  assign validSink_7_bits_decodeResult_vtype = shifterReg_7_0_bits_decodeResult_vtype;
  reg          shifterReg_7_0_bits_decodeResult_sWrite;
  assign validSink_7_bits_decodeResult_sWrite = shifterReg_7_0_bits_decodeResult_sWrite;
  reg          shifterReg_7_0_bits_decodeResult_crossRead;
  assign validSink_7_bits_decodeResult_crossRead = shifterReg_7_0_bits_decodeResult_crossRead;
  reg          shifterReg_7_0_bits_decodeResult_crossWrite;
  assign validSink_7_bits_decodeResult_crossWrite = shifterReg_7_0_bits_decodeResult_crossWrite;
  reg          shifterReg_7_0_bits_decodeResult_maskUnit;
  assign validSink_7_bits_decodeResult_maskUnit = shifterReg_7_0_bits_decodeResult_maskUnit;
  reg          shifterReg_7_0_bits_decodeResult_special;
  assign validSink_7_bits_decodeResult_special = shifterReg_7_0_bits_decodeResult_special;
  reg          shifterReg_7_0_bits_decodeResult_saturate;
  assign validSink_7_bits_decodeResult_saturate = shifterReg_7_0_bits_decodeResult_saturate;
  reg          shifterReg_7_0_bits_decodeResult_vwmacc;
  assign validSink_7_bits_decodeResult_vwmacc = shifterReg_7_0_bits_decodeResult_vwmacc;
  reg          shifterReg_7_0_bits_decodeResult_readOnly;
  assign validSink_7_bits_decodeResult_readOnly = shifterReg_7_0_bits_decodeResult_readOnly;
  reg          shifterReg_7_0_bits_decodeResult_maskSource;
  assign validSink_7_bits_decodeResult_maskSource = shifterReg_7_0_bits_decodeResult_maskSource;
  reg          shifterReg_7_0_bits_decodeResult_maskDestination;
  assign validSink_7_bits_decodeResult_maskDestination = shifterReg_7_0_bits_decodeResult_maskDestination;
  reg          shifterReg_7_0_bits_decodeResult_maskLogic;
  assign validSink_7_bits_decodeResult_maskLogic = shifterReg_7_0_bits_decodeResult_maskLogic;
  reg  [3:0]   shifterReg_7_0_bits_decodeResult_uop;
  assign validSink_7_bits_decodeResult_uop = shifterReg_7_0_bits_decodeResult_uop;
  reg          shifterReg_7_0_bits_decodeResult_iota;
  assign validSink_7_bits_decodeResult_iota = shifterReg_7_0_bits_decodeResult_iota;
  reg          shifterReg_7_0_bits_decodeResult_mv;
  assign validSink_7_bits_decodeResult_mv = shifterReg_7_0_bits_decodeResult_mv;
  reg          shifterReg_7_0_bits_decodeResult_extend;
  assign validSink_7_bits_decodeResult_extend = shifterReg_7_0_bits_decodeResult_extend;
  reg          shifterReg_7_0_bits_decodeResult_unOrderWrite;
  assign validSink_7_bits_decodeResult_unOrderWrite = shifterReg_7_0_bits_decodeResult_unOrderWrite;
  reg          shifterReg_7_0_bits_decodeResult_compress;
  assign validSink_7_bits_decodeResult_compress = shifterReg_7_0_bits_decodeResult_compress;
  reg          shifterReg_7_0_bits_decodeResult_gather16;
  assign validSink_7_bits_decodeResult_gather16 = shifterReg_7_0_bits_decodeResult_gather16;
  reg          shifterReg_7_0_bits_decodeResult_gather;
  assign validSink_7_bits_decodeResult_gather = shifterReg_7_0_bits_decodeResult_gather;
  reg          shifterReg_7_0_bits_decodeResult_slid;
  assign validSink_7_bits_decodeResult_slid = shifterReg_7_0_bits_decodeResult_slid;
  reg          shifterReg_7_0_bits_decodeResult_targetRd;
  assign validSink_7_bits_decodeResult_targetRd = shifterReg_7_0_bits_decodeResult_targetRd;
  reg          shifterReg_7_0_bits_decodeResult_widenReduce;
  assign validSink_7_bits_decodeResult_widenReduce = shifterReg_7_0_bits_decodeResult_widenReduce;
  reg          shifterReg_7_0_bits_decodeResult_red;
  assign validSink_7_bits_decodeResult_red = shifterReg_7_0_bits_decodeResult_red;
  reg          shifterReg_7_0_bits_decodeResult_nr;
  assign validSink_7_bits_decodeResult_nr = shifterReg_7_0_bits_decodeResult_nr;
  reg          shifterReg_7_0_bits_decodeResult_itype;
  assign validSink_7_bits_decodeResult_itype = shifterReg_7_0_bits_decodeResult_itype;
  reg          shifterReg_7_0_bits_decodeResult_unsigned1;
  assign validSink_7_bits_decodeResult_unsigned1 = shifterReg_7_0_bits_decodeResult_unsigned1;
  reg          shifterReg_7_0_bits_decodeResult_unsigned0;
  assign validSink_7_bits_decodeResult_unsigned0 = shifterReg_7_0_bits_decodeResult_unsigned0;
  reg          shifterReg_7_0_bits_decodeResult_other;
  assign validSink_7_bits_decodeResult_other = shifterReg_7_0_bits_decodeResult_other;
  reg          shifterReg_7_0_bits_decodeResult_multiCycle;
  assign validSink_7_bits_decodeResult_multiCycle = shifterReg_7_0_bits_decodeResult_multiCycle;
  reg          shifterReg_7_0_bits_decodeResult_divider;
  assign validSink_7_bits_decodeResult_divider = shifterReg_7_0_bits_decodeResult_divider;
  reg          shifterReg_7_0_bits_decodeResult_multiplier;
  assign validSink_7_bits_decodeResult_multiplier = shifterReg_7_0_bits_decodeResult_multiplier;
  reg          shifterReg_7_0_bits_decodeResult_shift;
  assign validSink_7_bits_decodeResult_shift = shifterReg_7_0_bits_decodeResult_shift;
  reg          shifterReg_7_0_bits_decodeResult_adder;
  assign validSink_7_bits_decodeResult_adder = shifterReg_7_0_bits_decodeResult_adder;
  reg          shifterReg_7_0_bits_decodeResult_logic;
  assign validSink_7_bits_decodeResult_logic = shifterReg_7_0_bits_decodeResult_logic;
  reg          shifterReg_7_0_bits_loadStore;
  assign validSink_7_bits_loadStore = shifterReg_7_0_bits_loadStore;
  reg          shifterReg_7_0_bits_issueInst;
  assign validSink_7_bits_issueInst = shifterReg_7_0_bits_issueInst;
  reg          shifterReg_7_0_bits_store;
  assign validSink_7_bits_store = shifterReg_7_0_bits_store;
  reg          shifterReg_7_0_bits_special;
  assign validSink_7_bits_special = shifterReg_7_0_bits_special;
  reg          shifterReg_7_0_bits_lsWholeReg;
  assign validSink_7_bits_lsWholeReg = shifterReg_7_0_bits_lsWholeReg;
  reg  [4:0]   shifterReg_7_0_bits_vs1;
  assign validSink_7_bits_vs1 = shifterReg_7_0_bits_vs1;
  reg  [4:0]   shifterReg_7_0_bits_vs2;
  assign validSink_7_bits_vs2 = shifterReg_7_0_bits_vs2;
  reg  [4:0]   shifterReg_7_0_bits_vd;
  assign validSink_7_bits_vd = shifterReg_7_0_bits_vd;
  reg  [1:0]   shifterReg_7_0_bits_loadStoreEEW;
  assign validSink_7_bits_loadStoreEEW = shifterReg_7_0_bits_loadStoreEEW;
  reg          shifterReg_7_0_bits_mask;
  assign validSink_7_bits_mask = shifterReg_7_0_bits_mask;
  reg  [2:0]   shifterReg_7_0_bits_segment;
  assign validSink_7_bits_segment = shifterReg_7_0_bits_segment;
  reg  [31:0]  shifterReg_7_0_bits_readFromScalar;
  assign validSink_7_bits_readFromScalar = shifterReg_7_0_bits_readFromScalar;
  reg  [11:0]  shifterReg_7_0_bits_csrInterface_vl;
  assign validSink_7_bits_csrInterface_vl = shifterReg_7_0_bits_csrInterface_vl;
  reg  [11:0]  shifterReg_7_0_bits_csrInterface_vStart;
  assign validSink_7_bits_csrInterface_vStart = shifterReg_7_0_bits_csrInterface_vStart;
  reg  [2:0]   shifterReg_7_0_bits_csrInterface_vlmul;
  assign validSink_7_bits_csrInterface_vlmul = shifterReg_7_0_bits_csrInterface_vlmul;
  reg  [1:0]   shifterReg_7_0_bits_csrInterface_vSew;
  assign validSink_7_bits_csrInterface_vSew = shifterReg_7_0_bits_csrInterface_vSew;
  reg  [1:0]   shifterReg_7_0_bits_csrInterface_vxrm;
  assign validSink_7_bits_csrInterface_vxrm = shifterReg_7_0_bits_csrInterface_vxrm;
  reg          shifterReg_7_0_bits_csrInterface_vta;
  assign validSink_7_bits_csrInterface_vta = shifterReg_7_0_bits_csrInterface_vta;
  reg          shifterReg_7_0_bits_csrInterface_vma;
  assign validSink_7_bits_csrInterface_vma = shifterReg_7_0_bits_csrInterface_vma;
  wire         shifterValid_7 = shifterReg_7_0_valid | validSource_7_valid;
  wire [1:0]   allLaneReady_lo_lo = {laneRequestSourceWire_1_ready, laneRequestSourceWire_0_ready};
  wire [1:0]   allLaneReady_lo_hi = {laneRequestSourceWire_3_ready, laneRequestSourceWire_2_ready};
  wire [3:0]   allLaneReady_lo = {allLaneReady_lo_hi, allLaneReady_lo_lo};
  wire [1:0]   allLaneReady_hi_lo = {laneRequestSourceWire_5_ready, laneRequestSourceWire_4_ready};
  wire [1:0]   allLaneReady_hi_hi = {laneRequestSourceWire_7_ready, laneRequestSourceWire_6_ready};
  wire [3:0]   allLaneReady_hi = {allLaneReady_hi_hi, allLaneReady_hi_lo};
  wire         allLaneReady = &{allLaneReady_hi, allLaneReady_lo};
  wire         completeIndexInstruction = (|(8'h1 << _GEN_2 & _lsu_lastReport)) & ~slots_3_state_idle;
  wire [1:0]   _GEN_3 = {slots_1_state_idle, slots_0_state_idle};
  wire [1:0]   freeOR_lo;
  assign freeOR_lo = _GEN_3;
  wire [1:0]   free_lo;
  assign free_lo = _GEN_3;
  wire [1:0]   _GEN_4 = {slots_3_state_idle, slots_2_state_idle};
  wire [1:0]   freeOR_hi;
  assign freeOR_hi = _GEN_4;
  wire [1:0]   free_hi;
  assign free_hi = _GEN_4;
  wire         freeOR = |{freeOR_hi, freeOR_lo};
  wire         slotReady = specialInstruction ? slots_3_state_idle : freeOR;
  wire         olderCheck_notSameLSB = slots_0_record_instructionIndex[1:0] != requestReg_bits_instructionIndex[1:0];
  wire         olderCheck_notSameLSB_1 = slots_1_record_instructionIndex[1:0] != requestReg_bits_instructionIndex[1:0];
  wire         olderCheck_notSameLSB_2 = slots_2_record_instructionIndex[1:0] != requestReg_bits_instructionIndex[1:0];
  wire         olderCheck_notSameLSB_3 = slots_3_record_instructionIndex[1:0] != requestReg_bits_instructionIndex[1:0];
  wire         olderCheck =
    (slots_0_state_idle | (slots_0_record_instructionIndex[1:0] < requestReg_bits_instructionIndex[1:0] ^ slots_0_record_instructionIndex[2] ^ requestReg_bits_instructionIndex[2]) & olderCheck_notSameLSB)
    & (slots_1_state_idle | (slots_1_record_instructionIndex[1:0] < requestReg_bits_instructionIndex[1:0] ^ slots_1_record_instructionIndex[2] ^ requestReg_bits_instructionIndex[2]) & olderCheck_notSameLSB_1)
    & (slots_2_state_idle | (slots_2_record_instructionIndex[1:0] < requestReg_bits_instructionIndex[1:0] ^ slots_2_record_instructionIndex[2] ^ requestReg_bits_instructionIndex[2]) & olderCheck_notSameLSB_2)
    & (slots_3_state_idle | (slots_3_record_instructionIndex[1:0] < requestReg_bits_instructionIndex[1:0] ^ slots_3_record_instructionIndex[2] ^ requestReg_bits_instructionIndex[2]) & olderCheck_notSameLSB_3);
  assign source1Select = requestReg_bits_decodeResult_gather ? _maskUnit_gatherData_bits : requestReg_bits_decodeResult_itype ? immSignExtend : source1Extend;
  assign laneRequestSourceWire_0_bits_readFromScalar = source1Select;
  assign laneRequestSourceWire_1_bits_readFromScalar = source1Select;
  assign laneRequestSourceWire_2_bits_readFromScalar = source1Select;
  assign laneRequestSourceWire_3_bits_readFromScalar = source1Select;
  assign laneRequestSourceWire_4_bits_readFromScalar = source1Select;
  assign laneRequestSourceWire_5_bits_readFromScalar = source1Select;
  assign laneRequestSourceWire_6_bits_readFromScalar = source1Select;
  assign laneRequestSourceWire_7_bits_readFromScalar = source1Select;
  wire         extendDataEEW = requestReg_bits_issue_vtype[3] - requestReg_bits_decodeResult_topUop[1];
  assign laneRequestSourceWire_0_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  assign laneRequestSourceWire_1_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  assign laneRequestSourceWire_2_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  assign laneRequestSourceWire_3_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  assign laneRequestSourceWire_4_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  assign laneRequestSourceWire_5_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  assign laneRequestSourceWire_6_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  assign laneRequestSourceWire_7_bits_loadStoreEEW = requestRegDequeue_bits_instruction[13:12];
  wire [2:0]   vSewSelect =
    isLoadStoreType
      ? {1'h0, requestRegDequeue_bits_instruction[13:12]}
      : requestReg_bits_decodeResult_nr | requestReg_bits_decodeResult_maskLogic ? 3'h2 : requestReg_bits_decodeResult_gather16 ? 3'h1 : requestReg_bits_decodeResult_extend ? {2'h0, extendDataEEW} : requestReg_bits_issue_vtype[5:3];
  wire [31:0]  evlForLane = requestReg_bits_decodeResult_nr ? {22'h0, {1'h0, requestRegDequeue_bits_instruction[17:15]} + 4'h1, 6'h0} : requestReg_bits_issue_vl;
  wire [1:0]   vSewForLsu = lsWholeReg ? 2'h2 : requestRegDequeue_bits_instruction[13:12];
  wire [31:0]  evlForLsu = lsWholeReg ? {22'h0, {1'h0, requestRegDequeue_bits_instruction[31:29]} + 4'h1, 6'h0} : requestReg_bits_issue_vl;
  assign laneRequestSourceWire_0_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_1_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_2_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_3_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_4_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_5_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_6_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_7_bits_vs1 = requestRegDequeue_bits_instruction[19:15];
  assign laneRequestSourceWire_0_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_1_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_2_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_3_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_4_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_5_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_6_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_7_bits_vd = requestRegDequeue_bits_instruction[11:7];
  assign laneRequestSourceWire_0_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_0_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSourceWire_0_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_1_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_2_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_3_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_4_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_5_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_6_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_7_bits_csrInterface_vSew = vSewSelect[1:0];
  assign laneRequestSourceWire_0_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_1_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_2_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_3_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_4_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_5_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_6_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_7_bits_csrInterface_vl = evlForLane[11:0];
  assign laneRequestSourceWire_1_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_1_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSourceWire_2_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_2_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSourceWire_3_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_3_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSourceWire_4_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_4_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSourceWire_5_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_5_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSourceWire_6_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_6_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSourceWire_7_bits_segment = requestReg_bits_decodeResult_nr ? requestRegDequeue_bits_instruction[17:15] : requestRegDequeue_bits_instruction[31:29];
  assign laneRequestSourceWire_7_bits_issueInst = ~noOffsetReadLoadStore & ~maskUnitInstruction;
  assign laneRequestSinkWire_0_ready = ~laneRequestSinkWire_0_bits_issueInst | _laneVec_0_laneRequest_ready;
  wire         sinkVec_tokenCheck;
  wire [4:0]   sinkVec_validSource_bits_vs = x13_0_bits_vs;
  wire [2:0]   sinkVec_validSource_bits_offset = x13_0_bits_offset;
  wire [2:0]   sinkVec_validSource_bits_instructionIndex = x13_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_1;
  wire [4:0]   sinkVec_validSource_1_bits_vs = x13_1_bits_vs;
  wire [2:0]   sinkVec_validSource_1_bits_offset = x13_1_bits_offset;
  wire [2:0]   sinkVec_validSource_1_bits_instructionIndex = x13_1_bits_instructionIndex;
  wire         sinkVec_0_ready;
  wire         sinkVec_queue_deq_ready = sinkVec_sinkWire_ready;
  wire         sinkVec_queue_deq_valid;
  wire [4:0]   sinkVec_queue_deq_bits_vs;
  wire         sinkVec_0_valid = sinkVec_sinkWire_valid;
  wire [1:0]   sinkVec_queue_deq_bits_readSource;
  wire [4:0]   sinkVec_0_bits_vs = sinkVec_sinkWire_bits_vs;
  wire [2:0]   sinkVec_queue_deq_bits_offset;
  wire [1:0]   sinkVec_0_bits_readSource = sinkVec_sinkWire_bits_readSource;
  wire [2:0]   sinkVec_queue_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_0_bits_offset = sinkVec_sinkWire_bits_offset;
  wire [2:0]   sinkVec_0_bits_instructionIndex = sinkVec_sinkWire_bits_instructionIndex;
  wire         sinkVec_validSink_valid;
  wire [4:0]   sinkVec_validSink_bits_vs;
  wire [1:0]   sinkVec_validSink_bits_readSource;
  wire [2:0]   sinkVec_validSink_bits_offset;
  wire [2:0]   sinkVec_validSink_bits_instructionIndex;
  assign sinkVec_sinkWire_valid = sinkVec_queue_deq_valid;
  assign sinkVec_sinkWire_bits_vs = sinkVec_queue_deq_bits_vs;
  assign sinkVec_sinkWire_bits_readSource = sinkVec_queue_deq_bits_readSource;
  assign sinkVec_sinkWire_bits_offset = sinkVec_queue_deq_bits_offset;
  assign sinkVec_sinkWire_bits_instructionIndex = sinkVec_queue_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_queue_enq_bits_offset;
  wire [2:0]   sinkVec_queue_enq_bits_instructionIndex;
  wire [5:0]   sinkVec_queue_dataIn_lo = {sinkVec_queue_enq_bits_offset, sinkVec_queue_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_enq_bits_vs;
  wire [1:0]   sinkVec_queue_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi = {sinkVec_queue_enq_bits_vs, sinkVec_queue_enq_bits_readSource};
  wire [12:0]  sinkVec_queue_dataIn = {sinkVec_queue_dataIn_hi, sinkVec_queue_dataIn_lo};
  wire [2:0]   sinkVec_queue_dataOut_instructionIndex = _sinkVec_queue_fifo_data_out[2:0];
  wire [2:0]   sinkVec_queue_dataOut_offset = _sinkVec_queue_fifo_data_out[5:3];
  wire [1:0]   sinkVec_queue_dataOut_readSource = _sinkVec_queue_fifo_data_out[7:6];
  wire [4:0]   sinkVec_queue_dataOut_vs = _sinkVec_queue_fifo_data_out[12:8];
  wire         sinkVec_queue_enq_ready = ~_sinkVec_queue_fifo_full;
  wire         sinkVec_queue_enq_valid;
  assign sinkVec_queue_deq_valid = ~_sinkVec_queue_fifo_empty | sinkVec_queue_enq_valid;
  assign sinkVec_queue_deq_bits_vs = _sinkVec_queue_fifo_empty ? sinkVec_queue_enq_bits_vs : sinkVec_queue_dataOut_vs;
  assign sinkVec_queue_deq_bits_readSource = _sinkVec_queue_fifo_empty ? sinkVec_queue_enq_bits_readSource : sinkVec_queue_dataOut_readSource;
  assign sinkVec_queue_deq_bits_offset = _sinkVec_queue_fifo_empty ? sinkVec_queue_enq_bits_offset : sinkVec_queue_dataOut_offset;
  assign sinkVec_queue_deq_bits_instructionIndex = _sinkVec_queue_fifo_empty ? sinkVec_queue_enq_bits_instructionIndex : sinkVec_queue_dataOut_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v;
  wire         sinkVec_releasePipe_pipe_out_valid = sinkVec_releasePipe_pipe_v;
  wire         x13_0_ready;
  wire         x13_0_valid;
  wire         sinkVec_validSource_valid = x13_0_ready & x13_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter;
  wire [2:0]   sinkVec_tokenCheck_counterChange = sinkVec_validSource_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck = ~(sinkVec_tokenCheck_counter[2]);
  assign x13_0_ready = sinkVec_tokenCheck;
  assign sinkVec_queue_enq_valid = sinkVec_validSink_valid;
  assign sinkVec_queue_enq_bits_vs = sinkVec_validSink_bits_vs;
  assign sinkVec_queue_enq_bits_readSource = sinkVec_validSink_bits_readSource;
  assign sinkVec_queue_enq_bits_offset = sinkVec_validSink_bits_offset;
  assign sinkVec_queue_enq_bits_instructionIndex = sinkVec_validSink_bits_instructionIndex;
  reg          sinkVec_shifterReg_0_valid;
  assign sinkVec_validSink_valid = sinkVec_shifterReg_0_valid;
  reg  [4:0]   sinkVec_shifterReg_0_bits_vs;
  assign sinkVec_validSink_bits_vs = sinkVec_shifterReg_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_0_bits_readSource;
  assign sinkVec_validSink_bits_readSource = sinkVec_shifterReg_0_bits_readSource;
  reg  [2:0]   sinkVec_shifterReg_0_bits_offset;
  assign sinkVec_validSink_bits_offset = sinkVec_shifterReg_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_0_bits_instructionIndex;
  assign sinkVec_validSink_bits_instructionIndex = sinkVec_shifterReg_0_bits_instructionIndex;
  wire         sinkVec_shifterValid = sinkVec_shifterReg_0_valid | sinkVec_validSource_valid;
  wire         sinkVec_1_ready;
  wire         sinkVec_queue_1_deq_ready = sinkVec_sinkWire_1_ready;
  wire         sinkVec_queue_1_deq_valid;
  wire [4:0]   sinkVec_queue_1_deq_bits_vs;
  wire         sinkVec_1_valid = sinkVec_sinkWire_1_valid;
  wire [1:0]   sinkVec_queue_1_deq_bits_readSource;
  wire [4:0]   sinkVec_1_bits_vs = sinkVec_sinkWire_1_bits_vs;
  wire [2:0]   sinkVec_queue_1_deq_bits_offset;
  wire [1:0]   sinkVec_1_bits_readSource = sinkVec_sinkWire_1_bits_readSource;
  wire [2:0]   sinkVec_queue_1_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_1_bits_offset = sinkVec_sinkWire_1_bits_offset;
  wire [2:0]   sinkVec_1_bits_instructionIndex = sinkVec_sinkWire_1_bits_instructionIndex;
  wire         sinkVec_validSink_1_valid;
  wire [4:0]   sinkVec_validSink_1_bits_vs;
  wire [1:0]   sinkVec_validSink_1_bits_readSource;
  wire [2:0]   sinkVec_validSink_1_bits_offset;
  wire [2:0]   sinkVec_validSink_1_bits_instructionIndex;
  assign sinkVec_sinkWire_1_valid = sinkVec_queue_1_deq_valid;
  assign sinkVec_sinkWire_1_bits_vs = sinkVec_queue_1_deq_bits_vs;
  assign sinkVec_sinkWire_1_bits_readSource = sinkVec_queue_1_deq_bits_readSource;
  assign sinkVec_sinkWire_1_bits_offset = sinkVec_queue_1_deq_bits_offset;
  assign sinkVec_sinkWire_1_bits_instructionIndex = sinkVec_queue_1_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_queue_1_enq_bits_offset;
  wire [2:0]   sinkVec_queue_1_enq_bits_instructionIndex;
  wire [5:0]   sinkVec_queue_dataIn_lo_1 = {sinkVec_queue_1_enq_bits_offset, sinkVec_queue_1_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_1_enq_bits_vs;
  wire [1:0]   sinkVec_queue_1_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_1 = {sinkVec_queue_1_enq_bits_vs, sinkVec_queue_1_enq_bits_readSource};
  wire [12:0]  sinkVec_queue_dataIn_1 = {sinkVec_queue_dataIn_hi_1, sinkVec_queue_dataIn_lo_1};
  wire [2:0]   sinkVec_queue_dataOut_1_instructionIndex = _sinkVec_queue_fifo_1_data_out[2:0];
  wire [2:0]   sinkVec_queue_dataOut_1_offset = _sinkVec_queue_fifo_1_data_out[5:3];
  wire [1:0]   sinkVec_queue_dataOut_1_readSource = _sinkVec_queue_fifo_1_data_out[7:6];
  wire [4:0]   sinkVec_queue_dataOut_1_vs = _sinkVec_queue_fifo_1_data_out[12:8];
  wire         sinkVec_queue_1_enq_ready = ~_sinkVec_queue_fifo_1_full;
  wire         sinkVec_queue_1_enq_valid;
  assign sinkVec_queue_1_deq_valid = ~_sinkVec_queue_fifo_1_empty | sinkVec_queue_1_enq_valid;
  assign sinkVec_queue_1_deq_bits_vs = _sinkVec_queue_fifo_1_empty ? sinkVec_queue_1_enq_bits_vs : sinkVec_queue_dataOut_1_vs;
  assign sinkVec_queue_1_deq_bits_readSource = _sinkVec_queue_fifo_1_empty ? sinkVec_queue_1_enq_bits_readSource : sinkVec_queue_dataOut_1_readSource;
  assign sinkVec_queue_1_deq_bits_offset = _sinkVec_queue_fifo_1_empty ? sinkVec_queue_1_enq_bits_offset : sinkVec_queue_dataOut_1_offset;
  assign sinkVec_queue_1_deq_bits_instructionIndex = _sinkVec_queue_fifo_1_empty ? sinkVec_queue_1_enq_bits_instructionIndex : sinkVec_queue_dataOut_1_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_1;
  wire         sinkVec_releasePipe_pipe_out_1_valid = sinkVec_releasePipe_pipe_v_1;
  wire         x13_1_ready;
  wire         x13_1_valid;
  wire         sinkVec_validSource_1_valid = x13_1_ready & x13_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_1;
  wire [2:0]   sinkVec_tokenCheck_counterChange_1 = sinkVec_validSource_1_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_1 = ~(sinkVec_tokenCheck_counter_1[2]);
  assign x13_1_ready = sinkVec_tokenCheck_1;
  assign sinkVec_queue_1_enq_valid = sinkVec_validSink_1_valid;
  assign sinkVec_queue_1_enq_bits_vs = sinkVec_validSink_1_bits_vs;
  assign sinkVec_queue_1_enq_bits_readSource = sinkVec_validSink_1_bits_readSource;
  assign sinkVec_queue_1_enq_bits_offset = sinkVec_validSink_1_bits_offset;
  assign sinkVec_queue_1_enq_bits_instructionIndex = sinkVec_validSink_1_bits_instructionIndex;
  reg          sinkVec_shifterReg_1_0_valid;
  assign sinkVec_validSink_1_valid = sinkVec_shifterReg_1_0_valid;
  reg  [4:0]   sinkVec_shifterReg_1_0_bits_vs;
  assign sinkVec_validSink_1_bits_vs = sinkVec_shifterReg_1_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_1_0_bits_readSource;
  assign sinkVec_validSink_1_bits_readSource = sinkVec_shifterReg_1_0_bits_readSource;
  reg  [2:0]   sinkVec_shifterReg_1_0_bits_offset;
  assign sinkVec_validSink_1_bits_offset = sinkVec_shifterReg_1_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_1_0_bits_instructionIndex;
  assign sinkVec_validSink_1_bits_instructionIndex = sinkVec_shifterReg_1_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_1 = sinkVec_shifterReg_1_0_valid | sinkVec_validSource_1_valid;
  assign sinkVec_sinkWire_ready = sinkVec_0_ready;
  assign sinkVec_sinkWire_1_ready = sinkVec_1_ready;
  reg          maskUnitFirst;
  wire         tryToRead = sinkVec_0_valid | sinkVec_1_valid;
  wire         sinkWire_valid = maskUnitFirst ? sinkVec_0_valid : sinkVec_1_valid;
  wire [4:0]   sinkWire_bits_vs = maskUnitFirst ? sinkVec_0_bits_vs : sinkVec_1_bits_vs;
  wire [1:0]   sinkWire_bits_readSource = maskUnitFirst ? sinkVec_0_bits_readSource : sinkVec_1_bits_readSource;
  wire [2:0]   sinkWire_bits_offset = maskUnitFirst ? sinkVec_0_bits_offset : sinkVec_1_bits_offset;
  wire [2:0]   sinkWire_bits_instructionIndex = maskUnitFirst ? sinkVec_0_bits_instructionIndex : sinkVec_1_bits_instructionIndex;
  wire         sinkWire_ready;
  assign sinkVec_1_ready = sinkWire_ready & ~maskUnitFirst;
  assign sinkVec_0_ready = sinkWire_ready & maskUnitFirst;
  reg          accessDataValid_pipe_v;
  reg          accessDataValid_pipe_pipe_v;
  wire         accessDataValid_pipe_pipe_out_valid = accessDataValid_pipe_pipe_v;
  wire         accessDataSource_valid = accessDataValid_pipe_pipe_out_valid;
  reg          shifterReg_8_0_valid;
  reg  [31:0]  shifterReg_8_0_bits;
  wire         shifterValid_8 = shifterReg_8_0_valid | accessDataSource_valid;
  reg          accessDataValid_pipe_v_1;
  reg          accessDataValid_pipe_pipe_v_1;
  wire         accessDataValid_pipe_pipe_out_1_valid = accessDataValid_pipe_pipe_v_1;
  wire         accessDataSource_1_valid = accessDataValid_pipe_pipe_out_1_valid;
  reg          shifterReg_9_0_valid;
  reg  [31:0]  shifterReg_9_0_bits;
  wire         shifterValid_9 = shifterReg_9_0_valid | accessDataSource_1_valid;
  wire         sinkVec_tokenCheck_2;
  wire [4:0]   sinkVec_validSource_2_bits_vd = x22_0_bits_vd;
  wire [2:0]   sinkVec_validSource_2_bits_offset = x22_0_bits_offset;
  wire [3:0]   sinkVec_validSource_2_bits_mask = x22_0_bits_mask;
  wire [31:0]  sinkVec_validSource_2_bits_data = x22_0_bits_data;
  wire [2:0]   sinkVec_validSource_2_bits_instructionIndex = x22_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_3;
  wire [4:0]   sinkVec_validSource_3_bits_vd = x22_1_bits_vd;
  wire [2:0]   sinkVec_validSource_3_bits_offset = x22_1_bits_offset;
  wire [3:0]   sinkVec_validSource_3_bits_mask = x22_1_bits_mask;
  wire [31:0]  sinkVec_validSource_3_bits_data = x22_1_bits_data;
  wire         sinkVec_validSource_3_bits_last = x22_1_bits_last;
  wire [2:0]   sinkVec_validSource_3_bits_instructionIndex = x22_1_bits_instructionIndex;
  wire         sinkVec_1_0_ready;
  wire         sinkVec_queue_2_deq_ready = sinkVec_sinkWire_2_ready;
  wire         sinkVec_queue_2_deq_valid;
  wire [4:0]   sinkVec_queue_2_deq_bits_vd;
  wire         sinkVec_1_0_valid = sinkVec_sinkWire_2_valid;
  wire [2:0]   sinkVec_queue_2_deq_bits_offset;
  wire [4:0]   sinkVec_1_0_bits_vd = sinkVec_sinkWire_2_bits_vd;
  wire [3:0]   sinkVec_queue_2_deq_bits_mask;
  wire [2:0]   sinkVec_1_0_bits_offset = sinkVec_sinkWire_2_bits_offset;
  wire [31:0]  sinkVec_queue_2_deq_bits_data;
  wire [3:0]   sinkVec_1_0_bits_mask = sinkVec_sinkWire_2_bits_mask;
  wire         sinkVec_queue_2_deq_bits_last;
  wire [31:0]  sinkVec_1_0_bits_data = sinkVec_sinkWire_2_bits_data;
  wire [2:0]   sinkVec_queue_2_deq_bits_instructionIndex;
  wire         sinkVec_1_0_bits_last = sinkVec_sinkWire_2_bits_last;
  wire [2:0]   sinkVec_1_0_bits_instructionIndex = sinkVec_sinkWire_2_bits_instructionIndex;
  wire         sinkVec_validSink_2_valid;
  wire [4:0]   sinkVec_validSink_2_bits_vd;
  wire [2:0]   sinkVec_validSink_2_bits_offset;
  wire [3:0]   sinkVec_validSink_2_bits_mask;
  wire [31:0]  sinkVec_validSink_2_bits_data;
  wire [2:0]   sinkVec_validSink_2_bits_instructionIndex;
  assign sinkVec_sinkWire_2_valid = sinkVec_queue_2_deq_valid;
  assign sinkVec_sinkWire_2_bits_vd = sinkVec_queue_2_deq_bits_vd;
  assign sinkVec_sinkWire_2_bits_offset = sinkVec_queue_2_deq_bits_offset;
  assign sinkVec_sinkWire_2_bits_mask = sinkVec_queue_2_deq_bits_mask;
  assign sinkVec_sinkWire_2_bits_data = sinkVec_queue_2_deq_bits_data;
  assign sinkVec_sinkWire_2_bits_last = sinkVec_queue_2_deq_bits_last;
  assign sinkVec_sinkWire_2_bits_instructionIndex = sinkVec_queue_2_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_2_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi = {sinkVec_queue_2_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_2_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_2 = {sinkVec_queue_dataIn_lo_hi, sinkVec_queue_2_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_2_enq_bits_vd;
  wire [2:0]   sinkVec_queue_2_enq_bits_offset;
  wire [7:0]   sinkVec_queue_dataIn_hi_hi = {sinkVec_queue_2_enq_bits_vd, sinkVec_queue_2_enq_bits_offset};
  wire [3:0]   sinkVec_queue_2_enq_bits_mask;
  wire [11:0]  sinkVec_queue_dataIn_hi_2 = {sinkVec_queue_dataIn_hi_hi, sinkVec_queue_2_enq_bits_mask};
  wire [47:0]  sinkVec_queue_dataIn_2 = {sinkVec_queue_dataIn_hi_2, sinkVec_queue_dataIn_lo_2};
  wire [2:0]   sinkVec_queue_dataOut_2_instructionIndex = _sinkVec_queue_fifo_2_data_out[2:0];
  wire         sinkVec_queue_dataOut_2_last = _sinkVec_queue_fifo_2_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_2_data = _sinkVec_queue_fifo_2_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_2_mask = _sinkVec_queue_fifo_2_data_out[39:36];
  wire [2:0]   sinkVec_queue_dataOut_2_offset = _sinkVec_queue_fifo_2_data_out[42:40];
  wire [4:0]   sinkVec_queue_dataOut_2_vd = _sinkVec_queue_fifo_2_data_out[47:43];
  wire         sinkVec_queue_2_enq_ready = ~_sinkVec_queue_fifo_2_full;
  wire         sinkVec_queue_2_enq_valid;
  assign sinkVec_queue_2_deq_valid = ~_sinkVec_queue_fifo_2_empty | sinkVec_queue_2_enq_valid;
  assign sinkVec_queue_2_deq_bits_vd = _sinkVec_queue_fifo_2_empty ? sinkVec_queue_2_enq_bits_vd : sinkVec_queue_dataOut_2_vd;
  assign sinkVec_queue_2_deq_bits_offset = _sinkVec_queue_fifo_2_empty ? sinkVec_queue_2_enq_bits_offset : sinkVec_queue_dataOut_2_offset;
  assign sinkVec_queue_2_deq_bits_mask = _sinkVec_queue_fifo_2_empty ? sinkVec_queue_2_enq_bits_mask : sinkVec_queue_dataOut_2_mask;
  assign sinkVec_queue_2_deq_bits_data = _sinkVec_queue_fifo_2_empty ? sinkVec_queue_2_enq_bits_data : sinkVec_queue_dataOut_2_data;
  assign sinkVec_queue_2_deq_bits_last = ~_sinkVec_queue_fifo_2_empty & sinkVec_queue_dataOut_2_last;
  assign sinkVec_queue_2_deq_bits_instructionIndex = _sinkVec_queue_fifo_2_empty ? sinkVec_queue_2_enq_bits_instructionIndex : sinkVec_queue_dataOut_2_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_2;
  wire         sinkVec_releasePipe_pipe_out_2_valid = sinkVec_releasePipe_pipe_v_2;
  wire         x22_0_ready;
  wire         x22_0_valid;
  wire         sinkVec_validSource_2_valid = x22_0_ready & x22_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_2;
  wire [2:0]   sinkVec_tokenCheck_counterChange_2 = sinkVec_validSource_2_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_2 = ~(sinkVec_tokenCheck_counter_2[2]);
  assign x22_0_ready = sinkVec_tokenCheck_2;
  assign sinkVec_queue_2_enq_valid = sinkVec_validSink_2_valid;
  assign sinkVec_queue_2_enq_bits_vd = sinkVec_validSink_2_bits_vd;
  assign sinkVec_queue_2_enq_bits_offset = sinkVec_validSink_2_bits_offset;
  assign sinkVec_queue_2_enq_bits_mask = sinkVec_validSink_2_bits_mask;
  assign sinkVec_queue_2_enq_bits_data = sinkVec_validSink_2_bits_data;
  assign sinkVec_queue_2_enq_bits_instructionIndex = sinkVec_validSink_2_bits_instructionIndex;
  reg          sinkVec_shifterReg_2_0_valid;
  assign sinkVec_validSink_2_valid = sinkVec_shifterReg_2_0_valid;
  reg  [4:0]   sinkVec_shifterReg_2_0_bits_vd;
  assign sinkVec_validSink_2_bits_vd = sinkVec_shifterReg_2_0_bits_vd;
  reg  [2:0]   sinkVec_shifterReg_2_0_bits_offset;
  assign sinkVec_validSink_2_bits_offset = sinkVec_shifterReg_2_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_2_0_bits_mask;
  assign sinkVec_validSink_2_bits_mask = sinkVec_shifterReg_2_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_2_0_bits_data;
  assign sinkVec_validSink_2_bits_data = sinkVec_shifterReg_2_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_2_0_bits_instructionIndex;
  assign sinkVec_validSink_2_bits_instructionIndex = sinkVec_shifterReg_2_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_2 = sinkVec_shifterReg_2_0_valid | sinkVec_validSource_2_valid;
  wire         sinkVec_1_1_ready;
  wire         sinkVec_queue_3_deq_ready = sinkVec_sinkWire_3_ready;
  wire         sinkVec_queue_3_deq_valid;
  wire [4:0]   sinkVec_queue_3_deq_bits_vd;
  wire         sinkVec_1_1_valid = sinkVec_sinkWire_3_valid;
  wire [2:0]   sinkVec_queue_3_deq_bits_offset;
  wire [4:0]   sinkVec_1_1_bits_vd = sinkVec_sinkWire_3_bits_vd;
  wire [3:0]   sinkVec_queue_3_deq_bits_mask;
  wire [2:0]   sinkVec_1_1_bits_offset = sinkVec_sinkWire_3_bits_offset;
  wire [31:0]  sinkVec_queue_3_deq_bits_data;
  wire [3:0]   sinkVec_1_1_bits_mask = sinkVec_sinkWire_3_bits_mask;
  wire         sinkVec_queue_3_deq_bits_last;
  wire [31:0]  sinkVec_1_1_bits_data = sinkVec_sinkWire_3_bits_data;
  wire [2:0]   sinkVec_queue_3_deq_bits_instructionIndex;
  wire         sinkVec_1_1_bits_last = sinkVec_sinkWire_3_bits_last;
  wire [2:0]   sinkVec_1_1_bits_instructionIndex = sinkVec_sinkWire_3_bits_instructionIndex;
  wire         sinkVec_validSink_3_valid;
  wire [4:0]   sinkVec_validSink_3_bits_vd;
  wire [2:0]   sinkVec_validSink_3_bits_offset;
  wire [3:0]   sinkVec_validSink_3_bits_mask;
  wire [31:0]  sinkVec_validSink_3_bits_data;
  wire         sinkVec_validSink_3_bits_last;
  wire [2:0]   sinkVec_validSink_3_bits_instructionIndex;
  assign sinkVec_sinkWire_3_valid = sinkVec_queue_3_deq_valid;
  assign sinkVec_sinkWire_3_bits_vd = sinkVec_queue_3_deq_bits_vd;
  assign sinkVec_sinkWire_3_bits_offset = sinkVec_queue_3_deq_bits_offset;
  assign sinkVec_sinkWire_3_bits_mask = sinkVec_queue_3_deq_bits_mask;
  assign sinkVec_sinkWire_3_bits_data = sinkVec_queue_3_deq_bits_data;
  assign sinkVec_sinkWire_3_bits_last = sinkVec_queue_3_deq_bits_last;
  assign sinkVec_sinkWire_3_bits_instructionIndex = sinkVec_queue_3_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_3_enq_bits_data;
  wire         sinkVec_queue_3_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_1 = {sinkVec_queue_3_enq_bits_data, sinkVec_queue_3_enq_bits_last};
  wire [2:0]   sinkVec_queue_3_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_3 = {sinkVec_queue_dataIn_lo_hi_1, sinkVec_queue_3_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_3_enq_bits_vd;
  wire [2:0]   sinkVec_queue_3_enq_bits_offset;
  wire [7:0]   sinkVec_queue_dataIn_hi_hi_1 = {sinkVec_queue_3_enq_bits_vd, sinkVec_queue_3_enq_bits_offset};
  wire [3:0]   sinkVec_queue_3_enq_bits_mask;
  wire [11:0]  sinkVec_queue_dataIn_hi_3 = {sinkVec_queue_dataIn_hi_hi_1, sinkVec_queue_3_enq_bits_mask};
  wire [47:0]  sinkVec_queue_dataIn_3 = {sinkVec_queue_dataIn_hi_3, sinkVec_queue_dataIn_lo_3};
  wire [2:0]   sinkVec_queue_dataOut_3_instructionIndex = _sinkVec_queue_fifo_3_data_out[2:0];
  wire         sinkVec_queue_dataOut_3_last = _sinkVec_queue_fifo_3_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_3_data = _sinkVec_queue_fifo_3_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_3_mask = _sinkVec_queue_fifo_3_data_out[39:36];
  wire [2:0]   sinkVec_queue_dataOut_3_offset = _sinkVec_queue_fifo_3_data_out[42:40];
  wire [4:0]   sinkVec_queue_dataOut_3_vd = _sinkVec_queue_fifo_3_data_out[47:43];
  wire         sinkVec_queue_3_enq_ready = ~_sinkVec_queue_fifo_3_full;
  wire         sinkVec_queue_3_enq_valid;
  assign sinkVec_queue_3_deq_valid = ~_sinkVec_queue_fifo_3_empty | sinkVec_queue_3_enq_valid;
  assign sinkVec_queue_3_deq_bits_vd = _sinkVec_queue_fifo_3_empty ? sinkVec_queue_3_enq_bits_vd : sinkVec_queue_dataOut_3_vd;
  assign sinkVec_queue_3_deq_bits_offset = _sinkVec_queue_fifo_3_empty ? sinkVec_queue_3_enq_bits_offset : sinkVec_queue_dataOut_3_offset;
  assign sinkVec_queue_3_deq_bits_mask = _sinkVec_queue_fifo_3_empty ? sinkVec_queue_3_enq_bits_mask : sinkVec_queue_dataOut_3_mask;
  assign sinkVec_queue_3_deq_bits_data = _sinkVec_queue_fifo_3_empty ? sinkVec_queue_3_enq_bits_data : sinkVec_queue_dataOut_3_data;
  assign sinkVec_queue_3_deq_bits_last = _sinkVec_queue_fifo_3_empty ? sinkVec_queue_3_enq_bits_last : sinkVec_queue_dataOut_3_last;
  assign sinkVec_queue_3_deq_bits_instructionIndex = _sinkVec_queue_fifo_3_empty ? sinkVec_queue_3_enq_bits_instructionIndex : sinkVec_queue_dataOut_3_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_3;
  wire         sinkVec_releasePipe_pipe_out_3_valid = sinkVec_releasePipe_pipe_v_3;
  wire         x22_1_ready;
  wire         x22_1_valid;
  wire         sinkVec_validSource_3_valid = x22_1_ready & x22_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_3;
  wire [2:0]   sinkVec_tokenCheck_counterChange_3 = sinkVec_validSource_3_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_3 = ~(sinkVec_tokenCheck_counter_3[2]);
  assign x22_1_ready = sinkVec_tokenCheck_3;
  assign sinkVec_queue_3_enq_valid = sinkVec_validSink_3_valid;
  assign sinkVec_queue_3_enq_bits_vd = sinkVec_validSink_3_bits_vd;
  assign sinkVec_queue_3_enq_bits_offset = sinkVec_validSink_3_bits_offset;
  assign sinkVec_queue_3_enq_bits_mask = sinkVec_validSink_3_bits_mask;
  assign sinkVec_queue_3_enq_bits_data = sinkVec_validSink_3_bits_data;
  assign sinkVec_queue_3_enq_bits_last = sinkVec_validSink_3_bits_last;
  assign sinkVec_queue_3_enq_bits_instructionIndex = sinkVec_validSink_3_bits_instructionIndex;
  reg          sinkVec_shifterReg_3_0_valid;
  assign sinkVec_validSink_3_valid = sinkVec_shifterReg_3_0_valid;
  reg  [4:0]   sinkVec_shifterReg_3_0_bits_vd;
  assign sinkVec_validSink_3_bits_vd = sinkVec_shifterReg_3_0_bits_vd;
  reg  [2:0]   sinkVec_shifterReg_3_0_bits_offset;
  assign sinkVec_validSink_3_bits_offset = sinkVec_shifterReg_3_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_3_0_bits_mask;
  assign sinkVec_validSink_3_bits_mask = sinkVec_shifterReg_3_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_3_0_bits_data;
  assign sinkVec_validSink_3_bits_data = sinkVec_shifterReg_3_0_bits_data;
  reg          sinkVec_shifterReg_3_0_bits_last;
  assign sinkVec_validSink_3_bits_last = sinkVec_shifterReg_3_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_3_0_bits_instructionIndex;
  assign sinkVec_validSink_3_bits_instructionIndex = sinkVec_shifterReg_3_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_3 = sinkVec_shifterReg_3_0_valid | sinkVec_validSource_3_valid;
  assign sinkVec_sinkWire_2_ready = sinkVec_1_0_ready;
  assign sinkVec_sinkWire_3_ready = sinkVec_1_1_ready;
  reg          maskUnitFirst_1;
  wire         tryToRead_1 = sinkVec_1_0_valid | sinkVec_1_1_valid;
  wire         sinkWire_1_valid = maskUnitFirst_1 ? sinkVec_1_0_valid : sinkVec_1_1_valid;
  wire [4:0]   sinkWire_1_bits_vd = maskUnitFirst_1 ? sinkVec_1_0_bits_vd : sinkVec_1_1_bits_vd;
  wire [2:0]   sinkWire_1_bits_offset = maskUnitFirst_1 ? sinkVec_1_0_bits_offset : sinkVec_1_1_bits_offset;
  wire [3:0]   sinkWire_1_bits_mask = maskUnitFirst_1 ? sinkVec_1_0_bits_mask : sinkVec_1_1_bits_mask;
  wire [31:0]  sinkWire_1_bits_data = maskUnitFirst_1 ? sinkVec_1_0_bits_data : sinkVec_1_1_bits_data;
  wire         sinkWire_1_bits_last = maskUnitFirst_1 ? sinkVec_1_0_bits_last : sinkVec_1_1_bits_last;
  wire [2:0]   sinkWire_1_bits_instructionIndex = maskUnitFirst_1 ? sinkVec_1_0_bits_instructionIndex : sinkVec_1_1_bits_instructionIndex;
  wire         sinkWire_1_ready;
  assign sinkVec_1_1_ready = sinkWire_1_ready & ~maskUnitFirst_1;
  assign sinkVec_1_0_ready = sinkWire_1_ready & maskUnitFirst_1;
  reg          view__writeRelease_0_pipe_v;
  wire         view__writeRelease_0_pipe_out_valid = view__writeRelease_0_pipe_v;
  reg          pipe_v;
  wire         pipe_out_valid = pipe_v;
  wire         _probeWire_writeQueueEnqVec_0_valid_T = x22_0_ready & _maskUnit_exeResp_0_valid;
  reg          instructionFinishedPipe_pipe_v;
  wire         instructionFinishedPipe_pipe_out_valid = instructionFinishedPipe_pipe_v;
  reg  [7:0]   instructionFinishedPipe_pipe_b;
  wire [7:0]   instructionFinishedPipe_pipe_out_bits = instructionFinishedPipe_pipe_b;
  wire         instructionFinished_0_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_bits);
  wire         instructionFinished_0_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_bits);
  wire         instructionFinished_0_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_bits);
  wire         instructionFinished_0_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_bits);
  assign vxsatReportVec_0 = _laneVec_0_vxsatReport[3:0];
  reg          pipe_v_1;
  reg  [31:0]  pipe_b_1;
  reg          pipe_pipe_v;
  wire         pipe_pipe_out_valid = pipe_pipe_v;
  reg  [31:0]  pipe_pipe_b;
  wire [31:0]  pipe_pipe_out_bits = pipe_pipe_b;
  reg          view__laneMaskSelect_0_pipe_v;
  reg  [5:0]   view__laneMaskSelect_0_pipe_b;
  reg          view__laneMaskSelect_0_pipe_pipe_v;
  wire         view__laneMaskSelect_0_pipe_pipe_out_valid = view__laneMaskSelect_0_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_0_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_0_pipe_pipe_out_bits = view__laneMaskSelect_0_pipe_pipe_b;
  reg          view__laneMaskSewSelect_0_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_0_pipe_b;
  reg          view__laneMaskSewSelect_0_pipe_pipe_v;
  wire         view__laneMaskSewSelect_0_pipe_pipe_out_valid = view__laneMaskSewSelect_0_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_0_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_0_pipe_pipe_out_bits = view__laneMaskSewSelect_0_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v;
  wire         lsuLastPipe_pipe_out_valid = lsuLastPipe_pipe_v;
  reg  [7:0]   lsuLastPipe_pipe_b;
  wire [7:0]   lsuLastPipe_pipe_out_bits = lsuLastPipe_pipe_b;
  reg          maskLastPipe_pipe_v;
  wire         maskLastPipe_pipe_out_valid = maskLastPipe_pipe_v;
  reg  [7:0]   maskLastPipe_pipe_b;
  wire [7:0]   maskLastPipe_pipe_out_bits = maskLastPipe_pipe_b;
  wire [6:0]   writeCounter = requestReg_bits_writeByte[11:5] + {6'h0, |(requestReg_bits_writeByte[4:0])};
  reg          pipe_v_2;
  wire         pipe_out_1_valid = pipe_v_2;
  reg  [6:0]   pipe_b_2;
  wire [6:0]   pipe_out_1_bits = pipe_b_2;
  assign laneRequestSinkWire_1_ready = ~laneRequestSinkWire_1_bits_issueInst | _laneVec_1_laneRequest_ready;
  wire         sinkVec_tokenCheck_4;
  wire [4:0]   sinkVec_validSource_4_bits_vs = x13_1_0_bits_vs;
  wire [2:0]   sinkVec_validSource_4_bits_offset = x13_1_0_bits_offset;
  wire [2:0]   sinkVec_validSource_4_bits_instructionIndex = x13_1_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_5;
  wire [4:0]   sinkVec_validSource_5_bits_vs = x13_1_1_bits_vs;
  wire [2:0]   sinkVec_validSource_5_bits_offset = x13_1_1_bits_offset;
  wire [2:0]   sinkVec_validSource_5_bits_instructionIndex = x13_1_1_bits_instructionIndex;
  wire         sinkVec_2_0_ready;
  wire         sinkVec_queue_4_deq_ready = sinkVec_sinkWire_4_ready;
  wire         sinkVec_queue_4_deq_valid;
  wire [4:0]   sinkVec_queue_4_deq_bits_vs;
  wire         sinkVec_2_0_valid = sinkVec_sinkWire_4_valid;
  wire [1:0]   sinkVec_queue_4_deq_bits_readSource;
  wire [4:0]   sinkVec_2_0_bits_vs = sinkVec_sinkWire_4_bits_vs;
  wire [2:0]   sinkVec_queue_4_deq_bits_offset;
  wire [1:0]   sinkVec_2_0_bits_readSource = sinkVec_sinkWire_4_bits_readSource;
  wire [2:0]   sinkVec_queue_4_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_2_0_bits_offset = sinkVec_sinkWire_4_bits_offset;
  wire [2:0]   sinkVec_2_0_bits_instructionIndex = sinkVec_sinkWire_4_bits_instructionIndex;
  wire         sinkVec_validSink_4_valid;
  wire [4:0]   sinkVec_validSink_4_bits_vs;
  wire [1:0]   sinkVec_validSink_4_bits_readSource;
  wire [2:0]   sinkVec_validSink_4_bits_offset;
  wire [2:0]   sinkVec_validSink_4_bits_instructionIndex;
  assign sinkVec_sinkWire_4_valid = sinkVec_queue_4_deq_valid;
  assign sinkVec_sinkWire_4_bits_vs = sinkVec_queue_4_deq_bits_vs;
  assign sinkVec_sinkWire_4_bits_readSource = sinkVec_queue_4_deq_bits_readSource;
  assign sinkVec_sinkWire_4_bits_offset = sinkVec_queue_4_deq_bits_offset;
  assign sinkVec_sinkWire_4_bits_instructionIndex = sinkVec_queue_4_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_queue_4_enq_bits_offset;
  wire [2:0]   sinkVec_queue_4_enq_bits_instructionIndex;
  wire [5:0]   sinkVec_queue_dataIn_lo_4 = {sinkVec_queue_4_enq_bits_offset, sinkVec_queue_4_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_4_enq_bits_vs;
  wire [1:0]   sinkVec_queue_4_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_4 = {sinkVec_queue_4_enq_bits_vs, sinkVec_queue_4_enq_bits_readSource};
  wire [12:0]  sinkVec_queue_dataIn_4 = {sinkVec_queue_dataIn_hi_4, sinkVec_queue_dataIn_lo_4};
  wire [2:0]   sinkVec_queue_dataOut_4_instructionIndex = _sinkVec_queue_fifo_4_data_out[2:0];
  wire [2:0]   sinkVec_queue_dataOut_4_offset = _sinkVec_queue_fifo_4_data_out[5:3];
  wire [1:0]   sinkVec_queue_dataOut_4_readSource = _sinkVec_queue_fifo_4_data_out[7:6];
  wire [4:0]   sinkVec_queue_dataOut_4_vs = _sinkVec_queue_fifo_4_data_out[12:8];
  wire         sinkVec_queue_4_enq_ready = ~_sinkVec_queue_fifo_4_full;
  wire         sinkVec_queue_4_enq_valid;
  assign sinkVec_queue_4_deq_valid = ~_sinkVec_queue_fifo_4_empty | sinkVec_queue_4_enq_valid;
  assign sinkVec_queue_4_deq_bits_vs = _sinkVec_queue_fifo_4_empty ? sinkVec_queue_4_enq_bits_vs : sinkVec_queue_dataOut_4_vs;
  assign sinkVec_queue_4_deq_bits_readSource = _sinkVec_queue_fifo_4_empty ? sinkVec_queue_4_enq_bits_readSource : sinkVec_queue_dataOut_4_readSource;
  assign sinkVec_queue_4_deq_bits_offset = _sinkVec_queue_fifo_4_empty ? sinkVec_queue_4_enq_bits_offset : sinkVec_queue_dataOut_4_offset;
  assign sinkVec_queue_4_deq_bits_instructionIndex = _sinkVec_queue_fifo_4_empty ? sinkVec_queue_4_enq_bits_instructionIndex : sinkVec_queue_dataOut_4_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_4;
  wire         sinkVec_releasePipe_pipe_out_4_valid = sinkVec_releasePipe_pipe_v_4;
  wire         x13_1_0_ready;
  wire         x13_1_0_valid;
  wire         sinkVec_validSource_4_valid = x13_1_0_ready & x13_1_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_4;
  wire [2:0]   sinkVec_tokenCheck_counterChange_4 = sinkVec_validSource_4_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_4 = ~(sinkVec_tokenCheck_counter_4[2]);
  assign x13_1_0_ready = sinkVec_tokenCheck_4;
  assign sinkVec_queue_4_enq_valid = sinkVec_validSink_4_valid;
  assign sinkVec_queue_4_enq_bits_vs = sinkVec_validSink_4_bits_vs;
  assign sinkVec_queue_4_enq_bits_readSource = sinkVec_validSink_4_bits_readSource;
  assign sinkVec_queue_4_enq_bits_offset = sinkVec_validSink_4_bits_offset;
  assign sinkVec_queue_4_enq_bits_instructionIndex = sinkVec_validSink_4_bits_instructionIndex;
  reg          sinkVec_shifterReg_4_0_valid;
  assign sinkVec_validSink_4_valid = sinkVec_shifterReg_4_0_valid;
  reg  [4:0]   sinkVec_shifterReg_4_0_bits_vs;
  assign sinkVec_validSink_4_bits_vs = sinkVec_shifterReg_4_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_4_0_bits_readSource;
  assign sinkVec_validSink_4_bits_readSource = sinkVec_shifterReg_4_0_bits_readSource;
  reg  [2:0]   sinkVec_shifterReg_4_0_bits_offset;
  assign sinkVec_validSink_4_bits_offset = sinkVec_shifterReg_4_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_4_0_bits_instructionIndex;
  assign sinkVec_validSink_4_bits_instructionIndex = sinkVec_shifterReg_4_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_4 = sinkVec_shifterReg_4_0_valid | sinkVec_validSource_4_valid;
  wire         sinkVec_2_1_ready;
  wire         sinkVec_queue_5_deq_ready = sinkVec_sinkWire_5_ready;
  wire         sinkVec_queue_5_deq_valid;
  wire [4:0]   sinkVec_queue_5_deq_bits_vs;
  wire         sinkVec_2_1_valid = sinkVec_sinkWire_5_valid;
  wire [1:0]   sinkVec_queue_5_deq_bits_readSource;
  wire [4:0]   sinkVec_2_1_bits_vs = sinkVec_sinkWire_5_bits_vs;
  wire [2:0]   sinkVec_queue_5_deq_bits_offset;
  wire [1:0]   sinkVec_2_1_bits_readSource = sinkVec_sinkWire_5_bits_readSource;
  wire [2:0]   sinkVec_queue_5_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_2_1_bits_offset = sinkVec_sinkWire_5_bits_offset;
  wire [2:0]   sinkVec_2_1_bits_instructionIndex = sinkVec_sinkWire_5_bits_instructionIndex;
  wire         sinkVec_validSink_5_valid;
  wire [4:0]   sinkVec_validSink_5_bits_vs;
  wire [1:0]   sinkVec_validSink_5_bits_readSource;
  wire [2:0]   sinkVec_validSink_5_bits_offset;
  wire [2:0]   sinkVec_validSink_5_bits_instructionIndex;
  assign sinkVec_sinkWire_5_valid = sinkVec_queue_5_deq_valid;
  assign sinkVec_sinkWire_5_bits_vs = sinkVec_queue_5_deq_bits_vs;
  assign sinkVec_sinkWire_5_bits_readSource = sinkVec_queue_5_deq_bits_readSource;
  assign sinkVec_sinkWire_5_bits_offset = sinkVec_queue_5_deq_bits_offset;
  assign sinkVec_sinkWire_5_bits_instructionIndex = sinkVec_queue_5_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_queue_5_enq_bits_offset;
  wire [2:0]   sinkVec_queue_5_enq_bits_instructionIndex;
  wire [5:0]   sinkVec_queue_dataIn_lo_5 = {sinkVec_queue_5_enq_bits_offset, sinkVec_queue_5_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_5_enq_bits_vs;
  wire [1:0]   sinkVec_queue_5_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_5 = {sinkVec_queue_5_enq_bits_vs, sinkVec_queue_5_enq_bits_readSource};
  wire [12:0]  sinkVec_queue_dataIn_5 = {sinkVec_queue_dataIn_hi_5, sinkVec_queue_dataIn_lo_5};
  wire [2:0]   sinkVec_queue_dataOut_5_instructionIndex = _sinkVec_queue_fifo_5_data_out[2:0];
  wire [2:0]   sinkVec_queue_dataOut_5_offset = _sinkVec_queue_fifo_5_data_out[5:3];
  wire [1:0]   sinkVec_queue_dataOut_5_readSource = _sinkVec_queue_fifo_5_data_out[7:6];
  wire [4:0]   sinkVec_queue_dataOut_5_vs = _sinkVec_queue_fifo_5_data_out[12:8];
  wire         sinkVec_queue_5_enq_ready = ~_sinkVec_queue_fifo_5_full;
  wire         sinkVec_queue_5_enq_valid;
  assign sinkVec_queue_5_deq_valid = ~_sinkVec_queue_fifo_5_empty | sinkVec_queue_5_enq_valid;
  assign sinkVec_queue_5_deq_bits_vs = _sinkVec_queue_fifo_5_empty ? sinkVec_queue_5_enq_bits_vs : sinkVec_queue_dataOut_5_vs;
  assign sinkVec_queue_5_deq_bits_readSource = _sinkVec_queue_fifo_5_empty ? sinkVec_queue_5_enq_bits_readSource : sinkVec_queue_dataOut_5_readSource;
  assign sinkVec_queue_5_deq_bits_offset = _sinkVec_queue_fifo_5_empty ? sinkVec_queue_5_enq_bits_offset : sinkVec_queue_dataOut_5_offset;
  assign sinkVec_queue_5_deq_bits_instructionIndex = _sinkVec_queue_fifo_5_empty ? sinkVec_queue_5_enq_bits_instructionIndex : sinkVec_queue_dataOut_5_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_5;
  wire         sinkVec_releasePipe_pipe_out_5_valid = sinkVec_releasePipe_pipe_v_5;
  wire         x13_1_1_ready;
  wire         x13_1_1_valid;
  wire         sinkVec_validSource_5_valid = x13_1_1_ready & x13_1_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_5;
  wire [2:0]   sinkVec_tokenCheck_counterChange_5 = sinkVec_validSource_5_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_5 = ~(sinkVec_tokenCheck_counter_5[2]);
  assign x13_1_1_ready = sinkVec_tokenCheck_5;
  assign sinkVec_queue_5_enq_valid = sinkVec_validSink_5_valid;
  assign sinkVec_queue_5_enq_bits_vs = sinkVec_validSink_5_bits_vs;
  assign sinkVec_queue_5_enq_bits_readSource = sinkVec_validSink_5_bits_readSource;
  assign sinkVec_queue_5_enq_bits_offset = sinkVec_validSink_5_bits_offset;
  assign sinkVec_queue_5_enq_bits_instructionIndex = sinkVec_validSink_5_bits_instructionIndex;
  reg          sinkVec_shifterReg_5_0_valid;
  assign sinkVec_validSink_5_valid = sinkVec_shifterReg_5_0_valid;
  reg  [4:0]   sinkVec_shifterReg_5_0_bits_vs;
  assign sinkVec_validSink_5_bits_vs = sinkVec_shifterReg_5_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_5_0_bits_readSource;
  assign sinkVec_validSink_5_bits_readSource = sinkVec_shifterReg_5_0_bits_readSource;
  reg  [2:0]   sinkVec_shifterReg_5_0_bits_offset;
  assign sinkVec_validSink_5_bits_offset = sinkVec_shifterReg_5_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_5_0_bits_instructionIndex;
  assign sinkVec_validSink_5_bits_instructionIndex = sinkVec_shifterReg_5_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_5 = sinkVec_shifterReg_5_0_valid | sinkVec_validSource_5_valid;
  assign sinkVec_sinkWire_4_ready = sinkVec_2_0_ready;
  assign sinkVec_sinkWire_5_ready = sinkVec_2_1_ready;
  reg          maskUnitFirst_2;
  wire         tryToRead_2 = sinkVec_2_0_valid | sinkVec_2_1_valid;
  wire         sinkWire_2_valid = maskUnitFirst_2 ? sinkVec_2_0_valid : sinkVec_2_1_valid;
  wire [4:0]   sinkWire_2_bits_vs = maskUnitFirst_2 ? sinkVec_2_0_bits_vs : sinkVec_2_1_bits_vs;
  wire [1:0]   sinkWire_2_bits_readSource = maskUnitFirst_2 ? sinkVec_2_0_bits_readSource : sinkVec_2_1_bits_readSource;
  wire [2:0]   sinkWire_2_bits_offset = maskUnitFirst_2 ? sinkVec_2_0_bits_offset : sinkVec_2_1_bits_offset;
  wire [2:0]   sinkWire_2_bits_instructionIndex = maskUnitFirst_2 ? sinkVec_2_0_bits_instructionIndex : sinkVec_2_1_bits_instructionIndex;
  wire         sinkWire_2_ready;
  assign sinkVec_2_1_ready = sinkWire_2_ready & ~maskUnitFirst_2;
  assign sinkVec_2_0_ready = sinkWire_2_ready & maskUnitFirst_2;
  reg          accessDataValid_pipe_v_2;
  reg          accessDataValid_pipe_pipe_v_2;
  wire         accessDataValid_pipe_pipe_out_2_valid = accessDataValid_pipe_pipe_v_2;
  wire         accessDataSource_2_valid = accessDataValid_pipe_pipe_out_2_valid;
  reg          shifterReg_10_0_valid;
  reg  [31:0]  shifterReg_10_0_bits;
  wire         shifterValid_10 = shifterReg_10_0_valid | accessDataSource_2_valid;
  reg          accessDataValid_pipe_v_3;
  reg          accessDataValid_pipe_pipe_v_3;
  wire         accessDataValid_pipe_pipe_out_3_valid = accessDataValid_pipe_pipe_v_3;
  wire         accessDataSource_3_valid = accessDataValid_pipe_pipe_out_3_valid;
  reg          shifterReg_11_0_valid;
  reg  [31:0]  shifterReg_11_0_bits;
  wire         shifterValid_11 = shifterReg_11_0_valid | accessDataSource_3_valid;
  wire         sinkVec_tokenCheck_6;
  wire [4:0]   sinkVec_validSource_6_bits_vd = x22_1_0_bits_vd;
  wire [2:0]   sinkVec_validSource_6_bits_offset = x22_1_0_bits_offset;
  wire [3:0]   sinkVec_validSource_6_bits_mask = x22_1_0_bits_mask;
  wire [31:0]  sinkVec_validSource_6_bits_data = x22_1_0_bits_data;
  wire [2:0]   sinkVec_validSource_6_bits_instructionIndex = x22_1_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_7;
  wire [4:0]   sinkVec_validSource_7_bits_vd = x22_1_1_bits_vd;
  wire [2:0]   sinkVec_validSource_7_bits_offset = x22_1_1_bits_offset;
  wire [3:0]   sinkVec_validSource_7_bits_mask = x22_1_1_bits_mask;
  wire [31:0]  sinkVec_validSource_7_bits_data = x22_1_1_bits_data;
  wire         sinkVec_validSource_7_bits_last = x22_1_1_bits_last;
  wire [2:0]   sinkVec_validSource_7_bits_instructionIndex = x22_1_1_bits_instructionIndex;
  wire         sinkVec_3_0_ready;
  wire         sinkVec_queue_6_deq_ready = sinkVec_sinkWire_6_ready;
  wire         sinkVec_queue_6_deq_valid;
  wire [4:0]   sinkVec_queue_6_deq_bits_vd;
  wire         sinkVec_3_0_valid = sinkVec_sinkWire_6_valid;
  wire [2:0]   sinkVec_queue_6_deq_bits_offset;
  wire [4:0]   sinkVec_3_0_bits_vd = sinkVec_sinkWire_6_bits_vd;
  wire [3:0]   sinkVec_queue_6_deq_bits_mask;
  wire [2:0]   sinkVec_3_0_bits_offset = sinkVec_sinkWire_6_bits_offset;
  wire [31:0]  sinkVec_queue_6_deq_bits_data;
  wire [3:0]   sinkVec_3_0_bits_mask = sinkVec_sinkWire_6_bits_mask;
  wire         sinkVec_queue_6_deq_bits_last;
  wire [31:0]  sinkVec_3_0_bits_data = sinkVec_sinkWire_6_bits_data;
  wire [2:0]   sinkVec_queue_6_deq_bits_instructionIndex;
  wire         sinkVec_3_0_bits_last = sinkVec_sinkWire_6_bits_last;
  wire [2:0]   sinkVec_3_0_bits_instructionIndex = sinkVec_sinkWire_6_bits_instructionIndex;
  wire         sinkVec_validSink_6_valid;
  wire [4:0]   sinkVec_validSink_6_bits_vd;
  wire [2:0]   sinkVec_validSink_6_bits_offset;
  wire [3:0]   sinkVec_validSink_6_bits_mask;
  wire [31:0]  sinkVec_validSink_6_bits_data;
  wire [2:0]   sinkVec_validSink_6_bits_instructionIndex;
  assign sinkVec_sinkWire_6_valid = sinkVec_queue_6_deq_valid;
  assign sinkVec_sinkWire_6_bits_vd = sinkVec_queue_6_deq_bits_vd;
  assign sinkVec_sinkWire_6_bits_offset = sinkVec_queue_6_deq_bits_offset;
  assign sinkVec_sinkWire_6_bits_mask = sinkVec_queue_6_deq_bits_mask;
  assign sinkVec_sinkWire_6_bits_data = sinkVec_queue_6_deq_bits_data;
  assign sinkVec_sinkWire_6_bits_last = sinkVec_queue_6_deq_bits_last;
  assign sinkVec_sinkWire_6_bits_instructionIndex = sinkVec_queue_6_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_6_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_2 = {sinkVec_queue_6_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_6_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_6 = {sinkVec_queue_dataIn_lo_hi_2, sinkVec_queue_6_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_6_enq_bits_vd;
  wire [2:0]   sinkVec_queue_6_enq_bits_offset;
  wire [7:0]   sinkVec_queue_dataIn_hi_hi_2 = {sinkVec_queue_6_enq_bits_vd, sinkVec_queue_6_enq_bits_offset};
  wire [3:0]   sinkVec_queue_6_enq_bits_mask;
  wire [11:0]  sinkVec_queue_dataIn_hi_6 = {sinkVec_queue_dataIn_hi_hi_2, sinkVec_queue_6_enq_bits_mask};
  wire [47:0]  sinkVec_queue_dataIn_6 = {sinkVec_queue_dataIn_hi_6, sinkVec_queue_dataIn_lo_6};
  wire [2:0]   sinkVec_queue_dataOut_6_instructionIndex = _sinkVec_queue_fifo_6_data_out[2:0];
  wire         sinkVec_queue_dataOut_6_last = _sinkVec_queue_fifo_6_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_6_data = _sinkVec_queue_fifo_6_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_6_mask = _sinkVec_queue_fifo_6_data_out[39:36];
  wire [2:0]   sinkVec_queue_dataOut_6_offset = _sinkVec_queue_fifo_6_data_out[42:40];
  wire [4:0]   sinkVec_queue_dataOut_6_vd = _sinkVec_queue_fifo_6_data_out[47:43];
  wire         sinkVec_queue_6_enq_ready = ~_sinkVec_queue_fifo_6_full;
  wire         sinkVec_queue_6_enq_valid;
  assign sinkVec_queue_6_deq_valid = ~_sinkVec_queue_fifo_6_empty | sinkVec_queue_6_enq_valid;
  assign sinkVec_queue_6_deq_bits_vd = _sinkVec_queue_fifo_6_empty ? sinkVec_queue_6_enq_bits_vd : sinkVec_queue_dataOut_6_vd;
  assign sinkVec_queue_6_deq_bits_offset = _sinkVec_queue_fifo_6_empty ? sinkVec_queue_6_enq_bits_offset : sinkVec_queue_dataOut_6_offset;
  assign sinkVec_queue_6_deq_bits_mask = _sinkVec_queue_fifo_6_empty ? sinkVec_queue_6_enq_bits_mask : sinkVec_queue_dataOut_6_mask;
  assign sinkVec_queue_6_deq_bits_data = _sinkVec_queue_fifo_6_empty ? sinkVec_queue_6_enq_bits_data : sinkVec_queue_dataOut_6_data;
  assign sinkVec_queue_6_deq_bits_last = ~_sinkVec_queue_fifo_6_empty & sinkVec_queue_dataOut_6_last;
  assign sinkVec_queue_6_deq_bits_instructionIndex = _sinkVec_queue_fifo_6_empty ? sinkVec_queue_6_enq_bits_instructionIndex : sinkVec_queue_dataOut_6_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_6;
  wire         sinkVec_releasePipe_pipe_out_6_valid = sinkVec_releasePipe_pipe_v_6;
  wire         x22_1_0_ready;
  wire         x22_1_0_valid;
  wire         sinkVec_validSource_6_valid = x22_1_0_ready & x22_1_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_6;
  wire [2:0]   sinkVec_tokenCheck_counterChange_6 = sinkVec_validSource_6_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_6 = ~(sinkVec_tokenCheck_counter_6[2]);
  assign x22_1_0_ready = sinkVec_tokenCheck_6;
  assign sinkVec_queue_6_enq_valid = sinkVec_validSink_6_valid;
  assign sinkVec_queue_6_enq_bits_vd = sinkVec_validSink_6_bits_vd;
  assign sinkVec_queue_6_enq_bits_offset = sinkVec_validSink_6_bits_offset;
  assign sinkVec_queue_6_enq_bits_mask = sinkVec_validSink_6_bits_mask;
  assign sinkVec_queue_6_enq_bits_data = sinkVec_validSink_6_bits_data;
  assign sinkVec_queue_6_enq_bits_instructionIndex = sinkVec_validSink_6_bits_instructionIndex;
  reg          sinkVec_shifterReg_6_0_valid;
  assign sinkVec_validSink_6_valid = sinkVec_shifterReg_6_0_valid;
  reg  [4:0]   sinkVec_shifterReg_6_0_bits_vd;
  assign sinkVec_validSink_6_bits_vd = sinkVec_shifterReg_6_0_bits_vd;
  reg  [2:0]   sinkVec_shifterReg_6_0_bits_offset;
  assign sinkVec_validSink_6_bits_offset = sinkVec_shifterReg_6_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_6_0_bits_mask;
  assign sinkVec_validSink_6_bits_mask = sinkVec_shifterReg_6_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_6_0_bits_data;
  assign sinkVec_validSink_6_bits_data = sinkVec_shifterReg_6_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_6_0_bits_instructionIndex;
  assign sinkVec_validSink_6_bits_instructionIndex = sinkVec_shifterReg_6_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_6 = sinkVec_shifterReg_6_0_valid | sinkVec_validSource_6_valid;
  wire         sinkVec_3_1_ready;
  wire         sinkVec_queue_7_deq_ready = sinkVec_sinkWire_7_ready;
  wire         sinkVec_queue_7_deq_valid;
  wire [4:0]   sinkVec_queue_7_deq_bits_vd;
  wire         sinkVec_3_1_valid = sinkVec_sinkWire_7_valid;
  wire [2:0]   sinkVec_queue_7_deq_bits_offset;
  wire [4:0]   sinkVec_3_1_bits_vd = sinkVec_sinkWire_7_bits_vd;
  wire [3:0]   sinkVec_queue_7_deq_bits_mask;
  wire [2:0]   sinkVec_3_1_bits_offset = sinkVec_sinkWire_7_bits_offset;
  wire [31:0]  sinkVec_queue_7_deq_bits_data;
  wire [3:0]   sinkVec_3_1_bits_mask = sinkVec_sinkWire_7_bits_mask;
  wire         sinkVec_queue_7_deq_bits_last;
  wire [31:0]  sinkVec_3_1_bits_data = sinkVec_sinkWire_7_bits_data;
  wire [2:0]   sinkVec_queue_7_deq_bits_instructionIndex;
  wire         sinkVec_3_1_bits_last = sinkVec_sinkWire_7_bits_last;
  wire [2:0]   sinkVec_3_1_bits_instructionIndex = sinkVec_sinkWire_7_bits_instructionIndex;
  wire         sinkVec_validSink_7_valid;
  wire [4:0]   sinkVec_validSink_7_bits_vd;
  wire [2:0]   sinkVec_validSink_7_bits_offset;
  wire [3:0]   sinkVec_validSink_7_bits_mask;
  wire [31:0]  sinkVec_validSink_7_bits_data;
  wire         sinkVec_validSink_7_bits_last;
  wire [2:0]   sinkVec_validSink_7_bits_instructionIndex;
  assign sinkVec_sinkWire_7_valid = sinkVec_queue_7_deq_valid;
  assign sinkVec_sinkWire_7_bits_vd = sinkVec_queue_7_deq_bits_vd;
  assign sinkVec_sinkWire_7_bits_offset = sinkVec_queue_7_deq_bits_offset;
  assign sinkVec_sinkWire_7_bits_mask = sinkVec_queue_7_deq_bits_mask;
  assign sinkVec_sinkWire_7_bits_data = sinkVec_queue_7_deq_bits_data;
  assign sinkVec_sinkWire_7_bits_last = sinkVec_queue_7_deq_bits_last;
  assign sinkVec_sinkWire_7_bits_instructionIndex = sinkVec_queue_7_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_7_enq_bits_data;
  wire         sinkVec_queue_7_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_3 = {sinkVec_queue_7_enq_bits_data, sinkVec_queue_7_enq_bits_last};
  wire [2:0]   sinkVec_queue_7_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_7 = {sinkVec_queue_dataIn_lo_hi_3, sinkVec_queue_7_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_7_enq_bits_vd;
  wire [2:0]   sinkVec_queue_7_enq_bits_offset;
  wire [7:0]   sinkVec_queue_dataIn_hi_hi_3 = {sinkVec_queue_7_enq_bits_vd, sinkVec_queue_7_enq_bits_offset};
  wire [3:0]   sinkVec_queue_7_enq_bits_mask;
  wire [11:0]  sinkVec_queue_dataIn_hi_7 = {sinkVec_queue_dataIn_hi_hi_3, sinkVec_queue_7_enq_bits_mask};
  wire [47:0]  sinkVec_queue_dataIn_7 = {sinkVec_queue_dataIn_hi_7, sinkVec_queue_dataIn_lo_7};
  wire [2:0]   sinkVec_queue_dataOut_7_instructionIndex = _sinkVec_queue_fifo_7_data_out[2:0];
  wire         sinkVec_queue_dataOut_7_last = _sinkVec_queue_fifo_7_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_7_data = _sinkVec_queue_fifo_7_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_7_mask = _sinkVec_queue_fifo_7_data_out[39:36];
  wire [2:0]   sinkVec_queue_dataOut_7_offset = _sinkVec_queue_fifo_7_data_out[42:40];
  wire [4:0]   sinkVec_queue_dataOut_7_vd = _sinkVec_queue_fifo_7_data_out[47:43];
  wire         sinkVec_queue_7_enq_ready = ~_sinkVec_queue_fifo_7_full;
  wire         sinkVec_queue_7_enq_valid;
  assign sinkVec_queue_7_deq_valid = ~_sinkVec_queue_fifo_7_empty | sinkVec_queue_7_enq_valid;
  assign sinkVec_queue_7_deq_bits_vd = _sinkVec_queue_fifo_7_empty ? sinkVec_queue_7_enq_bits_vd : sinkVec_queue_dataOut_7_vd;
  assign sinkVec_queue_7_deq_bits_offset = _sinkVec_queue_fifo_7_empty ? sinkVec_queue_7_enq_bits_offset : sinkVec_queue_dataOut_7_offset;
  assign sinkVec_queue_7_deq_bits_mask = _sinkVec_queue_fifo_7_empty ? sinkVec_queue_7_enq_bits_mask : sinkVec_queue_dataOut_7_mask;
  assign sinkVec_queue_7_deq_bits_data = _sinkVec_queue_fifo_7_empty ? sinkVec_queue_7_enq_bits_data : sinkVec_queue_dataOut_7_data;
  assign sinkVec_queue_7_deq_bits_last = _sinkVec_queue_fifo_7_empty ? sinkVec_queue_7_enq_bits_last : sinkVec_queue_dataOut_7_last;
  assign sinkVec_queue_7_deq_bits_instructionIndex = _sinkVec_queue_fifo_7_empty ? sinkVec_queue_7_enq_bits_instructionIndex : sinkVec_queue_dataOut_7_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_7;
  wire         sinkVec_releasePipe_pipe_out_7_valid = sinkVec_releasePipe_pipe_v_7;
  wire         x22_1_1_ready;
  wire         x22_1_1_valid;
  wire         sinkVec_validSource_7_valid = x22_1_1_ready & x22_1_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_7;
  wire [2:0]   sinkVec_tokenCheck_counterChange_7 = sinkVec_validSource_7_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_7 = ~(sinkVec_tokenCheck_counter_7[2]);
  assign x22_1_1_ready = sinkVec_tokenCheck_7;
  assign sinkVec_queue_7_enq_valid = sinkVec_validSink_7_valid;
  assign sinkVec_queue_7_enq_bits_vd = sinkVec_validSink_7_bits_vd;
  assign sinkVec_queue_7_enq_bits_offset = sinkVec_validSink_7_bits_offset;
  assign sinkVec_queue_7_enq_bits_mask = sinkVec_validSink_7_bits_mask;
  assign sinkVec_queue_7_enq_bits_data = sinkVec_validSink_7_bits_data;
  assign sinkVec_queue_7_enq_bits_last = sinkVec_validSink_7_bits_last;
  assign sinkVec_queue_7_enq_bits_instructionIndex = sinkVec_validSink_7_bits_instructionIndex;
  reg          sinkVec_shifterReg_7_0_valid;
  assign sinkVec_validSink_7_valid = sinkVec_shifterReg_7_0_valid;
  reg  [4:0]   sinkVec_shifterReg_7_0_bits_vd;
  assign sinkVec_validSink_7_bits_vd = sinkVec_shifterReg_7_0_bits_vd;
  reg  [2:0]   sinkVec_shifterReg_7_0_bits_offset;
  assign sinkVec_validSink_7_bits_offset = sinkVec_shifterReg_7_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_7_0_bits_mask;
  assign sinkVec_validSink_7_bits_mask = sinkVec_shifterReg_7_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_7_0_bits_data;
  assign sinkVec_validSink_7_bits_data = sinkVec_shifterReg_7_0_bits_data;
  reg          sinkVec_shifterReg_7_0_bits_last;
  assign sinkVec_validSink_7_bits_last = sinkVec_shifterReg_7_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_7_0_bits_instructionIndex;
  assign sinkVec_validSink_7_bits_instructionIndex = sinkVec_shifterReg_7_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_7 = sinkVec_shifterReg_7_0_valid | sinkVec_validSource_7_valid;
  assign sinkVec_sinkWire_6_ready = sinkVec_3_0_ready;
  assign sinkVec_sinkWire_7_ready = sinkVec_3_1_ready;
  reg          maskUnitFirst_3;
  wire         tryToRead_3 = sinkVec_3_0_valid | sinkVec_3_1_valid;
  wire         sinkWire_3_valid = maskUnitFirst_3 ? sinkVec_3_0_valid : sinkVec_3_1_valid;
  wire [4:0]   sinkWire_3_bits_vd = maskUnitFirst_3 ? sinkVec_3_0_bits_vd : sinkVec_3_1_bits_vd;
  wire [2:0]   sinkWire_3_bits_offset = maskUnitFirst_3 ? sinkVec_3_0_bits_offset : sinkVec_3_1_bits_offset;
  wire [3:0]   sinkWire_3_bits_mask = maskUnitFirst_3 ? sinkVec_3_0_bits_mask : sinkVec_3_1_bits_mask;
  wire [31:0]  sinkWire_3_bits_data = maskUnitFirst_3 ? sinkVec_3_0_bits_data : sinkVec_3_1_bits_data;
  wire         sinkWire_3_bits_last = maskUnitFirst_3 ? sinkVec_3_0_bits_last : sinkVec_3_1_bits_last;
  wire [2:0]   sinkWire_3_bits_instructionIndex = maskUnitFirst_3 ? sinkVec_3_0_bits_instructionIndex : sinkVec_3_1_bits_instructionIndex;
  wire         sinkWire_3_ready;
  assign sinkVec_3_1_ready = sinkWire_3_ready & ~maskUnitFirst_3;
  assign sinkVec_3_0_ready = sinkWire_3_ready & maskUnitFirst_3;
  reg          view__writeRelease_1_pipe_v;
  wire         view__writeRelease_1_pipe_out_valid = view__writeRelease_1_pipe_v;
  reg          pipe_v_3;
  wire         pipe_out_2_valid = pipe_v_3;
  wire         _probeWire_writeQueueEnqVec_1_valid_T = x22_1_0_ready & _maskUnit_exeResp_1_valid;
  reg          instructionFinishedPipe_pipe_v_1;
  wire         instructionFinishedPipe_pipe_out_1_valid = instructionFinishedPipe_pipe_v_1;
  reg  [7:0]   instructionFinishedPipe_pipe_b_1;
  wire [7:0]   instructionFinishedPipe_pipe_out_1_bits = instructionFinishedPipe_pipe_b_1;
  wire         instructionFinished_1_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_1_bits);
  wire         instructionFinished_1_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_1_bits);
  wire         instructionFinished_1_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_1_bits);
  wire         instructionFinished_1_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_1_bits);
  assign vxsatReportVec_1 = _laneVec_1_vxsatReport[3:0];
  reg          pipe_v_4;
  reg  [31:0]  pipe_b_4;
  reg          pipe_pipe_v_1;
  wire         pipe_pipe_out_1_valid = pipe_pipe_v_1;
  reg  [31:0]  pipe_pipe_b_1;
  wire [31:0]  pipe_pipe_out_1_bits = pipe_pipe_b_1;
  reg          view__laneMaskSelect_1_pipe_v;
  reg  [5:0]   view__laneMaskSelect_1_pipe_b;
  reg          view__laneMaskSelect_1_pipe_pipe_v;
  wire         view__laneMaskSelect_1_pipe_pipe_out_valid = view__laneMaskSelect_1_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_1_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_1_pipe_pipe_out_bits = view__laneMaskSelect_1_pipe_pipe_b;
  reg          view__laneMaskSewSelect_1_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_1_pipe_b;
  reg          view__laneMaskSewSelect_1_pipe_pipe_v;
  wire         view__laneMaskSewSelect_1_pipe_pipe_out_valid = view__laneMaskSewSelect_1_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_1_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_1_pipe_pipe_out_bits = view__laneMaskSewSelect_1_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v_1;
  wire         lsuLastPipe_pipe_out_1_valid = lsuLastPipe_pipe_v_1;
  reg  [7:0]   lsuLastPipe_pipe_b_1;
  wire [7:0]   lsuLastPipe_pipe_out_1_bits = lsuLastPipe_pipe_b_1;
  reg          maskLastPipe_pipe_v_1;
  wire         maskLastPipe_pipe_out_1_valid = maskLastPipe_pipe_v_1;
  reg  [7:0]   maskLastPipe_pipe_b_1;
  wire [7:0]   maskLastPipe_pipe_out_1_bits = maskLastPipe_pipe_b_1;
  wire [6:0]   writeCounter_1 = requestReg_bits_writeByte[11:5] + {6'h0, requestReg_bits_writeByte[4:0] > 5'h4};
  reg          pipe_v_5;
  wire         pipe_out_3_valid = pipe_v_5;
  reg  [6:0]   pipe_b_5;
  wire [6:0]   pipe_out_3_bits = pipe_b_5;
  assign laneRequestSinkWire_2_ready = ~laneRequestSinkWire_2_bits_issueInst | _laneVec_2_laneRequest_ready;
  wire         sinkVec_tokenCheck_8;
  wire [4:0]   sinkVec_validSource_8_bits_vs = x13_2_0_bits_vs;
  wire [2:0]   sinkVec_validSource_8_bits_offset = x13_2_0_bits_offset;
  wire [2:0]   sinkVec_validSource_8_bits_instructionIndex = x13_2_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_9;
  wire [4:0]   sinkVec_validSource_9_bits_vs = x13_2_1_bits_vs;
  wire [2:0]   sinkVec_validSource_9_bits_offset = x13_2_1_bits_offset;
  wire [2:0]   sinkVec_validSource_9_bits_instructionIndex = x13_2_1_bits_instructionIndex;
  wire         sinkVec_4_0_ready;
  wire         sinkVec_queue_8_deq_ready = sinkVec_sinkWire_8_ready;
  wire         sinkVec_queue_8_deq_valid;
  wire [4:0]   sinkVec_queue_8_deq_bits_vs;
  wire         sinkVec_4_0_valid = sinkVec_sinkWire_8_valid;
  wire [1:0]   sinkVec_queue_8_deq_bits_readSource;
  wire [4:0]   sinkVec_4_0_bits_vs = sinkVec_sinkWire_8_bits_vs;
  wire [2:0]   sinkVec_queue_8_deq_bits_offset;
  wire [1:0]   sinkVec_4_0_bits_readSource = sinkVec_sinkWire_8_bits_readSource;
  wire [2:0]   sinkVec_queue_8_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_4_0_bits_offset = sinkVec_sinkWire_8_bits_offset;
  wire [2:0]   sinkVec_4_0_bits_instructionIndex = sinkVec_sinkWire_8_bits_instructionIndex;
  wire         sinkVec_validSink_8_valid;
  wire [4:0]   sinkVec_validSink_8_bits_vs;
  wire [1:0]   sinkVec_validSink_8_bits_readSource;
  wire [2:0]   sinkVec_validSink_8_bits_offset;
  wire [2:0]   sinkVec_validSink_8_bits_instructionIndex;
  assign sinkVec_sinkWire_8_valid = sinkVec_queue_8_deq_valid;
  assign sinkVec_sinkWire_8_bits_vs = sinkVec_queue_8_deq_bits_vs;
  assign sinkVec_sinkWire_8_bits_readSource = sinkVec_queue_8_deq_bits_readSource;
  assign sinkVec_sinkWire_8_bits_offset = sinkVec_queue_8_deq_bits_offset;
  assign sinkVec_sinkWire_8_bits_instructionIndex = sinkVec_queue_8_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_queue_8_enq_bits_offset;
  wire [2:0]   sinkVec_queue_8_enq_bits_instructionIndex;
  wire [5:0]   sinkVec_queue_dataIn_lo_8 = {sinkVec_queue_8_enq_bits_offset, sinkVec_queue_8_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_8_enq_bits_vs;
  wire [1:0]   sinkVec_queue_8_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_8 = {sinkVec_queue_8_enq_bits_vs, sinkVec_queue_8_enq_bits_readSource};
  wire [12:0]  sinkVec_queue_dataIn_8 = {sinkVec_queue_dataIn_hi_8, sinkVec_queue_dataIn_lo_8};
  wire [2:0]   sinkVec_queue_dataOut_8_instructionIndex = _sinkVec_queue_fifo_8_data_out[2:0];
  wire [2:0]   sinkVec_queue_dataOut_8_offset = _sinkVec_queue_fifo_8_data_out[5:3];
  wire [1:0]   sinkVec_queue_dataOut_8_readSource = _sinkVec_queue_fifo_8_data_out[7:6];
  wire [4:0]   sinkVec_queue_dataOut_8_vs = _sinkVec_queue_fifo_8_data_out[12:8];
  wire         sinkVec_queue_8_enq_ready = ~_sinkVec_queue_fifo_8_full;
  wire         sinkVec_queue_8_enq_valid;
  assign sinkVec_queue_8_deq_valid = ~_sinkVec_queue_fifo_8_empty | sinkVec_queue_8_enq_valid;
  assign sinkVec_queue_8_deq_bits_vs = _sinkVec_queue_fifo_8_empty ? sinkVec_queue_8_enq_bits_vs : sinkVec_queue_dataOut_8_vs;
  assign sinkVec_queue_8_deq_bits_readSource = _sinkVec_queue_fifo_8_empty ? sinkVec_queue_8_enq_bits_readSource : sinkVec_queue_dataOut_8_readSource;
  assign sinkVec_queue_8_deq_bits_offset = _sinkVec_queue_fifo_8_empty ? sinkVec_queue_8_enq_bits_offset : sinkVec_queue_dataOut_8_offset;
  assign sinkVec_queue_8_deq_bits_instructionIndex = _sinkVec_queue_fifo_8_empty ? sinkVec_queue_8_enq_bits_instructionIndex : sinkVec_queue_dataOut_8_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_8;
  wire         sinkVec_releasePipe_pipe_out_8_valid = sinkVec_releasePipe_pipe_v_8;
  wire         x13_2_0_ready;
  wire         x13_2_0_valid;
  wire         sinkVec_validSource_8_valid = x13_2_0_ready & x13_2_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_8;
  wire [2:0]   sinkVec_tokenCheck_counterChange_8 = sinkVec_validSource_8_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_8 = ~(sinkVec_tokenCheck_counter_8[2]);
  assign x13_2_0_ready = sinkVec_tokenCheck_8;
  assign sinkVec_queue_8_enq_valid = sinkVec_validSink_8_valid;
  assign sinkVec_queue_8_enq_bits_vs = sinkVec_validSink_8_bits_vs;
  assign sinkVec_queue_8_enq_bits_readSource = sinkVec_validSink_8_bits_readSource;
  assign sinkVec_queue_8_enq_bits_offset = sinkVec_validSink_8_bits_offset;
  assign sinkVec_queue_8_enq_bits_instructionIndex = sinkVec_validSink_8_bits_instructionIndex;
  reg          sinkVec_shifterReg_8_0_valid;
  assign sinkVec_validSink_8_valid = sinkVec_shifterReg_8_0_valid;
  reg  [4:0]   sinkVec_shifterReg_8_0_bits_vs;
  assign sinkVec_validSink_8_bits_vs = sinkVec_shifterReg_8_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_8_0_bits_readSource;
  assign sinkVec_validSink_8_bits_readSource = sinkVec_shifterReg_8_0_bits_readSource;
  reg  [2:0]   sinkVec_shifterReg_8_0_bits_offset;
  assign sinkVec_validSink_8_bits_offset = sinkVec_shifterReg_8_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_8_0_bits_instructionIndex;
  assign sinkVec_validSink_8_bits_instructionIndex = sinkVec_shifterReg_8_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_8 = sinkVec_shifterReg_8_0_valid | sinkVec_validSource_8_valid;
  wire         sinkVec_4_1_ready;
  wire         sinkVec_queue_9_deq_ready = sinkVec_sinkWire_9_ready;
  wire         sinkVec_queue_9_deq_valid;
  wire [4:0]   sinkVec_queue_9_deq_bits_vs;
  wire         sinkVec_4_1_valid = sinkVec_sinkWire_9_valid;
  wire [1:0]   sinkVec_queue_9_deq_bits_readSource;
  wire [4:0]   sinkVec_4_1_bits_vs = sinkVec_sinkWire_9_bits_vs;
  wire [2:0]   sinkVec_queue_9_deq_bits_offset;
  wire [1:0]   sinkVec_4_1_bits_readSource = sinkVec_sinkWire_9_bits_readSource;
  wire [2:0]   sinkVec_queue_9_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_4_1_bits_offset = sinkVec_sinkWire_9_bits_offset;
  wire [2:0]   sinkVec_4_1_bits_instructionIndex = sinkVec_sinkWire_9_bits_instructionIndex;
  wire         sinkVec_validSink_9_valid;
  wire [4:0]   sinkVec_validSink_9_bits_vs;
  wire [1:0]   sinkVec_validSink_9_bits_readSource;
  wire [2:0]   sinkVec_validSink_9_bits_offset;
  wire [2:0]   sinkVec_validSink_9_bits_instructionIndex;
  assign sinkVec_sinkWire_9_valid = sinkVec_queue_9_deq_valid;
  assign sinkVec_sinkWire_9_bits_vs = sinkVec_queue_9_deq_bits_vs;
  assign sinkVec_sinkWire_9_bits_readSource = sinkVec_queue_9_deq_bits_readSource;
  assign sinkVec_sinkWire_9_bits_offset = sinkVec_queue_9_deq_bits_offset;
  assign sinkVec_sinkWire_9_bits_instructionIndex = sinkVec_queue_9_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_queue_9_enq_bits_offset;
  wire [2:0]   sinkVec_queue_9_enq_bits_instructionIndex;
  wire [5:0]   sinkVec_queue_dataIn_lo_9 = {sinkVec_queue_9_enq_bits_offset, sinkVec_queue_9_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_9_enq_bits_vs;
  wire [1:0]   sinkVec_queue_9_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_9 = {sinkVec_queue_9_enq_bits_vs, sinkVec_queue_9_enq_bits_readSource};
  wire [12:0]  sinkVec_queue_dataIn_9 = {sinkVec_queue_dataIn_hi_9, sinkVec_queue_dataIn_lo_9};
  wire [2:0]   sinkVec_queue_dataOut_9_instructionIndex = _sinkVec_queue_fifo_9_data_out[2:0];
  wire [2:0]   sinkVec_queue_dataOut_9_offset = _sinkVec_queue_fifo_9_data_out[5:3];
  wire [1:0]   sinkVec_queue_dataOut_9_readSource = _sinkVec_queue_fifo_9_data_out[7:6];
  wire [4:0]   sinkVec_queue_dataOut_9_vs = _sinkVec_queue_fifo_9_data_out[12:8];
  wire         sinkVec_queue_9_enq_ready = ~_sinkVec_queue_fifo_9_full;
  wire         sinkVec_queue_9_enq_valid;
  assign sinkVec_queue_9_deq_valid = ~_sinkVec_queue_fifo_9_empty | sinkVec_queue_9_enq_valid;
  assign sinkVec_queue_9_deq_bits_vs = _sinkVec_queue_fifo_9_empty ? sinkVec_queue_9_enq_bits_vs : sinkVec_queue_dataOut_9_vs;
  assign sinkVec_queue_9_deq_bits_readSource = _sinkVec_queue_fifo_9_empty ? sinkVec_queue_9_enq_bits_readSource : sinkVec_queue_dataOut_9_readSource;
  assign sinkVec_queue_9_deq_bits_offset = _sinkVec_queue_fifo_9_empty ? sinkVec_queue_9_enq_bits_offset : sinkVec_queue_dataOut_9_offset;
  assign sinkVec_queue_9_deq_bits_instructionIndex = _sinkVec_queue_fifo_9_empty ? sinkVec_queue_9_enq_bits_instructionIndex : sinkVec_queue_dataOut_9_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_9;
  wire         sinkVec_releasePipe_pipe_out_9_valid = sinkVec_releasePipe_pipe_v_9;
  wire         x13_2_1_ready;
  wire         x13_2_1_valid;
  wire         sinkVec_validSource_9_valid = x13_2_1_ready & x13_2_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_9;
  wire [2:0]   sinkVec_tokenCheck_counterChange_9 = sinkVec_validSource_9_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_9 = ~(sinkVec_tokenCheck_counter_9[2]);
  assign x13_2_1_ready = sinkVec_tokenCheck_9;
  assign sinkVec_queue_9_enq_valid = sinkVec_validSink_9_valid;
  assign sinkVec_queue_9_enq_bits_vs = sinkVec_validSink_9_bits_vs;
  assign sinkVec_queue_9_enq_bits_readSource = sinkVec_validSink_9_bits_readSource;
  assign sinkVec_queue_9_enq_bits_offset = sinkVec_validSink_9_bits_offset;
  assign sinkVec_queue_9_enq_bits_instructionIndex = sinkVec_validSink_9_bits_instructionIndex;
  reg          sinkVec_shifterReg_9_0_valid;
  assign sinkVec_validSink_9_valid = sinkVec_shifterReg_9_0_valid;
  reg  [4:0]   sinkVec_shifterReg_9_0_bits_vs;
  assign sinkVec_validSink_9_bits_vs = sinkVec_shifterReg_9_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_9_0_bits_readSource;
  assign sinkVec_validSink_9_bits_readSource = sinkVec_shifterReg_9_0_bits_readSource;
  reg  [2:0]   sinkVec_shifterReg_9_0_bits_offset;
  assign sinkVec_validSink_9_bits_offset = sinkVec_shifterReg_9_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_9_0_bits_instructionIndex;
  assign sinkVec_validSink_9_bits_instructionIndex = sinkVec_shifterReg_9_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_9 = sinkVec_shifterReg_9_0_valid | sinkVec_validSource_9_valid;
  assign sinkVec_sinkWire_8_ready = sinkVec_4_0_ready;
  assign sinkVec_sinkWire_9_ready = sinkVec_4_1_ready;
  reg          maskUnitFirst_4;
  wire         tryToRead_4 = sinkVec_4_0_valid | sinkVec_4_1_valid;
  wire         sinkWire_4_valid = maskUnitFirst_4 ? sinkVec_4_0_valid : sinkVec_4_1_valid;
  wire [4:0]   sinkWire_4_bits_vs = maskUnitFirst_4 ? sinkVec_4_0_bits_vs : sinkVec_4_1_bits_vs;
  wire [1:0]   sinkWire_4_bits_readSource = maskUnitFirst_4 ? sinkVec_4_0_bits_readSource : sinkVec_4_1_bits_readSource;
  wire [2:0]   sinkWire_4_bits_offset = maskUnitFirst_4 ? sinkVec_4_0_bits_offset : sinkVec_4_1_bits_offset;
  wire [2:0]   sinkWire_4_bits_instructionIndex = maskUnitFirst_4 ? sinkVec_4_0_bits_instructionIndex : sinkVec_4_1_bits_instructionIndex;
  wire         sinkWire_4_ready;
  assign sinkVec_4_1_ready = sinkWire_4_ready & ~maskUnitFirst_4;
  assign sinkVec_4_0_ready = sinkWire_4_ready & maskUnitFirst_4;
  reg          accessDataValid_pipe_v_4;
  reg          accessDataValid_pipe_pipe_v_4;
  wire         accessDataValid_pipe_pipe_out_4_valid = accessDataValid_pipe_pipe_v_4;
  wire         accessDataSource_4_valid = accessDataValid_pipe_pipe_out_4_valid;
  reg          shifterReg_12_0_valid;
  reg  [31:0]  shifterReg_12_0_bits;
  wire         shifterValid_12 = shifterReg_12_0_valid | accessDataSource_4_valid;
  reg          accessDataValid_pipe_v_5;
  reg          accessDataValid_pipe_pipe_v_5;
  wire         accessDataValid_pipe_pipe_out_5_valid = accessDataValid_pipe_pipe_v_5;
  wire         accessDataSource_5_valid = accessDataValid_pipe_pipe_out_5_valid;
  reg          shifterReg_13_0_valid;
  reg  [31:0]  shifterReg_13_0_bits;
  wire         shifterValid_13 = shifterReg_13_0_valid | accessDataSource_5_valid;
  wire         sinkVec_tokenCheck_10;
  wire [4:0]   sinkVec_validSource_10_bits_vd = x22_2_0_bits_vd;
  wire [2:0]   sinkVec_validSource_10_bits_offset = x22_2_0_bits_offset;
  wire [3:0]   sinkVec_validSource_10_bits_mask = x22_2_0_bits_mask;
  wire [31:0]  sinkVec_validSource_10_bits_data = x22_2_0_bits_data;
  wire [2:0]   sinkVec_validSource_10_bits_instructionIndex = x22_2_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_11;
  wire [4:0]   sinkVec_validSource_11_bits_vd = x22_2_1_bits_vd;
  wire [2:0]   sinkVec_validSource_11_bits_offset = x22_2_1_bits_offset;
  wire [3:0]   sinkVec_validSource_11_bits_mask = x22_2_1_bits_mask;
  wire [31:0]  sinkVec_validSource_11_bits_data = x22_2_1_bits_data;
  wire         sinkVec_validSource_11_bits_last = x22_2_1_bits_last;
  wire [2:0]   sinkVec_validSource_11_bits_instructionIndex = x22_2_1_bits_instructionIndex;
  wire         sinkVec_5_0_ready;
  wire         sinkVec_queue_10_deq_ready = sinkVec_sinkWire_10_ready;
  wire         sinkVec_queue_10_deq_valid;
  wire [4:0]   sinkVec_queue_10_deq_bits_vd;
  wire         sinkVec_5_0_valid = sinkVec_sinkWire_10_valid;
  wire [2:0]   sinkVec_queue_10_deq_bits_offset;
  wire [4:0]   sinkVec_5_0_bits_vd = sinkVec_sinkWire_10_bits_vd;
  wire [3:0]   sinkVec_queue_10_deq_bits_mask;
  wire [2:0]   sinkVec_5_0_bits_offset = sinkVec_sinkWire_10_bits_offset;
  wire [31:0]  sinkVec_queue_10_deq_bits_data;
  wire [3:0]   sinkVec_5_0_bits_mask = sinkVec_sinkWire_10_bits_mask;
  wire         sinkVec_queue_10_deq_bits_last;
  wire [31:0]  sinkVec_5_0_bits_data = sinkVec_sinkWire_10_bits_data;
  wire [2:0]   sinkVec_queue_10_deq_bits_instructionIndex;
  wire         sinkVec_5_0_bits_last = sinkVec_sinkWire_10_bits_last;
  wire [2:0]   sinkVec_5_0_bits_instructionIndex = sinkVec_sinkWire_10_bits_instructionIndex;
  wire         sinkVec_validSink_10_valid;
  wire [4:0]   sinkVec_validSink_10_bits_vd;
  wire [2:0]   sinkVec_validSink_10_bits_offset;
  wire [3:0]   sinkVec_validSink_10_bits_mask;
  wire [31:0]  sinkVec_validSink_10_bits_data;
  wire [2:0]   sinkVec_validSink_10_bits_instructionIndex;
  assign sinkVec_sinkWire_10_valid = sinkVec_queue_10_deq_valid;
  assign sinkVec_sinkWire_10_bits_vd = sinkVec_queue_10_deq_bits_vd;
  assign sinkVec_sinkWire_10_bits_offset = sinkVec_queue_10_deq_bits_offset;
  assign sinkVec_sinkWire_10_bits_mask = sinkVec_queue_10_deq_bits_mask;
  assign sinkVec_sinkWire_10_bits_data = sinkVec_queue_10_deq_bits_data;
  assign sinkVec_sinkWire_10_bits_last = sinkVec_queue_10_deq_bits_last;
  assign sinkVec_sinkWire_10_bits_instructionIndex = sinkVec_queue_10_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_10_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_4 = {sinkVec_queue_10_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_10_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_10 = {sinkVec_queue_dataIn_lo_hi_4, sinkVec_queue_10_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_10_enq_bits_vd;
  wire [2:0]   sinkVec_queue_10_enq_bits_offset;
  wire [7:0]   sinkVec_queue_dataIn_hi_hi_4 = {sinkVec_queue_10_enq_bits_vd, sinkVec_queue_10_enq_bits_offset};
  wire [3:0]   sinkVec_queue_10_enq_bits_mask;
  wire [11:0]  sinkVec_queue_dataIn_hi_10 = {sinkVec_queue_dataIn_hi_hi_4, sinkVec_queue_10_enq_bits_mask};
  wire [47:0]  sinkVec_queue_dataIn_10 = {sinkVec_queue_dataIn_hi_10, sinkVec_queue_dataIn_lo_10};
  wire [2:0]   sinkVec_queue_dataOut_10_instructionIndex = _sinkVec_queue_fifo_10_data_out[2:0];
  wire         sinkVec_queue_dataOut_10_last = _sinkVec_queue_fifo_10_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_10_data = _sinkVec_queue_fifo_10_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_10_mask = _sinkVec_queue_fifo_10_data_out[39:36];
  wire [2:0]   sinkVec_queue_dataOut_10_offset = _sinkVec_queue_fifo_10_data_out[42:40];
  wire [4:0]   sinkVec_queue_dataOut_10_vd = _sinkVec_queue_fifo_10_data_out[47:43];
  wire         sinkVec_queue_10_enq_ready = ~_sinkVec_queue_fifo_10_full;
  wire         sinkVec_queue_10_enq_valid;
  assign sinkVec_queue_10_deq_valid = ~_sinkVec_queue_fifo_10_empty | sinkVec_queue_10_enq_valid;
  assign sinkVec_queue_10_deq_bits_vd = _sinkVec_queue_fifo_10_empty ? sinkVec_queue_10_enq_bits_vd : sinkVec_queue_dataOut_10_vd;
  assign sinkVec_queue_10_deq_bits_offset = _sinkVec_queue_fifo_10_empty ? sinkVec_queue_10_enq_bits_offset : sinkVec_queue_dataOut_10_offset;
  assign sinkVec_queue_10_deq_bits_mask = _sinkVec_queue_fifo_10_empty ? sinkVec_queue_10_enq_bits_mask : sinkVec_queue_dataOut_10_mask;
  assign sinkVec_queue_10_deq_bits_data = _sinkVec_queue_fifo_10_empty ? sinkVec_queue_10_enq_bits_data : sinkVec_queue_dataOut_10_data;
  assign sinkVec_queue_10_deq_bits_last = ~_sinkVec_queue_fifo_10_empty & sinkVec_queue_dataOut_10_last;
  assign sinkVec_queue_10_deq_bits_instructionIndex = _sinkVec_queue_fifo_10_empty ? sinkVec_queue_10_enq_bits_instructionIndex : sinkVec_queue_dataOut_10_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_10;
  wire         sinkVec_releasePipe_pipe_out_10_valid = sinkVec_releasePipe_pipe_v_10;
  wire         x22_2_0_ready;
  wire         x22_2_0_valid;
  wire         sinkVec_validSource_10_valid = x22_2_0_ready & x22_2_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_10;
  wire [2:0]   sinkVec_tokenCheck_counterChange_10 = sinkVec_validSource_10_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_10 = ~(sinkVec_tokenCheck_counter_10[2]);
  assign x22_2_0_ready = sinkVec_tokenCheck_10;
  assign sinkVec_queue_10_enq_valid = sinkVec_validSink_10_valid;
  assign sinkVec_queue_10_enq_bits_vd = sinkVec_validSink_10_bits_vd;
  assign sinkVec_queue_10_enq_bits_offset = sinkVec_validSink_10_bits_offset;
  assign sinkVec_queue_10_enq_bits_mask = sinkVec_validSink_10_bits_mask;
  assign sinkVec_queue_10_enq_bits_data = sinkVec_validSink_10_bits_data;
  assign sinkVec_queue_10_enq_bits_instructionIndex = sinkVec_validSink_10_bits_instructionIndex;
  reg          sinkVec_shifterReg_10_0_valid;
  assign sinkVec_validSink_10_valid = sinkVec_shifterReg_10_0_valid;
  reg  [4:0]   sinkVec_shifterReg_10_0_bits_vd;
  assign sinkVec_validSink_10_bits_vd = sinkVec_shifterReg_10_0_bits_vd;
  reg  [2:0]   sinkVec_shifterReg_10_0_bits_offset;
  assign sinkVec_validSink_10_bits_offset = sinkVec_shifterReg_10_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_10_0_bits_mask;
  assign sinkVec_validSink_10_bits_mask = sinkVec_shifterReg_10_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_10_0_bits_data;
  assign sinkVec_validSink_10_bits_data = sinkVec_shifterReg_10_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_10_0_bits_instructionIndex;
  assign sinkVec_validSink_10_bits_instructionIndex = sinkVec_shifterReg_10_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_10 = sinkVec_shifterReg_10_0_valid | sinkVec_validSource_10_valid;
  wire         sinkVec_5_1_ready;
  wire         sinkVec_queue_11_deq_ready = sinkVec_sinkWire_11_ready;
  wire         sinkVec_queue_11_deq_valid;
  wire [4:0]   sinkVec_queue_11_deq_bits_vd;
  wire         sinkVec_5_1_valid = sinkVec_sinkWire_11_valid;
  wire [2:0]   sinkVec_queue_11_deq_bits_offset;
  wire [4:0]   sinkVec_5_1_bits_vd = sinkVec_sinkWire_11_bits_vd;
  wire [3:0]   sinkVec_queue_11_deq_bits_mask;
  wire [2:0]   sinkVec_5_1_bits_offset = sinkVec_sinkWire_11_bits_offset;
  wire [31:0]  sinkVec_queue_11_deq_bits_data;
  wire [3:0]   sinkVec_5_1_bits_mask = sinkVec_sinkWire_11_bits_mask;
  wire         sinkVec_queue_11_deq_bits_last;
  wire [31:0]  sinkVec_5_1_bits_data = sinkVec_sinkWire_11_bits_data;
  wire [2:0]   sinkVec_queue_11_deq_bits_instructionIndex;
  wire         sinkVec_5_1_bits_last = sinkVec_sinkWire_11_bits_last;
  wire [2:0]   sinkVec_5_1_bits_instructionIndex = sinkVec_sinkWire_11_bits_instructionIndex;
  wire         sinkVec_validSink_11_valid;
  wire [4:0]   sinkVec_validSink_11_bits_vd;
  wire [2:0]   sinkVec_validSink_11_bits_offset;
  wire [3:0]   sinkVec_validSink_11_bits_mask;
  wire [31:0]  sinkVec_validSink_11_bits_data;
  wire         sinkVec_validSink_11_bits_last;
  wire [2:0]   sinkVec_validSink_11_bits_instructionIndex;
  assign sinkVec_sinkWire_11_valid = sinkVec_queue_11_deq_valid;
  assign sinkVec_sinkWire_11_bits_vd = sinkVec_queue_11_deq_bits_vd;
  assign sinkVec_sinkWire_11_bits_offset = sinkVec_queue_11_deq_bits_offset;
  assign sinkVec_sinkWire_11_bits_mask = sinkVec_queue_11_deq_bits_mask;
  assign sinkVec_sinkWire_11_bits_data = sinkVec_queue_11_deq_bits_data;
  assign sinkVec_sinkWire_11_bits_last = sinkVec_queue_11_deq_bits_last;
  assign sinkVec_sinkWire_11_bits_instructionIndex = sinkVec_queue_11_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_11_enq_bits_data;
  wire         sinkVec_queue_11_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_5 = {sinkVec_queue_11_enq_bits_data, sinkVec_queue_11_enq_bits_last};
  wire [2:0]   sinkVec_queue_11_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_11 = {sinkVec_queue_dataIn_lo_hi_5, sinkVec_queue_11_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_11_enq_bits_vd;
  wire [2:0]   sinkVec_queue_11_enq_bits_offset;
  wire [7:0]   sinkVec_queue_dataIn_hi_hi_5 = {sinkVec_queue_11_enq_bits_vd, sinkVec_queue_11_enq_bits_offset};
  wire [3:0]   sinkVec_queue_11_enq_bits_mask;
  wire [11:0]  sinkVec_queue_dataIn_hi_11 = {sinkVec_queue_dataIn_hi_hi_5, sinkVec_queue_11_enq_bits_mask};
  wire [47:0]  sinkVec_queue_dataIn_11 = {sinkVec_queue_dataIn_hi_11, sinkVec_queue_dataIn_lo_11};
  wire [2:0]   sinkVec_queue_dataOut_11_instructionIndex = _sinkVec_queue_fifo_11_data_out[2:0];
  wire         sinkVec_queue_dataOut_11_last = _sinkVec_queue_fifo_11_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_11_data = _sinkVec_queue_fifo_11_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_11_mask = _sinkVec_queue_fifo_11_data_out[39:36];
  wire [2:0]   sinkVec_queue_dataOut_11_offset = _sinkVec_queue_fifo_11_data_out[42:40];
  wire [4:0]   sinkVec_queue_dataOut_11_vd = _sinkVec_queue_fifo_11_data_out[47:43];
  wire         sinkVec_queue_11_enq_ready = ~_sinkVec_queue_fifo_11_full;
  wire         sinkVec_queue_11_enq_valid;
  assign sinkVec_queue_11_deq_valid = ~_sinkVec_queue_fifo_11_empty | sinkVec_queue_11_enq_valid;
  assign sinkVec_queue_11_deq_bits_vd = _sinkVec_queue_fifo_11_empty ? sinkVec_queue_11_enq_bits_vd : sinkVec_queue_dataOut_11_vd;
  assign sinkVec_queue_11_deq_bits_offset = _sinkVec_queue_fifo_11_empty ? sinkVec_queue_11_enq_bits_offset : sinkVec_queue_dataOut_11_offset;
  assign sinkVec_queue_11_deq_bits_mask = _sinkVec_queue_fifo_11_empty ? sinkVec_queue_11_enq_bits_mask : sinkVec_queue_dataOut_11_mask;
  assign sinkVec_queue_11_deq_bits_data = _sinkVec_queue_fifo_11_empty ? sinkVec_queue_11_enq_bits_data : sinkVec_queue_dataOut_11_data;
  assign sinkVec_queue_11_deq_bits_last = _sinkVec_queue_fifo_11_empty ? sinkVec_queue_11_enq_bits_last : sinkVec_queue_dataOut_11_last;
  assign sinkVec_queue_11_deq_bits_instructionIndex = _sinkVec_queue_fifo_11_empty ? sinkVec_queue_11_enq_bits_instructionIndex : sinkVec_queue_dataOut_11_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_11;
  wire         sinkVec_releasePipe_pipe_out_11_valid = sinkVec_releasePipe_pipe_v_11;
  wire         x22_2_1_ready;
  wire         x22_2_1_valid;
  wire         sinkVec_validSource_11_valid = x22_2_1_ready & x22_2_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_11;
  wire [2:0]   sinkVec_tokenCheck_counterChange_11 = sinkVec_validSource_11_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_11 = ~(sinkVec_tokenCheck_counter_11[2]);
  assign x22_2_1_ready = sinkVec_tokenCheck_11;
  assign sinkVec_queue_11_enq_valid = sinkVec_validSink_11_valid;
  assign sinkVec_queue_11_enq_bits_vd = sinkVec_validSink_11_bits_vd;
  assign sinkVec_queue_11_enq_bits_offset = sinkVec_validSink_11_bits_offset;
  assign sinkVec_queue_11_enq_bits_mask = sinkVec_validSink_11_bits_mask;
  assign sinkVec_queue_11_enq_bits_data = sinkVec_validSink_11_bits_data;
  assign sinkVec_queue_11_enq_bits_last = sinkVec_validSink_11_bits_last;
  assign sinkVec_queue_11_enq_bits_instructionIndex = sinkVec_validSink_11_bits_instructionIndex;
  reg          sinkVec_shifterReg_11_0_valid;
  assign sinkVec_validSink_11_valid = sinkVec_shifterReg_11_0_valid;
  reg  [4:0]   sinkVec_shifterReg_11_0_bits_vd;
  assign sinkVec_validSink_11_bits_vd = sinkVec_shifterReg_11_0_bits_vd;
  reg  [2:0]   sinkVec_shifterReg_11_0_bits_offset;
  assign sinkVec_validSink_11_bits_offset = sinkVec_shifterReg_11_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_11_0_bits_mask;
  assign sinkVec_validSink_11_bits_mask = sinkVec_shifterReg_11_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_11_0_bits_data;
  assign sinkVec_validSink_11_bits_data = sinkVec_shifterReg_11_0_bits_data;
  reg          sinkVec_shifterReg_11_0_bits_last;
  assign sinkVec_validSink_11_bits_last = sinkVec_shifterReg_11_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_11_0_bits_instructionIndex;
  assign sinkVec_validSink_11_bits_instructionIndex = sinkVec_shifterReg_11_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_11 = sinkVec_shifterReg_11_0_valid | sinkVec_validSource_11_valid;
  assign sinkVec_sinkWire_10_ready = sinkVec_5_0_ready;
  assign sinkVec_sinkWire_11_ready = sinkVec_5_1_ready;
  reg          maskUnitFirst_5;
  wire         tryToRead_5 = sinkVec_5_0_valid | sinkVec_5_1_valid;
  wire         sinkWire_5_valid = maskUnitFirst_5 ? sinkVec_5_0_valid : sinkVec_5_1_valid;
  wire [4:0]   sinkWire_5_bits_vd = maskUnitFirst_5 ? sinkVec_5_0_bits_vd : sinkVec_5_1_bits_vd;
  wire [2:0]   sinkWire_5_bits_offset = maskUnitFirst_5 ? sinkVec_5_0_bits_offset : sinkVec_5_1_bits_offset;
  wire [3:0]   sinkWire_5_bits_mask = maskUnitFirst_5 ? sinkVec_5_0_bits_mask : sinkVec_5_1_bits_mask;
  wire [31:0]  sinkWire_5_bits_data = maskUnitFirst_5 ? sinkVec_5_0_bits_data : sinkVec_5_1_bits_data;
  wire         sinkWire_5_bits_last = maskUnitFirst_5 ? sinkVec_5_0_bits_last : sinkVec_5_1_bits_last;
  wire [2:0]   sinkWire_5_bits_instructionIndex = maskUnitFirst_5 ? sinkVec_5_0_bits_instructionIndex : sinkVec_5_1_bits_instructionIndex;
  wire         sinkWire_5_ready;
  assign sinkVec_5_1_ready = sinkWire_5_ready & ~maskUnitFirst_5;
  assign sinkVec_5_0_ready = sinkWire_5_ready & maskUnitFirst_5;
  reg          view__writeRelease_2_pipe_v;
  wire         view__writeRelease_2_pipe_out_valid = view__writeRelease_2_pipe_v;
  reg          pipe_v_6;
  wire         pipe_out_4_valid = pipe_v_6;
  wire         _probeWire_writeQueueEnqVec_2_valid_T = x22_2_0_ready & _maskUnit_exeResp_2_valid;
  reg          instructionFinishedPipe_pipe_v_2;
  wire         instructionFinishedPipe_pipe_out_2_valid = instructionFinishedPipe_pipe_v_2;
  reg  [7:0]   instructionFinishedPipe_pipe_b_2;
  wire [7:0]   instructionFinishedPipe_pipe_out_2_bits = instructionFinishedPipe_pipe_b_2;
  wire         instructionFinished_2_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_2_bits);
  wire         instructionFinished_2_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_2_bits);
  wire         instructionFinished_2_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_2_bits);
  wire         instructionFinished_2_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_2_bits);
  assign vxsatReportVec_2 = _laneVec_2_vxsatReport[3:0];
  reg          pipe_v_7;
  reg  [31:0]  pipe_b_7;
  reg          pipe_pipe_v_2;
  wire         pipe_pipe_out_2_valid = pipe_pipe_v_2;
  reg  [31:0]  pipe_pipe_b_2;
  wire [31:0]  pipe_pipe_out_2_bits = pipe_pipe_b_2;
  reg          view__laneMaskSelect_2_pipe_v;
  reg  [5:0]   view__laneMaskSelect_2_pipe_b;
  reg          view__laneMaskSelect_2_pipe_pipe_v;
  wire         view__laneMaskSelect_2_pipe_pipe_out_valid = view__laneMaskSelect_2_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_2_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_2_pipe_pipe_out_bits = view__laneMaskSelect_2_pipe_pipe_b;
  reg          view__laneMaskSewSelect_2_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_2_pipe_b;
  reg          view__laneMaskSewSelect_2_pipe_pipe_v;
  wire         view__laneMaskSewSelect_2_pipe_pipe_out_valid = view__laneMaskSewSelect_2_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_2_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_2_pipe_pipe_out_bits = view__laneMaskSewSelect_2_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v_2;
  wire         lsuLastPipe_pipe_out_2_valid = lsuLastPipe_pipe_v_2;
  reg  [7:0]   lsuLastPipe_pipe_b_2;
  wire [7:0]   lsuLastPipe_pipe_out_2_bits = lsuLastPipe_pipe_b_2;
  reg          maskLastPipe_pipe_v_2;
  wire         maskLastPipe_pipe_out_2_valid = maskLastPipe_pipe_v_2;
  reg  [7:0]   maskLastPipe_pipe_b_2;
  wire [7:0]   maskLastPipe_pipe_out_2_bits = maskLastPipe_pipe_b_2;
  wire [6:0]   writeCounter_2 = requestReg_bits_writeByte[11:5] + {6'h0, requestReg_bits_writeByte[4:0] > 5'h8};
  reg          pipe_v_8;
  wire         pipe_out_5_valid = pipe_v_8;
  reg  [6:0]   pipe_b_8;
  wire [6:0]   pipe_out_5_bits = pipe_b_8;
  assign laneRequestSinkWire_3_ready = ~laneRequestSinkWire_3_bits_issueInst | _laneVec_3_laneRequest_ready;
  wire         sinkVec_tokenCheck_12;
  wire [4:0]   sinkVec_validSource_12_bits_vs = x13_3_0_bits_vs;
  wire [2:0]   sinkVec_validSource_12_bits_offset = x13_3_0_bits_offset;
  wire [2:0]   sinkVec_validSource_12_bits_instructionIndex = x13_3_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_13;
  wire [4:0]   sinkVec_validSource_13_bits_vs = x13_3_1_bits_vs;
  wire [2:0]   sinkVec_validSource_13_bits_offset = x13_3_1_bits_offset;
  wire [2:0]   sinkVec_validSource_13_bits_instructionIndex = x13_3_1_bits_instructionIndex;
  wire         sinkVec_6_0_ready;
  wire         sinkVec_queue_12_deq_ready = sinkVec_sinkWire_12_ready;
  wire         sinkVec_queue_12_deq_valid;
  wire [4:0]   sinkVec_queue_12_deq_bits_vs;
  wire         sinkVec_6_0_valid = sinkVec_sinkWire_12_valid;
  wire [1:0]   sinkVec_queue_12_deq_bits_readSource;
  wire [4:0]   sinkVec_6_0_bits_vs = sinkVec_sinkWire_12_bits_vs;
  wire [2:0]   sinkVec_queue_12_deq_bits_offset;
  wire [1:0]   sinkVec_6_0_bits_readSource = sinkVec_sinkWire_12_bits_readSource;
  wire [2:0]   sinkVec_queue_12_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_6_0_bits_offset = sinkVec_sinkWire_12_bits_offset;
  wire [2:0]   sinkVec_6_0_bits_instructionIndex = sinkVec_sinkWire_12_bits_instructionIndex;
  wire         sinkVec_validSink_12_valid;
  wire [4:0]   sinkVec_validSink_12_bits_vs;
  wire [1:0]   sinkVec_validSink_12_bits_readSource;
  wire [2:0]   sinkVec_validSink_12_bits_offset;
  wire [2:0]   sinkVec_validSink_12_bits_instructionIndex;
  assign sinkVec_sinkWire_12_valid = sinkVec_queue_12_deq_valid;
  assign sinkVec_sinkWire_12_bits_vs = sinkVec_queue_12_deq_bits_vs;
  assign sinkVec_sinkWire_12_bits_readSource = sinkVec_queue_12_deq_bits_readSource;
  assign sinkVec_sinkWire_12_bits_offset = sinkVec_queue_12_deq_bits_offset;
  assign sinkVec_sinkWire_12_bits_instructionIndex = sinkVec_queue_12_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_queue_12_enq_bits_offset;
  wire [2:0]   sinkVec_queue_12_enq_bits_instructionIndex;
  wire [5:0]   sinkVec_queue_dataIn_lo_12 = {sinkVec_queue_12_enq_bits_offset, sinkVec_queue_12_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_12_enq_bits_vs;
  wire [1:0]   sinkVec_queue_12_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_12 = {sinkVec_queue_12_enq_bits_vs, sinkVec_queue_12_enq_bits_readSource};
  wire [12:0]  sinkVec_queue_dataIn_12 = {sinkVec_queue_dataIn_hi_12, sinkVec_queue_dataIn_lo_12};
  wire [2:0]   sinkVec_queue_dataOut_12_instructionIndex = _sinkVec_queue_fifo_12_data_out[2:0];
  wire [2:0]   sinkVec_queue_dataOut_12_offset = _sinkVec_queue_fifo_12_data_out[5:3];
  wire [1:0]   sinkVec_queue_dataOut_12_readSource = _sinkVec_queue_fifo_12_data_out[7:6];
  wire [4:0]   sinkVec_queue_dataOut_12_vs = _sinkVec_queue_fifo_12_data_out[12:8];
  wire         sinkVec_queue_12_enq_ready = ~_sinkVec_queue_fifo_12_full;
  wire         sinkVec_queue_12_enq_valid;
  assign sinkVec_queue_12_deq_valid = ~_sinkVec_queue_fifo_12_empty | sinkVec_queue_12_enq_valid;
  assign sinkVec_queue_12_deq_bits_vs = _sinkVec_queue_fifo_12_empty ? sinkVec_queue_12_enq_bits_vs : sinkVec_queue_dataOut_12_vs;
  assign sinkVec_queue_12_deq_bits_readSource = _sinkVec_queue_fifo_12_empty ? sinkVec_queue_12_enq_bits_readSource : sinkVec_queue_dataOut_12_readSource;
  assign sinkVec_queue_12_deq_bits_offset = _sinkVec_queue_fifo_12_empty ? sinkVec_queue_12_enq_bits_offset : sinkVec_queue_dataOut_12_offset;
  assign sinkVec_queue_12_deq_bits_instructionIndex = _sinkVec_queue_fifo_12_empty ? sinkVec_queue_12_enq_bits_instructionIndex : sinkVec_queue_dataOut_12_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_12;
  wire         sinkVec_releasePipe_pipe_out_12_valid = sinkVec_releasePipe_pipe_v_12;
  wire         x13_3_0_ready;
  wire         x13_3_0_valid;
  wire         sinkVec_validSource_12_valid = x13_3_0_ready & x13_3_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_12;
  wire [2:0]   sinkVec_tokenCheck_counterChange_12 = sinkVec_validSource_12_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_12 = ~(sinkVec_tokenCheck_counter_12[2]);
  assign x13_3_0_ready = sinkVec_tokenCheck_12;
  assign sinkVec_queue_12_enq_valid = sinkVec_validSink_12_valid;
  assign sinkVec_queue_12_enq_bits_vs = sinkVec_validSink_12_bits_vs;
  assign sinkVec_queue_12_enq_bits_readSource = sinkVec_validSink_12_bits_readSource;
  assign sinkVec_queue_12_enq_bits_offset = sinkVec_validSink_12_bits_offset;
  assign sinkVec_queue_12_enq_bits_instructionIndex = sinkVec_validSink_12_bits_instructionIndex;
  reg          sinkVec_shifterReg_12_0_valid;
  assign sinkVec_validSink_12_valid = sinkVec_shifterReg_12_0_valid;
  reg  [4:0]   sinkVec_shifterReg_12_0_bits_vs;
  assign sinkVec_validSink_12_bits_vs = sinkVec_shifterReg_12_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_12_0_bits_readSource;
  assign sinkVec_validSink_12_bits_readSource = sinkVec_shifterReg_12_0_bits_readSource;
  reg  [2:0]   sinkVec_shifterReg_12_0_bits_offset;
  assign sinkVec_validSink_12_bits_offset = sinkVec_shifterReg_12_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_12_0_bits_instructionIndex;
  assign sinkVec_validSink_12_bits_instructionIndex = sinkVec_shifterReg_12_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_12 = sinkVec_shifterReg_12_0_valid | sinkVec_validSource_12_valid;
  wire         sinkVec_6_1_ready;
  wire         sinkVec_queue_13_deq_ready = sinkVec_sinkWire_13_ready;
  wire         sinkVec_queue_13_deq_valid;
  wire [4:0]   sinkVec_queue_13_deq_bits_vs;
  wire         sinkVec_6_1_valid = sinkVec_sinkWire_13_valid;
  wire [1:0]   sinkVec_queue_13_deq_bits_readSource;
  wire [4:0]   sinkVec_6_1_bits_vs = sinkVec_sinkWire_13_bits_vs;
  wire [2:0]   sinkVec_queue_13_deq_bits_offset;
  wire [1:0]   sinkVec_6_1_bits_readSource = sinkVec_sinkWire_13_bits_readSource;
  wire [2:0]   sinkVec_queue_13_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_6_1_bits_offset = sinkVec_sinkWire_13_bits_offset;
  wire [2:0]   sinkVec_6_1_bits_instructionIndex = sinkVec_sinkWire_13_bits_instructionIndex;
  wire         sinkVec_validSink_13_valid;
  wire [4:0]   sinkVec_validSink_13_bits_vs;
  wire [1:0]   sinkVec_validSink_13_bits_readSource;
  wire [2:0]   sinkVec_validSink_13_bits_offset;
  wire [2:0]   sinkVec_validSink_13_bits_instructionIndex;
  assign sinkVec_sinkWire_13_valid = sinkVec_queue_13_deq_valid;
  assign sinkVec_sinkWire_13_bits_vs = sinkVec_queue_13_deq_bits_vs;
  assign sinkVec_sinkWire_13_bits_readSource = sinkVec_queue_13_deq_bits_readSource;
  assign sinkVec_sinkWire_13_bits_offset = sinkVec_queue_13_deq_bits_offset;
  assign sinkVec_sinkWire_13_bits_instructionIndex = sinkVec_queue_13_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_queue_13_enq_bits_offset;
  wire [2:0]   sinkVec_queue_13_enq_bits_instructionIndex;
  wire [5:0]   sinkVec_queue_dataIn_lo_13 = {sinkVec_queue_13_enq_bits_offset, sinkVec_queue_13_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_13_enq_bits_vs;
  wire [1:0]   sinkVec_queue_13_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_13 = {sinkVec_queue_13_enq_bits_vs, sinkVec_queue_13_enq_bits_readSource};
  wire [12:0]  sinkVec_queue_dataIn_13 = {sinkVec_queue_dataIn_hi_13, sinkVec_queue_dataIn_lo_13};
  wire [2:0]   sinkVec_queue_dataOut_13_instructionIndex = _sinkVec_queue_fifo_13_data_out[2:0];
  wire [2:0]   sinkVec_queue_dataOut_13_offset = _sinkVec_queue_fifo_13_data_out[5:3];
  wire [1:0]   sinkVec_queue_dataOut_13_readSource = _sinkVec_queue_fifo_13_data_out[7:6];
  wire [4:0]   sinkVec_queue_dataOut_13_vs = _sinkVec_queue_fifo_13_data_out[12:8];
  wire         sinkVec_queue_13_enq_ready = ~_sinkVec_queue_fifo_13_full;
  wire         sinkVec_queue_13_enq_valid;
  assign sinkVec_queue_13_deq_valid = ~_sinkVec_queue_fifo_13_empty | sinkVec_queue_13_enq_valid;
  assign sinkVec_queue_13_deq_bits_vs = _sinkVec_queue_fifo_13_empty ? sinkVec_queue_13_enq_bits_vs : sinkVec_queue_dataOut_13_vs;
  assign sinkVec_queue_13_deq_bits_readSource = _sinkVec_queue_fifo_13_empty ? sinkVec_queue_13_enq_bits_readSource : sinkVec_queue_dataOut_13_readSource;
  assign sinkVec_queue_13_deq_bits_offset = _sinkVec_queue_fifo_13_empty ? sinkVec_queue_13_enq_bits_offset : sinkVec_queue_dataOut_13_offset;
  assign sinkVec_queue_13_deq_bits_instructionIndex = _sinkVec_queue_fifo_13_empty ? sinkVec_queue_13_enq_bits_instructionIndex : sinkVec_queue_dataOut_13_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_13;
  wire         sinkVec_releasePipe_pipe_out_13_valid = sinkVec_releasePipe_pipe_v_13;
  wire         x13_3_1_ready;
  wire         x13_3_1_valid;
  wire         sinkVec_validSource_13_valid = x13_3_1_ready & x13_3_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_13;
  wire [2:0]   sinkVec_tokenCheck_counterChange_13 = sinkVec_validSource_13_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_13 = ~(sinkVec_tokenCheck_counter_13[2]);
  assign x13_3_1_ready = sinkVec_tokenCheck_13;
  assign sinkVec_queue_13_enq_valid = sinkVec_validSink_13_valid;
  assign sinkVec_queue_13_enq_bits_vs = sinkVec_validSink_13_bits_vs;
  assign sinkVec_queue_13_enq_bits_readSource = sinkVec_validSink_13_bits_readSource;
  assign sinkVec_queue_13_enq_bits_offset = sinkVec_validSink_13_bits_offset;
  assign sinkVec_queue_13_enq_bits_instructionIndex = sinkVec_validSink_13_bits_instructionIndex;
  reg          sinkVec_shifterReg_13_0_valid;
  assign sinkVec_validSink_13_valid = sinkVec_shifterReg_13_0_valid;
  reg  [4:0]   sinkVec_shifterReg_13_0_bits_vs;
  assign sinkVec_validSink_13_bits_vs = sinkVec_shifterReg_13_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_13_0_bits_readSource;
  assign sinkVec_validSink_13_bits_readSource = sinkVec_shifterReg_13_0_bits_readSource;
  reg  [2:0]   sinkVec_shifterReg_13_0_bits_offset;
  assign sinkVec_validSink_13_bits_offset = sinkVec_shifterReg_13_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_13_0_bits_instructionIndex;
  assign sinkVec_validSink_13_bits_instructionIndex = sinkVec_shifterReg_13_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_13 = sinkVec_shifterReg_13_0_valid | sinkVec_validSource_13_valid;
  assign sinkVec_sinkWire_12_ready = sinkVec_6_0_ready;
  assign sinkVec_sinkWire_13_ready = sinkVec_6_1_ready;
  reg          maskUnitFirst_6;
  wire         tryToRead_6 = sinkVec_6_0_valid | sinkVec_6_1_valid;
  wire         sinkWire_6_valid = maskUnitFirst_6 ? sinkVec_6_0_valid : sinkVec_6_1_valid;
  wire [4:0]   sinkWire_6_bits_vs = maskUnitFirst_6 ? sinkVec_6_0_bits_vs : sinkVec_6_1_bits_vs;
  wire [1:0]   sinkWire_6_bits_readSource = maskUnitFirst_6 ? sinkVec_6_0_bits_readSource : sinkVec_6_1_bits_readSource;
  wire [2:0]   sinkWire_6_bits_offset = maskUnitFirst_6 ? sinkVec_6_0_bits_offset : sinkVec_6_1_bits_offset;
  wire [2:0]   sinkWire_6_bits_instructionIndex = maskUnitFirst_6 ? sinkVec_6_0_bits_instructionIndex : sinkVec_6_1_bits_instructionIndex;
  wire         sinkWire_6_ready;
  assign sinkVec_6_1_ready = sinkWire_6_ready & ~maskUnitFirst_6;
  assign sinkVec_6_0_ready = sinkWire_6_ready & maskUnitFirst_6;
  reg          accessDataValid_pipe_v_6;
  reg          accessDataValid_pipe_pipe_v_6;
  wire         accessDataValid_pipe_pipe_out_6_valid = accessDataValid_pipe_pipe_v_6;
  wire         accessDataSource_6_valid = accessDataValid_pipe_pipe_out_6_valid;
  reg          shifterReg_14_0_valid;
  reg  [31:0]  shifterReg_14_0_bits;
  wire         shifterValid_14 = shifterReg_14_0_valid | accessDataSource_6_valid;
  reg          accessDataValid_pipe_v_7;
  reg          accessDataValid_pipe_pipe_v_7;
  wire         accessDataValid_pipe_pipe_out_7_valid = accessDataValid_pipe_pipe_v_7;
  wire         accessDataSource_7_valid = accessDataValid_pipe_pipe_out_7_valid;
  reg          shifterReg_15_0_valid;
  reg  [31:0]  shifterReg_15_0_bits;
  wire         shifterValid_15 = shifterReg_15_0_valid | accessDataSource_7_valid;
  wire         sinkVec_tokenCheck_14;
  wire [4:0]   sinkVec_validSource_14_bits_vd = x22_3_0_bits_vd;
  wire [2:0]   sinkVec_validSource_14_bits_offset = x22_3_0_bits_offset;
  wire [3:0]   sinkVec_validSource_14_bits_mask = x22_3_0_bits_mask;
  wire [31:0]  sinkVec_validSource_14_bits_data = x22_3_0_bits_data;
  wire [2:0]   sinkVec_validSource_14_bits_instructionIndex = x22_3_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_15;
  wire [4:0]   sinkVec_validSource_15_bits_vd = x22_3_1_bits_vd;
  wire [2:0]   sinkVec_validSource_15_bits_offset = x22_3_1_bits_offset;
  wire [3:0]   sinkVec_validSource_15_bits_mask = x22_3_1_bits_mask;
  wire [31:0]  sinkVec_validSource_15_bits_data = x22_3_1_bits_data;
  wire         sinkVec_validSource_15_bits_last = x22_3_1_bits_last;
  wire [2:0]   sinkVec_validSource_15_bits_instructionIndex = x22_3_1_bits_instructionIndex;
  wire         sinkVec_7_0_ready;
  wire         sinkVec_queue_14_deq_ready = sinkVec_sinkWire_14_ready;
  wire         sinkVec_queue_14_deq_valid;
  wire [4:0]   sinkVec_queue_14_deq_bits_vd;
  wire         sinkVec_7_0_valid = sinkVec_sinkWire_14_valid;
  wire [2:0]   sinkVec_queue_14_deq_bits_offset;
  wire [4:0]   sinkVec_7_0_bits_vd = sinkVec_sinkWire_14_bits_vd;
  wire [3:0]   sinkVec_queue_14_deq_bits_mask;
  wire [2:0]   sinkVec_7_0_bits_offset = sinkVec_sinkWire_14_bits_offset;
  wire [31:0]  sinkVec_queue_14_deq_bits_data;
  wire [3:0]   sinkVec_7_0_bits_mask = sinkVec_sinkWire_14_bits_mask;
  wire         sinkVec_queue_14_deq_bits_last;
  wire [31:0]  sinkVec_7_0_bits_data = sinkVec_sinkWire_14_bits_data;
  wire [2:0]   sinkVec_queue_14_deq_bits_instructionIndex;
  wire         sinkVec_7_0_bits_last = sinkVec_sinkWire_14_bits_last;
  wire [2:0]   sinkVec_7_0_bits_instructionIndex = sinkVec_sinkWire_14_bits_instructionIndex;
  wire         sinkVec_validSink_14_valid;
  wire [4:0]   sinkVec_validSink_14_bits_vd;
  wire [2:0]   sinkVec_validSink_14_bits_offset;
  wire [3:0]   sinkVec_validSink_14_bits_mask;
  wire [31:0]  sinkVec_validSink_14_bits_data;
  wire [2:0]   sinkVec_validSink_14_bits_instructionIndex;
  assign sinkVec_sinkWire_14_valid = sinkVec_queue_14_deq_valid;
  assign sinkVec_sinkWire_14_bits_vd = sinkVec_queue_14_deq_bits_vd;
  assign sinkVec_sinkWire_14_bits_offset = sinkVec_queue_14_deq_bits_offset;
  assign sinkVec_sinkWire_14_bits_mask = sinkVec_queue_14_deq_bits_mask;
  assign sinkVec_sinkWire_14_bits_data = sinkVec_queue_14_deq_bits_data;
  assign sinkVec_sinkWire_14_bits_last = sinkVec_queue_14_deq_bits_last;
  assign sinkVec_sinkWire_14_bits_instructionIndex = sinkVec_queue_14_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_14_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_6 = {sinkVec_queue_14_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_14_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_14 = {sinkVec_queue_dataIn_lo_hi_6, sinkVec_queue_14_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_14_enq_bits_vd;
  wire [2:0]   sinkVec_queue_14_enq_bits_offset;
  wire [7:0]   sinkVec_queue_dataIn_hi_hi_6 = {sinkVec_queue_14_enq_bits_vd, sinkVec_queue_14_enq_bits_offset};
  wire [3:0]   sinkVec_queue_14_enq_bits_mask;
  wire [11:0]  sinkVec_queue_dataIn_hi_14 = {sinkVec_queue_dataIn_hi_hi_6, sinkVec_queue_14_enq_bits_mask};
  wire [47:0]  sinkVec_queue_dataIn_14 = {sinkVec_queue_dataIn_hi_14, sinkVec_queue_dataIn_lo_14};
  wire [2:0]   sinkVec_queue_dataOut_14_instructionIndex = _sinkVec_queue_fifo_14_data_out[2:0];
  wire         sinkVec_queue_dataOut_14_last = _sinkVec_queue_fifo_14_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_14_data = _sinkVec_queue_fifo_14_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_14_mask = _sinkVec_queue_fifo_14_data_out[39:36];
  wire [2:0]   sinkVec_queue_dataOut_14_offset = _sinkVec_queue_fifo_14_data_out[42:40];
  wire [4:0]   sinkVec_queue_dataOut_14_vd = _sinkVec_queue_fifo_14_data_out[47:43];
  wire         sinkVec_queue_14_enq_ready = ~_sinkVec_queue_fifo_14_full;
  wire         sinkVec_queue_14_enq_valid;
  assign sinkVec_queue_14_deq_valid = ~_sinkVec_queue_fifo_14_empty | sinkVec_queue_14_enq_valid;
  assign sinkVec_queue_14_deq_bits_vd = _sinkVec_queue_fifo_14_empty ? sinkVec_queue_14_enq_bits_vd : sinkVec_queue_dataOut_14_vd;
  assign sinkVec_queue_14_deq_bits_offset = _sinkVec_queue_fifo_14_empty ? sinkVec_queue_14_enq_bits_offset : sinkVec_queue_dataOut_14_offset;
  assign sinkVec_queue_14_deq_bits_mask = _sinkVec_queue_fifo_14_empty ? sinkVec_queue_14_enq_bits_mask : sinkVec_queue_dataOut_14_mask;
  assign sinkVec_queue_14_deq_bits_data = _sinkVec_queue_fifo_14_empty ? sinkVec_queue_14_enq_bits_data : sinkVec_queue_dataOut_14_data;
  assign sinkVec_queue_14_deq_bits_last = ~_sinkVec_queue_fifo_14_empty & sinkVec_queue_dataOut_14_last;
  assign sinkVec_queue_14_deq_bits_instructionIndex = _sinkVec_queue_fifo_14_empty ? sinkVec_queue_14_enq_bits_instructionIndex : sinkVec_queue_dataOut_14_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_14;
  wire         sinkVec_releasePipe_pipe_out_14_valid = sinkVec_releasePipe_pipe_v_14;
  wire         x22_3_0_ready;
  wire         x22_3_0_valid;
  wire         sinkVec_validSource_14_valid = x22_3_0_ready & x22_3_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_14;
  wire [2:0]   sinkVec_tokenCheck_counterChange_14 = sinkVec_validSource_14_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_14 = ~(sinkVec_tokenCheck_counter_14[2]);
  assign x22_3_0_ready = sinkVec_tokenCheck_14;
  assign sinkVec_queue_14_enq_valid = sinkVec_validSink_14_valid;
  assign sinkVec_queue_14_enq_bits_vd = sinkVec_validSink_14_bits_vd;
  assign sinkVec_queue_14_enq_bits_offset = sinkVec_validSink_14_bits_offset;
  assign sinkVec_queue_14_enq_bits_mask = sinkVec_validSink_14_bits_mask;
  assign sinkVec_queue_14_enq_bits_data = sinkVec_validSink_14_bits_data;
  assign sinkVec_queue_14_enq_bits_instructionIndex = sinkVec_validSink_14_bits_instructionIndex;
  reg          sinkVec_shifterReg_14_0_valid;
  assign sinkVec_validSink_14_valid = sinkVec_shifterReg_14_0_valid;
  reg  [4:0]   sinkVec_shifterReg_14_0_bits_vd;
  assign sinkVec_validSink_14_bits_vd = sinkVec_shifterReg_14_0_bits_vd;
  reg  [2:0]   sinkVec_shifterReg_14_0_bits_offset;
  assign sinkVec_validSink_14_bits_offset = sinkVec_shifterReg_14_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_14_0_bits_mask;
  assign sinkVec_validSink_14_bits_mask = sinkVec_shifterReg_14_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_14_0_bits_data;
  assign sinkVec_validSink_14_bits_data = sinkVec_shifterReg_14_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_14_0_bits_instructionIndex;
  assign sinkVec_validSink_14_bits_instructionIndex = sinkVec_shifterReg_14_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_14 = sinkVec_shifterReg_14_0_valid | sinkVec_validSource_14_valid;
  wire         sinkVec_7_1_ready;
  wire         sinkVec_queue_15_deq_ready = sinkVec_sinkWire_15_ready;
  wire         sinkVec_queue_15_deq_valid;
  wire [4:0]   sinkVec_queue_15_deq_bits_vd;
  wire         sinkVec_7_1_valid = sinkVec_sinkWire_15_valid;
  wire [2:0]   sinkVec_queue_15_deq_bits_offset;
  wire [4:0]   sinkVec_7_1_bits_vd = sinkVec_sinkWire_15_bits_vd;
  wire [3:0]   sinkVec_queue_15_deq_bits_mask;
  wire [2:0]   sinkVec_7_1_bits_offset = sinkVec_sinkWire_15_bits_offset;
  wire [31:0]  sinkVec_queue_15_deq_bits_data;
  wire [3:0]   sinkVec_7_1_bits_mask = sinkVec_sinkWire_15_bits_mask;
  wire         sinkVec_queue_15_deq_bits_last;
  wire [31:0]  sinkVec_7_1_bits_data = sinkVec_sinkWire_15_bits_data;
  wire [2:0]   sinkVec_queue_15_deq_bits_instructionIndex;
  wire         sinkVec_7_1_bits_last = sinkVec_sinkWire_15_bits_last;
  wire [2:0]   sinkVec_7_1_bits_instructionIndex = sinkVec_sinkWire_15_bits_instructionIndex;
  wire         sinkVec_validSink_15_valid;
  wire [4:0]   sinkVec_validSink_15_bits_vd;
  wire [2:0]   sinkVec_validSink_15_bits_offset;
  wire [3:0]   sinkVec_validSink_15_bits_mask;
  wire [31:0]  sinkVec_validSink_15_bits_data;
  wire         sinkVec_validSink_15_bits_last;
  wire [2:0]   sinkVec_validSink_15_bits_instructionIndex;
  assign sinkVec_sinkWire_15_valid = sinkVec_queue_15_deq_valid;
  assign sinkVec_sinkWire_15_bits_vd = sinkVec_queue_15_deq_bits_vd;
  assign sinkVec_sinkWire_15_bits_offset = sinkVec_queue_15_deq_bits_offset;
  assign sinkVec_sinkWire_15_bits_mask = sinkVec_queue_15_deq_bits_mask;
  assign sinkVec_sinkWire_15_bits_data = sinkVec_queue_15_deq_bits_data;
  assign sinkVec_sinkWire_15_bits_last = sinkVec_queue_15_deq_bits_last;
  assign sinkVec_sinkWire_15_bits_instructionIndex = sinkVec_queue_15_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_15_enq_bits_data;
  wire         sinkVec_queue_15_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_7 = {sinkVec_queue_15_enq_bits_data, sinkVec_queue_15_enq_bits_last};
  wire [2:0]   sinkVec_queue_15_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_15 = {sinkVec_queue_dataIn_lo_hi_7, sinkVec_queue_15_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_15_enq_bits_vd;
  wire [2:0]   sinkVec_queue_15_enq_bits_offset;
  wire [7:0]   sinkVec_queue_dataIn_hi_hi_7 = {sinkVec_queue_15_enq_bits_vd, sinkVec_queue_15_enq_bits_offset};
  wire [3:0]   sinkVec_queue_15_enq_bits_mask;
  wire [11:0]  sinkVec_queue_dataIn_hi_15 = {sinkVec_queue_dataIn_hi_hi_7, sinkVec_queue_15_enq_bits_mask};
  wire [47:0]  sinkVec_queue_dataIn_15 = {sinkVec_queue_dataIn_hi_15, sinkVec_queue_dataIn_lo_15};
  wire [2:0]   sinkVec_queue_dataOut_15_instructionIndex = _sinkVec_queue_fifo_15_data_out[2:0];
  wire         sinkVec_queue_dataOut_15_last = _sinkVec_queue_fifo_15_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_15_data = _sinkVec_queue_fifo_15_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_15_mask = _sinkVec_queue_fifo_15_data_out[39:36];
  wire [2:0]   sinkVec_queue_dataOut_15_offset = _sinkVec_queue_fifo_15_data_out[42:40];
  wire [4:0]   sinkVec_queue_dataOut_15_vd = _sinkVec_queue_fifo_15_data_out[47:43];
  wire         sinkVec_queue_15_enq_ready = ~_sinkVec_queue_fifo_15_full;
  wire         sinkVec_queue_15_enq_valid;
  assign sinkVec_queue_15_deq_valid = ~_sinkVec_queue_fifo_15_empty | sinkVec_queue_15_enq_valid;
  assign sinkVec_queue_15_deq_bits_vd = _sinkVec_queue_fifo_15_empty ? sinkVec_queue_15_enq_bits_vd : sinkVec_queue_dataOut_15_vd;
  assign sinkVec_queue_15_deq_bits_offset = _sinkVec_queue_fifo_15_empty ? sinkVec_queue_15_enq_bits_offset : sinkVec_queue_dataOut_15_offset;
  assign sinkVec_queue_15_deq_bits_mask = _sinkVec_queue_fifo_15_empty ? sinkVec_queue_15_enq_bits_mask : sinkVec_queue_dataOut_15_mask;
  assign sinkVec_queue_15_deq_bits_data = _sinkVec_queue_fifo_15_empty ? sinkVec_queue_15_enq_bits_data : sinkVec_queue_dataOut_15_data;
  assign sinkVec_queue_15_deq_bits_last = _sinkVec_queue_fifo_15_empty ? sinkVec_queue_15_enq_bits_last : sinkVec_queue_dataOut_15_last;
  assign sinkVec_queue_15_deq_bits_instructionIndex = _sinkVec_queue_fifo_15_empty ? sinkVec_queue_15_enq_bits_instructionIndex : sinkVec_queue_dataOut_15_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_15;
  wire         sinkVec_releasePipe_pipe_out_15_valid = sinkVec_releasePipe_pipe_v_15;
  wire         x22_3_1_ready;
  wire         x22_3_1_valid;
  wire         sinkVec_validSource_15_valid = x22_3_1_ready & x22_3_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_15;
  wire [2:0]   sinkVec_tokenCheck_counterChange_15 = sinkVec_validSource_15_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_15 = ~(sinkVec_tokenCheck_counter_15[2]);
  assign x22_3_1_ready = sinkVec_tokenCheck_15;
  assign sinkVec_queue_15_enq_valid = sinkVec_validSink_15_valid;
  assign sinkVec_queue_15_enq_bits_vd = sinkVec_validSink_15_bits_vd;
  assign sinkVec_queue_15_enq_bits_offset = sinkVec_validSink_15_bits_offset;
  assign sinkVec_queue_15_enq_bits_mask = sinkVec_validSink_15_bits_mask;
  assign sinkVec_queue_15_enq_bits_data = sinkVec_validSink_15_bits_data;
  assign sinkVec_queue_15_enq_bits_last = sinkVec_validSink_15_bits_last;
  assign sinkVec_queue_15_enq_bits_instructionIndex = sinkVec_validSink_15_bits_instructionIndex;
  reg          sinkVec_shifterReg_15_0_valid;
  assign sinkVec_validSink_15_valid = sinkVec_shifterReg_15_0_valid;
  reg  [4:0]   sinkVec_shifterReg_15_0_bits_vd;
  assign sinkVec_validSink_15_bits_vd = sinkVec_shifterReg_15_0_bits_vd;
  reg  [2:0]   sinkVec_shifterReg_15_0_bits_offset;
  assign sinkVec_validSink_15_bits_offset = sinkVec_shifterReg_15_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_15_0_bits_mask;
  assign sinkVec_validSink_15_bits_mask = sinkVec_shifterReg_15_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_15_0_bits_data;
  assign sinkVec_validSink_15_bits_data = sinkVec_shifterReg_15_0_bits_data;
  reg          sinkVec_shifterReg_15_0_bits_last;
  assign sinkVec_validSink_15_bits_last = sinkVec_shifterReg_15_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_15_0_bits_instructionIndex;
  assign sinkVec_validSink_15_bits_instructionIndex = sinkVec_shifterReg_15_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_15 = sinkVec_shifterReg_15_0_valid | sinkVec_validSource_15_valid;
  assign sinkVec_sinkWire_14_ready = sinkVec_7_0_ready;
  assign sinkVec_sinkWire_15_ready = sinkVec_7_1_ready;
  reg          maskUnitFirst_7;
  wire         tryToRead_7 = sinkVec_7_0_valid | sinkVec_7_1_valid;
  wire         sinkWire_7_valid = maskUnitFirst_7 ? sinkVec_7_0_valid : sinkVec_7_1_valid;
  wire [4:0]   sinkWire_7_bits_vd = maskUnitFirst_7 ? sinkVec_7_0_bits_vd : sinkVec_7_1_bits_vd;
  wire [2:0]   sinkWire_7_bits_offset = maskUnitFirst_7 ? sinkVec_7_0_bits_offset : sinkVec_7_1_bits_offset;
  wire [3:0]   sinkWire_7_bits_mask = maskUnitFirst_7 ? sinkVec_7_0_bits_mask : sinkVec_7_1_bits_mask;
  wire [31:0]  sinkWire_7_bits_data = maskUnitFirst_7 ? sinkVec_7_0_bits_data : sinkVec_7_1_bits_data;
  wire         sinkWire_7_bits_last = maskUnitFirst_7 ? sinkVec_7_0_bits_last : sinkVec_7_1_bits_last;
  wire [2:0]   sinkWire_7_bits_instructionIndex = maskUnitFirst_7 ? sinkVec_7_0_bits_instructionIndex : sinkVec_7_1_bits_instructionIndex;
  wire         sinkWire_7_ready;
  assign sinkVec_7_1_ready = sinkWire_7_ready & ~maskUnitFirst_7;
  assign sinkVec_7_0_ready = sinkWire_7_ready & maskUnitFirst_7;
  reg          view__writeRelease_3_pipe_v;
  wire         view__writeRelease_3_pipe_out_valid = view__writeRelease_3_pipe_v;
  reg          pipe_v_9;
  wire         pipe_out_6_valid = pipe_v_9;
  wire         _probeWire_writeQueueEnqVec_3_valid_T = x22_3_0_ready & _maskUnit_exeResp_3_valid;
  reg          instructionFinishedPipe_pipe_v_3;
  wire         instructionFinishedPipe_pipe_out_3_valid = instructionFinishedPipe_pipe_v_3;
  reg  [7:0]   instructionFinishedPipe_pipe_b_3;
  wire [7:0]   instructionFinishedPipe_pipe_out_3_bits = instructionFinishedPipe_pipe_b_3;
  wire         instructionFinished_3_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_3_bits);
  wire         instructionFinished_3_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_3_bits);
  wire         instructionFinished_3_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_3_bits);
  wire         instructionFinished_3_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_3_bits);
  assign vxsatReportVec_3 = _laneVec_3_vxsatReport[3:0];
  reg          pipe_v_10;
  reg  [31:0]  pipe_b_10;
  reg          pipe_pipe_v_3;
  wire         pipe_pipe_out_3_valid = pipe_pipe_v_3;
  reg  [31:0]  pipe_pipe_b_3;
  wire [31:0]  pipe_pipe_out_3_bits = pipe_pipe_b_3;
  reg          view__laneMaskSelect_3_pipe_v;
  reg  [5:0]   view__laneMaskSelect_3_pipe_b;
  reg          view__laneMaskSelect_3_pipe_pipe_v;
  wire         view__laneMaskSelect_3_pipe_pipe_out_valid = view__laneMaskSelect_3_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_3_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_3_pipe_pipe_out_bits = view__laneMaskSelect_3_pipe_pipe_b;
  reg          view__laneMaskSewSelect_3_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_3_pipe_b;
  reg          view__laneMaskSewSelect_3_pipe_pipe_v;
  wire         view__laneMaskSewSelect_3_pipe_pipe_out_valid = view__laneMaskSewSelect_3_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_3_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_3_pipe_pipe_out_bits = view__laneMaskSewSelect_3_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v_3;
  wire         lsuLastPipe_pipe_out_3_valid = lsuLastPipe_pipe_v_3;
  reg  [7:0]   lsuLastPipe_pipe_b_3;
  wire [7:0]   lsuLastPipe_pipe_out_3_bits = lsuLastPipe_pipe_b_3;
  reg          maskLastPipe_pipe_v_3;
  wire         maskLastPipe_pipe_out_3_valid = maskLastPipe_pipe_v_3;
  reg  [7:0]   maskLastPipe_pipe_b_3;
  wire [7:0]   maskLastPipe_pipe_out_3_bits = maskLastPipe_pipe_b_3;
  wire [6:0]   writeCounter_3 = requestReg_bits_writeByte[11:5] + {6'h0, requestReg_bits_writeByte[4:0] > 5'hC};
  reg          pipe_v_11;
  wire         pipe_out_7_valid = pipe_v_11;
  reg  [6:0]   pipe_b_11;
  wire [6:0]   pipe_out_7_bits = pipe_b_11;
  assign laneRequestSinkWire_4_ready = ~laneRequestSinkWire_4_bits_issueInst | _laneVec_4_laneRequest_ready;
  wire         sinkVec_tokenCheck_16;
  wire [4:0]   sinkVec_validSource_16_bits_vs = x13_4_0_bits_vs;
  wire [2:0]   sinkVec_validSource_16_bits_offset = x13_4_0_bits_offset;
  wire [2:0]   sinkVec_validSource_16_bits_instructionIndex = x13_4_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_17;
  wire [4:0]   sinkVec_validSource_17_bits_vs = x13_4_1_bits_vs;
  wire [2:0]   sinkVec_validSource_17_bits_offset = x13_4_1_bits_offset;
  wire [2:0]   sinkVec_validSource_17_bits_instructionIndex = x13_4_1_bits_instructionIndex;
  wire         sinkVec_8_0_ready;
  wire         sinkVec_queue_16_deq_ready = sinkVec_sinkWire_16_ready;
  wire         sinkVec_queue_16_deq_valid;
  wire [4:0]   sinkVec_queue_16_deq_bits_vs;
  wire         sinkVec_8_0_valid = sinkVec_sinkWire_16_valid;
  wire [1:0]   sinkVec_queue_16_deq_bits_readSource;
  wire [4:0]   sinkVec_8_0_bits_vs = sinkVec_sinkWire_16_bits_vs;
  wire [2:0]   sinkVec_queue_16_deq_bits_offset;
  wire [1:0]   sinkVec_8_0_bits_readSource = sinkVec_sinkWire_16_bits_readSource;
  wire [2:0]   sinkVec_queue_16_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_8_0_bits_offset = sinkVec_sinkWire_16_bits_offset;
  wire [2:0]   sinkVec_8_0_bits_instructionIndex = sinkVec_sinkWire_16_bits_instructionIndex;
  wire         sinkVec_validSink_16_valid;
  wire [4:0]   sinkVec_validSink_16_bits_vs;
  wire [1:0]   sinkVec_validSink_16_bits_readSource;
  wire [2:0]   sinkVec_validSink_16_bits_offset;
  wire [2:0]   sinkVec_validSink_16_bits_instructionIndex;
  assign sinkVec_sinkWire_16_valid = sinkVec_queue_16_deq_valid;
  assign sinkVec_sinkWire_16_bits_vs = sinkVec_queue_16_deq_bits_vs;
  assign sinkVec_sinkWire_16_bits_readSource = sinkVec_queue_16_deq_bits_readSource;
  assign sinkVec_sinkWire_16_bits_offset = sinkVec_queue_16_deq_bits_offset;
  assign sinkVec_sinkWire_16_bits_instructionIndex = sinkVec_queue_16_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_queue_16_enq_bits_offset;
  wire [2:0]   sinkVec_queue_16_enq_bits_instructionIndex;
  wire [5:0]   sinkVec_queue_dataIn_lo_16 = {sinkVec_queue_16_enq_bits_offset, sinkVec_queue_16_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_16_enq_bits_vs;
  wire [1:0]   sinkVec_queue_16_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_16 = {sinkVec_queue_16_enq_bits_vs, sinkVec_queue_16_enq_bits_readSource};
  wire [12:0]  sinkVec_queue_dataIn_16 = {sinkVec_queue_dataIn_hi_16, sinkVec_queue_dataIn_lo_16};
  wire [2:0]   sinkVec_queue_dataOut_16_instructionIndex = _sinkVec_queue_fifo_16_data_out[2:0];
  wire [2:0]   sinkVec_queue_dataOut_16_offset = _sinkVec_queue_fifo_16_data_out[5:3];
  wire [1:0]   sinkVec_queue_dataOut_16_readSource = _sinkVec_queue_fifo_16_data_out[7:6];
  wire [4:0]   sinkVec_queue_dataOut_16_vs = _sinkVec_queue_fifo_16_data_out[12:8];
  wire         sinkVec_queue_16_enq_ready = ~_sinkVec_queue_fifo_16_full;
  wire         sinkVec_queue_16_enq_valid;
  assign sinkVec_queue_16_deq_valid = ~_sinkVec_queue_fifo_16_empty | sinkVec_queue_16_enq_valid;
  assign sinkVec_queue_16_deq_bits_vs = _sinkVec_queue_fifo_16_empty ? sinkVec_queue_16_enq_bits_vs : sinkVec_queue_dataOut_16_vs;
  assign sinkVec_queue_16_deq_bits_readSource = _sinkVec_queue_fifo_16_empty ? sinkVec_queue_16_enq_bits_readSource : sinkVec_queue_dataOut_16_readSource;
  assign sinkVec_queue_16_deq_bits_offset = _sinkVec_queue_fifo_16_empty ? sinkVec_queue_16_enq_bits_offset : sinkVec_queue_dataOut_16_offset;
  assign sinkVec_queue_16_deq_bits_instructionIndex = _sinkVec_queue_fifo_16_empty ? sinkVec_queue_16_enq_bits_instructionIndex : sinkVec_queue_dataOut_16_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_16;
  wire         sinkVec_releasePipe_pipe_out_16_valid = sinkVec_releasePipe_pipe_v_16;
  wire         x13_4_0_ready;
  wire         x13_4_0_valid;
  wire         sinkVec_validSource_16_valid = x13_4_0_ready & x13_4_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_16;
  wire [2:0]   sinkVec_tokenCheck_counterChange_16 = sinkVec_validSource_16_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_16 = ~(sinkVec_tokenCheck_counter_16[2]);
  assign x13_4_0_ready = sinkVec_tokenCheck_16;
  assign sinkVec_queue_16_enq_valid = sinkVec_validSink_16_valid;
  assign sinkVec_queue_16_enq_bits_vs = sinkVec_validSink_16_bits_vs;
  assign sinkVec_queue_16_enq_bits_readSource = sinkVec_validSink_16_bits_readSource;
  assign sinkVec_queue_16_enq_bits_offset = sinkVec_validSink_16_bits_offset;
  assign sinkVec_queue_16_enq_bits_instructionIndex = sinkVec_validSink_16_bits_instructionIndex;
  reg          sinkVec_shifterReg_16_0_valid;
  assign sinkVec_validSink_16_valid = sinkVec_shifterReg_16_0_valid;
  reg  [4:0]   sinkVec_shifterReg_16_0_bits_vs;
  assign sinkVec_validSink_16_bits_vs = sinkVec_shifterReg_16_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_16_0_bits_readSource;
  assign sinkVec_validSink_16_bits_readSource = sinkVec_shifterReg_16_0_bits_readSource;
  reg  [2:0]   sinkVec_shifterReg_16_0_bits_offset;
  assign sinkVec_validSink_16_bits_offset = sinkVec_shifterReg_16_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_16_0_bits_instructionIndex;
  assign sinkVec_validSink_16_bits_instructionIndex = sinkVec_shifterReg_16_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_16 = sinkVec_shifterReg_16_0_valid | sinkVec_validSource_16_valid;
  wire         sinkVec_8_1_ready;
  wire         sinkVec_queue_17_deq_ready = sinkVec_sinkWire_17_ready;
  wire         sinkVec_queue_17_deq_valid;
  wire [4:0]   sinkVec_queue_17_deq_bits_vs;
  wire         sinkVec_8_1_valid = sinkVec_sinkWire_17_valid;
  wire [1:0]   sinkVec_queue_17_deq_bits_readSource;
  wire [4:0]   sinkVec_8_1_bits_vs = sinkVec_sinkWire_17_bits_vs;
  wire [2:0]   sinkVec_queue_17_deq_bits_offset;
  wire [1:0]   sinkVec_8_1_bits_readSource = sinkVec_sinkWire_17_bits_readSource;
  wire [2:0]   sinkVec_queue_17_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_8_1_bits_offset = sinkVec_sinkWire_17_bits_offset;
  wire [2:0]   sinkVec_8_1_bits_instructionIndex = sinkVec_sinkWire_17_bits_instructionIndex;
  wire         sinkVec_validSink_17_valid;
  wire [4:0]   sinkVec_validSink_17_bits_vs;
  wire [1:0]   sinkVec_validSink_17_bits_readSource;
  wire [2:0]   sinkVec_validSink_17_bits_offset;
  wire [2:0]   sinkVec_validSink_17_bits_instructionIndex;
  assign sinkVec_sinkWire_17_valid = sinkVec_queue_17_deq_valid;
  assign sinkVec_sinkWire_17_bits_vs = sinkVec_queue_17_deq_bits_vs;
  assign sinkVec_sinkWire_17_bits_readSource = sinkVec_queue_17_deq_bits_readSource;
  assign sinkVec_sinkWire_17_bits_offset = sinkVec_queue_17_deq_bits_offset;
  assign sinkVec_sinkWire_17_bits_instructionIndex = sinkVec_queue_17_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_queue_17_enq_bits_offset;
  wire [2:0]   sinkVec_queue_17_enq_bits_instructionIndex;
  wire [5:0]   sinkVec_queue_dataIn_lo_17 = {sinkVec_queue_17_enq_bits_offset, sinkVec_queue_17_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_17_enq_bits_vs;
  wire [1:0]   sinkVec_queue_17_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_17 = {sinkVec_queue_17_enq_bits_vs, sinkVec_queue_17_enq_bits_readSource};
  wire [12:0]  sinkVec_queue_dataIn_17 = {sinkVec_queue_dataIn_hi_17, sinkVec_queue_dataIn_lo_17};
  wire [2:0]   sinkVec_queue_dataOut_17_instructionIndex = _sinkVec_queue_fifo_17_data_out[2:0];
  wire [2:0]   sinkVec_queue_dataOut_17_offset = _sinkVec_queue_fifo_17_data_out[5:3];
  wire [1:0]   sinkVec_queue_dataOut_17_readSource = _sinkVec_queue_fifo_17_data_out[7:6];
  wire [4:0]   sinkVec_queue_dataOut_17_vs = _sinkVec_queue_fifo_17_data_out[12:8];
  wire         sinkVec_queue_17_enq_ready = ~_sinkVec_queue_fifo_17_full;
  wire         sinkVec_queue_17_enq_valid;
  assign sinkVec_queue_17_deq_valid = ~_sinkVec_queue_fifo_17_empty | sinkVec_queue_17_enq_valid;
  assign sinkVec_queue_17_deq_bits_vs = _sinkVec_queue_fifo_17_empty ? sinkVec_queue_17_enq_bits_vs : sinkVec_queue_dataOut_17_vs;
  assign sinkVec_queue_17_deq_bits_readSource = _sinkVec_queue_fifo_17_empty ? sinkVec_queue_17_enq_bits_readSource : sinkVec_queue_dataOut_17_readSource;
  assign sinkVec_queue_17_deq_bits_offset = _sinkVec_queue_fifo_17_empty ? sinkVec_queue_17_enq_bits_offset : sinkVec_queue_dataOut_17_offset;
  assign sinkVec_queue_17_deq_bits_instructionIndex = _sinkVec_queue_fifo_17_empty ? sinkVec_queue_17_enq_bits_instructionIndex : sinkVec_queue_dataOut_17_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_17;
  wire         sinkVec_releasePipe_pipe_out_17_valid = sinkVec_releasePipe_pipe_v_17;
  wire         x13_4_1_ready;
  wire         x13_4_1_valid;
  wire         sinkVec_validSource_17_valid = x13_4_1_ready & x13_4_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_17;
  wire [2:0]   sinkVec_tokenCheck_counterChange_17 = sinkVec_validSource_17_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_17 = ~(sinkVec_tokenCheck_counter_17[2]);
  assign x13_4_1_ready = sinkVec_tokenCheck_17;
  assign sinkVec_queue_17_enq_valid = sinkVec_validSink_17_valid;
  assign sinkVec_queue_17_enq_bits_vs = sinkVec_validSink_17_bits_vs;
  assign sinkVec_queue_17_enq_bits_readSource = sinkVec_validSink_17_bits_readSource;
  assign sinkVec_queue_17_enq_bits_offset = sinkVec_validSink_17_bits_offset;
  assign sinkVec_queue_17_enq_bits_instructionIndex = sinkVec_validSink_17_bits_instructionIndex;
  reg          sinkVec_shifterReg_17_0_valid;
  assign sinkVec_validSink_17_valid = sinkVec_shifterReg_17_0_valid;
  reg  [4:0]   sinkVec_shifterReg_17_0_bits_vs;
  assign sinkVec_validSink_17_bits_vs = sinkVec_shifterReg_17_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_17_0_bits_readSource;
  assign sinkVec_validSink_17_bits_readSource = sinkVec_shifterReg_17_0_bits_readSource;
  reg  [2:0]   sinkVec_shifterReg_17_0_bits_offset;
  assign sinkVec_validSink_17_bits_offset = sinkVec_shifterReg_17_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_17_0_bits_instructionIndex;
  assign sinkVec_validSink_17_bits_instructionIndex = sinkVec_shifterReg_17_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_17 = sinkVec_shifterReg_17_0_valid | sinkVec_validSource_17_valid;
  assign sinkVec_sinkWire_16_ready = sinkVec_8_0_ready;
  assign sinkVec_sinkWire_17_ready = sinkVec_8_1_ready;
  reg          maskUnitFirst_8;
  wire         tryToRead_8 = sinkVec_8_0_valid | sinkVec_8_1_valid;
  wire         sinkWire_8_valid = maskUnitFirst_8 ? sinkVec_8_0_valid : sinkVec_8_1_valid;
  wire [4:0]   sinkWire_8_bits_vs = maskUnitFirst_8 ? sinkVec_8_0_bits_vs : sinkVec_8_1_bits_vs;
  wire [1:0]   sinkWire_8_bits_readSource = maskUnitFirst_8 ? sinkVec_8_0_bits_readSource : sinkVec_8_1_bits_readSource;
  wire [2:0]   sinkWire_8_bits_offset = maskUnitFirst_8 ? sinkVec_8_0_bits_offset : sinkVec_8_1_bits_offset;
  wire [2:0]   sinkWire_8_bits_instructionIndex = maskUnitFirst_8 ? sinkVec_8_0_bits_instructionIndex : sinkVec_8_1_bits_instructionIndex;
  wire         sinkWire_8_ready;
  assign sinkVec_8_1_ready = sinkWire_8_ready & ~maskUnitFirst_8;
  assign sinkVec_8_0_ready = sinkWire_8_ready & maskUnitFirst_8;
  reg          accessDataValid_pipe_v_8;
  reg          accessDataValid_pipe_pipe_v_8;
  wire         accessDataValid_pipe_pipe_out_8_valid = accessDataValid_pipe_pipe_v_8;
  wire         accessDataSource_8_valid = accessDataValid_pipe_pipe_out_8_valid;
  reg          shifterReg_16_0_valid;
  reg  [31:0]  shifterReg_16_0_bits;
  wire         shifterValid_16 = shifterReg_16_0_valid | accessDataSource_8_valid;
  reg          accessDataValid_pipe_v_9;
  reg          accessDataValid_pipe_pipe_v_9;
  wire         accessDataValid_pipe_pipe_out_9_valid = accessDataValid_pipe_pipe_v_9;
  wire         accessDataSource_9_valid = accessDataValid_pipe_pipe_out_9_valid;
  reg          shifterReg_17_0_valid;
  reg  [31:0]  shifterReg_17_0_bits;
  wire         shifterValid_17 = shifterReg_17_0_valid | accessDataSource_9_valid;
  wire         sinkVec_tokenCheck_18;
  wire [4:0]   sinkVec_validSource_18_bits_vd = x22_4_0_bits_vd;
  wire [2:0]   sinkVec_validSource_18_bits_offset = x22_4_0_bits_offset;
  wire [3:0]   sinkVec_validSource_18_bits_mask = x22_4_0_bits_mask;
  wire [31:0]  sinkVec_validSource_18_bits_data = x22_4_0_bits_data;
  wire [2:0]   sinkVec_validSource_18_bits_instructionIndex = x22_4_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_19;
  wire [4:0]   sinkVec_validSource_19_bits_vd = x22_4_1_bits_vd;
  wire [2:0]   sinkVec_validSource_19_bits_offset = x22_4_1_bits_offset;
  wire [3:0]   sinkVec_validSource_19_bits_mask = x22_4_1_bits_mask;
  wire [31:0]  sinkVec_validSource_19_bits_data = x22_4_1_bits_data;
  wire         sinkVec_validSource_19_bits_last = x22_4_1_bits_last;
  wire [2:0]   sinkVec_validSource_19_bits_instructionIndex = x22_4_1_bits_instructionIndex;
  wire         sinkVec_9_0_ready;
  wire         sinkVec_queue_18_deq_ready = sinkVec_sinkWire_18_ready;
  wire         sinkVec_queue_18_deq_valid;
  wire [4:0]   sinkVec_queue_18_deq_bits_vd;
  wire         sinkVec_9_0_valid = sinkVec_sinkWire_18_valid;
  wire [2:0]   sinkVec_queue_18_deq_bits_offset;
  wire [4:0]   sinkVec_9_0_bits_vd = sinkVec_sinkWire_18_bits_vd;
  wire [3:0]   sinkVec_queue_18_deq_bits_mask;
  wire [2:0]   sinkVec_9_0_bits_offset = sinkVec_sinkWire_18_bits_offset;
  wire [31:0]  sinkVec_queue_18_deq_bits_data;
  wire [3:0]   sinkVec_9_0_bits_mask = sinkVec_sinkWire_18_bits_mask;
  wire         sinkVec_queue_18_deq_bits_last;
  wire [31:0]  sinkVec_9_0_bits_data = sinkVec_sinkWire_18_bits_data;
  wire [2:0]   sinkVec_queue_18_deq_bits_instructionIndex;
  wire         sinkVec_9_0_bits_last = sinkVec_sinkWire_18_bits_last;
  wire [2:0]   sinkVec_9_0_bits_instructionIndex = sinkVec_sinkWire_18_bits_instructionIndex;
  wire         sinkVec_validSink_18_valid;
  wire [4:0]   sinkVec_validSink_18_bits_vd;
  wire [2:0]   sinkVec_validSink_18_bits_offset;
  wire [3:0]   sinkVec_validSink_18_bits_mask;
  wire [31:0]  sinkVec_validSink_18_bits_data;
  wire [2:0]   sinkVec_validSink_18_bits_instructionIndex;
  assign sinkVec_sinkWire_18_valid = sinkVec_queue_18_deq_valid;
  assign sinkVec_sinkWire_18_bits_vd = sinkVec_queue_18_deq_bits_vd;
  assign sinkVec_sinkWire_18_bits_offset = sinkVec_queue_18_deq_bits_offset;
  assign sinkVec_sinkWire_18_bits_mask = sinkVec_queue_18_deq_bits_mask;
  assign sinkVec_sinkWire_18_bits_data = sinkVec_queue_18_deq_bits_data;
  assign sinkVec_sinkWire_18_bits_last = sinkVec_queue_18_deq_bits_last;
  assign sinkVec_sinkWire_18_bits_instructionIndex = sinkVec_queue_18_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_18_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_8 = {sinkVec_queue_18_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_18_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_18 = {sinkVec_queue_dataIn_lo_hi_8, sinkVec_queue_18_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_18_enq_bits_vd;
  wire [2:0]   sinkVec_queue_18_enq_bits_offset;
  wire [7:0]   sinkVec_queue_dataIn_hi_hi_8 = {sinkVec_queue_18_enq_bits_vd, sinkVec_queue_18_enq_bits_offset};
  wire [3:0]   sinkVec_queue_18_enq_bits_mask;
  wire [11:0]  sinkVec_queue_dataIn_hi_18 = {sinkVec_queue_dataIn_hi_hi_8, sinkVec_queue_18_enq_bits_mask};
  wire [47:0]  sinkVec_queue_dataIn_18 = {sinkVec_queue_dataIn_hi_18, sinkVec_queue_dataIn_lo_18};
  wire [2:0]   sinkVec_queue_dataOut_18_instructionIndex = _sinkVec_queue_fifo_18_data_out[2:0];
  wire         sinkVec_queue_dataOut_18_last = _sinkVec_queue_fifo_18_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_18_data = _sinkVec_queue_fifo_18_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_18_mask = _sinkVec_queue_fifo_18_data_out[39:36];
  wire [2:0]   sinkVec_queue_dataOut_18_offset = _sinkVec_queue_fifo_18_data_out[42:40];
  wire [4:0]   sinkVec_queue_dataOut_18_vd = _sinkVec_queue_fifo_18_data_out[47:43];
  wire         sinkVec_queue_18_enq_ready = ~_sinkVec_queue_fifo_18_full;
  wire         sinkVec_queue_18_enq_valid;
  assign sinkVec_queue_18_deq_valid = ~_sinkVec_queue_fifo_18_empty | sinkVec_queue_18_enq_valid;
  assign sinkVec_queue_18_deq_bits_vd = _sinkVec_queue_fifo_18_empty ? sinkVec_queue_18_enq_bits_vd : sinkVec_queue_dataOut_18_vd;
  assign sinkVec_queue_18_deq_bits_offset = _sinkVec_queue_fifo_18_empty ? sinkVec_queue_18_enq_bits_offset : sinkVec_queue_dataOut_18_offset;
  assign sinkVec_queue_18_deq_bits_mask = _sinkVec_queue_fifo_18_empty ? sinkVec_queue_18_enq_bits_mask : sinkVec_queue_dataOut_18_mask;
  assign sinkVec_queue_18_deq_bits_data = _sinkVec_queue_fifo_18_empty ? sinkVec_queue_18_enq_bits_data : sinkVec_queue_dataOut_18_data;
  assign sinkVec_queue_18_deq_bits_last = ~_sinkVec_queue_fifo_18_empty & sinkVec_queue_dataOut_18_last;
  assign sinkVec_queue_18_deq_bits_instructionIndex = _sinkVec_queue_fifo_18_empty ? sinkVec_queue_18_enq_bits_instructionIndex : sinkVec_queue_dataOut_18_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_18;
  wire         sinkVec_releasePipe_pipe_out_18_valid = sinkVec_releasePipe_pipe_v_18;
  wire         x22_4_0_ready;
  wire         x22_4_0_valid;
  wire         sinkVec_validSource_18_valid = x22_4_0_ready & x22_4_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_18;
  wire [2:0]   sinkVec_tokenCheck_counterChange_18 = sinkVec_validSource_18_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_18 = ~(sinkVec_tokenCheck_counter_18[2]);
  assign x22_4_0_ready = sinkVec_tokenCheck_18;
  assign sinkVec_queue_18_enq_valid = sinkVec_validSink_18_valid;
  assign sinkVec_queue_18_enq_bits_vd = sinkVec_validSink_18_bits_vd;
  assign sinkVec_queue_18_enq_bits_offset = sinkVec_validSink_18_bits_offset;
  assign sinkVec_queue_18_enq_bits_mask = sinkVec_validSink_18_bits_mask;
  assign sinkVec_queue_18_enq_bits_data = sinkVec_validSink_18_bits_data;
  assign sinkVec_queue_18_enq_bits_instructionIndex = sinkVec_validSink_18_bits_instructionIndex;
  reg          sinkVec_shifterReg_18_0_valid;
  assign sinkVec_validSink_18_valid = sinkVec_shifterReg_18_0_valid;
  reg  [4:0]   sinkVec_shifterReg_18_0_bits_vd;
  assign sinkVec_validSink_18_bits_vd = sinkVec_shifterReg_18_0_bits_vd;
  reg  [2:0]   sinkVec_shifterReg_18_0_bits_offset;
  assign sinkVec_validSink_18_bits_offset = sinkVec_shifterReg_18_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_18_0_bits_mask;
  assign sinkVec_validSink_18_bits_mask = sinkVec_shifterReg_18_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_18_0_bits_data;
  assign sinkVec_validSink_18_bits_data = sinkVec_shifterReg_18_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_18_0_bits_instructionIndex;
  assign sinkVec_validSink_18_bits_instructionIndex = sinkVec_shifterReg_18_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_18 = sinkVec_shifterReg_18_0_valid | sinkVec_validSource_18_valid;
  wire         sinkVec_9_1_ready;
  wire         sinkVec_queue_19_deq_ready = sinkVec_sinkWire_19_ready;
  wire         sinkVec_queue_19_deq_valid;
  wire [4:0]   sinkVec_queue_19_deq_bits_vd;
  wire         sinkVec_9_1_valid = sinkVec_sinkWire_19_valid;
  wire [2:0]   sinkVec_queue_19_deq_bits_offset;
  wire [4:0]   sinkVec_9_1_bits_vd = sinkVec_sinkWire_19_bits_vd;
  wire [3:0]   sinkVec_queue_19_deq_bits_mask;
  wire [2:0]   sinkVec_9_1_bits_offset = sinkVec_sinkWire_19_bits_offset;
  wire [31:0]  sinkVec_queue_19_deq_bits_data;
  wire [3:0]   sinkVec_9_1_bits_mask = sinkVec_sinkWire_19_bits_mask;
  wire         sinkVec_queue_19_deq_bits_last;
  wire [31:0]  sinkVec_9_1_bits_data = sinkVec_sinkWire_19_bits_data;
  wire [2:0]   sinkVec_queue_19_deq_bits_instructionIndex;
  wire         sinkVec_9_1_bits_last = sinkVec_sinkWire_19_bits_last;
  wire [2:0]   sinkVec_9_1_bits_instructionIndex = sinkVec_sinkWire_19_bits_instructionIndex;
  wire         sinkVec_validSink_19_valid;
  wire [4:0]   sinkVec_validSink_19_bits_vd;
  wire [2:0]   sinkVec_validSink_19_bits_offset;
  wire [3:0]   sinkVec_validSink_19_bits_mask;
  wire [31:0]  sinkVec_validSink_19_bits_data;
  wire         sinkVec_validSink_19_bits_last;
  wire [2:0]   sinkVec_validSink_19_bits_instructionIndex;
  assign sinkVec_sinkWire_19_valid = sinkVec_queue_19_deq_valid;
  assign sinkVec_sinkWire_19_bits_vd = sinkVec_queue_19_deq_bits_vd;
  assign sinkVec_sinkWire_19_bits_offset = sinkVec_queue_19_deq_bits_offset;
  assign sinkVec_sinkWire_19_bits_mask = sinkVec_queue_19_deq_bits_mask;
  assign sinkVec_sinkWire_19_bits_data = sinkVec_queue_19_deq_bits_data;
  assign sinkVec_sinkWire_19_bits_last = sinkVec_queue_19_deq_bits_last;
  assign sinkVec_sinkWire_19_bits_instructionIndex = sinkVec_queue_19_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_19_enq_bits_data;
  wire         sinkVec_queue_19_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_9 = {sinkVec_queue_19_enq_bits_data, sinkVec_queue_19_enq_bits_last};
  wire [2:0]   sinkVec_queue_19_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_19 = {sinkVec_queue_dataIn_lo_hi_9, sinkVec_queue_19_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_19_enq_bits_vd;
  wire [2:0]   sinkVec_queue_19_enq_bits_offset;
  wire [7:0]   sinkVec_queue_dataIn_hi_hi_9 = {sinkVec_queue_19_enq_bits_vd, sinkVec_queue_19_enq_bits_offset};
  wire [3:0]   sinkVec_queue_19_enq_bits_mask;
  wire [11:0]  sinkVec_queue_dataIn_hi_19 = {sinkVec_queue_dataIn_hi_hi_9, sinkVec_queue_19_enq_bits_mask};
  wire [47:0]  sinkVec_queue_dataIn_19 = {sinkVec_queue_dataIn_hi_19, sinkVec_queue_dataIn_lo_19};
  wire [2:0]   sinkVec_queue_dataOut_19_instructionIndex = _sinkVec_queue_fifo_19_data_out[2:0];
  wire         sinkVec_queue_dataOut_19_last = _sinkVec_queue_fifo_19_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_19_data = _sinkVec_queue_fifo_19_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_19_mask = _sinkVec_queue_fifo_19_data_out[39:36];
  wire [2:0]   sinkVec_queue_dataOut_19_offset = _sinkVec_queue_fifo_19_data_out[42:40];
  wire [4:0]   sinkVec_queue_dataOut_19_vd = _sinkVec_queue_fifo_19_data_out[47:43];
  wire         sinkVec_queue_19_enq_ready = ~_sinkVec_queue_fifo_19_full;
  wire         sinkVec_queue_19_enq_valid;
  assign sinkVec_queue_19_deq_valid = ~_sinkVec_queue_fifo_19_empty | sinkVec_queue_19_enq_valid;
  assign sinkVec_queue_19_deq_bits_vd = _sinkVec_queue_fifo_19_empty ? sinkVec_queue_19_enq_bits_vd : sinkVec_queue_dataOut_19_vd;
  assign sinkVec_queue_19_deq_bits_offset = _sinkVec_queue_fifo_19_empty ? sinkVec_queue_19_enq_bits_offset : sinkVec_queue_dataOut_19_offset;
  assign sinkVec_queue_19_deq_bits_mask = _sinkVec_queue_fifo_19_empty ? sinkVec_queue_19_enq_bits_mask : sinkVec_queue_dataOut_19_mask;
  assign sinkVec_queue_19_deq_bits_data = _sinkVec_queue_fifo_19_empty ? sinkVec_queue_19_enq_bits_data : sinkVec_queue_dataOut_19_data;
  assign sinkVec_queue_19_deq_bits_last = _sinkVec_queue_fifo_19_empty ? sinkVec_queue_19_enq_bits_last : sinkVec_queue_dataOut_19_last;
  assign sinkVec_queue_19_deq_bits_instructionIndex = _sinkVec_queue_fifo_19_empty ? sinkVec_queue_19_enq_bits_instructionIndex : sinkVec_queue_dataOut_19_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_19;
  wire         sinkVec_releasePipe_pipe_out_19_valid = sinkVec_releasePipe_pipe_v_19;
  wire         x22_4_1_ready;
  wire         x22_4_1_valid;
  wire         sinkVec_validSource_19_valid = x22_4_1_ready & x22_4_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_19;
  wire [2:0]   sinkVec_tokenCheck_counterChange_19 = sinkVec_validSource_19_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_19 = ~(sinkVec_tokenCheck_counter_19[2]);
  assign x22_4_1_ready = sinkVec_tokenCheck_19;
  assign sinkVec_queue_19_enq_valid = sinkVec_validSink_19_valid;
  assign sinkVec_queue_19_enq_bits_vd = sinkVec_validSink_19_bits_vd;
  assign sinkVec_queue_19_enq_bits_offset = sinkVec_validSink_19_bits_offset;
  assign sinkVec_queue_19_enq_bits_mask = sinkVec_validSink_19_bits_mask;
  assign sinkVec_queue_19_enq_bits_data = sinkVec_validSink_19_bits_data;
  assign sinkVec_queue_19_enq_bits_last = sinkVec_validSink_19_bits_last;
  assign sinkVec_queue_19_enq_bits_instructionIndex = sinkVec_validSink_19_bits_instructionIndex;
  reg          sinkVec_shifterReg_19_0_valid;
  assign sinkVec_validSink_19_valid = sinkVec_shifterReg_19_0_valid;
  reg  [4:0]   sinkVec_shifterReg_19_0_bits_vd;
  assign sinkVec_validSink_19_bits_vd = sinkVec_shifterReg_19_0_bits_vd;
  reg  [2:0]   sinkVec_shifterReg_19_0_bits_offset;
  assign sinkVec_validSink_19_bits_offset = sinkVec_shifterReg_19_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_19_0_bits_mask;
  assign sinkVec_validSink_19_bits_mask = sinkVec_shifterReg_19_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_19_0_bits_data;
  assign sinkVec_validSink_19_bits_data = sinkVec_shifterReg_19_0_bits_data;
  reg          sinkVec_shifterReg_19_0_bits_last;
  assign sinkVec_validSink_19_bits_last = sinkVec_shifterReg_19_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_19_0_bits_instructionIndex;
  assign sinkVec_validSink_19_bits_instructionIndex = sinkVec_shifterReg_19_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_19 = sinkVec_shifterReg_19_0_valid | sinkVec_validSource_19_valid;
  assign sinkVec_sinkWire_18_ready = sinkVec_9_0_ready;
  assign sinkVec_sinkWire_19_ready = sinkVec_9_1_ready;
  reg          maskUnitFirst_9;
  wire         tryToRead_9 = sinkVec_9_0_valid | sinkVec_9_1_valid;
  wire         sinkWire_9_valid = maskUnitFirst_9 ? sinkVec_9_0_valid : sinkVec_9_1_valid;
  wire [4:0]   sinkWire_9_bits_vd = maskUnitFirst_9 ? sinkVec_9_0_bits_vd : sinkVec_9_1_bits_vd;
  wire [2:0]   sinkWire_9_bits_offset = maskUnitFirst_9 ? sinkVec_9_0_bits_offset : sinkVec_9_1_bits_offset;
  wire [3:0]   sinkWire_9_bits_mask = maskUnitFirst_9 ? sinkVec_9_0_bits_mask : sinkVec_9_1_bits_mask;
  wire [31:0]  sinkWire_9_bits_data = maskUnitFirst_9 ? sinkVec_9_0_bits_data : sinkVec_9_1_bits_data;
  wire         sinkWire_9_bits_last = maskUnitFirst_9 ? sinkVec_9_0_bits_last : sinkVec_9_1_bits_last;
  wire [2:0]   sinkWire_9_bits_instructionIndex = maskUnitFirst_9 ? sinkVec_9_0_bits_instructionIndex : sinkVec_9_1_bits_instructionIndex;
  wire         sinkWire_9_ready;
  assign sinkVec_9_1_ready = sinkWire_9_ready & ~maskUnitFirst_9;
  assign sinkVec_9_0_ready = sinkWire_9_ready & maskUnitFirst_9;
  reg          view__writeRelease_4_pipe_v;
  wire         view__writeRelease_4_pipe_out_valid = view__writeRelease_4_pipe_v;
  reg          pipe_v_12;
  wire         pipe_out_8_valid = pipe_v_12;
  wire         _probeWire_writeQueueEnqVec_4_valid_T = x22_4_0_ready & _maskUnit_exeResp_4_valid;
  reg          instructionFinishedPipe_pipe_v_4;
  wire         instructionFinishedPipe_pipe_out_4_valid = instructionFinishedPipe_pipe_v_4;
  reg  [7:0]   instructionFinishedPipe_pipe_b_4;
  wire [7:0]   instructionFinishedPipe_pipe_out_4_bits = instructionFinishedPipe_pipe_b_4;
  wire         instructionFinished_4_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_4_bits);
  wire         instructionFinished_4_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_4_bits);
  wire         instructionFinished_4_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_4_bits);
  wire         instructionFinished_4_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_4_bits);
  assign vxsatReportVec_4 = _laneVec_4_vxsatReport[3:0];
  reg          pipe_v_13;
  reg  [31:0]  pipe_b_13;
  reg          pipe_pipe_v_4;
  wire         pipe_pipe_out_4_valid = pipe_pipe_v_4;
  reg  [31:0]  pipe_pipe_b_4;
  wire [31:0]  pipe_pipe_out_4_bits = pipe_pipe_b_4;
  reg          view__laneMaskSelect_4_pipe_v;
  reg  [5:0]   view__laneMaskSelect_4_pipe_b;
  reg          view__laneMaskSelect_4_pipe_pipe_v;
  wire         view__laneMaskSelect_4_pipe_pipe_out_valid = view__laneMaskSelect_4_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_4_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_4_pipe_pipe_out_bits = view__laneMaskSelect_4_pipe_pipe_b;
  reg          view__laneMaskSewSelect_4_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_4_pipe_b;
  reg          view__laneMaskSewSelect_4_pipe_pipe_v;
  wire         view__laneMaskSewSelect_4_pipe_pipe_out_valid = view__laneMaskSewSelect_4_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_4_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_4_pipe_pipe_out_bits = view__laneMaskSewSelect_4_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v_4;
  wire         lsuLastPipe_pipe_out_4_valid = lsuLastPipe_pipe_v_4;
  reg  [7:0]   lsuLastPipe_pipe_b_4;
  wire [7:0]   lsuLastPipe_pipe_out_4_bits = lsuLastPipe_pipe_b_4;
  reg          maskLastPipe_pipe_v_4;
  wire         maskLastPipe_pipe_out_4_valid = maskLastPipe_pipe_v_4;
  reg  [7:0]   maskLastPipe_pipe_b_4;
  wire [7:0]   maskLastPipe_pipe_out_4_bits = maskLastPipe_pipe_b_4;
  wire [6:0]   writeCounter_4 = requestReg_bits_writeByte[11:5] + {6'h0, requestReg_bits_writeByte[4:0] > 5'h10};
  reg          pipe_v_14;
  wire         pipe_out_9_valid = pipe_v_14;
  reg  [6:0]   pipe_b_14;
  wire [6:0]   pipe_out_9_bits = pipe_b_14;
  assign laneRequestSinkWire_5_ready = ~laneRequestSinkWire_5_bits_issueInst | _laneVec_5_laneRequest_ready;
  wire         sinkVec_tokenCheck_20;
  wire [4:0]   sinkVec_validSource_20_bits_vs = x13_5_0_bits_vs;
  wire [2:0]   sinkVec_validSource_20_bits_offset = x13_5_0_bits_offset;
  wire [2:0]   sinkVec_validSource_20_bits_instructionIndex = x13_5_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_21;
  wire [4:0]   sinkVec_validSource_21_bits_vs = x13_5_1_bits_vs;
  wire [2:0]   sinkVec_validSource_21_bits_offset = x13_5_1_bits_offset;
  wire [2:0]   sinkVec_validSource_21_bits_instructionIndex = x13_5_1_bits_instructionIndex;
  wire         sinkVec_10_0_ready;
  wire         sinkVec_queue_20_deq_ready = sinkVec_sinkWire_20_ready;
  wire         sinkVec_queue_20_deq_valid;
  wire [4:0]   sinkVec_queue_20_deq_bits_vs;
  wire         sinkVec_10_0_valid = sinkVec_sinkWire_20_valid;
  wire [1:0]   sinkVec_queue_20_deq_bits_readSource;
  wire [4:0]   sinkVec_10_0_bits_vs = sinkVec_sinkWire_20_bits_vs;
  wire [2:0]   sinkVec_queue_20_deq_bits_offset;
  wire [1:0]   sinkVec_10_0_bits_readSource = sinkVec_sinkWire_20_bits_readSource;
  wire [2:0]   sinkVec_queue_20_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_10_0_bits_offset = sinkVec_sinkWire_20_bits_offset;
  wire [2:0]   sinkVec_10_0_bits_instructionIndex = sinkVec_sinkWire_20_bits_instructionIndex;
  wire         sinkVec_validSink_20_valid;
  wire [4:0]   sinkVec_validSink_20_bits_vs;
  wire [1:0]   sinkVec_validSink_20_bits_readSource;
  wire [2:0]   sinkVec_validSink_20_bits_offset;
  wire [2:0]   sinkVec_validSink_20_bits_instructionIndex;
  assign sinkVec_sinkWire_20_valid = sinkVec_queue_20_deq_valid;
  assign sinkVec_sinkWire_20_bits_vs = sinkVec_queue_20_deq_bits_vs;
  assign sinkVec_sinkWire_20_bits_readSource = sinkVec_queue_20_deq_bits_readSource;
  assign sinkVec_sinkWire_20_bits_offset = sinkVec_queue_20_deq_bits_offset;
  assign sinkVec_sinkWire_20_bits_instructionIndex = sinkVec_queue_20_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_queue_20_enq_bits_offset;
  wire [2:0]   sinkVec_queue_20_enq_bits_instructionIndex;
  wire [5:0]   sinkVec_queue_dataIn_lo_20 = {sinkVec_queue_20_enq_bits_offset, sinkVec_queue_20_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_20_enq_bits_vs;
  wire [1:0]   sinkVec_queue_20_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_20 = {sinkVec_queue_20_enq_bits_vs, sinkVec_queue_20_enq_bits_readSource};
  wire [12:0]  sinkVec_queue_dataIn_20 = {sinkVec_queue_dataIn_hi_20, sinkVec_queue_dataIn_lo_20};
  wire [2:0]   sinkVec_queue_dataOut_20_instructionIndex = _sinkVec_queue_fifo_20_data_out[2:0];
  wire [2:0]   sinkVec_queue_dataOut_20_offset = _sinkVec_queue_fifo_20_data_out[5:3];
  wire [1:0]   sinkVec_queue_dataOut_20_readSource = _sinkVec_queue_fifo_20_data_out[7:6];
  wire [4:0]   sinkVec_queue_dataOut_20_vs = _sinkVec_queue_fifo_20_data_out[12:8];
  wire         sinkVec_queue_20_enq_ready = ~_sinkVec_queue_fifo_20_full;
  wire         sinkVec_queue_20_enq_valid;
  assign sinkVec_queue_20_deq_valid = ~_sinkVec_queue_fifo_20_empty | sinkVec_queue_20_enq_valid;
  assign sinkVec_queue_20_deq_bits_vs = _sinkVec_queue_fifo_20_empty ? sinkVec_queue_20_enq_bits_vs : sinkVec_queue_dataOut_20_vs;
  assign sinkVec_queue_20_deq_bits_readSource = _sinkVec_queue_fifo_20_empty ? sinkVec_queue_20_enq_bits_readSource : sinkVec_queue_dataOut_20_readSource;
  assign sinkVec_queue_20_deq_bits_offset = _sinkVec_queue_fifo_20_empty ? sinkVec_queue_20_enq_bits_offset : sinkVec_queue_dataOut_20_offset;
  assign sinkVec_queue_20_deq_bits_instructionIndex = _sinkVec_queue_fifo_20_empty ? sinkVec_queue_20_enq_bits_instructionIndex : sinkVec_queue_dataOut_20_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_20;
  wire         sinkVec_releasePipe_pipe_out_20_valid = sinkVec_releasePipe_pipe_v_20;
  wire         x13_5_0_ready;
  wire         x13_5_0_valid;
  wire         sinkVec_validSource_20_valid = x13_5_0_ready & x13_5_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_20;
  wire [2:0]   sinkVec_tokenCheck_counterChange_20 = sinkVec_validSource_20_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_20 = ~(sinkVec_tokenCheck_counter_20[2]);
  assign x13_5_0_ready = sinkVec_tokenCheck_20;
  assign sinkVec_queue_20_enq_valid = sinkVec_validSink_20_valid;
  assign sinkVec_queue_20_enq_bits_vs = sinkVec_validSink_20_bits_vs;
  assign sinkVec_queue_20_enq_bits_readSource = sinkVec_validSink_20_bits_readSource;
  assign sinkVec_queue_20_enq_bits_offset = sinkVec_validSink_20_bits_offset;
  assign sinkVec_queue_20_enq_bits_instructionIndex = sinkVec_validSink_20_bits_instructionIndex;
  reg          sinkVec_shifterReg_20_0_valid;
  assign sinkVec_validSink_20_valid = sinkVec_shifterReg_20_0_valid;
  reg  [4:0]   sinkVec_shifterReg_20_0_bits_vs;
  assign sinkVec_validSink_20_bits_vs = sinkVec_shifterReg_20_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_20_0_bits_readSource;
  assign sinkVec_validSink_20_bits_readSource = sinkVec_shifterReg_20_0_bits_readSource;
  reg  [2:0]   sinkVec_shifterReg_20_0_bits_offset;
  assign sinkVec_validSink_20_bits_offset = sinkVec_shifterReg_20_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_20_0_bits_instructionIndex;
  assign sinkVec_validSink_20_bits_instructionIndex = sinkVec_shifterReg_20_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_20 = sinkVec_shifterReg_20_0_valid | sinkVec_validSource_20_valid;
  wire         sinkVec_10_1_ready;
  wire         sinkVec_queue_21_deq_ready = sinkVec_sinkWire_21_ready;
  wire         sinkVec_queue_21_deq_valid;
  wire [4:0]   sinkVec_queue_21_deq_bits_vs;
  wire         sinkVec_10_1_valid = sinkVec_sinkWire_21_valid;
  wire [1:0]   sinkVec_queue_21_deq_bits_readSource;
  wire [4:0]   sinkVec_10_1_bits_vs = sinkVec_sinkWire_21_bits_vs;
  wire [2:0]   sinkVec_queue_21_deq_bits_offset;
  wire [1:0]   sinkVec_10_1_bits_readSource = sinkVec_sinkWire_21_bits_readSource;
  wire [2:0]   sinkVec_queue_21_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_10_1_bits_offset = sinkVec_sinkWire_21_bits_offset;
  wire [2:0]   sinkVec_10_1_bits_instructionIndex = sinkVec_sinkWire_21_bits_instructionIndex;
  wire         sinkVec_validSink_21_valid;
  wire [4:0]   sinkVec_validSink_21_bits_vs;
  wire [1:0]   sinkVec_validSink_21_bits_readSource;
  wire [2:0]   sinkVec_validSink_21_bits_offset;
  wire [2:0]   sinkVec_validSink_21_bits_instructionIndex;
  assign sinkVec_sinkWire_21_valid = sinkVec_queue_21_deq_valid;
  assign sinkVec_sinkWire_21_bits_vs = sinkVec_queue_21_deq_bits_vs;
  assign sinkVec_sinkWire_21_bits_readSource = sinkVec_queue_21_deq_bits_readSource;
  assign sinkVec_sinkWire_21_bits_offset = sinkVec_queue_21_deq_bits_offset;
  assign sinkVec_sinkWire_21_bits_instructionIndex = sinkVec_queue_21_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_queue_21_enq_bits_offset;
  wire [2:0]   sinkVec_queue_21_enq_bits_instructionIndex;
  wire [5:0]   sinkVec_queue_dataIn_lo_21 = {sinkVec_queue_21_enq_bits_offset, sinkVec_queue_21_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_21_enq_bits_vs;
  wire [1:0]   sinkVec_queue_21_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_21 = {sinkVec_queue_21_enq_bits_vs, sinkVec_queue_21_enq_bits_readSource};
  wire [12:0]  sinkVec_queue_dataIn_21 = {sinkVec_queue_dataIn_hi_21, sinkVec_queue_dataIn_lo_21};
  wire [2:0]   sinkVec_queue_dataOut_21_instructionIndex = _sinkVec_queue_fifo_21_data_out[2:0];
  wire [2:0]   sinkVec_queue_dataOut_21_offset = _sinkVec_queue_fifo_21_data_out[5:3];
  wire [1:0]   sinkVec_queue_dataOut_21_readSource = _sinkVec_queue_fifo_21_data_out[7:6];
  wire [4:0]   sinkVec_queue_dataOut_21_vs = _sinkVec_queue_fifo_21_data_out[12:8];
  wire         sinkVec_queue_21_enq_ready = ~_sinkVec_queue_fifo_21_full;
  wire         sinkVec_queue_21_enq_valid;
  assign sinkVec_queue_21_deq_valid = ~_sinkVec_queue_fifo_21_empty | sinkVec_queue_21_enq_valid;
  assign sinkVec_queue_21_deq_bits_vs = _sinkVec_queue_fifo_21_empty ? sinkVec_queue_21_enq_bits_vs : sinkVec_queue_dataOut_21_vs;
  assign sinkVec_queue_21_deq_bits_readSource = _sinkVec_queue_fifo_21_empty ? sinkVec_queue_21_enq_bits_readSource : sinkVec_queue_dataOut_21_readSource;
  assign sinkVec_queue_21_deq_bits_offset = _sinkVec_queue_fifo_21_empty ? sinkVec_queue_21_enq_bits_offset : sinkVec_queue_dataOut_21_offset;
  assign sinkVec_queue_21_deq_bits_instructionIndex = _sinkVec_queue_fifo_21_empty ? sinkVec_queue_21_enq_bits_instructionIndex : sinkVec_queue_dataOut_21_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_21;
  wire         sinkVec_releasePipe_pipe_out_21_valid = sinkVec_releasePipe_pipe_v_21;
  wire         x13_5_1_ready;
  wire         x13_5_1_valid;
  wire         sinkVec_validSource_21_valid = x13_5_1_ready & x13_5_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_21;
  wire [2:0]   sinkVec_tokenCheck_counterChange_21 = sinkVec_validSource_21_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_21 = ~(sinkVec_tokenCheck_counter_21[2]);
  assign x13_5_1_ready = sinkVec_tokenCheck_21;
  assign sinkVec_queue_21_enq_valid = sinkVec_validSink_21_valid;
  assign sinkVec_queue_21_enq_bits_vs = sinkVec_validSink_21_bits_vs;
  assign sinkVec_queue_21_enq_bits_readSource = sinkVec_validSink_21_bits_readSource;
  assign sinkVec_queue_21_enq_bits_offset = sinkVec_validSink_21_bits_offset;
  assign sinkVec_queue_21_enq_bits_instructionIndex = sinkVec_validSink_21_bits_instructionIndex;
  reg          sinkVec_shifterReg_21_0_valid;
  assign sinkVec_validSink_21_valid = sinkVec_shifterReg_21_0_valid;
  reg  [4:0]   sinkVec_shifterReg_21_0_bits_vs;
  assign sinkVec_validSink_21_bits_vs = sinkVec_shifterReg_21_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_21_0_bits_readSource;
  assign sinkVec_validSink_21_bits_readSource = sinkVec_shifterReg_21_0_bits_readSource;
  reg  [2:0]   sinkVec_shifterReg_21_0_bits_offset;
  assign sinkVec_validSink_21_bits_offset = sinkVec_shifterReg_21_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_21_0_bits_instructionIndex;
  assign sinkVec_validSink_21_bits_instructionIndex = sinkVec_shifterReg_21_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_21 = sinkVec_shifterReg_21_0_valid | sinkVec_validSource_21_valid;
  assign sinkVec_sinkWire_20_ready = sinkVec_10_0_ready;
  assign sinkVec_sinkWire_21_ready = sinkVec_10_1_ready;
  reg          maskUnitFirst_10;
  wire         tryToRead_10 = sinkVec_10_0_valid | sinkVec_10_1_valid;
  wire         sinkWire_10_valid = maskUnitFirst_10 ? sinkVec_10_0_valid : sinkVec_10_1_valid;
  wire [4:0]   sinkWire_10_bits_vs = maskUnitFirst_10 ? sinkVec_10_0_bits_vs : sinkVec_10_1_bits_vs;
  wire [1:0]   sinkWire_10_bits_readSource = maskUnitFirst_10 ? sinkVec_10_0_bits_readSource : sinkVec_10_1_bits_readSource;
  wire [2:0]   sinkWire_10_bits_offset = maskUnitFirst_10 ? sinkVec_10_0_bits_offset : sinkVec_10_1_bits_offset;
  wire [2:0]   sinkWire_10_bits_instructionIndex = maskUnitFirst_10 ? sinkVec_10_0_bits_instructionIndex : sinkVec_10_1_bits_instructionIndex;
  wire         sinkWire_10_ready;
  assign sinkVec_10_1_ready = sinkWire_10_ready & ~maskUnitFirst_10;
  assign sinkVec_10_0_ready = sinkWire_10_ready & maskUnitFirst_10;
  reg          accessDataValid_pipe_v_10;
  reg          accessDataValid_pipe_pipe_v_10;
  wire         accessDataValid_pipe_pipe_out_10_valid = accessDataValid_pipe_pipe_v_10;
  wire         accessDataSource_10_valid = accessDataValid_pipe_pipe_out_10_valid;
  reg          shifterReg_18_0_valid;
  reg  [31:0]  shifterReg_18_0_bits;
  wire         shifterValid_18 = shifterReg_18_0_valid | accessDataSource_10_valid;
  reg          accessDataValid_pipe_v_11;
  reg          accessDataValid_pipe_pipe_v_11;
  wire         accessDataValid_pipe_pipe_out_11_valid = accessDataValid_pipe_pipe_v_11;
  wire         accessDataSource_11_valid = accessDataValid_pipe_pipe_out_11_valid;
  reg          shifterReg_19_0_valid;
  reg  [31:0]  shifterReg_19_0_bits;
  wire         shifterValid_19 = shifterReg_19_0_valid | accessDataSource_11_valid;
  wire         sinkVec_tokenCheck_22;
  wire [4:0]   sinkVec_validSource_22_bits_vd = x22_5_0_bits_vd;
  wire [2:0]   sinkVec_validSource_22_bits_offset = x22_5_0_bits_offset;
  wire [3:0]   sinkVec_validSource_22_bits_mask = x22_5_0_bits_mask;
  wire [31:0]  sinkVec_validSource_22_bits_data = x22_5_0_bits_data;
  wire [2:0]   sinkVec_validSource_22_bits_instructionIndex = x22_5_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_23;
  wire [4:0]   sinkVec_validSource_23_bits_vd = x22_5_1_bits_vd;
  wire [2:0]   sinkVec_validSource_23_bits_offset = x22_5_1_bits_offset;
  wire [3:0]   sinkVec_validSource_23_bits_mask = x22_5_1_bits_mask;
  wire [31:0]  sinkVec_validSource_23_bits_data = x22_5_1_bits_data;
  wire         sinkVec_validSource_23_bits_last = x22_5_1_bits_last;
  wire [2:0]   sinkVec_validSource_23_bits_instructionIndex = x22_5_1_bits_instructionIndex;
  wire         sinkVec_11_0_ready;
  wire         sinkVec_queue_22_deq_ready = sinkVec_sinkWire_22_ready;
  wire         sinkVec_queue_22_deq_valid;
  wire [4:0]   sinkVec_queue_22_deq_bits_vd;
  wire         sinkVec_11_0_valid = sinkVec_sinkWire_22_valid;
  wire [2:0]   sinkVec_queue_22_deq_bits_offset;
  wire [4:0]   sinkVec_11_0_bits_vd = sinkVec_sinkWire_22_bits_vd;
  wire [3:0]   sinkVec_queue_22_deq_bits_mask;
  wire [2:0]   sinkVec_11_0_bits_offset = sinkVec_sinkWire_22_bits_offset;
  wire [31:0]  sinkVec_queue_22_deq_bits_data;
  wire [3:0]   sinkVec_11_0_bits_mask = sinkVec_sinkWire_22_bits_mask;
  wire         sinkVec_queue_22_deq_bits_last;
  wire [31:0]  sinkVec_11_0_bits_data = sinkVec_sinkWire_22_bits_data;
  wire [2:0]   sinkVec_queue_22_deq_bits_instructionIndex;
  wire         sinkVec_11_0_bits_last = sinkVec_sinkWire_22_bits_last;
  wire [2:0]   sinkVec_11_0_bits_instructionIndex = sinkVec_sinkWire_22_bits_instructionIndex;
  wire         sinkVec_validSink_22_valid;
  wire [4:0]   sinkVec_validSink_22_bits_vd;
  wire [2:0]   sinkVec_validSink_22_bits_offset;
  wire [3:0]   sinkVec_validSink_22_bits_mask;
  wire [31:0]  sinkVec_validSink_22_bits_data;
  wire [2:0]   sinkVec_validSink_22_bits_instructionIndex;
  assign sinkVec_sinkWire_22_valid = sinkVec_queue_22_deq_valid;
  assign sinkVec_sinkWire_22_bits_vd = sinkVec_queue_22_deq_bits_vd;
  assign sinkVec_sinkWire_22_bits_offset = sinkVec_queue_22_deq_bits_offset;
  assign sinkVec_sinkWire_22_bits_mask = sinkVec_queue_22_deq_bits_mask;
  assign sinkVec_sinkWire_22_bits_data = sinkVec_queue_22_deq_bits_data;
  assign sinkVec_sinkWire_22_bits_last = sinkVec_queue_22_deq_bits_last;
  assign sinkVec_sinkWire_22_bits_instructionIndex = sinkVec_queue_22_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_22_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_10 = {sinkVec_queue_22_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_22_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_22 = {sinkVec_queue_dataIn_lo_hi_10, sinkVec_queue_22_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_22_enq_bits_vd;
  wire [2:0]   sinkVec_queue_22_enq_bits_offset;
  wire [7:0]   sinkVec_queue_dataIn_hi_hi_10 = {sinkVec_queue_22_enq_bits_vd, sinkVec_queue_22_enq_bits_offset};
  wire [3:0]   sinkVec_queue_22_enq_bits_mask;
  wire [11:0]  sinkVec_queue_dataIn_hi_22 = {sinkVec_queue_dataIn_hi_hi_10, sinkVec_queue_22_enq_bits_mask};
  wire [47:0]  sinkVec_queue_dataIn_22 = {sinkVec_queue_dataIn_hi_22, sinkVec_queue_dataIn_lo_22};
  wire [2:0]   sinkVec_queue_dataOut_22_instructionIndex = _sinkVec_queue_fifo_22_data_out[2:0];
  wire         sinkVec_queue_dataOut_22_last = _sinkVec_queue_fifo_22_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_22_data = _sinkVec_queue_fifo_22_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_22_mask = _sinkVec_queue_fifo_22_data_out[39:36];
  wire [2:0]   sinkVec_queue_dataOut_22_offset = _sinkVec_queue_fifo_22_data_out[42:40];
  wire [4:0]   sinkVec_queue_dataOut_22_vd = _sinkVec_queue_fifo_22_data_out[47:43];
  wire         sinkVec_queue_22_enq_ready = ~_sinkVec_queue_fifo_22_full;
  wire         sinkVec_queue_22_enq_valid;
  assign sinkVec_queue_22_deq_valid = ~_sinkVec_queue_fifo_22_empty | sinkVec_queue_22_enq_valid;
  assign sinkVec_queue_22_deq_bits_vd = _sinkVec_queue_fifo_22_empty ? sinkVec_queue_22_enq_bits_vd : sinkVec_queue_dataOut_22_vd;
  assign sinkVec_queue_22_deq_bits_offset = _sinkVec_queue_fifo_22_empty ? sinkVec_queue_22_enq_bits_offset : sinkVec_queue_dataOut_22_offset;
  assign sinkVec_queue_22_deq_bits_mask = _sinkVec_queue_fifo_22_empty ? sinkVec_queue_22_enq_bits_mask : sinkVec_queue_dataOut_22_mask;
  assign sinkVec_queue_22_deq_bits_data = _sinkVec_queue_fifo_22_empty ? sinkVec_queue_22_enq_bits_data : sinkVec_queue_dataOut_22_data;
  assign sinkVec_queue_22_deq_bits_last = ~_sinkVec_queue_fifo_22_empty & sinkVec_queue_dataOut_22_last;
  assign sinkVec_queue_22_deq_bits_instructionIndex = _sinkVec_queue_fifo_22_empty ? sinkVec_queue_22_enq_bits_instructionIndex : sinkVec_queue_dataOut_22_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_22;
  wire         sinkVec_releasePipe_pipe_out_22_valid = sinkVec_releasePipe_pipe_v_22;
  wire         x22_5_0_ready;
  wire         x22_5_0_valid;
  wire         sinkVec_validSource_22_valid = x22_5_0_ready & x22_5_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_22;
  wire [2:0]   sinkVec_tokenCheck_counterChange_22 = sinkVec_validSource_22_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_22 = ~(sinkVec_tokenCheck_counter_22[2]);
  assign x22_5_0_ready = sinkVec_tokenCheck_22;
  assign sinkVec_queue_22_enq_valid = sinkVec_validSink_22_valid;
  assign sinkVec_queue_22_enq_bits_vd = sinkVec_validSink_22_bits_vd;
  assign sinkVec_queue_22_enq_bits_offset = sinkVec_validSink_22_bits_offset;
  assign sinkVec_queue_22_enq_bits_mask = sinkVec_validSink_22_bits_mask;
  assign sinkVec_queue_22_enq_bits_data = sinkVec_validSink_22_bits_data;
  assign sinkVec_queue_22_enq_bits_instructionIndex = sinkVec_validSink_22_bits_instructionIndex;
  reg          sinkVec_shifterReg_22_0_valid;
  assign sinkVec_validSink_22_valid = sinkVec_shifterReg_22_0_valid;
  reg  [4:0]   sinkVec_shifterReg_22_0_bits_vd;
  assign sinkVec_validSink_22_bits_vd = sinkVec_shifterReg_22_0_bits_vd;
  reg  [2:0]   sinkVec_shifterReg_22_0_bits_offset;
  assign sinkVec_validSink_22_bits_offset = sinkVec_shifterReg_22_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_22_0_bits_mask;
  assign sinkVec_validSink_22_bits_mask = sinkVec_shifterReg_22_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_22_0_bits_data;
  assign sinkVec_validSink_22_bits_data = sinkVec_shifterReg_22_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_22_0_bits_instructionIndex;
  assign sinkVec_validSink_22_bits_instructionIndex = sinkVec_shifterReg_22_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_22 = sinkVec_shifterReg_22_0_valid | sinkVec_validSource_22_valid;
  wire         sinkVec_11_1_ready;
  wire         sinkVec_queue_23_deq_ready = sinkVec_sinkWire_23_ready;
  wire         sinkVec_queue_23_deq_valid;
  wire [4:0]   sinkVec_queue_23_deq_bits_vd;
  wire         sinkVec_11_1_valid = sinkVec_sinkWire_23_valid;
  wire [2:0]   sinkVec_queue_23_deq_bits_offset;
  wire [4:0]   sinkVec_11_1_bits_vd = sinkVec_sinkWire_23_bits_vd;
  wire [3:0]   sinkVec_queue_23_deq_bits_mask;
  wire [2:0]   sinkVec_11_1_bits_offset = sinkVec_sinkWire_23_bits_offset;
  wire [31:0]  sinkVec_queue_23_deq_bits_data;
  wire [3:0]   sinkVec_11_1_bits_mask = sinkVec_sinkWire_23_bits_mask;
  wire         sinkVec_queue_23_deq_bits_last;
  wire [31:0]  sinkVec_11_1_bits_data = sinkVec_sinkWire_23_bits_data;
  wire [2:0]   sinkVec_queue_23_deq_bits_instructionIndex;
  wire         sinkVec_11_1_bits_last = sinkVec_sinkWire_23_bits_last;
  wire [2:0]   sinkVec_11_1_bits_instructionIndex = sinkVec_sinkWire_23_bits_instructionIndex;
  wire         sinkVec_validSink_23_valid;
  wire [4:0]   sinkVec_validSink_23_bits_vd;
  wire [2:0]   sinkVec_validSink_23_bits_offset;
  wire [3:0]   sinkVec_validSink_23_bits_mask;
  wire [31:0]  sinkVec_validSink_23_bits_data;
  wire         sinkVec_validSink_23_bits_last;
  wire [2:0]   sinkVec_validSink_23_bits_instructionIndex;
  assign sinkVec_sinkWire_23_valid = sinkVec_queue_23_deq_valid;
  assign sinkVec_sinkWire_23_bits_vd = sinkVec_queue_23_deq_bits_vd;
  assign sinkVec_sinkWire_23_bits_offset = sinkVec_queue_23_deq_bits_offset;
  assign sinkVec_sinkWire_23_bits_mask = sinkVec_queue_23_deq_bits_mask;
  assign sinkVec_sinkWire_23_bits_data = sinkVec_queue_23_deq_bits_data;
  assign sinkVec_sinkWire_23_bits_last = sinkVec_queue_23_deq_bits_last;
  assign sinkVec_sinkWire_23_bits_instructionIndex = sinkVec_queue_23_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_23_enq_bits_data;
  wire         sinkVec_queue_23_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_11 = {sinkVec_queue_23_enq_bits_data, sinkVec_queue_23_enq_bits_last};
  wire [2:0]   sinkVec_queue_23_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_23 = {sinkVec_queue_dataIn_lo_hi_11, sinkVec_queue_23_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_23_enq_bits_vd;
  wire [2:0]   sinkVec_queue_23_enq_bits_offset;
  wire [7:0]   sinkVec_queue_dataIn_hi_hi_11 = {sinkVec_queue_23_enq_bits_vd, sinkVec_queue_23_enq_bits_offset};
  wire [3:0]   sinkVec_queue_23_enq_bits_mask;
  wire [11:0]  sinkVec_queue_dataIn_hi_23 = {sinkVec_queue_dataIn_hi_hi_11, sinkVec_queue_23_enq_bits_mask};
  wire [47:0]  sinkVec_queue_dataIn_23 = {sinkVec_queue_dataIn_hi_23, sinkVec_queue_dataIn_lo_23};
  wire [2:0]   sinkVec_queue_dataOut_23_instructionIndex = _sinkVec_queue_fifo_23_data_out[2:0];
  wire         sinkVec_queue_dataOut_23_last = _sinkVec_queue_fifo_23_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_23_data = _sinkVec_queue_fifo_23_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_23_mask = _sinkVec_queue_fifo_23_data_out[39:36];
  wire [2:0]   sinkVec_queue_dataOut_23_offset = _sinkVec_queue_fifo_23_data_out[42:40];
  wire [4:0]   sinkVec_queue_dataOut_23_vd = _sinkVec_queue_fifo_23_data_out[47:43];
  wire         sinkVec_queue_23_enq_ready = ~_sinkVec_queue_fifo_23_full;
  wire         sinkVec_queue_23_enq_valid;
  assign sinkVec_queue_23_deq_valid = ~_sinkVec_queue_fifo_23_empty | sinkVec_queue_23_enq_valid;
  assign sinkVec_queue_23_deq_bits_vd = _sinkVec_queue_fifo_23_empty ? sinkVec_queue_23_enq_bits_vd : sinkVec_queue_dataOut_23_vd;
  assign sinkVec_queue_23_deq_bits_offset = _sinkVec_queue_fifo_23_empty ? sinkVec_queue_23_enq_bits_offset : sinkVec_queue_dataOut_23_offset;
  assign sinkVec_queue_23_deq_bits_mask = _sinkVec_queue_fifo_23_empty ? sinkVec_queue_23_enq_bits_mask : sinkVec_queue_dataOut_23_mask;
  assign sinkVec_queue_23_deq_bits_data = _sinkVec_queue_fifo_23_empty ? sinkVec_queue_23_enq_bits_data : sinkVec_queue_dataOut_23_data;
  assign sinkVec_queue_23_deq_bits_last = _sinkVec_queue_fifo_23_empty ? sinkVec_queue_23_enq_bits_last : sinkVec_queue_dataOut_23_last;
  assign sinkVec_queue_23_deq_bits_instructionIndex = _sinkVec_queue_fifo_23_empty ? sinkVec_queue_23_enq_bits_instructionIndex : sinkVec_queue_dataOut_23_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_23;
  wire         sinkVec_releasePipe_pipe_out_23_valid = sinkVec_releasePipe_pipe_v_23;
  wire         x22_5_1_ready;
  wire         x22_5_1_valid;
  wire         sinkVec_validSource_23_valid = x22_5_1_ready & x22_5_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_23;
  wire [2:0]   sinkVec_tokenCheck_counterChange_23 = sinkVec_validSource_23_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_23 = ~(sinkVec_tokenCheck_counter_23[2]);
  assign x22_5_1_ready = sinkVec_tokenCheck_23;
  assign sinkVec_queue_23_enq_valid = sinkVec_validSink_23_valid;
  assign sinkVec_queue_23_enq_bits_vd = sinkVec_validSink_23_bits_vd;
  assign sinkVec_queue_23_enq_bits_offset = sinkVec_validSink_23_bits_offset;
  assign sinkVec_queue_23_enq_bits_mask = sinkVec_validSink_23_bits_mask;
  assign sinkVec_queue_23_enq_bits_data = sinkVec_validSink_23_bits_data;
  assign sinkVec_queue_23_enq_bits_last = sinkVec_validSink_23_bits_last;
  assign sinkVec_queue_23_enq_bits_instructionIndex = sinkVec_validSink_23_bits_instructionIndex;
  reg          sinkVec_shifterReg_23_0_valid;
  assign sinkVec_validSink_23_valid = sinkVec_shifterReg_23_0_valid;
  reg  [4:0]   sinkVec_shifterReg_23_0_bits_vd;
  assign sinkVec_validSink_23_bits_vd = sinkVec_shifterReg_23_0_bits_vd;
  reg  [2:0]   sinkVec_shifterReg_23_0_bits_offset;
  assign sinkVec_validSink_23_bits_offset = sinkVec_shifterReg_23_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_23_0_bits_mask;
  assign sinkVec_validSink_23_bits_mask = sinkVec_shifterReg_23_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_23_0_bits_data;
  assign sinkVec_validSink_23_bits_data = sinkVec_shifterReg_23_0_bits_data;
  reg          sinkVec_shifterReg_23_0_bits_last;
  assign sinkVec_validSink_23_bits_last = sinkVec_shifterReg_23_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_23_0_bits_instructionIndex;
  assign sinkVec_validSink_23_bits_instructionIndex = sinkVec_shifterReg_23_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_23 = sinkVec_shifterReg_23_0_valid | sinkVec_validSource_23_valid;
  assign sinkVec_sinkWire_22_ready = sinkVec_11_0_ready;
  assign sinkVec_sinkWire_23_ready = sinkVec_11_1_ready;
  reg          maskUnitFirst_11;
  wire         tryToRead_11 = sinkVec_11_0_valid | sinkVec_11_1_valid;
  wire         sinkWire_11_valid = maskUnitFirst_11 ? sinkVec_11_0_valid : sinkVec_11_1_valid;
  wire [4:0]   sinkWire_11_bits_vd = maskUnitFirst_11 ? sinkVec_11_0_bits_vd : sinkVec_11_1_bits_vd;
  wire [2:0]   sinkWire_11_bits_offset = maskUnitFirst_11 ? sinkVec_11_0_bits_offset : sinkVec_11_1_bits_offset;
  wire [3:0]   sinkWire_11_bits_mask = maskUnitFirst_11 ? sinkVec_11_0_bits_mask : sinkVec_11_1_bits_mask;
  wire [31:0]  sinkWire_11_bits_data = maskUnitFirst_11 ? sinkVec_11_0_bits_data : sinkVec_11_1_bits_data;
  wire         sinkWire_11_bits_last = maskUnitFirst_11 ? sinkVec_11_0_bits_last : sinkVec_11_1_bits_last;
  wire [2:0]   sinkWire_11_bits_instructionIndex = maskUnitFirst_11 ? sinkVec_11_0_bits_instructionIndex : sinkVec_11_1_bits_instructionIndex;
  wire         sinkWire_11_ready;
  assign sinkVec_11_1_ready = sinkWire_11_ready & ~maskUnitFirst_11;
  assign sinkVec_11_0_ready = sinkWire_11_ready & maskUnitFirst_11;
  reg          view__writeRelease_5_pipe_v;
  wire         view__writeRelease_5_pipe_out_valid = view__writeRelease_5_pipe_v;
  reg          pipe_v_15;
  wire         pipe_out_10_valid = pipe_v_15;
  wire         _probeWire_writeQueueEnqVec_5_valid_T = x22_5_0_ready & _maskUnit_exeResp_5_valid;
  reg          instructionFinishedPipe_pipe_v_5;
  wire         instructionFinishedPipe_pipe_out_5_valid = instructionFinishedPipe_pipe_v_5;
  reg  [7:0]   instructionFinishedPipe_pipe_b_5;
  wire [7:0]   instructionFinishedPipe_pipe_out_5_bits = instructionFinishedPipe_pipe_b_5;
  wire         instructionFinished_5_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_5_bits);
  wire         instructionFinished_5_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_5_bits);
  wire         instructionFinished_5_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_5_bits);
  wire         instructionFinished_5_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_5_bits);
  assign vxsatReportVec_5 = _laneVec_5_vxsatReport[3:0];
  reg          pipe_v_16;
  reg  [31:0]  pipe_b_16;
  reg          pipe_pipe_v_5;
  wire         pipe_pipe_out_5_valid = pipe_pipe_v_5;
  reg  [31:0]  pipe_pipe_b_5;
  wire [31:0]  pipe_pipe_out_5_bits = pipe_pipe_b_5;
  reg          view__laneMaskSelect_5_pipe_v;
  reg  [5:0]   view__laneMaskSelect_5_pipe_b;
  reg          view__laneMaskSelect_5_pipe_pipe_v;
  wire         view__laneMaskSelect_5_pipe_pipe_out_valid = view__laneMaskSelect_5_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_5_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_5_pipe_pipe_out_bits = view__laneMaskSelect_5_pipe_pipe_b;
  reg          view__laneMaskSewSelect_5_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_5_pipe_b;
  reg          view__laneMaskSewSelect_5_pipe_pipe_v;
  wire         view__laneMaskSewSelect_5_pipe_pipe_out_valid = view__laneMaskSewSelect_5_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_5_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_5_pipe_pipe_out_bits = view__laneMaskSewSelect_5_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v_5;
  wire         lsuLastPipe_pipe_out_5_valid = lsuLastPipe_pipe_v_5;
  reg  [7:0]   lsuLastPipe_pipe_b_5;
  wire [7:0]   lsuLastPipe_pipe_out_5_bits = lsuLastPipe_pipe_b_5;
  reg          maskLastPipe_pipe_v_5;
  wire         maskLastPipe_pipe_out_5_valid = maskLastPipe_pipe_v_5;
  reg  [7:0]   maskLastPipe_pipe_b_5;
  wire [7:0]   maskLastPipe_pipe_out_5_bits = maskLastPipe_pipe_b_5;
  wire [6:0]   writeCounter_5 = requestReg_bits_writeByte[11:5] + {6'h0, requestReg_bits_writeByte[4:0] > 5'h14};
  reg          pipe_v_17;
  wire         pipe_out_11_valid = pipe_v_17;
  reg  [6:0]   pipe_b_17;
  wire [6:0]   pipe_out_11_bits = pipe_b_17;
  assign laneRequestSinkWire_6_ready = ~laneRequestSinkWire_6_bits_issueInst | _laneVec_6_laneRequest_ready;
  wire         sinkVec_tokenCheck_24;
  wire [4:0]   sinkVec_validSource_24_bits_vs = x13_6_0_bits_vs;
  wire [2:0]   sinkVec_validSource_24_bits_offset = x13_6_0_bits_offset;
  wire [2:0]   sinkVec_validSource_24_bits_instructionIndex = x13_6_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_25;
  wire [4:0]   sinkVec_validSource_25_bits_vs = x13_6_1_bits_vs;
  wire [2:0]   sinkVec_validSource_25_bits_offset = x13_6_1_bits_offset;
  wire [2:0]   sinkVec_validSource_25_bits_instructionIndex = x13_6_1_bits_instructionIndex;
  wire         sinkVec_12_0_ready;
  wire         sinkVec_queue_24_deq_ready = sinkVec_sinkWire_24_ready;
  wire         sinkVec_queue_24_deq_valid;
  wire [4:0]   sinkVec_queue_24_deq_bits_vs;
  wire         sinkVec_12_0_valid = sinkVec_sinkWire_24_valid;
  wire [1:0]   sinkVec_queue_24_deq_bits_readSource;
  wire [4:0]   sinkVec_12_0_bits_vs = sinkVec_sinkWire_24_bits_vs;
  wire [2:0]   sinkVec_queue_24_deq_bits_offset;
  wire [1:0]   sinkVec_12_0_bits_readSource = sinkVec_sinkWire_24_bits_readSource;
  wire [2:0]   sinkVec_queue_24_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_12_0_bits_offset = sinkVec_sinkWire_24_bits_offset;
  wire [2:0]   sinkVec_12_0_bits_instructionIndex = sinkVec_sinkWire_24_bits_instructionIndex;
  wire         sinkVec_validSink_24_valid;
  wire [4:0]   sinkVec_validSink_24_bits_vs;
  wire [1:0]   sinkVec_validSink_24_bits_readSource;
  wire [2:0]   sinkVec_validSink_24_bits_offset;
  wire [2:0]   sinkVec_validSink_24_bits_instructionIndex;
  assign sinkVec_sinkWire_24_valid = sinkVec_queue_24_deq_valid;
  assign sinkVec_sinkWire_24_bits_vs = sinkVec_queue_24_deq_bits_vs;
  assign sinkVec_sinkWire_24_bits_readSource = sinkVec_queue_24_deq_bits_readSource;
  assign sinkVec_sinkWire_24_bits_offset = sinkVec_queue_24_deq_bits_offset;
  assign sinkVec_sinkWire_24_bits_instructionIndex = sinkVec_queue_24_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_queue_24_enq_bits_offset;
  wire [2:0]   sinkVec_queue_24_enq_bits_instructionIndex;
  wire [5:0]   sinkVec_queue_dataIn_lo_24 = {sinkVec_queue_24_enq_bits_offset, sinkVec_queue_24_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_24_enq_bits_vs;
  wire [1:0]   sinkVec_queue_24_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_24 = {sinkVec_queue_24_enq_bits_vs, sinkVec_queue_24_enq_bits_readSource};
  wire [12:0]  sinkVec_queue_dataIn_24 = {sinkVec_queue_dataIn_hi_24, sinkVec_queue_dataIn_lo_24};
  wire [2:0]   sinkVec_queue_dataOut_24_instructionIndex = _sinkVec_queue_fifo_24_data_out[2:0];
  wire [2:0]   sinkVec_queue_dataOut_24_offset = _sinkVec_queue_fifo_24_data_out[5:3];
  wire [1:0]   sinkVec_queue_dataOut_24_readSource = _sinkVec_queue_fifo_24_data_out[7:6];
  wire [4:0]   sinkVec_queue_dataOut_24_vs = _sinkVec_queue_fifo_24_data_out[12:8];
  wire         sinkVec_queue_24_enq_ready = ~_sinkVec_queue_fifo_24_full;
  wire         sinkVec_queue_24_enq_valid;
  assign sinkVec_queue_24_deq_valid = ~_sinkVec_queue_fifo_24_empty | sinkVec_queue_24_enq_valid;
  assign sinkVec_queue_24_deq_bits_vs = _sinkVec_queue_fifo_24_empty ? sinkVec_queue_24_enq_bits_vs : sinkVec_queue_dataOut_24_vs;
  assign sinkVec_queue_24_deq_bits_readSource = _sinkVec_queue_fifo_24_empty ? sinkVec_queue_24_enq_bits_readSource : sinkVec_queue_dataOut_24_readSource;
  assign sinkVec_queue_24_deq_bits_offset = _sinkVec_queue_fifo_24_empty ? sinkVec_queue_24_enq_bits_offset : sinkVec_queue_dataOut_24_offset;
  assign sinkVec_queue_24_deq_bits_instructionIndex = _sinkVec_queue_fifo_24_empty ? sinkVec_queue_24_enq_bits_instructionIndex : sinkVec_queue_dataOut_24_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_24;
  wire         sinkVec_releasePipe_pipe_out_24_valid = sinkVec_releasePipe_pipe_v_24;
  wire         x13_6_0_ready;
  wire         x13_6_0_valid;
  wire         sinkVec_validSource_24_valid = x13_6_0_ready & x13_6_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_24;
  wire [2:0]   sinkVec_tokenCheck_counterChange_24 = sinkVec_validSource_24_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_24 = ~(sinkVec_tokenCheck_counter_24[2]);
  assign x13_6_0_ready = sinkVec_tokenCheck_24;
  assign sinkVec_queue_24_enq_valid = sinkVec_validSink_24_valid;
  assign sinkVec_queue_24_enq_bits_vs = sinkVec_validSink_24_bits_vs;
  assign sinkVec_queue_24_enq_bits_readSource = sinkVec_validSink_24_bits_readSource;
  assign sinkVec_queue_24_enq_bits_offset = sinkVec_validSink_24_bits_offset;
  assign sinkVec_queue_24_enq_bits_instructionIndex = sinkVec_validSink_24_bits_instructionIndex;
  reg          sinkVec_shifterReg_24_0_valid;
  assign sinkVec_validSink_24_valid = sinkVec_shifterReg_24_0_valid;
  reg  [4:0]   sinkVec_shifterReg_24_0_bits_vs;
  assign sinkVec_validSink_24_bits_vs = sinkVec_shifterReg_24_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_24_0_bits_readSource;
  assign sinkVec_validSink_24_bits_readSource = sinkVec_shifterReg_24_0_bits_readSource;
  reg  [2:0]   sinkVec_shifterReg_24_0_bits_offset;
  assign sinkVec_validSink_24_bits_offset = sinkVec_shifterReg_24_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_24_0_bits_instructionIndex;
  assign sinkVec_validSink_24_bits_instructionIndex = sinkVec_shifterReg_24_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_24 = sinkVec_shifterReg_24_0_valid | sinkVec_validSource_24_valid;
  wire         sinkVec_12_1_ready;
  wire         sinkVec_queue_25_deq_ready = sinkVec_sinkWire_25_ready;
  wire         sinkVec_queue_25_deq_valid;
  wire [4:0]   sinkVec_queue_25_deq_bits_vs;
  wire         sinkVec_12_1_valid = sinkVec_sinkWire_25_valid;
  wire [1:0]   sinkVec_queue_25_deq_bits_readSource;
  wire [4:0]   sinkVec_12_1_bits_vs = sinkVec_sinkWire_25_bits_vs;
  wire [2:0]   sinkVec_queue_25_deq_bits_offset;
  wire [1:0]   sinkVec_12_1_bits_readSource = sinkVec_sinkWire_25_bits_readSource;
  wire [2:0]   sinkVec_queue_25_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_12_1_bits_offset = sinkVec_sinkWire_25_bits_offset;
  wire [2:0]   sinkVec_12_1_bits_instructionIndex = sinkVec_sinkWire_25_bits_instructionIndex;
  wire         sinkVec_validSink_25_valid;
  wire [4:0]   sinkVec_validSink_25_bits_vs;
  wire [1:0]   sinkVec_validSink_25_bits_readSource;
  wire [2:0]   sinkVec_validSink_25_bits_offset;
  wire [2:0]   sinkVec_validSink_25_bits_instructionIndex;
  assign sinkVec_sinkWire_25_valid = sinkVec_queue_25_deq_valid;
  assign sinkVec_sinkWire_25_bits_vs = sinkVec_queue_25_deq_bits_vs;
  assign sinkVec_sinkWire_25_bits_readSource = sinkVec_queue_25_deq_bits_readSource;
  assign sinkVec_sinkWire_25_bits_offset = sinkVec_queue_25_deq_bits_offset;
  assign sinkVec_sinkWire_25_bits_instructionIndex = sinkVec_queue_25_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_queue_25_enq_bits_offset;
  wire [2:0]   sinkVec_queue_25_enq_bits_instructionIndex;
  wire [5:0]   sinkVec_queue_dataIn_lo_25 = {sinkVec_queue_25_enq_bits_offset, sinkVec_queue_25_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_25_enq_bits_vs;
  wire [1:0]   sinkVec_queue_25_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_25 = {sinkVec_queue_25_enq_bits_vs, sinkVec_queue_25_enq_bits_readSource};
  wire [12:0]  sinkVec_queue_dataIn_25 = {sinkVec_queue_dataIn_hi_25, sinkVec_queue_dataIn_lo_25};
  wire [2:0]   sinkVec_queue_dataOut_25_instructionIndex = _sinkVec_queue_fifo_25_data_out[2:0];
  wire [2:0]   sinkVec_queue_dataOut_25_offset = _sinkVec_queue_fifo_25_data_out[5:3];
  wire [1:0]   sinkVec_queue_dataOut_25_readSource = _sinkVec_queue_fifo_25_data_out[7:6];
  wire [4:0]   sinkVec_queue_dataOut_25_vs = _sinkVec_queue_fifo_25_data_out[12:8];
  wire         sinkVec_queue_25_enq_ready = ~_sinkVec_queue_fifo_25_full;
  wire         sinkVec_queue_25_enq_valid;
  assign sinkVec_queue_25_deq_valid = ~_sinkVec_queue_fifo_25_empty | sinkVec_queue_25_enq_valid;
  assign sinkVec_queue_25_deq_bits_vs = _sinkVec_queue_fifo_25_empty ? sinkVec_queue_25_enq_bits_vs : sinkVec_queue_dataOut_25_vs;
  assign sinkVec_queue_25_deq_bits_readSource = _sinkVec_queue_fifo_25_empty ? sinkVec_queue_25_enq_bits_readSource : sinkVec_queue_dataOut_25_readSource;
  assign sinkVec_queue_25_deq_bits_offset = _sinkVec_queue_fifo_25_empty ? sinkVec_queue_25_enq_bits_offset : sinkVec_queue_dataOut_25_offset;
  assign sinkVec_queue_25_deq_bits_instructionIndex = _sinkVec_queue_fifo_25_empty ? sinkVec_queue_25_enq_bits_instructionIndex : sinkVec_queue_dataOut_25_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_25;
  wire         sinkVec_releasePipe_pipe_out_25_valid = sinkVec_releasePipe_pipe_v_25;
  wire         x13_6_1_ready;
  wire         x13_6_1_valid;
  wire         sinkVec_validSource_25_valid = x13_6_1_ready & x13_6_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_25;
  wire [2:0]   sinkVec_tokenCheck_counterChange_25 = sinkVec_validSource_25_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_25 = ~(sinkVec_tokenCheck_counter_25[2]);
  assign x13_6_1_ready = sinkVec_tokenCheck_25;
  assign sinkVec_queue_25_enq_valid = sinkVec_validSink_25_valid;
  assign sinkVec_queue_25_enq_bits_vs = sinkVec_validSink_25_bits_vs;
  assign sinkVec_queue_25_enq_bits_readSource = sinkVec_validSink_25_bits_readSource;
  assign sinkVec_queue_25_enq_bits_offset = sinkVec_validSink_25_bits_offset;
  assign sinkVec_queue_25_enq_bits_instructionIndex = sinkVec_validSink_25_bits_instructionIndex;
  reg          sinkVec_shifterReg_25_0_valid;
  assign sinkVec_validSink_25_valid = sinkVec_shifterReg_25_0_valid;
  reg  [4:0]   sinkVec_shifterReg_25_0_bits_vs;
  assign sinkVec_validSink_25_bits_vs = sinkVec_shifterReg_25_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_25_0_bits_readSource;
  assign sinkVec_validSink_25_bits_readSource = sinkVec_shifterReg_25_0_bits_readSource;
  reg  [2:0]   sinkVec_shifterReg_25_0_bits_offset;
  assign sinkVec_validSink_25_bits_offset = sinkVec_shifterReg_25_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_25_0_bits_instructionIndex;
  assign sinkVec_validSink_25_bits_instructionIndex = sinkVec_shifterReg_25_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_25 = sinkVec_shifterReg_25_0_valid | sinkVec_validSource_25_valid;
  assign sinkVec_sinkWire_24_ready = sinkVec_12_0_ready;
  assign sinkVec_sinkWire_25_ready = sinkVec_12_1_ready;
  reg          maskUnitFirst_12;
  wire         tryToRead_12 = sinkVec_12_0_valid | sinkVec_12_1_valid;
  wire         sinkWire_12_valid = maskUnitFirst_12 ? sinkVec_12_0_valid : sinkVec_12_1_valid;
  wire [4:0]   sinkWire_12_bits_vs = maskUnitFirst_12 ? sinkVec_12_0_bits_vs : sinkVec_12_1_bits_vs;
  wire [1:0]   sinkWire_12_bits_readSource = maskUnitFirst_12 ? sinkVec_12_0_bits_readSource : sinkVec_12_1_bits_readSource;
  wire [2:0]   sinkWire_12_bits_offset = maskUnitFirst_12 ? sinkVec_12_0_bits_offset : sinkVec_12_1_bits_offset;
  wire [2:0]   sinkWire_12_bits_instructionIndex = maskUnitFirst_12 ? sinkVec_12_0_bits_instructionIndex : sinkVec_12_1_bits_instructionIndex;
  wire         sinkWire_12_ready;
  assign sinkVec_12_1_ready = sinkWire_12_ready & ~maskUnitFirst_12;
  assign sinkVec_12_0_ready = sinkWire_12_ready & maskUnitFirst_12;
  reg          accessDataValid_pipe_v_12;
  reg          accessDataValid_pipe_pipe_v_12;
  wire         accessDataValid_pipe_pipe_out_12_valid = accessDataValid_pipe_pipe_v_12;
  wire         accessDataSource_12_valid = accessDataValid_pipe_pipe_out_12_valid;
  reg          shifterReg_20_0_valid;
  reg  [31:0]  shifterReg_20_0_bits;
  wire         shifterValid_20 = shifterReg_20_0_valid | accessDataSource_12_valid;
  reg          accessDataValid_pipe_v_13;
  reg          accessDataValid_pipe_pipe_v_13;
  wire         accessDataValid_pipe_pipe_out_13_valid = accessDataValid_pipe_pipe_v_13;
  wire         accessDataSource_13_valid = accessDataValid_pipe_pipe_out_13_valid;
  reg          shifterReg_21_0_valid;
  reg  [31:0]  shifterReg_21_0_bits;
  wire         shifterValid_21 = shifterReg_21_0_valid | accessDataSource_13_valid;
  wire         sinkVec_tokenCheck_26;
  wire [4:0]   sinkVec_validSource_26_bits_vd = x22_6_0_bits_vd;
  wire [2:0]   sinkVec_validSource_26_bits_offset = x22_6_0_bits_offset;
  wire [3:0]   sinkVec_validSource_26_bits_mask = x22_6_0_bits_mask;
  wire [31:0]  sinkVec_validSource_26_bits_data = x22_6_0_bits_data;
  wire [2:0]   sinkVec_validSource_26_bits_instructionIndex = x22_6_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_27;
  wire [4:0]   sinkVec_validSource_27_bits_vd = x22_6_1_bits_vd;
  wire [2:0]   sinkVec_validSource_27_bits_offset = x22_6_1_bits_offset;
  wire [3:0]   sinkVec_validSource_27_bits_mask = x22_6_1_bits_mask;
  wire [31:0]  sinkVec_validSource_27_bits_data = x22_6_1_bits_data;
  wire         sinkVec_validSource_27_bits_last = x22_6_1_bits_last;
  wire [2:0]   sinkVec_validSource_27_bits_instructionIndex = x22_6_1_bits_instructionIndex;
  wire         sinkVec_13_0_ready;
  wire         sinkVec_queue_26_deq_ready = sinkVec_sinkWire_26_ready;
  wire         sinkVec_queue_26_deq_valid;
  wire [4:0]   sinkVec_queue_26_deq_bits_vd;
  wire         sinkVec_13_0_valid = sinkVec_sinkWire_26_valid;
  wire [2:0]   sinkVec_queue_26_deq_bits_offset;
  wire [4:0]   sinkVec_13_0_bits_vd = sinkVec_sinkWire_26_bits_vd;
  wire [3:0]   sinkVec_queue_26_deq_bits_mask;
  wire [2:0]   sinkVec_13_0_bits_offset = sinkVec_sinkWire_26_bits_offset;
  wire [31:0]  sinkVec_queue_26_deq_bits_data;
  wire [3:0]   sinkVec_13_0_bits_mask = sinkVec_sinkWire_26_bits_mask;
  wire         sinkVec_queue_26_deq_bits_last;
  wire [31:0]  sinkVec_13_0_bits_data = sinkVec_sinkWire_26_bits_data;
  wire [2:0]   sinkVec_queue_26_deq_bits_instructionIndex;
  wire         sinkVec_13_0_bits_last = sinkVec_sinkWire_26_bits_last;
  wire [2:0]   sinkVec_13_0_bits_instructionIndex = sinkVec_sinkWire_26_bits_instructionIndex;
  wire         sinkVec_validSink_26_valid;
  wire [4:0]   sinkVec_validSink_26_bits_vd;
  wire [2:0]   sinkVec_validSink_26_bits_offset;
  wire [3:0]   sinkVec_validSink_26_bits_mask;
  wire [31:0]  sinkVec_validSink_26_bits_data;
  wire [2:0]   sinkVec_validSink_26_bits_instructionIndex;
  assign sinkVec_sinkWire_26_valid = sinkVec_queue_26_deq_valid;
  assign sinkVec_sinkWire_26_bits_vd = sinkVec_queue_26_deq_bits_vd;
  assign sinkVec_sinkWire_26_bits_offset = sinkVec_queue_26_deq_bits_offset;
  assign sinkVec_sinkWire_26_bits_mask = sinkVec_queue_26_deq_bits_mask;
  assign sinkVec_sinkWire_26_bits_data = sinkVec_queue_26_deq_bits_data;
  assign sinkVec_sinkWire_26_bits_last = sinkVec_queue_26_deq_bits_last;
  assign sinkVec_sinkWire_26_bits_instructionIndex = sinkVec_queue_26_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_26_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_12 = {sinkVec_queue_26_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_26_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_26 = {sinkVec_queue_dataIn_lo_hi_12, sinkVec_queue_26_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_26_enq_bits_vd;
  wire [2:0]   sinkVec_queue_26_enq_bits_offset;
  wire [7:0]   sinkVec_queue_dataIn_hi_hi_12 = {sinkVec_queue_26_enq_bits_vd, sinkVec_queue_26_enq_bits_offset};
  wire [3:0]   sinkVec_queue_26_enq_bits_mask;
  wire [11:0]  sinkVec_queue_dataIn_hi_26 = {sinkVec_queue_dataIn_hi_hi_12, sinkVec_queue_26_enq_bits_mask};
  wire [47:0]  sinkVec_queue_dataIn_26 = {sinkVec_queue_dataIn_hi_26, sinkVec_queue_dataIn_lo_26};
  wire [2:0]   sinkVec_queue_dataOut_26_instructionIndex = _sinkVec_queue_fifo_26_data_out[2:0];
  wire         sinkVec_queue_dataOut_26_last = _sinkVec_queue_fifo_26_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_26_data = _sinkVec_queue_fifo_26_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_26_mask = _sinkVec_queue_fifo_26_data_out[39:36];
  wire [2:0]   sinkVec_queue_dataOut_26_offset = _sinkVec_queue_fifo_26_data_out[42:40];
  wire [4:0]   sinkVec_queue_dataOut_26_vd = _sinkVec_queue_fifo_26_data_out[47:43];
  wire         sinkVec_queue_26_enq_ready = ~_sinkVec_queue_fifo_26_full;
  wire         sinkVec_queue_26_enq_valid;
  assign sinkVec_queue_26_deq_valid = ~_sinkVec_queue_fifo_26_empty | sinkVec_queue_26_enq_valid;
  assign sinkVec_queue_26_deq_bits_vd = _sinkVec_queue_fifo_26_empty ? sinkVec_queue_26_enq_bits_vd : sinkVec_queue_dataOut_26_vd;
  assign sinkVec_queue_26_deq_bits_offset = _sinkVec_queue_fifo_26_empty ? sinkVec_queue_26_enq_bits_offset : sinkVec_queue_dataOut_26_offset;
  assign sinkVec_queue_26_deq_bits_mask = _sinkVec_queue_fifo_26_empty ? sinkVec_queue_26_enq_bits_mask : sinkVec_queue_dataOut_26_mask;
  assign sinkVec_queue_26_deq_bits_data = _sinkVec_queue_fifo_26_empty ? sinkVec_queue_26_enq_bits_data : sinkVec_queue_dataOut_26_data;
  assign sinkVec_queue_26_deq_bits_last = ~_sinkVec_queue_fifo_26_empty & sinkVec_queue_dataOut_26_last;
  assign sinkVec_queue_26_deq_bits_instructionIndex = _sinkVec_queue_fifo_26_empty ? sinkVec_queue_26_enq_bits_instructionIndex : sinkVec_queue_dataOut_26_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_26;
  wire         sinkVec_releasePipe_pipe_out_26_valid = sinkVec_releasePipe_pipe_v_26;
  wire         x22_6_0_ready;
  wire         x22_6_0_valid;
  wire         sinkVec_validSource_26_valid = x22_6_0_ready & x22_6_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_26;
  wire [2:0]   sinkVec_tokenCheck_counterChange_26 = sinkVec_validSource_26_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_26 = ~(sinkVec_tokenCheck_counter_26[2]);
  assign x22_6_0_ready = sinkVec_tokenCheck_26;
  assign sinkVec_queue_26_enq_valid = sinkVec_validSink_26_valid;
  assign sinkVec_queue_26_enq_bits_vd = sinkVec_validSink_26_bits_vd;
  assign sinkVec_queue_26_enq_bits_offset = sinkVec_validSink_26_bits_offset;
  assign sinkVec_queue_26_enq_bits_mask = sinkVec_validSink_26_bits_mask;
  assign sinkVec_queue_26_enq_bits_data = sinkVec_validSink_26_bits_data;
  assign sinkVec_queue_26_enq_bits_instructionIndex = sinkVec_validSink_26_bits_instructionIndex;
  reg          sinkVec_shifterReg_26_0_valid;
  assign sinkVec_validSink_26_valid = sinkVec_shifterReg_26_0_valid;
  reg  [4:0]   sinkVec_shifterReg_26_0_bits_vd;
  assign sinkVec_validSink_26_bits_vd = sinkVec_shifterReg_26_0_bits_vd;
  reg  [2:0]   sinkVec_shifterReg_26_0_bits_offset;
  assign sinkVec_validSink_26_bits_offset = sinkVec_shifterReg_26_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_26_0_bits_mask;
  assign sinkVec_validSink_26_bits_mask = sinkVec_shifterReg_26_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_26_0_bits_data;
  assign sinkVec_validSink_26_bits_data = sinkVec_shifterReg_26_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_26_0_bits_instructionIndex;
  assign sinkVec_validSink_26_bits_instructionIndex = sinkVec_shifterReg_26_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_26 = sinkVec_shifterReg_26_0_valid | sinkVec_validSource_26_valid;
  wire         sinkVec_13_1_ready;
  wire         sinkVec_queue_27_deq_ready = sinkVec_sinkWire_27_ready;
  wire         sinkVec_queue_27_deq_valid;
  wire [4:0]   sinkVec_queue_27_deq_bits_vd;
  wire         sinkVec_13_1_valid = sinkVec_sinkWire_27_valid;
  wire [2:0]   sinkVec_queue_27_deq_bits_offset;
  wire [4:0]   sinkVec_13_1_bits_vd = sinkVec_sinkWire_27_bits_vd;
  wire [3:0]   sinkVec_queue_27_deq_bits_mask;
  wire [2:0]   sinkVec_13_1_bits_offset = sinkVec_sinkWire_27_bits_offset;
  wire [31:0]  sinkVec_queue_27_deq_bits_data;
  wire [3:0]   sinkVec_13_1_bits_mask = sinkVec_sinkWire_27_bits_mask;
  wire         sinkVec_queue_27_deq_bits_last;
  wire [31:0]  sinkVec_13_1_bits_data = sinkVec_sinkWire_27_bits_data;
  wire [2:0]   sinkVec_queue_27_deq_bits_instructionIndex;
  wire         sinkVec_13_1_bits_last = sinkVec_sinkWire_27_bits_last;
  wire [2:0]   sinkVec_13_1_bits_instructionIndex = sinkVec_sinkWire_27_bits_instructionIndex;
  wire         sinkVec_validSink_27_valid;
  wire [4:0]   sinkVec_validSink_27_bits_vd;
  wire [2:0]   sinkVec_validSink_27_bits_offset;
  wire [3:0]   sinkVec_validSink_27_bits_mask;
  wire [31:0]  sinkVec_validSink_27_bits_data;
  wire         sinkVec_validSink_27_bits_last;
  wire [2:0]   sinkVec_validSink_27_bits_instructionIndex;
  assign sinkVec_sinkWire_27_valid = sinkVec_queue_27_deq_valid;
  assign sinkVec_sinkWire_27_bits_vd = sinkVec_queue_27_deq_bits_vd;
  assign sinkVec_sinkWire_27_bits_offset = sinkVec_queue_27_deq_bits_offset;
  assign sinkVec_sinkWire_27_bits_mask = sinkVec_queue_27_deq_bits_mask;
  assign sinkVec_sinkWire_27_bits_data = sinkVec_queue_27_deq_bits_data;
  assign sinkVec_sinkWire_27_bits_last = sinkVec_queue_27_deq_bits_last;
  assign sinkVec_sinkWire_27_bits_instructionIndex = sinkVec_queue_27_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_27_enq_bits_data;
  wire         sinkVec_queue_27_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_13 = {sinkVec_queue_27_enq_bits_data, sinkVec_queue_27_enq_bits_last};
  wire [2:0]   sinkVec_queue_27_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_27 = {sinkVec_queue_dataIn_lo_hi_13, sinkVec_queue_27_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_27_enq_bits_vd;
  wire [2:0]   sinkVec_queue_27_enq_bits_offset;
  wire [7:0]   sinkVec_queue_dataIn_hi_hi_13 = {sinkVec_queue_27_enq_bits_vd, sinkVec_queue_27_enq_bits_offset};
  wire [3:0]   sinkVec_queue_27_enq_bits_mask;
  wire [11:0]  sinkVec_queue_dataIn_hi_27 = {sinkVec_queue_dataIn_hi_hi_13, sinkVec_queue_27_enq_bits_mask};
  wire [47:0]  sinkVec_queue_dataIn_27 = {sinkVec_queue_dataIn_hi_27, sinkVec_queue_dataIn_lo_27};
  wire [2:0]   sinkVec_queue_dataOut_27_instructionIndex = _sinkVec_queue_fifo_27_data_out[2:0];
  wire         sinkVec_queue_dataOut_27_last = _sinkVec_queue_fifo_27_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_27_data = _sinkVec_queue_fifo_27_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_27_mask = _sinkVec_queue_fifo_27_data_out[39:36];
  wire [2:0]   sinkVec_queue_dataOut_27_offset = _sinkVec_queue_fifo_27_data_out[42:40];
  wire [4:0]   sinkVec_queue_dataOut_27_vd = _sinkVec_queue_fifo_27_data_out[47:43];
  wire         sinkVec_queue_27_enq_ready = ~_sinkVec_queue_fifo_27_full;
  wire         sinkVec_queue_27_enq_valid;
  assign sinkVec_queue_27_deq_valid = ~_sinkVec_queue_fifo_27_empty | sinkVec_queue_27_enq_valid;
  assign sinkVec_queue_27_deq_bits_vd = _sinkVec_queue_fifo_27_empty ? sinkVec_queue_27_enq_bits_vd : sinkVec_queue_dataOut_27_vd;
  assign sinkVec_queue_27_deq_bits_offset = _sinkVec_queue_fifo_27_empty ? sinkVec_queue_27_enq_bits_offset : sinkVec_queue_dataOut_27_offset;
  assign sinkVec_queue_27_deq_bits_mask = _sinkVec_queue_fifo_27_empty ? sinkVec_queue_27_enq_bits_mask : sinkVec_queue_dataOut_27_mask;
  assign sinkVec_queue_27_deq_bits_data = _sinkVec_queue_fifo_27_empty ? sinkVec_queue_27_enq_bits_data : sinkVec_queue_dataOut_27_data;
  assign sinkVec_queue_27_deq_bits_last = _sinkVec_queue_fifo_27_empty ? sinkVec_queue_27_enq_bits_last : sinkVec_queue_dataOut_27_last;
  assign sinkVec_queue_27_deq_bits_instructionIndex = _sinkVec_queue_fifo_27_empty ? sinkVec_queue_27_enq_bits_instructionIndex : sinkVec_queue_dataOut_27_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_27;
  wire         sinkVec_releasePipe_pipe_out_27_valid = sinkVec_releasePipe_pipe_v_27;
  wire         x22_6_1_ready;
  wire         x22_6_1_valid;
  wire         sinkVec_validSource_27_valid = x22_6_1_ready & x22_6_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_27;
  wire [2:0]   sinkVec_tokenCheck_counterChange_27 = sinkVec_validSource_27_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_27 = ~(sinkVec_tokenCheck_counter_27[2]);
  assign x22_6_1_ready = sinkVec_tokenCheck_27;
  assign sinkVec_queue_27_enq_valid = sinkVec_validSink_27_valid;
  assign sinkVec_queue_27_enq_bits_vd = sinkVec_validSink_27_bits_vd;
  assign sinkVec_queue_27_enq_bits_offset = sinkVec_validSink_27_bits_offset;
  assign sinkVec_queue_27_enq_bits_mask = sinkVec_validSink_27_bits_mask;
  assign sinkVec_queue_27_enq_bits_data = sinkVec_validSink_27_bits_data;
  assign sinkVec_queue_27_enq_bits_last = sinkVec_validSink_27_bits_last;
  assign sinkVec_queue_27_enq_bits_instructionIndex = sinkVec_validSink_27_bits_instructionIndex;
  reg          sinkVec_shifterReg_27_0_valid;
  assign sinkVec_validSink_27_valid = sinkVec_shifterReg_27_0_valid;
  reg  [4:0]   sinkVec_shifterReg_27_0_bits_vd;
  assign sinkVec_validSink_27_bits_vd = sinkVec_shifterReg_27_0_bits_vd;
  reg  [2:0]   sinkVec_shifterReg_27_0_bits_offset;
  assign sinkVec_validSink_27_bits_offset = sinkVec_shifterReg_27_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_27_0_bits_mask;
  assign sinkVec_validSink_27_bits_mask = sinkVec_shifterReg_27_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_27_0_bits_data;
  assign sinkVec_validSink_27_bits_data = sinkVec_shifterReg_27_0_bits_data;
  reg          sinkVec_shifterReg_27_0_bits_last;
  assign sinkVec_validSink_27_bits_last = sinkVec_shifterReg_27_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_27_0_bits_instructionIndex;
  assign sinkVec_validSink_27_bits_instructionIndex = sinkVec_shifterReg_27_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_27 = sinkVec_shifterReg_27_0_valid | sinkVec_validSource_27_valid;
  assign sinkVec_sinkWire_26_ready = sinkVec_13_0_ready;
  assign sinkVec_sinkWire_27_ready = sinkVec_13_1_ready;
  reg          maskUnitFirst_13;
  wire         tryToRead_13 = sinkVec_13_0_valid | sinkVec_13_1_valid;
  wire         sinkWire_13_valid = maskUnitFirst_13 ? sinkVec_13_0_valid : sinkVec_13_1_valid;
  wire [4:0]   sinkWire_13_bits_vd = maskUnitFirst_13 ? sinkVec_13_0_bits_vd : sinkVec_13_1_bits_vd;
  wire [2:0]   sinkWire_13_bits_offset = maskUnitFirst_13 ? sinkVec_13_0_bits_offset : sinkVec_13_1_bits_offset;
  wire [3:0]   sinkWire_13_bits_mask = maskUnitFirst_13 ? sinkVec_13_0_bits_mask : sinkVec_13_1_bits_mask;
  wire [31:0]  sinkWire_13_bits_data = maskUnitFirst_13 ? sinkVec_13_0_bits_data : sinkVec_13_1_bits_data;
  wire         sinkWire_13_bits_last = maskUnitFirst_13 ? sinkVec_13_0_bits_last : sinkVec_13_1_bits_last;
  wire [2:0]   sinkWire_13_bits_instructionIndex = maskUnitFirst_13 ? sinkVec_13_0_bits_instructionIndex : sinkVec_13_1_bits_instructionIndex;
  wire         sinkWire_13_ready;
  assign sinkVec_13_1_ready = sinkWire_13_ready & ~maskUnitFirst_13;
  assign sinkVec_13_0_ready = sinkWire_13_ready & maskUnitFirst_13;
  reg          view__writeRelease_6_pipe_v;
  wire         view__writeRelease_6_pipe_out_valid = view__writeRelease_6_pipe_v;
  reg          pipe_v_18;
  wire         pipe_out_12_valid = pipe_v_18;
  wire         _probeWire_writeQueueEnqVec_6_valid_T = x22_6_0_ready & _maskUnit_exeResp_6_valid;
  reg          instructionFinishedPipe_pipe_v_6;
  wire         instructionFinishedPipe_pipe_out_6_valid = instructionFinishedPipe_pipe_v_6;
  reg  [7:0]   instructionFinishedPipe_pipe_b_6;
  wire [7:0]   instructionFinishedPipe_pipe_out_6_bits = instructionFinishedPipe_pipe_b_6;
  wire         instructionFinished_6_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_6_bits);
  wire         instructionFinished_6_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_6_bits);
  wire         instructionFinished_6_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_6_bits);
  wire         instructionFinished_6_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_6_bits);
  assign vxsatReportVec_6 = _laneVec_6_vxsatReport[3:0];
  reg          pipe_v_19;
  reg  [31:0]  pipe_b_19;
  reg          pipe_pipe_v_6;
  wire         pipe_pipe_out_6_valid = pipe_pipe_v_6;
  reg  [31:0]  pipe_pipe_b_6;
  wire [31:0]  pipe_pipe_out_6_bits = pipe_pipe_b_6;
  reg          view__laneMaskSelect_6_pipe_v;
  reg  [5:0]   view__laneMaskSelect_6_pipe_b;
  reg          view__laneMaskSelect_6_pipe_pipe_v;
  wire         view__laneMaskSelect_6_pipe_pipe_out_valid = view__laneMaskSelect_6_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_6_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_6_pipe_pipe_out_bits = view__laneMaskSelect_6_pipe_pipe_b;
  reg          view__laneMaskSewSelect_6_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_6_pipe_b;
  reg          view__laneMaskSewSelect_6_pipe_pipe_v;
  wire         view__laneMaskSewSelect_6_pipe_pipe_out_valid = view__laneMaskSewSelect_6_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_6_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_6_pipe_pipe_out_bits = view__laneMaskSewSelect_6_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v_6;
  wire         lsuLastPipe_pipe_out_6_valid = lsuLastPipe_pipe_v_6;
  reg  [7:0]   lsuLastPipe_pipe_b_6;
  wire [7:0]   lsuLastPipe_pipe_out_6_bits = lsuLastPipe_pipe_b_6;
  reg          maskLastPipe_pipe_v_6;
  wire         maskLastPipe_pipe_out_6_valid = maskLastPipe_pipe_v_6;
  reg  [7:0]   maskLastPipe_pipe_b_6;
  wire [7:0]   maskLastPipe_pipe_out_6_bits = maskLastPipe_pipe_b_6;
  wire [6:0]   writeCounter_6 = requestReg_bits_writeByte[11:5] + {6'h0, requestReg_bits_writeByte[4:0] > 5'h18};
  reg          pipe_v_20;
  wire         pipe_out_13_valid = pipe_v_20;
  reg  [6:0]   pipe_b_20;
  wire [6:0]   pipe_out_13_bits = pipe_b_20;
  assign laneRequestSinkWire_7_ready = ~laneRequestSinkWire_7_bits_issueInst | _laneVec_7_laneRequest_ready;
  wire         sinkVec_tokenCheck_28;
  wire [4:0]   sinkVec_validSource_28_bits_vs = x13_7_0_bits_vs;
  wire [2:0]   sinkVec_validSource_28_bits_offset = x13_7_0_bits_offset;
  wire [2:0]   sinkVec_validSource_28_bits_instructionIndex = x13_7_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_29;
  wire [4:0]   sinkVec_validSource_29_bits_vs = x13_7_1_bits_vs;
  wire [2:0]   sinkVec_validSource_29_bits_offset = x13_7_1_bits_offset;
  wire [2:0]   sinkVec_validSource_29_bits_instructionIndex = x13_7_1_bits_instructionIndex;
  wire         sinkVec_14_0_ready;
  wire         sinkVec_queue_28_deq_ready = sinkVec_sinkWire_28_ready;
  wire         sinkVec_queue_28_deq_valid;
  wire [4:0]   sinkVec_queue_28_deq_bits_vs;
  wire         sinkVec_14_0_valid = sinkVec_sinkWire_28_valid;
  wire [1:0]   sinkVec_queue_28_deq_bits_readSource;
  wire [4:0]   sinkVec_14_0_bits_vs = sinkVec_sinkWire_28_bits_vs;
  wire [2:0]   sinkVec_queue_28_deq_bits_offset;
  wire [1:0]   sinkVec_14_0_bits_readSource = sinkVec_sinkWire_28_bits_readSource;
  wire [2:0]   sinkVec_queue_28_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_14_0_bits_offset = sinkVec_sinkWire_28_bits_offset;
  wire [2:0]   sinkVec_14_0_bits_instructionIndex = sinkVec_sinkWire_28_bits_instructionIndex;
  wire         sinkVec_validSink_28_valid;
  wire [4:0]   sinkVec_validSink_28_bits_vs;
  wire [1:0]   sinkVec_validSink_28_bits_readSource;
  wire [2:0]   sinkVec_validSink_28_bits_offset;
  wire [2:0]   sinkVec_validSink_28_bits_instructionIndex;
  assign sinkVec_sinkWire_28_valid = sinkVec_queue_28_deq_valid;
  assign sinkVec_sinkWire_28_bits_vs = sinkVec_queue_28_deq_bits_vs;
  assign sinkVec_sinkWire_28_bits_readSource = sinkVec_queue_28_deq_bits_readSource;
  assign sinkVec_sinkWire_28_bits_offset = sinkVec_queue_28_deq_bits_offset;
  assign sinkVec_sinkWire_28_bits_instructionIndex = sinkVec_queue_28_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_queue_28_enq_bits_offset;
  wire [2:0]   sinkVec_queue_28_enq_bits_instructionIndex;
  wire [5:0]   sinkVec_queue_dataIn_lo_28 = {sinkVec_queue_28_enq_bits_offset, sinkVec_queue_28_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_28_enq_bits_vs;
  wire [1:0]   sinkVec_queue_28_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_28 = {sinkVec_queue_28_enq_bits_vs, sinkVec_queue_28_enq_bits_readSource};
  wire [12:0]  sinkVec_queue_dataIn_28 = {sinkVec_queue_dataIn_hi_28, sinkVec_queue_dataIn_lo_28};
  wire [2:0]   sinkVec_queue_dataOut_28_instructionIndex = _sinkVec_queue_fifo_28_data_out[2:0];
  wire [2:0]   sinkVec_queue_dataOut_28_offset = _sinkVec_queue_fifo_28_data_out[5:3];
  wire [1:0]   sinkVec_queue_dataOut_28_readSource = _sinkVec_queue_fifo_28_data_out[7:6];
  wire [4:0]   sinkVec_queue_dataOut_28_vs = _sinkVec_queue_fifo_28_data_out[12:8];
  wire         sinkVec_queue_28_enq_ready = ~_sinkVec_queue_fifo_28_full;
  wire         sinkVec_queue_28_enq_valid;
  assign sinkVec_queue_28_deq_valid = ~_sinkVec_queue_fifo_28_empty | sinkVec_queue_28_enq_valid;
  assign sinkVec_queue_28_deq_bits_vs = _sinkVec_queue_fifo_28_empty ? sinkVec_queue_28_enq_bits_vs : sinkVec_queue_dataOut_28_vs;
  assign sinkVec_queue_28_deq_bits_readSource = _sinkVec_queue_fifo_28_empty ? sinkVec_queue_28_enq_bits_readSource : sinkVec_queue_dataOut_28_readSource;
  assign sinkVec_queue_28_deq_bits_offset = _sinkVec_queue_fifo_28_empty ? sinkVec_queue_28_enq_bits_offset : sinkVec_queue_dataOut_28_offset;
  assign sinkVec_queue_28_deq_bits_instructionIndex = _sinkVec_queue_fifo_28_empty ? sinkVec_queue_28_enq_bits_instructionIndex : sinkVec_queue_dataOut_28_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_28;
  wire         sinkVec_releasePipe_pipe_out_28_valid = sinkVec_releasePipe_pipe_v_28;
  wire         x13_7_0_ready;
  wire         x13_7_0_valid;
  wire         sinkVec_validSource_28_valid = x13_7_0_ready & x13_7_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_28;
  wire [2:0]   sinkVec_tokenCheck_counterChange_28 = sinkVec_validSource_28_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_28 = ~(sinkVec_tokenCheck_counter_28[2]);
  assign x13_7_0_ready = sinkVec_tokenCheck_28;
  assign sinkVec_queue_28_enq_valid = sinkVec_validSink_28_valid;
  assign sinkVec_queue_28_enq_bits_vs = sinkVec_validSink_28_bits_vs;
  assign sinkVec_queue_28_enq_bits_readSource = sinkVec_validSink_28_bits_readSource;
  assign sinkVec_queue_28_enq_bits_offset = sinkVec_validSink_28_bits_offset;
  assign sinkVec_queue_28_enq_bits_instructionIndex = sinkVec_validSink_28_bits_instructionIndex;
  reg          sinkVec_shifterReg_28_0_valid;
  assign sinkVec_validSink_28_valid = sinkVec_shifterReg_28_0_valid;
  reg  [4:0]   sinkVec_shifterReg_28_0_bits_vs;
  assign sinkVec_validSink_28_bits_vs = sinkVec_shifterReg_28_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_28_0_bits_readSource;
  assign sinkVec_validSink_28_bits_readSource = sinkVec_shifterReg_28_0_bits_readSource;
  reg  [2:0]   sinkVec_shifterReg_28_0_bits_offset;
  assign sinkVec_validSink_28_bits_offset = sinkVec_shifterReg_28_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_28_0_bits_instructionIndex;
  assign sinkVec_validSink_28_bits_instructionIndex = sinkVec_shifterReg_28_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_28 = sinkVec_shifterReg_28_0_valid | sinkVec_validSource_28_valid;
  wire         sinkVec_14_1_ready;
  wire         sinkVec_queue_29_deq_ready = sinkVec_sinkWire_29_ready;
  wire         sinkVec_queue_29_deq_valid;
  wire [4:0]   sinkVec_queue_29_deq_bits_vs;
  wire         sinkVec_14_1_valid = sinkVec_sinkWire_29_valid;
  wire [1:0]   sinkVec_queue_29_deq_bits_readSource;
  wire [4:0]   sinkVec_14_1_bits_vs = sinkVec_sinkWire_29_bits_vs;
  wire [2:0]   sinkVec_queue_29_deq_bits_offset;
  wire [1:0]   sinkVec_14_1_bits_readSource = sinkVec_sinkWire_29_bits_readSource;
  wire [2:0]   sinkVec_queue_29_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_14_1_bits_offset = sinkVec_sinkWire_29_bits_offset;
  wire [2:0]   sinkVec_14_1_bits_instructionIndex = sinkVec_sinkWire_29_bits_instructionIndex;
  wire         sinkVec_validSink_29_valid;
  wire [4:0]   sinkVec_validSink_29_bits_vs;
  wire [1:0]   sinkVec_validSink_29_bits_readSource;
  wire [2:0]   sinkVec_validSink_29_bits_offset;
  wire [2:0]   sinkVec_validSink_29_bits_instructionIndex;
  assign sinkVec_sinkWire_29_valid = sinkVec_queue_29_deq_valid;
  assign sinkVec_sinkWire_29_bits_vs = sinkVec_queue_29_deq_bits_vs;
  assign sinkVec_sinkWire_29_bits_readSource = sinkVec_queue_29_deq_bits_readSource;
  assign sinkVec_sinkWire_29_bits_offset = sinkVec_queue_29_deq_bits_offset;
  assign sinkVec_sinkWire_29_bits_instructionIndex = sinkVec_queue_29_deq_bits_instructionIndex;
  wire [2:0]   sinkVec_queue_29_enq_bits_offset;
  wire [2:0]   sinkVec_queue_29_enq_bits_instructionIndex;
  wire [5:0]   sinkVec_queue_dataIn_lo_29 = {sinkVec_queue_29_enq_bits_offset, sinkVec_queue_29_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_29_enq_bits_vs;
  wire [1:0]   sinkVec_queue_29_enq_bits_readSource;
  wire [6:0]   sinkVec_queue_dataIn_hi_29 = {sinkVec_queue_29_enq_bits_vs, sinkVec_queue_29_enq_bits_readSource};
  wire [12:0]  sinkVec_queue_dataIn_29 = {sinkVec_queue_dataIn_hi_29, sinkVec_queue_dataIn_lo_29};
  wire [2:0]   sinkVec_queue_dataOut_29_instructionIndex = _sinkVec_queue_fifo_29_data_out[2:0];
  wire [2:0]   sinkVec_queue_dataOut_29_offset = _sinkVec_queue_fifo_29_data_out[5:3];
  wire [1:0]   sinkVec_queue_dataOut_29_readSource = _sinkVec_queue_fifo_29_data_out[7:6];
  wire [4:0]   sinkVec_queue_dataOut_29_vs = _sinkVec_queue_fifo_29_data_out[12:8];
  wire         sinkVec_queue_29_enq_ready = ~_sinkVec_queue_fifo_29_full;
  wire         sinkVec_queue_29_enq_valid;
  assign sinkVec_queue_29_deq_valid = ~_sinkVec_queue_fifo_29_empty | sinkVec_queue_29_enq_valid;
  assign sinkVec_queue_29_deq_bits_vs = _sinkVec_queue_fifo_29_empty ? sinkVec_queue_29_enq_bits_vs : sinkVec_queue_dataOut_29_vs;
  assign sinkVec_queue_29_deq_bits_readSource = _sinkVec_queue_fifo_29_empty ? sinkVec_queue_29_enq_bits_readSource : sinkVec_queue_dataOut_29_readSource;
  assign sinkVec_queue_29_deq_bits_offset = _sinkVec_queue_fifo_29_empty ? sinkVec_queue_29_enq_bits_offset : sinkVec_queue_dataOut_29_offset;
  assign sinkVec_queue_29_deq_bits_instructionIndex = _sinkVec_queue_fifo_29_empty ? sinkVec_queue_29_enq_bits_instructionIndex : sinkVec_queue_dataOut_29_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_29;
  wire         sinkVec_releasePipe_pipe_out_29_valid = sinkVec_releasePipe_pipe_v_29;
  wire         x13_7_1_ready;
  wire         x13_7_1_valid;
  wire         sinkVec_validSource_29_valid = x13_7_1_ready & x13_7_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_29;
  wire [2:0]   sinkVec_tokenCheck_counterChange_29 = sinkVec_validSource_29_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_29 = ~(sinkVec_tokenCheck_counter_29[2]);
  assign x13_7_1_ready = sinkVec_tokenCheck_29;
  assign sinkVec_queue_29_enq_valid = sinkVec_validSink_29_valid;
  assign sinkVec_queue_29_enq_bits_vs = sinkVec_validSink_29_bits_vs;
  assign sinkVec_queue_29_enq_bits_readSource = sinkVec_validSink_29_bits_readSource;
  assign sinkVec_queue_29_enq_bits_offset = sinkVec_validSink_29_bits_offset;
  assign sinkVec_queue_29_enq_bits_instructionIndex = sinkVec_validSink_29_bits_instructionIndex;
  reg          sinkVec_shifterReg_29_0_valid;
  assign sinkVec_validSink_29_valid = sinkVec_shifterReg_29_0_valid;
  reg  [4:0]   sinkVec_shifterReg_29_0_bits_vs;
  assign sinkVec_validSink_29_bits_vs = sinkVec_shifterReg_29_0_bits_vs;
  reg  [1:0]   sinkVec_shifterReg_29_0_bits_readSource;
  assign sinkVec_validSink_29_bits_readSource = sinkVec_shifterReg_29_0_bits_readSource;
  reg  [2:0]   sinkVec_shifterReg_29_0_bits_offset;
  assign sinkVec_validSink_29_bits_offset = sinkVec_shifterReg_29_0_bits_offset;
  reg  [2:0]   sinkVec_shifterReg_29_0_bits_instructionIndex;
  assign sinkVec_validSink_29_bits_instructionIndex = sinkVec_shifterReg_29_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_29 = sinkVec_shifterReg_29_0_valid | sinkVec_validSource_29_valid;
  assign sinkVec_sinkWire_28_ready = sinkVec_14_0_ready;
  assign sinkVec_sinkWire_29_ready = sinkVec_14_1_ready;
  reg          maskUnitFirst_14;
  wire         tryToRead_14 = sinkVec_14_0_valid | sinkVec_14_1_valid;
  wire         sinkWire_14_valid = maskUnitFirst_14 ? sinkVec_14_0_valid : sinkVec_14_1_valid;
  wire [4:0]   sinkWire_14_bits_vs = maskUnitFirst_14 ? sinkVec_14_0_bits_vs : sinkVec_14_1_bits_vs;
  wire [1:0]   sinkWire_14_bits_readSource = maskUnitFirst_14 ? sinkVec_14_0_bits_readSource : sinkVec_14_1_bits_readSource;
  wire [2:0]   sinkWire_14_bits_offset = maskUnitFirst_14 ? sinkVec_14_0_bits_offset : sinkVec_14_1_bits_offset;
  wire [2:0]   sinkWire_14_bits_instructionIndex = maskUnitFirst_14 ? sinkVec_14_0_bits_instructionIndex : sinkVec_14_1_bits_instructionIndex;
  wire         sinkWire_14_ready;
  assign sinkVec_14_1_ready = sinkWire_14_ready & ~maskUnitFirst_14;
  assign sinkVec_14_0_ready = sinkWire_14_ready & maskUnitFirst_14;
  reg          accessDataValid_pipe_v_14;
  reg          accessDataValid_pipe_pipe_v_14;
  wire         accessDataValid_pipe_pipe_out_14_valid = accessDataValid_pipe_pipe_v_14;
  wire         accessDataSource_14_valid = accessDataValid_pipe_pipe_out_14_valid;
  reg          shifterReg_22_0_valid;
  reg  [31:0]  shifterReg_22_0_bits;
  wire         shifterValid_22 = shifterReg_22_0_valid | accessDataSource_14_valid;
  reg          accessDataValid_pipe_v_15;
  reg          accessDataValid_pipe_pipe_v_15;
  wire         accessDataValid_pipe_pipe_out_15_valid = accessDataValid_pipe_pipe_v_15;
  wire         accessDataSource_15_valid = accessDataValid_pipe_pipe_out_15_valid;
  reg          shifterReg_23_0_valid;
  reg  [31:0]  shifterReg_23_0_bits;
  wire         shifterValid_23 = shifterReg_23_0_valid | accessDataSource_15_valid;
  wire         sinkVec_tokenCheck_30;
  wire [4:0]   sinkVec_validSource_30_bits_vd = x22_7_0_bits_vd;
  wire [2:0]   sinkVec_validSource_30_bits_offset = x22_7_0_bits_offset;
  wire [3:0]   sinkVec_validSource_30_bits_mask = x22_7_0_bits_mask;
  wire [31:0]  sinkVec_validSource_30_bits_data = x22_7_0_bits_data;
  wire [2:0]   sinkVec_validSource_30_bits_instructionIndex = x22_7_0_bits_instructionIndex;
  wire         sinkVec_tokenCheck_31;
  wire [4:0]   sinkVec_validSource_31_bits_vd = x22_7_1_bits_vd;
  wire [2:0]   sinkVec_validSource_31_bits_offset = x22_7_1_bits_offset;
  wire [3:0]   sinkVec_validSource_31_bits_mask = x22_7_1_bits_mask;
  wire [31:0]  sinkVec_validSource_31_bits_data = x22_7_1_bits_data;
  wire         sinkVec_validSource_31_bits_last = x22_7_1_bits_last;
  wire [2:0]   sinkVec_validSource_31_bits_instructionIndex = x22_7_1_bits_instructionIndex;
  wire         sinkVec_15_0_ready;
  wire         sinkVec_queue_30_deq_ready = sinkVec_sinkWire_30_ready;
  wire         sinkVec_queue_30_deq_valid;
  wire [4:0]   sinkVec_queue_30_deq_bits_vd;
  wire         sinkVec_15_0_valid = sinkVec_sinkWire_30_valid;
  wire [2:0]   sinkVec_queue_30_deq_bits_offset;
  wire [4:0]   sinkVec_15_0_bits_vd = sinkVec_sinkWire_30_bits_vd;
  wire [3:0]   sinkVec_queue_30_deq_bits_mask;
  wire [2:0]   sinkVec_15_0_bits_offset = sinkVec_sinkWire_30_bits_offset;
  wire [31:0]  sinkVec_queue_30_deq_bits_data;
  wire [3:0]   sinkVec_15_0_bits_mask = sinkVec_sinkWire_30_bits_mask;
  wire         sinkVec_queue_30_deq_bits_last;
  wire [31:0]  sinkVec_15_0_bits_data = sinkVec_sinkWire_30_bits_data;
  wire [2:0]   sinkVec_queue_30_deq_bits_instructionIndex;
  wire         sinkVec_15_0_bits_last = sinkVec_sinkWire_30_bits_last;
  wire [2:0]   sinkVec_15_0_bits_instructionIndex = sinkVec_sinkWire_30_bits_instructionIndex;
  wire         sinkVec_validSink_30_valid;
  wire [4:0]   sinkVec_validSink_30_bits_vd;
  wire [2:0]   sinkVec_validSink_30_bits_offset;
  wire [3:0]   sinkVec_validSink_30_bits_mask;
  wire [31:0]  sinkVec_validSink_30_bits_data;
  wire [2:0]   sinkVec_validSink_30_bits_instructionIndex;
  assign sinkVec_sinkWire_30_valid = sinkVec_queue_30_deq_valid;
  assign sinkVec_sinkWire_30_bits_vd = sinkVec_queue_30_deq_bits_vd;
  assign sinkVec_sinkWire_30_bits_offset = sinkVec_queue_30_deq_bits_offset;
  assign sinkVec_sinkWire_30_bits_mask = sinkVec_queue_30_deq_bits_mask;
  assign sinkVec_sinkWire_30_bits_data = sinkVec_queue_30_deq_bits_data;
  assign sinkVec_sinkWire_30_bits_last = sinkVec_queue_30_deq_bits_last;
  assign sinkVec_sinkWire_30_bits_instructionIndex = sinkVec_queue_30_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_30_enq_bits_data;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_14 = {sinkVec_queue_30_enq_bits_data, 1'h0};
  wire [2:0]   sinkVec_queue_30_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_30 = {sinkVec_queue_dataIn_lo_hi_14, sinkVec_queue_30_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_30_enq_bits_vd;
  wire [2:0]   sinkVec_queue_30_enq_bits_offset;
  wire [7:0]   sinkVec_queue_dataIn_hi_hi_14 = {sinkVec_queue_30_enq_bits_vd, sinkVec_queue_30_enq_bits_offset};
  wire [3:0]   sinkVec_queue_30_enq_bits_mask;
  wire [11:0]  sinkVec_queue_dataIn_hi_30 = {sinkVec_queue_dataIn_hi_hi_14, sinkVec_queue_30_enq_bits_mask};
  wire [47:0]  sinkVec_queue_dataIn_30 = {sinkVec_queue_dataIn_hi_30, sinkVec_queue_dataIn_lo_30};
  wire [2:0]   sinkVec_queue_dataOut_30_instructionIndex = _sinkVec_queue_fifo_30_data_out[2:0];
  wire         sinkVec_queue_dataOut_30_last = _sinkVec_queue_fifo_30_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_30_data = _sinkVec_queue_fifo_30_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_30_mask = _sinkVec_queue_fifo_30_data_out[39:36];
  wire [2:0]   sinkVec_queue_dataOut_30_offset = _sinkVec_queue_fifo_30_data_out[42:40];
  wire [4:0]   sinkVec_queue_dataOut_30_vd = _sinkVec_queue_fifo_30_data_out[47:43];
  wire         sinkVec_queue_30_enq_ready = ~_sinkVec_queue_fifo_30_full;
  wire         sinkVec_queue_30_enq_valid;
  assign sinkVec_queue_30_deq_valid = ~_sinkVec_queue_fifo_30_empty | sinkVec_queue_30_enq_valid;
  assign sinkVec_queue_30_deq_bits_vd = _sinkVec_queue_fifo_30_empty ? sinkVec_queue_30_enq_bits_vd : sinkVec_queue_dataOut_30_vd;
  assign sinkVec_queue_30_deq_bits_offset = _sinkVec_queue_fifo_30_empty ? sinkVec_queue_30_enq_bits_offset : sinkVec_queue_dataOut_30_offset;
  assign sinkVec_queue_30_deq_bits_mask = _sinkVec_queue_fifo_30_empty ? sinkVec_queue_30_enq_bits_mask : sinkVec_queue_dataOut_30_mask;
  assign sinkVec_queue_30_deq_bits_data = _sinkVec_queue_fifo_30_empty ? sinkVec_queue_30_enq_bits_data : sinkVec_queue_dataOut_30_data;
  assign sinkVec_queue_30_deq_bits_last = ~_sinkVec_queue_fifo_30_empty & sinkVec_queue_dataOut_30_last;
  assign sinkVec_queue_30_deq_bits_instructionIndex = _sinkVec_queue_fifo_30_empty ? sinkVec_queue_30_enq_bits_instructionIndex : sinkVec_queue_dataOut_30_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_30;
  wire         sinkVec_releasePipe_pipe_out_30_valid = sinkVec_releasePipe_pipe_v_30;
  wire         x22_7_0_ready;
  wire         x22_7_0_valid;
  wire         sinkVec_validSource_30_valid = x22_7_0_ready & x22_7_0_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_30;
  wire [2:0]   sinkVec_tokenCheck_counterChange_30 = sinkVec_validSource_30_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_30 = ~(sinkVec_tokenCheck_counter_30[2]);
  assign x22_7_0_ready = sinkVec_tokenCheck_30;
  assign sinkVec_queue_30_enq_valid = sinkVec_validSink_30_valid;
  assign sinkVec_queue_30_enq_bits_vd = sinkVec_validSink_30_bits_vd;
  assign sinkVec_queue_30_enq_bits_offset = sinkVec_validSink_30_bits_offset;
  assign sinkVec_queue_30_enq_bits_mask = sinkVec_validSink_30_bits_mask;
  assign sinkVec_queue_30_enq_bits_data = sinkVec_validSink_30_bits_data;
  assign sinkVec_queue_30_enq_bits_instructionIndex = sinkVec_validSink_30_bits_instructionIndex;
  reg          sinkVec_shifterReg_30_0_valid;
  assign sinkVec_validSink_30_valid = sinkVec_shifterReg_30_0_valid;
  reg  [4:0]   sinkVec_shifterReg_30_0_bits_vd;
  assign sinkVec_validSink_30_bits_vd = sinkVec_shifterReg_30_0_bits_vd;
  reg  [2:0]   sinkVec_shifterReg_30_0_bits_offset;
  assign sinkVec_validSink_30_bits_offset = sinkVec_shifterReg_30_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_30_0_bits_mask;
  assign sinkVec_validSink_30_bits_mask = sinkVec_shifterReg_30_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_30_0_bits_data;
  assign sinkVec_validSink_30_bits_data = sinkVec_shifterReg_30_0_bits_data;
  reg  [2:0]   sinkVec_shifterReg_30_0_bits_instructionIndex;
  assign sinkVec_validSink_30_bits_instructionIndex = sinkVec_shifterReg_30_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_30 = sinkVec_shifterReg_30_0_valid | sinkVec_validSource_30_valid;
  wire         sinkVec_15_1_ready;
  wire         sinkVec_queue_31_deq_ready = sinkVec_sinkWire_31_ready;
  wire         sinkVec_queue_31_deq_valid;
  wire [4:0]   sinkVec_queue_31_deq_bits_vd;
  wire         sinkVec_15_1_valid = sinkVec_sinkWire_31_valid;
  wire [2:0]   sinkVec_queue_31_deq_bits_offset;
  wire [4:0]   sinkVec_15_1_bits_vd = sinkVec_sinkWire_31_bits_vd;
  wire [3:0]   sinkVec_queue_31_deq_bits_mask;
  wire [2:0]   sinkVec_15_1_bits_offset = sinkVec_sinkWire_31_bits_offset;
  wire [31:0]  sinkVec_queue_31_deq_bits_data;
  wire [3:0]   sinkVec_15_1_bits_mask = sinkVec_sinkWire_31_bits_mask;
  wire         sinkVec_queue_31_deq_bits_last;
  wire [31:0]  sinkVec_15_1_bits_data = sinkVec_sinkWire_31_bits_data;
  wire [2:0]   sinkVec_queue_31_deq_bits_instructionIndex;
  wire         sinkVec_15_1_bits_last = sinkVec_sinkWire_31_bits_last;
  wire [2:0]   sinkVec_15_1_bits_instructionIndex = sinkVec_sinkWire_31_bits_instructionIndex;
  wire         sinkVec_validSink_31_valid;
  wire [4:0]   sinkVec_validSink_31_bits_vd;
  wire [2:0]   sinkVec_validSink_31_bits_offset;
  wire [3:0]   sinkVec_validSink_31_bits_mask;
  wire [31:0]  sinkVec_validSink_31_bits_data;
  wire         sinkVec_validSink_31_bits_last;
  wire [2:0]   sinkVec_validSink_31_bits_instructionIndex;
  assign sinkVec_sinkWire_31_valid = sinkVec_queue_31_deq_valid;
  assign sinkVec_sinkWire_31_bits_vd = sinkVec_queue_31_deq_bits_vd;
  assign sinkVec_sinkWire_31_bits_offset = sinkVec_queue_31_deq_bits_offset;
  assign sinkVec_sinkWire_31_bits_mask = sinkVec_queue_31_deq_bits_mask;
  assign sinkVec_sinkWire_31_bits_data = sinkVec_queue_31_deq_bits_data;
  assign sinkVec_sinkWire_31_bits_last = sinkVec_queue_31_deq_bits_last;
  assign sinkVec_sinkWire_31_bits_instructionIndex = sinkVec_queue_31_deq_bits_instructionIndex;
  wire [31:0]  sinkVec_queue_31_enq_bits_data;
  wire         sinkVec_queue_31_enq_bits_last;
  wire [32:0]  sinkVec_queue_dataIn_lo_hi_15 = {sinkVec_queue_31_enq_bits_data, sinkVec_queue_31_enq_bits_last};
  wire [2:0]   sinkVec_queue_31_enq_bits_instructionIndex;
  wire [35:0]  sinkVec_queue_dataIn_lo_31 = {sinkVec_queue_dataIn_lo_hi_15, sinkVec_queue_31_enq_bits_instructionIndex};
  wire [4:0]   sinkVec_queue_31_enq_bits_vd;
  wire [2:0]   sinkVec_queue_31_enq_bits_offset;
  wire [7:0]   sinkVec_queue_dataIn_hi_hi_15 = {sinkVec_queue_31_enq_bits_vd, sinkVec_queue_31_enq_bits_offset};
  wire [3:0]   sinkVec_queue_31_enq_bits_mask;
  wire [11:0]  sinkVec_queue_dataIn_hi_31 = {sinkVec_queue_dataIn_hi_hi_15, sinkVec_queue_31_enq_bits_mask};
  wire [47:0]  sinkVec_queue_dataIn_31 = {sinkVec_queue_dataIn_hi_31, sinkVec_queue_dataIn_lo_31};
  wire [2:0]   sinkVec_queue_dataOut_31_instructionIndex = _sinkVec_queue_fifo_31_data_out[2:0];
  wire         sinkVec_queue_dataOut_31_last = _sinkVec_queue_fifo_31_data_out[3];
  wire [31:0]  sinkVec_queue_dataOut_31_data = _sinkVec_queue_fifo_31_data_out[35:4];
  wire [3:0]   sinkVec_queue_dataOut_31_mask = _sinkVec_queue_fifo_31_data_out[39:36];
  wire [2:0]   sinkVec_queue_dataOut_31_offset = _sinkVec_queue_fifo_31_data_out[42:40];
  wire [4:0]   sinkVec_queue_dataOut_31_vd = _sinkVec_queue_fifo_31_data_out[47:43];
  wire         sinkVec_queue_31_enq_ready = ~_sinkVec_queue_fifo_31_full;
  wire         sinkVec_queue_31_enq_valid;
  assign sinkVec_queue_31_deq_valid = ~_sinkVec_queue_fifo_31_empty | sinkVec_queue_31_enq_valid;
  assign sinkVec_queue_31_deq_bits_vd = _sinkVec_queue_fifo_31_empty ? sinkVec_queue_31_enq_bits_vd : sinkVec_queue_dataOut_31_vd;
  assign sinkVec_queue_31_deq_bits_offset = _sinkVec_queue_fifo_31_empty ? sinkVec_queue_31_enq_bits_offset : sinkVec_queue_dataOut_31_offset;
  assign sinkVec_queue_31_deq_bits_mask = _sinkVec_queue_fifo_31_empty ? sinkVec_queue_31_enq_bits_mask : sinkVec_queue_dataOut_31_mask;
  assign sinkVec_queue_31_deq_bits_data = _sinkVec_queue_fifo_31_empty ? sinkVec_queue_31_enq_bits_data : sinkVec_queue_dataOut_31_data;
  assign sinkVec_queue_31_deq_bits_last = _sinkVec_queue_fifo_31_empty ? sinkVec_queue_31_enq_bits_last : sinkVec_queue_dataOut_31_last;
  assign sinkVec_queue_31_deq_bits_instructionIndex = _sinkVec_queue_fifo_31_empty ? sinkVec_queue_31_enq_bits_instructionIndex : sinkVec_queue_dataOut_31_instructionIndex;
  reg          sinkVec_releasePipe_pipe_v_31;
  wire         sinkVec_releasePipe_pipe_out_31_valid = sinkVec_releasePipe_pipe_v_31;
  wire         x22_7_1_ready;
  wire         x22_7_1_valid;
  wire         sinkVec_validSource_31_valid = x22_7_1_ready & x22_7_1_valid;
  reg  [2:0]   sinkVec_tokenCheck_counter_31;
  wire [2:0]   sinkVec_tokenCheck_counterChange_31 = sinkVec_validSource_31_valid ? 3'h1 : 3'h7;
  assign sinkVec_tokenCheck_31 = ~(sinkVec_tokenCheck_counter_31[2]);
  assign x22_7_1_ready = sinkVec_tokenCheck_31;
  assign sinkVec_queue_31_enq_valid = sinkVec_validSink_31_valid;
  assign sinkVec_queue_31_enq_bits_vd = sinkVec_validSink_31_bits_vd;
  assign sinkVec_queue_31_enq_bits_offset = sinkVec_validSink_31_bits_offset;
  assign sinkVec_queue_31_enq_bits_mask = sinkVec_validSink_31_bits_mask;
  assign sinkVec_queue_31_enq_bits_data = sinkVec_validSink_31_bits_data;
  assign sinkVec_queue_31_enq_bits_last = sinkVec_validSink_31_bits_last;
  assign sinkVec_queue_31_enq_bits_instructionIndex = sinkVec_validSink_31_bits_instructionIndex;
  reg          sinkVec_shifterReg_31_0_valid;
  assign sinkVec_validSink_31_valid = sinkVec_shifterReg_31_0_valid;
  reg  [4:0]   sinkVec_shifterReg_31_0_bits_vd;
  assign sinkVec_validSink_31_bits_vd = sinkVec_shifterReg_31_0_bits_vd;
  reg  [2:0]   sinkVec_shifterReg_31_0_bits_offset;
  assign sinkVec_validSink_31_bits_offset = sinkVec_shifterReg_31_0_bits_offset;
  reg  [3:0]   sinkVec_shifterReg_31_0_bits_mask;
  assign sinkVec_validSink_31_bits_mask = sinkVec_shifterReg_31_0_bits_mask;
  reg  [31:0]  sinkVec_shifterReg_31_0_bits_data;
  assign sinkVec_validSink_31_bits_data = sinkVec_shifterReg_31_0_bits_data;
  reg          sinkVec_shifterReg_31_0_bits_last;
  assign sinkVec_validSink_31_bits_last = sinkVec_shifterReg_31_0_bits_last;
  reg  [2:0]   sinkVec_shifterReg_31_0_bits_instructionIndex;
  assign sinkVec_validSink_31_bits_instructionIndex = sinkVec_shifterReg_31_0_bits_instructionIndex;
  wire         sinkVec_shifterValid_31 = sinkVec_shifterReg_31_0_valid | sinkVec_validSource_31_valid;
  assign sinkVec_sinkWire_30_ready = sinkVec_15_0_ready;
  assign sinkVec_sinkWire_31_ready = sinkVec_15_1_ready;
  reg          maskUnitFirst_15;
  wire         tryToRead_15 = sinkVec_15_0_valid | sinkVec_15_1_valid;
  wire         sinkWire_15_valid = maskUnitFirst_15 ? sinkVec_15_0_valid : sinkVec_15_1_valid;
  wire [4:0]   sinkWire_15_bits_vd = maskUnitFirst_15 ? sinkVec_15_0_bits_vd : sinkVec_15_1_bits_vd;
  wire [2:0]   sinkWire_15_bits_offset = maskUnitFirst_15 ? sinkVec_15_0_bits_offset : sinkVec_15_1_bits_offset;
  wire [3:0]   sinkWire_15_bits_mask = maskUnitFirst_15 ? sinkVec_15_0_bits_mask : sinkVec_15_1_bits_mask;
  wire [31:0]  sinkWire_15_bits_data = maskUnitFirst_15 ? sinkVec_15_0_bits_data : sinkVec_15_1_bits_data;
  wire         sinkWire_15_bits_last = maskUnitFirst_15 ? sinkVec_15_0_bits_last : sinkVec_15_1_bits_last;
  wire [2:0]   sinkWire_15_bits_instructionIndex = maskUnitFirst_15 ? sinkVec_15_0_bits_instructionIndex : sinkVec_15_1_bits_instructionIndex;
  wire         sinkWire_15_ready;
  assign sinkVec_15_1_ready = sinkWire_15_ready & ~maskUnitFirst_15;
  assign sinkVec_15_0_ready = sinkWire_15_ready & maskUnitFirst_15;
  reg          view__writeRelease_7_pipe_v;
  wire         view__writeRelease_7_pipe_out_valid = view__writeRelease_7_pipe_v;
  reg          pipe_v_21;
  wire         pipe_out_14_valid = pipe_v_21;
  wire         _probeWire_writeQueueEnqVec_7_valid_T = x22_7_0_ready & _maskUnit_exeResp_7_valid;
  reg          instructionFinishedPipe_pipe_v_7;
  wire         instructionFinishedPipe_pipe_out_7_valid = instructionFinishedPipe_pipe_v_7;
  reg  [7:0]   instructionFinishedPipe_pipe_b_7;
  wire [7:0]   instructionFinishedPipe_pipe_out_7_bits = instructionFinishedPipe_pipe_b_7;
  wire         instructionFinished_7_0 = |(8'h1 << _GEN & instructionFinishedPipe_pipe_out_7_bits);
  wire         instructionFinished_7_1 = |(8'h1 << _GEN_0 & instructionFinishedPipe_pipe_out_7_bits);
  wire         instructionFinished_7_2 = |(8'h1 << _GEN_1 & instructionFinishedPipe_pipe_out_7_bits);
  wire         instructionFinished_7_3 = |(8'h1 << _GEN_2 & instructionFinishedPipe_pipe_out_7_bits);
  assign vxsatReportVec_7 = _laneVec_7_vxsatReport[3:0];
  reg          pipe_v_22;
  reg  [31:0]  pipe_b_22;
  reg          pipe_pipe_v_7;
  wire         pipe_pipe_out_7_valid = pipe_pipe_v_7;
  reg  [31:0]  pipe_pipe_b_7;
  wire [31:0]  pipe_pipe_out_7_bits = pipe_pipe_b_7;
  reg          view__laneMaskSelect_7_pipe_v;
  reg  [5:0]   view__laneMaskSelect_7_pipe_b;
  reg          view__laneMaskSelect_7_pipe_pipe_v;
  wire         view__laneMaskSelect_7_pipe_pipe_out_valid = view__laneMaskSelect_7_pipe_pipe_v;
  reg  [5:0]   view__laneMaskSelect_7_pipe_pipe_b;
  wire [5:0]   view__laneMaskSelect_7_pipe_pipe_out_bits = view__laneMaskSelect_7_pipe_pipe_b;
  reg          view__laneMaskSewSelect_7_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_7_pipe_b;
  reg          view__laneMaskSewSelect_7_pipe_pipe_v;
  wire         view__laneMaskSewSelect_7_pipe_pipe_out_valid = view__laneMaskSewSelect_7_pipe_pipe_v;
  reg  [1:0]   view__laneMaskSewSelect_7_pipe_pipe_b;
  wire [1:0]   view__laneMaskSewSelect_7_pipe_pipe_out_bits = view__laneMaskSewSelect_7_pipe_pipe_b;
  reg          lsuLastPipe_pipe_v_7;
  wire         lsuLastPipe_pipe_out_7_valid = lsuLastPipe_pipe_v_7;
  reg  [7:0]   lsuLastPipe_pipe_b_7;
  wire [7:0]   lsuLastPipe_pipe_out_7_bits = lsuLastPipe_pipe_b_7;
  reg          maskLastPipe_pipe_v_7;
  wire         maskLastPipe_pipe_out_7_valid = maskLastPipe_pipe_v_7;
  reg  [7:0]   maskLastPipe_pipe_b_7;
  wire [7:0]   maskLastPipe_pipe_out_7_bits = maskLastPipe_pipe_b_7;
  wire [6:0]   writeCounter_7 = requestReg_bits_writeByte[11:5] + {6'h0, requestReg_bits_writeByte[4:0] > 5'h1C};
  reg          pipe_v_23;
  wire         pipe_out_15_valid = pipe_v_23;
  reg  [6:0]   pipe_b_23;
  wire [6:0]   pipe_out_15_bits = pipe_b_23;
  reg          pipe_v_24;
  wire         pipe_out_16_valid = pipe_v_24;
  reg          shifterReg_24_0_valid;
  reg  [31:0]  shifterReg_24_0_bits_data;
  wire         shifterValid_24 = shifterReg_24_0_valid | _laneVec_0_readBusPort_0_deq_valid;
  reg          pipe_v_25;
  wire         pipe_out_17_valid = pipe_v_25;
  reg          shifterReg_25_0_valid;
  reg  [31:0]  shifterReg_25_0_bits_data;
  reg  [1:0]   shifterReg_25_0_bits_mask;
  reg  [2:0]   shifterReg_25_0_bits_instructionIndex;
  reg  [6:0]   shifterReg_25_0_bits_counter;
  wire         shifterValid_25 = shifterReg_25_0_valid | _laneVec_0_writeBusPort_0_deq_valid;
  reg          pipe_v_26;
  wire         pipe_out_18_valid = pipe_v_26;
  reg          shifterReg_26_0_valid;
  reg  [31:0]  shifterReg_26_0_bits_data;
  wire         shifterValid_26 = shifterReg_26_0_valid | _laneVec_1_readBusPort_0_deq_valid;
  reg          pipe_v_27;
  wire         pipe_out_19_valid = pipe_v_27;
  reg          shifterReg_27_0_valid;
  reg  [31:0]  shifterReg_27_0_bits_data;
  reg  [1:0]   shifterReg_27_0_bits_mask;
  reg  [2:0]   shifterReg_27_0_bits_instructionIndex;
  reg  [6:0]   shifterReg_27_0_bits_counter;
  wire         shifterValid_27 = shifterReg_27_0_valid | _laneVec_0_writeBusPort_1_deq_valid;
  reg          pipe_v_28;
  wire         pipe_out_20_valid = pipe_v_28;
  reg          shifterReg_28_0_valid;
  reg  [31:0]  shifterReg_28_0_bits_data;
  wire         shifterValid_28 = shifterReg_28_0_valid | _laneVec_2_readBusPort_0_deq_valid;
  reg          pipe_v_29;
  wire         pipe_out_21_valid = pipe_v_29;
  reg          shifterReg_29_0_valid;
  reg  [31:0]  shifterReg_29_0_bits_data;
  reg  [1:0]   shifterReg_29_0_bits_mask;
  reg  [2:0]   shifterReg_29_0_bits_instructionIndex;
  reg  [6:0]   shifterReg_29_0_bits_counter;
  wire         shifterValid_29 = shifterReg_29_0_valid | _laneVec_1_writeBusPort_0_deq_valid;
  reg          pipe_v_30;
  wire         pipe_out_22_valid = pipe_v_30;
  reg          shifterReg_30_0_valid;
  reg  [31:0]  shifterReg_30_0_bits_data;
  wire         shifterValid_30 = shifterReg_30_0_valid | _laneVec_3_readBusPort_0_deq_valid;
  reg          pipe_v_31;
  wire         pipe_out_23_valid = pipe_v_31;
  reg          shifterReg_31_0_valid;
  reg  [31:0]  shifterReg_31_0_bits_data;
  reg  [1:0]   shifterReg_31_0_bits_mask;
  reg  [2:0]   shifterReg_31_0_bits_instructionIndex;
  reg  [6:0]   shifterReg_31_0_bits_counter;
  wire         shifterValid_31 = shifterReg_31_0_valid | _laneVec_1_writeBusPort_1_deq_valid;
  reg          pipe_v_32;
  wire         pipe_out_24_valid = pipe_v_32;
  reg          shifterReg_32_0_valid;
  reg  [31:0]  shifterReg_32_0_bits_data;
  wire         shifterValid_32 = shifterReg_32_0_valid | _laneVec_4_readBusPort_0_deq_valid;
  reg          pipe_v_33;
  wire         pipe_out_25_valid = pipe_v_33;
  reg          shifterReg_33_0_valid;
  reg  [31:0]  shifterReg_33_0_bits_data;
  reg  [1:0]   shifterReg_33_0_bits_mask;
  reg  [2:0]   shifterReg_33_0_bits_instructionIndex;
  reg  [6:0]   shifterReg_33_0_bits_counter;
  wire         shifterValid_33 = shifterReg_33_0_valid | _laneVec_2_writeBusPort_0_deq_valid;
  reg          pipe_v_34;
  wire         pipe_out_26_valid = pipe_v_34;
  reg          shifterReg_34_0_valid;
  reg  [31:0]  shifterReg_34_0_bits_data;
  wire         shifterValid_34 = shifterReg_34_0_valid | _laneVec_5_readBusPort_0_deq_valid;
  reg          pipe_v_35;
  wire         pipe_out_27_valid = pipe_v_35;
  reg          shifterReg_35_0_valid;
  reg  [31:0]  shifterReg_35_0_bits_data;
  reg  [1:0]   shifterReg_35_0_bits_mask;
  reg  [2:0]   shifterReg_35_0_bits_instructionIndex;
  reg  [6:0]   shifterReg_35_0_bits_counter;
  wire         shifterValid_35 = shifterReg_35_0_valid | _laneVec_2_writeBusPort_1_deq_valid;
  reg          pipe_v_36;
  wire         pipe_out_28_valid = pipe_v_36;
  reg          shifterReg_36_0_valid;
  reg  [31:0]  shifterReg_36_0_bits_data;
  wire         shifterValid_36 = shifterReg_36_0_valid | _laneVec_6_readBusPort_0_deq_valid;
  reg          pipe_v_37;
  wire         pipe_out_29_valid = pipe_v_37;
  reg          shifterReg_37_0_valid;
  reg  [31:0]  shifterReg_37_0_bits_data;
  reg  [1:0]   shifterReg_37_0_bits_mask;
  reg  [2:0]   shifterReg_37_0_bits_instructionIndex;
  reg  [6:0]   shifterReg_37_0_bits_counter;
  wire         shifterValid_37 = shifterReg_37_0_valid | _laneVec_3_writeBusPort_0_deq_valid;
  reg          pipe_v_38;
  wire         pipe_out_30_valid = pipe_v_38;
  reg          shifterReg_38_0_valid;
  reg  [31:0]  shifterReg_38_0_bits_data;
  wire         shifterValid_38 = shifterReg_38_0_valid | _laneVec_7_readBusPort_0_deq_valid;
  reg          pipe_v_39;
  wire         pipe_out_31_valid = pipe_v_39;
  reg          shifterReg_39_0_valid;
  reg  [31:0]  shifterReg_39_0_bits_data;
  reg  [1:0]   shifterReg_39_0_bits_mask;
  reg  [2:0]   shifterReg_39_0_bits_instructionIndex;
  reg  [6:0]   shifterReg_39_0_bits_counter;
  wire         shifterValid_39 = shifterReg_39_0_valid | _laneVec_3_writeBusPort_1_deq_valid;
  reg          pipe_v_40;
  wire         pipe_out_32_valid = pipe_v_40;
  reg          shifterReg_40_0_valid;
  reg  [31:0]  shifterReg_40_0_bits_data;
  wire         shifterValid_40 = shifterReg_40_0_valid | _laneVec_0_readBusPort_1_deq_valid;
  reg          pipe_v_41;
  wire         pipe_out_33_valid = pipe_v_41;
  reg          shifterReg_41_0_valid;
  reg  [31:0]  shifterReg_41_0_bits_data;
  reg  [1:0]   shifterReg_41_0_bits_mask;
  reg  [2:0]   shifterReg_41_0_bits_instructionIndex;
  reg  [6:0]   shifterReg_41_0_bits_counter;
  wire         shifterValid_41 = shifterReg_41_0_valid | _laneVec_4_writeBusPort_0_deq_valid;
  reg          pipe_v_42;
  wire         pipe_out_34_valid = pipe_v_42;
  reg          shifterReg_42_0_valid;
  reg  [31:0]  shifterReg_42_0_bits_data;
  wire         shifterValid_42 = shifterReg_42_0_valid | _laneVec_1_readBusPort_1_deq_valid;
  reg          pipe_v_43;
  wire         pipe_out_35_valid = pipe_v_43;
  reg          shifterReg_43_0_valid;
  reg  [31:0]  shifterReg_43_0_bits_data;
  reg  [1:0]   shifterReg_43_0_bits_mask;
  reg  [2:0]   shifterReg_43_0_bits_instructionIndex;
  reg  [6:0]   shifterReg_43_0_bits_counter;
  wire         shifterValid_43 = shifterReg_43_0_valid | _laneVec_4_writeBusPort_1_deq_valid;
  reg          pipe_v_44;
  wire         pipe_out_36_valid = pipe_v_44;
  reg          shifterReg_44_0_valid;
  reg  [31:0]  shifterReg_44_0_bits_data;
  wire         shifterValid_44 = shifterReg_44_0_valid | _laneVec_2_readBusPort_1_deq_valid;
  reg          pipe_v_45;
  wire         pipe_out_37_valid = pipe_v_45;
  reg          shifterReg_45_0_valid;
  reg  [31:0]  shifterReg_45_0_bits_data;
  reg  [1:0]   shifterReg_45_0_bits_mask;
  reg  [2:0]   shifterReg_45_0_bits_instructionIndex;
  reg  [6:0]   shifterReg_45_0_bits_counter;
  wire         shifterValid_45 = shifterReg_45_0_valid | _laneVec_5_writeBusPort_0_deq_valid;
  reg          pipe_v_46;
  wire         pipe_out_38_valid = pipe_v_46;
  reg          shifterReg_46_0_valid;
  reg  [31:0]  shifterReg_46_0_bits_data;
  wire         shifterValid_46 = shifterReg_46_0_valid | _laneVec_3_readBusPort_1_deq_valid;
  reg          pipe_v_47;
  wire         pipe_out_39_valid = pipe_v_47;
  reg          shifterReg_47_0_valid;
  reg  [31:0]  shifterReg_47_0_bits_data;
  reg  [1:0]   shifterReg_47_0_bits_mask;
  reg  [2:0]   shifterReg_47_0_bits_instructionIndex;
  reg  [6:0]   shifterReg_47_0_bits_counter;
  wire         shifterValid_47 = shifterReg_47_0_valid | _laneVec_5_writeBusPort_1_deq_valid;
  reg          pipe_v_48;
  wire         pipe_out_40_valid = pipe_v_48;
  reg          shifterReg_48_0_valid;
  reg  [31:0]  shifterReg_48_0_bits_data;
  wire         shifterValid_48 = shifterReg_48_0_valid | _laneVec_4_readBusPort_1_deq_valid;
  reg          pipe_v_49;
  wire         pipe_out_41_valid = pipe_v_49;
  reg          shifterReg_49_0_valid;
  reg  [31:0]  shifterReg_49_0_bits_data;
  reg  [1:0]   shifterReg_49_0_bits_mask;
  reg  [2:0]   shifterReg_49_0_bits_instructionIndex;
  reg  [6:0]   shifterReg_49_0_bits_counter;
  wire         shifterValid_49 = shifterReg_49_0_valid | _laneVec_6_writeBusPort_0_deq_valid;
  reg          pipe_v_50;
  wire         pipe_out_42_valid = pipe_v_50;
  reg          shifterReg_50_0_valid;
  reg  [31:0]  shifterReg_50_0_bits_data;
  wire         shifterValid_50 = shifterReg_50_0_valid | _laneVec_5_readBusPort_1_deq_valid;
  reg          pipe_v_51;
  wire         pipe_out_43_valid = pipe_v_51;
  reg          shifterReg_51_0_valid;
  reg  [31:0]  shifterReg_51_0_bits_data;
  reg  [1:0]   shifterReg_51_0_bits_mask;
  reg  [2:0]   shifterReg_51_0_bits_instructionIndex;
  reg  [6:0]   shifterReg_51_0_bits_counter;
  wire         shifterValid_51 = shifterReg_51_0_valid | _laneVec_6_writeBusPort_1_deq_valid;
  reg          pipe_v_52;
  wire         pipe_out_44_valid = pipe_v_52;
  reg          shifterReg_52_0_valid;
  reg  [31:0]  shifterReg_52_0_bits_data;
  wire         shifterValid_52 = shifterReg_52_0_valid | _laneVec_6_readBusPort_1_deq_valid;
  reg          pipe_v_53;
  wire         pipe_out_45_valid = pipe_v_53;
  reg          shifterReg_53_0_valid;
  reg  [31:0]  shifterReg_53_0_bits_data;
  reg  [1:0]   shifterReg_53_0_bits_mask;
  reg  [2:0]   shifterReg_53_0_bits_instructionIndex;
  reg  [6:0]   shifterReg_53_0_bits_counter;
  wire         shifterValid_53 = shifterReg_53_0_valid | _laneVec_7_writeBusPort_0_deq_valid;
  reg          pipe_v_54;
  wire         pipe_out_46_valid = pipe_v_54;
  reg          shifterReg_54_0_valid;
  reg  [31:0]  shifterReg_54_0_bits_data;
  wire         shifterValid_54 = shifterReg_54_0_valid | _laneVec_7_readBusPort_1_deq_valid;
  reg          pipe_v_55;
  wire         pipe_out_47_valid = pipe_v_55;
  reg          shifterReg_55_0_valid;
  reg  [31:0]  shifterReg_55_0_bits_data;
  reg  [1:0]   shifterReg_55_0_bits_mask;
  reg  [2:0]   shifterReg_55_0_bits_instructionIndex;
  reg  [6:0]   shifterReg_55_0_bits_counter;
  wire         shifterValid_55 = shifterReg_55_0_valid | _laneVec_7_writeBusPort_1_deq_valid;
  wire [3:0]   free = {free_hi, free_lo};
  wire         allSlotFree = &free;
  wire [1:0]   existMaskType_lo = {~slots_1_state_idle & slots_1_record_maskType, ~slots_0_state_idle & slots_0_record_maskType};
  wire [1:0]   existMaskType_hi = {~slots_3_state_idle & slots_3_record_maskType, ~slots_2_state_idle & slots_2_record_maskType};
  wire         existMaskType = |{existMaskType_hi, existMaskType_lo};
  wire [2:0]   _free1H_T_2 = free[2:0] | {free[1:0], 1'h0};
  wire [3:0]   free1H = {~(_free1H_T_2 | {_free1H_T_2[0], 2'h0}), 1'h1} & free;
  wire [3:0]   slotToEnqueue = specialInstruction ? 4'h8 : free1H;
  wire         instructionIndexFree =
    (slots_0_state_idle | slots_0_record_instructionIndex[1:0] != requestReg_bits_instructionIndex[1:0]) & (slots_1_state_idle | slots_1_record_instructionIndex[1:0] != requestReg_bits_instructionIndex[1:0])
    & (slots_2_state_idle | slots_2_record_instructionIndex[1:0] != requestReg_bits_instructionIndex[1:0]) & (slots_3_state_idle | slots_3_record_instructionIndex[1:0] != requestReg_bits_instructionIndex[1:0]);
  wire         executionReady = (~isLoadStoreType | _lsu_request_ready) & (noOffsetReadLoadStore | allLaneReady);
  assign requestRegDequeue_ready = executionReady & slotReady & (~gatherNeedRead | _maskUnit_gatherData_valid) & _tokenManager_issueAllow & instructionIndexFree & olderCheck;
  wire [3:0]   instructionToSlotOH = maskUnit_gatherData_ready ? slotToEnqueue : 4'h0;
  wire         slotCommit_0 = slots_0_state_wMaskUnitLast & slots_0_state_wLast & slots_0_state_wVRFWrite & ~slots_0_state_sCommit & slots_0_record_instructionIndex == responseCounter;
  wire         slotCommit_1 = slots_1_state_wMaskUnitLast & slots_1_state_wLast & slots_1_state_wVRFWrite & ~slots_1_state_sCommit & slots_1_record_instructionIndex == responseCounter;
  wire         slotCommit_2 = slots_2_state_wMaskUnitLast & slots_2_state_wLast & slots_2_state_wVRFWrite & ~slots_2_state_sCommit & slots_2_record_instructionIndex == responseCounter;
  assign slotCommit_3 = slots_3_state_wMaskUnitLast & slots_3_state_wLast & slots_3_state_wVRFWrite & ~slots_3_state_sCommit & slots_3_record_instructionIndex == responseCounter;
  assign lastSlotCommit = slotCommit_3;
  wire [1:0]   _GEN_5 = {slotCommit_1, slotCommit_0};
  wire [1:0]   retire_lo;
  assign retire_lo = _GEN_5;
  wire [1:0]   view__retire_csr_bits_vxsat_lo;
  assign view__retire_csr_bits_vxsat_lo = _GEN_5;
  wire [1:0]   view__retire_mem_valid_lo;
  assign view__retire_mem_valid_lo = _GEN_5;
  wire [1:0]   _GEN_6 = {slotCommit_3, slotCommit_2};
  wire [1:0]   retire_hi;
  assign retire_hi = _GEN_6;
  wire [1:0]   view__retire_csr_bits_vxsat_hi;
  assign view__retire_csr_bits_vxsat_hi = _GEN_6;
  wire [1:0]   view__retire_mem_valid_hi;
  assign view__retire_mem_valid_hi = _GEN_6;
  wire         retire_1 = |{retire_hi, retire_lo};
  wire [1:0]   view__retire_csr_bits_vxsat_lo_1 = {slots_1_vxsat, slots_0_vxsat};
  wire [1:0]   view__retire_csr_bits_vxsat_hi_1 = {slots_3_vxsat, slots_2_vxsat};
  wire [31:0]  retire_csr_bits_vxsat_0 = {31'h0, |({view__retire_csr_bits_vxsat_hi, view__retire_csr_bits_vxsat_lo} & {view__retire_csr_bits_vxsat_hi_1, view__retire_csr_bits_vxsat_lo_1})};
  wire [1:0]   view__retire_mem_valid_lo_1 = {slots_1_record_isLoadStore, slots_0_record_isLoadStore};
  wire [1:0]   view__retire_mem_valid_hi_1 = {slots_3_record_isLoadStore, slots_2_record_isLoadStore};
  wire         retire_mem_valid_0 = |({view__retire_mem_valid_hi, view__retire_mem_valid_lo} & {view__retire_mem_valid_hi_1, view__retire_mem_valid_lo_1});
  wire [31:0]  accessDataSource_bits;
  wire [31:0]  accessDataSource_1_bits;
  wire [31:0]  accessDataSource_2_bits;
  wire [31:0]  accessDataSource_3_bits;
  wire [31:0]  accessDataSource_4_bits;
  wire [31:0]  accessDataSource_5_bits;
  wire [31:0]  accessDataSource_6_bits;
  wire [31:0]  accessDataSource_7_bits;
  wire [31:0]  accessDataSource_8_bits;
  wire [31:0]  accessDataSource_9_bits;
  wire [31:0]  accessDataSource_10_bits;
  wire [31:0]  accessDataSource_11_bits;
  wire [31:0]  accessDataSource_12_bits;
  wire [31:0]  accessDataSource_13_bits;
  wire [31:0]  accessDataSource_14_bits;
  wire [31:0]  accessDataSource_15_bits;
  always @(posedge clock) begin
    if (reset) begin
      instructionCounter <= 3'h0;
      responseCounter <= 3'h0;
      requestReg_valid <= 1'h0;
      requestReg_bits_issue_instruction <= 32'h0;
      requestReg_bits_issue_rs1Data <= 32'h0;
      requestReg_bits_issue_rs2Data <= 32'h0;
      requestReg_bits_issue_vtype <= 32'h0;
      requestReg_bits_issue_vl <= 32'h0;
      requestReg_bits_issue_vstart <= 32'h0;
      requestReg_bits_issue_vcsr <= 32'h0;
      requestReg_bits_decodeResult_specialSlot <= 1'h0;
      requestReg_bits_decodeResult_topUop <= 5'h0;
      requestReg_bits_decodeResult_popCount <= 1'h0;
      requestReg_bits_decodeResult_ffo <= 1'h0;
      requestReg_bits_decodeResult_average <= 1'h0;
      requestReg_bits_decodeResult_reverse <= 1'h0;
      requestReg_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      requestReg_bits_decodeResult_scheduler <= 1'h0;
      requestReg_bits_decodeResult_sReadVD <= 1'h0;
      requestReg_bits_decodeResult_vtype <= 1'h0;
      requestReg_bits_decodeResult_sWrite <= 1'h0;
      requestReg_bits_decodeResult_crossRead <= 1'h0;
      requestReg_bits_decodeResult_crossWrite <= 1'h0;
      requestReg_bits_decodeResult_maskUnit <= 1'h0;
      requestReg_bits_decodeResult_special <= 1'h0;
      requestReg_bits_decodeResult_saturate <= 1'h0;
      requestReg_bits_decodeResult_vwmacc <= 1'h0;
      requestReg_bits_decodeResult_readOnly <= 1'h0;
      requestReg_bits_decodeResult_maskSource <= 1'h0;
      requestReg_bits_decodeResult_maskDestination <= 1'h0;
      requestReg_bits_decodeResult_maskLogic <= 1'h0;
      requestReg_bits_decodeResult_uop <= 4'h0;
      requestReg_bits_decodeResult_iota <= 1'h0;
      requestReg_bits_decodeResult_mv <= 1'h0;
      requestReg_bits_decodeResult_extend <= 1'h0;
      requestReg_bits_decodeResult_unOrderWrite <= 1'h0;
      requestReg_bits_decodeResult_compress <= 1'h0;
      requestReg_bits_decodeResult_gather16 <= 1'h0;
      requestReg_bits_decodeResult_gather <= 1'h0;
      requestReg_bits_decodeResult_slid <= 1'h0;
      requestReg_bits_decodeResult_targetRd <= 1'h0;
      requestReg_bits_decodeResult_widenReduce <= 1'h0;
      requestReg_bits_decodeResult_red <= 1'h0;
      requestReg_bits_decodeResult_nr <= 1'h0;
      requestReg_bits_decodeResult_itype <= 1'h0;
      requestReg_bits_decodeResult_unsigned1 <= 1'h0;
      requestReg_bits_decodeResult_unsigned0 <= 1'h0;
      requestReg_bits_decodeResult_other <= 1'h0;
      requestReg_bits_decodeResult_multiCycle <= 1'h0;
      requestReg_bits_decodeResult_divider <= 1'h0;
      requestReg_bits_decodeResult_multiplier <= 1'h0;
      requestReg_bits_decodeResult_shift <= 1'h0;
      requestReg_bits_decodeResult_adder <= 1'h0;
      requestReg_bits_decodeResult_logic <= 1'h0;
      requestReg_bits_instructionIndex <= 3'h0;
      requestReg_bits_vdIsV0 <= 1'h0;
      requestReg_bits_writeByte <= 12'h0;
      slots_0_record_instructionIndex <= 3'h7;
      slots_0_record_isLoadStore <= 1'h1;
      slots_0_record_maskType <= 1'h1;
      slots_0_state_wLast <= 1'h1;
      slots_0_state_idle <= 1'h1;
      slots_0_state_wMaskUnitLast <= 1'h1;
      slots_0_state_wVRFWrite <= 1'h1;
      slots_0_state_sCommit <= 1'h1;
      slots_0_endTag_0 <= 1'h1;
      slots_0_endTag_1 <= 1'h1;
      slots_0_endTag_2 <= 1'h1;
      slots_0_endTag_3 <= 1'h1;
      slots_0_endTag_4 <= 1'h1;
      slots_0_endTag_5 <= 1'h1;
      slots_0_endTag_6 <= 1'h1;
      slots_0_endTag_7 <= 1'h1;
      slots_0_endTag_8 <= 1'h1;
      slots_0_vxsat <= 1'h1;
      slots_1_record_instructionIndex <= 3'h7;
      slots_1_record_isLoadStore <= 1'h1;
      slots_1_record_maskType <= 1'h1;
      slots_1_state_wLast <= 1'h1;
      slots_1_state_idle <= 1'h1;
      slots_1_state_wMaskUnitLast <= 1'h1;
      slots_1_state_wVRFWrite <= 1'h1;
      slots_1_state_sCommit <= 1'h1;
      slots_1_endTag_0 <= 1'h1;
      slots_1_endTag_1 <= 1'h1;
      slots_1_endTag_2 <= 1'h1;
      slots_1_endTag_3 <= 1'h1;
      slots_1_endTag_4 <= 1'h1;
      slots_1_endTag_5 <= 1'h1;
      slots_1_endTag_6 <= 1'h1;
      slots_1_endTag_7 <= 1'h1;
      slots_1_endTag_8 <= 1'h1;
      slots_1_vxsat <= 1'h1;
      slots_2_record_instructionIndex <= 3'h7;
      slots_2_record_isLoadStore <= 1'h1;
      slots_2_record_maskType <= 1'h1;
      slots_2_state_wLast <= 1'h1;
      slots_2_state_idle <= 1'h1;
      slots_2_state_wMaskUnitLast <= 1'h1;
      slots_2_state_wVRFWrite <= 1'h1;
      slots_2_state_sCommit <= 1'h1;
      slots_2_endTag_0 <= 1'h1;
      slots_2_endTag_1 <= 1'h1;
      slots_2_endTag_2 <= 1'h1;
      slots_2_endTag_3 <= 1'h1;
      slots_2_endTag_4 <= 1'h1;
      slots_2_endTag_5 <= 1'h1;
      slots_2_endTag_6 <= 1'h1;
      slots_2_endTag_7 <= 1'h1;
      slots_2_endTag_8 <= 1'h1;
      slots_2_vxsat <= 1'h1;
      slots_3_record_instructionIndex <= 3'h7;
      slots_3_record_isLoadStore <= 1'h1;
      slots_3_record_maskType <= 1'h1;
      slots_3_state_wLast <= 1'h1;
      slots_3_state_idle <= 1'h1;
      slots_3_state_wMaskUnitLast <= 1'h1;
      slots_3_state_wVRFWrite <= 1'h1;
      slots_3_state_sCommit <= 1'h1;
      slots_3_endTag_0 <= 1'h1;
      slots_3_endTag_1 <= 1'h1;
      slots_3_endTag_2 <= 1'h1;
      slots_3_endTag_3 <= 1'h1;
      slots_3_endTag_4 <= 1'h1;
      slots_3_endTag_5 <= 1'h1;
      slots_3_endTag_6 <= 1'h1;
      slots_3_endTag_7 <= 1'h1;
      slots_3_endTag_8 <= 1'h1;
      slots_3_vxsat <= 1'h1;
      slots_writeRD <= 1'h0;
      slots_vd <= 5'h0;
      releasePipe_pipe_v <= 1'h0;
      tokenCheck_counter <= 3'h0;
      shifterReg_0_valid <= 1'h0;
      shifterReg_0_bits_instructionIndex <= 3'h0;
      shifterReg_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_0_bits_decodeResult_average <= 1'h0;
      shifterReg_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_0_bits_decodeResult_special <= 1'h0;
      shifterReg_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_0_bits_decodeResult_red <= 1'h0;
      shifterReg_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_0_bits_decodeResult_other <= 1'h0;
      shifterReg_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_0_bits_loadStore <= 1'h0;
      shifterReg_0_bits_issueInst <= 1'h0;
      shifterReg_0_bits_store <= 1'h0;
      shifterReg_0_bits_special <= 1'h0;
      shifterReg_0_bits_lsWholeReg <= 1'h0;
      shifterReg_0_bits_vs1 <= 5'h0;
      shifterReg_0_bits_vs2 <= 5'h0;
      shifterReg_0_bits_vd <= 5'h0;
      shifterReg_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_0_bits_mask <= 1'h0;
      shifterReg_0_bits_segment <= 3'h0;
      shifterReg_0_bits_readFromScalar <= 32'h0;
      shifterReg_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_0_bits_csrInterface_vma <= 1'h0;
      releasePipe_pipe_v_1 <= 1'h0;
      tokenCheck_counter_1 <= 3'h0;
      shifterReg_1_0_valid <= 1'h0;
      shifterReg_1_0_bits_instructionIndex <= 3'h0;
      shifterReg_1_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_1_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_1_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_1_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_1_0_bits_decodeResult_average <= 1'h0;
      shifterReg_1_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_1_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_1_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_1_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_1_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_1_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_1_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_1_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_1_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_1_0_bits_decodeResult_special <= 1'h0;
      shifterReg_1_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_1_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_1_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_1_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_1_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_1_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_1_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_1_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_1_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_1_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_1_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_1_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_1_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_1_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_1_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_1_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_1_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_1_0_bits_decodeResult_red <= 1'h0;
      shifterReg_1_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_1_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_1_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_1_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_1_0_bits_decodeResult_other <= 1'h0;
      shifterReg_1_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_1_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_1_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_1_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_1_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_1_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_1_0_bits_loadStore <= 1'h0;
      shifterReg_1_0_bits_issueInst <= 1'h0;
      shifterReg_1_0_bits_store <= 1'h0;
      shifterReg_1_0_bits_special <= 1'h0;
      shifterReg_1_0_bits_lsWholeReg <= 1'h0;
      shifterReg_1_0_bits_vs1 <= 5'h0;
      shifterReg_1_0_bits_vs2 <= 5'h0;
      shifterReg_1_0_bits_vd <= 5'h0;
      shifterReg_1_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_1_0_bits_mask <= 1'h0;
      shifterReg_1_0_bits_segment <= 3'h0;
      shifterReg_1_0_bits_readFromScalar <= 32'h0;
      shifterReg_1_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_1_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_1_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_1_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_1_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_1_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_1_0_bits_csrInterface_vma <= 1'h0;
      releasePipe_pipe_v_2 <= 1'h0;
      tokenCheck_counter_2 <= 3'h0;
      shifterReg_2_0_valid <= 1'h0;
      shifterReg_2_0_bits_instructionIndex <= 3'h0;
      shifterReg_2_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_2_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_2_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_2_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_2_0_bits_decodeResult_average <= 1'h0;
      shifterReg_2_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_2_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_2_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_2_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_2_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_2_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_2_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_2_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_2_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_2_0_bits_decodeResult_special <= 1'h0;
      shifterReg_2_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_2_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_2_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_2_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_2_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_2_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_2_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_2_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_2_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_2_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_2_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_2_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_2_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_2_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_2_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_2_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_2_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_2_0_bits_decodeResult_red <= 1'h0;
      shifterReg_2_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_2_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_2_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_2_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_2_0_bits_decodeResult_other <= 1'h0;
      shifterReg_2_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_2_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_2_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_2_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_2_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_2_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_2_0_bits_loadStore <= 1'h0;
      shifterReg_2_0_bits_issueInst <= 1'h0;
      shifterReg_2_0_bits_store <= 1'h0;
      shifterReg_2_0_bits_special <= 1'h0;
      shifterReg_2_0_bits_lsWholeReg <= 1'h0;
      shifterReg_2_0_bits_vs1 <= 5'h0;
      shifterReg_2_0_bits_vs2 <= 5'h0;
      shifterReg_2_0_bits_vd <= 5'h0;
      shifterReg_2_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_2_0_bits_mask <= 1'h0;
      shifterReg_2_0_bits_segment <= 3'h0;
      shifterReg_2_0_bits_readFromScalar <= 32'h0;
      shifterReg_2_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_2_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_2_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_2_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_2_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_2_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_2_0_bits_csrInterface_vma <= 1'h0;
      releasePipe_pipe_v_3 <= 1'h0;
      tokenCheck_counter_3 <= 3'h0;
      shifterReg_3_0_valid <= 1'h0;
      shifterReg_3_0_bits_instructionIndex <= 3'h0;
      shifterReg_3_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_3_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_3_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_3_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_3_0_bits_decodeResult_average <= 1'h0;
      shifterReg_3_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_3_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_3_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_3_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_3_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_3_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_3_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_3_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_3_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_3_0_bits_decodeResult_special <= 1'h0;
      shifterReg_3_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_3_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_3_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_3_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_3_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_3_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_3_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_3_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_3_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_3_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_3_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_3_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_3_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_3_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_3_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_3_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_3_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_3_0_bits_decodeResult_red <= 1'h0;
      shifterReg_3_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_3_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_3_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_3_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_3_0_bits_decodeResult_other <= 1'h0;
      shifterReg_3_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_3_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_3_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_3_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_3_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_3_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_3_0_bits_loadStore <= 1'h0;
      shifterReg_3_0_bits_issueInst <= 1'h0;
      shifterReg_3_0_bits_store <= 1'h0;
      shifterReg_3_0_bits_special <= 1'h0;
      shifterReg_3_0_bits_lsWholeReg <= 1'h0;
      shifterReg_3_0_bits_vs1 <= 5'h0;
      shifterReg_3_0_bits_vs2 <= 5'h0;
      shifterReg_3_0_bits_vd <= 5'h0;
      shifterReg_3_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_3_0_bits_mask <= 1'h0;
      shifterReg_3_0_bits_segment <= 3'h0;
      shifterReg_3_0_bits_readFromScalar <= 32'h0;
      shifterReg_3_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_3_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_3_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_3_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_3_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_3_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_3_0_bits_csrInterface_vma <= 1'h0;
      releasePipe_pipe_v_4 <= 1'h0;
      tokenCheck_counter_4 <= 3'h0;
      shifterReg_4_0_valid <= 1'h0;
      shifterReg_4_0_bits_instructionIndex <= 3'h0;
      shifterReg_4_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_4_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_4_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_4_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_4_0_bits_decodeResult_average <= 1'h0;
      shifterReg_4_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_4_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_4_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_4_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_4_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_4_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_4_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_4_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_4_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_4_0_bits_decodeResult_special <= 1'h0;
      shifterReg_4_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_4_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_4_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_4_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_4_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_4_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_4_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_4_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_4_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_4_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_4_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_4_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_4_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_4_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_4_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_4_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_4_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_4_0_bits_decodeResult_red <= 1'h0;
      shifterReg_4_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_4_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_4_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_4_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_4_0_bits_decodeResult_other <= 1'h0;
      shifterReg_4_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_4_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_4_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_4_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_4_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_4_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_4_0_bits_loadStore <= 1'h0;
      shifterReg_4_0_bits_issueInst <= 1'h0;
      shifterReg_4_0_bits_store <= 1'h0;
      shifterReg_4_0_bits_special <= 1'h0;
      shifterReg_4_0_bits_lsWholeReg <= 1'h0;
      shifterReg_4_0_bits_vs1 <= 5'h0;
      shifterReg_4_0_bits_vs2 <= 5'h0;
      shifterReg_4_0_bits_vd <= 5'h0;
      shifterReg_4_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_4_0_bits_mask <= 1'h0;
      shifterReg_4_0_bits_segment <= 3'h0;
      shifterReg_4_0_bits_readFromScalar <= 32'h0;
      shifterReg_4_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_4_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_4_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_4_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_4_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_4_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_4_0_bits_csrInterface_vma <= 1'h0;
      releasePipe_pipe_v_5 <= 1'h0;
      tokenCheck_counter_5 <= 3'h0;
      shifterReg_5_0_valid <= 1'h0;
      shifterReg_5_0_bits_instructionIndex <= 3'h0;
      shifterReg_5_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_5_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_5_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_5_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_5_0_bits_decodeResult_average <= 1'h0;
      shifterReg_5_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_5_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_5_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_5_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_5_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_5_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_5_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_5_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_5_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_5_0_bits_decodeResult_special <= 1'h0;
      shifterReg_5_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_5_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_5_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_5_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_5_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_5_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_5_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_5_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_5_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_5_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_5_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_5_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_5_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_5_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_5_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_5_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_5_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_5_0_bits_decodeResult_red <= 1'h0;
      shifterReg_5_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_5_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_5_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_5_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_5_0_bits_decodeResult_other <= 1'h0;
      shifterReg_5_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_5_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_5_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_5_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_5_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_5_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_5_0_bits_loadStore <= 1'h0;
      shifterReg_5_0_bits_issueInst <= 1'h0;
      shifterReg_5_0_bits_store <= 1'h0;
      shifterReg_5_0_bits_special <= 1'h0;
      shifterReg_5_0_bits_lsWholeReg <= 1'h0;
      shifterReg_5_0_bits_vs1 <= 5'h0;
      shifterReg_5_0_bits_vs2 <= 5'h0;
      shifterReg_5_0_bits_vd <= 5'h0;
      shifterReg_5_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_5_0_bits_mask <= 1'h0;
      shifterReg_5_0_bits_segment <= 3'h0;
      shifterReg_5_0_bits_readFromScalar <= 32'h0;
      shifterReg_5_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_5_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_5_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_5_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_5_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_5_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_5_0_bits_csrInterface_vma <= 1'h0;
      releasePipe_pipe_v_6 <= 1'h0;
      tokenCheck_counter_6 <= 3'h0;
      shifterReg_6_0_valid <= 1'h0;
      shifterReg_6_0_bits_instructionIndex <= 3'h0;
      shifterReg_6_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_6_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_6_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_6_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_6_0_bits_decodeResult_average <= 1'h0;
      shifterReg_6_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_6_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_6_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_6_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_6_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_6_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_6_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_6_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_6_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_6_0_bits_decodeResult_special <= 1'h0;
      shifterReg_6_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_6_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_6_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_6_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_6_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_6_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_6_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_6_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_6_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_6_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_6_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_6_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_6_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_6_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_6_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_6_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_6_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_6_0_bits_decodeResult_red <= 1'h0;
      shifterReg_6_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_6_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_6_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_6_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_6_0_bits_decodeResult_other <= 1'h0;
      shifterReg_6_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_6_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_6_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_6_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_6_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_6_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_6_0_bits_loadStore <= 1'h0;
      shifterReg_6_0_bits_issueInst <= 1'h0;
      shifterReg_6_0_bits_store <= 1'h0;
      shifterReg_6_0_bits_special <= 1'h0;
      shifterReg_6_0_bits_lsWholeReg <= 1'h0;
      shifterReg_6_0_bits_vs1 <= 5'h0;
      shifterReg_6_0_bits_vs2 <= 5'h0;
      shifterReg_6_0_bits_vd <= 5'h0;
      shifterReg_6_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_6_0_bits_mask <= 1'h0;
      shifterReg_6_0_bits_segment <= 3'h0;
      shifterReg_6_0_bits_readFromScalar <= 32'h0;
      shifterReg_6_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_6_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_6_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_6_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_6_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_6_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_6_0_bits_csrInterface_vma <= 1'h0;
      releasePipe_pipe_v_7 <= 1'h0;
      tokenCheck_counter_7 <= 3'h0;
      shifterReg_7_0_valid <= 1'h0;
      shifterReg_7_0_bits_instructionIndex <= 3'h0;
      shifterReg_7_0_bits_decodeResult_specialSlot <= 1'h0;
      shifterReg_7_0_bits_decodeResult_topUop <= 5'h0;
      shifterReg_7_0_bits_decodeResult_popCount <= 1'h0;
      shifterReg_7_0_bits_decodeResult_ffo <= 1'h0;
      shifterReg_7_0_bits_decodeResult_average <= 1'h0;
      shifterReg_7_0_bits_decodeResult_reverse <= 1'h0;
      shifterReg_7_0_bits_decodeResult_dontNeedExecuteInLane <= 1'h0;
      shifterReg_7_0_bits_decodeResult_scheduler <= 1'h0;
      shifterReg_7_0_bits_decodeResult_sReadVD <= 1'h0;
      shifterReg_7_0_bits_decodeResult_vtype <= 1'h0;
      shifterReg_7_0_bits_decodeResult_sWrite <= 1'h0;
      shifterReg_7_0_bits_decodeResult_crossRead <= 1'h0;
      shifterReg_7_0_bits_decodeResult_crossWrite <= 1'h0;
      shifterReg_7_0_bits_decodeResult_maskUnit <= 1'h0;
      shifterReg_7_0_bits_decodeResult_special <= 1'h0;
      shifterReg_7_0_bits_decodeResult_saturate <= 1'h0;
      shifterReg_7_0_bits_decodeResult_vwmacc <= 1'h0;
      shifterReg_7_0_bits_decodeResult_readOnly <= 1'h0;
      shifterReg_7_0_bits_decodeResult_maskSource <= 1'h0;
      shifterReg_7_0_bits_decodeResult_maskDestination <= 1'h0;
      shifterReg_7_0_bits_decodeResult_maskLogic <= 1'h0;
      shifterReg_7_0_bits_decodeResult_uop <= 4'h0;
      shifterReg_7_0_bits_decodeResult_iota <= 1'h0;
      shifterReg_7_0_bits_decodeResult_mv <= 1'h0;
      shifterReg_7_0_bits_decodeResult_extend <= 1'h0;
      shifterReg_7_0_bits_decodeResult_unOrderWrite <= 1'h0;
      shifterReg_7_0_bits_decodeResult_compress <= 1'h0;
      shifterReg_7_0_bits_decodeResult_gather16 <= 1'h0;
      shifterReg_7_0_bits_decodeResult_gather <= 1'h0;
      shifterReg_7_0_bits_decodeResult_slid <= 1'h0;
      shifterReg_7_0_bits_decodeResult_targetRd <= 1'h0;
      shifterReg_7_0_bits_decodeResult_widenReduce <= 1'h0;
      shifterReg_7_0_bits_decodeResult_red <= 1'h0;
      shifterReg_7_0_bits_decodeResult_nr <= 1'h0;
      shifterReg_7_0_bits_decodeResult_itype <= 1'h0;
      shifterReg_7_0_bits_decodeResult_unsigned1 <= 1'h0;
      shifterReg_7_0_bits_decodeResult_unsigned0 <= 1'h0;
      shifterReg_7_0_bits_decodeResult_other <= 1'h0;
      shifterReg_7_0_bits_decodeResult_multiCycle <= 1'h0;
      shifterReg_7_0_bits_decodeResult_divider <= 1'h0;
      shifterReg_7_0_bits_decodeResult_multiplier <= 1'h0;
      shifterReg_7_0_bits_decodeResult_shift <= 1'h0;
      shifterReg_7_0_bits_decodeResult_adder <= 1'h0;
      shifterReg_7_0_bits_decodeResult_logic <= 1'h0;
      shifterReg_7_0_bits_loadStore <= 1'h0;
      shifterReg_7_0_bits_issueInst <= 1'h0;
      shifterReg_7_0_bits_store <= 1'h0;
      shifterReg_7_0_bits_special <= 1'h0;
      shifterReg_7_0_bits_lsWholeReg <= 1'h0;
      shifterReg_7_0_bits_vs1 <= 5'h0;
      shifterReg_7_0_bits_vs2 <= 5'h0;
      shifterReg_7_0_bits_vd <= 5'h0;
      shifterReg_7_0_bits_loadStoreEEW <= 2'h0;
      shifterReg_7_0_bits_mask <= 1'h0;
      shifterReg_7_0_bits_segment <= 3'h0;
      shifterReg_7_0_bits_readFromScalar <= 32'h0;
      shifterReg_7_0_bits_csrInterface_vl <= 12'h0;
      shifterReg_7_0_bits_csrInterface_vStart <= 12'h0;
      shifterReg_7_0_bits_csrInterface_vlmul <= 3'h0;
      shifterReg_7_0_bits_csrInterface_vSew <= 2'h0;
      shifterReg_7_0_bits_csrInterface_vxrm <= 2'h0;
      shifterReg_7_0_bits_csrInterface_vta <= 1'h0;
      shifterReg_7_0_bits_csrInterface_vma <= 1'h0;
      sinkVec_releasePipe_pipe_v <= 1'h0;
      sinkVec_tokenCheck_counter <= 3'h0;
      sinkVec_shifterReg_0_valid <= 1'h0;
      sinkVec_shifterReg_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_1 <= 1'h0;
      sinkVec_tokenCheck_counter_1 <= 3'h0;
      sinkVec_shifterReg_1_0_valid <= 1'h0;
      sinkVec_shifterReg_1_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_1_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_1_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_1_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst <= 1'h0;
      accessDataValid_pipe_v <= 1'h0;
      accessDataValid_pipe_pipe_v <= 1'h0;
      shifterReg_8_0_valid <= 1'h0;
      shifterReg_8_0_bits <= 32'h0;
      accessDataValid_pipe_v_1 <= 1'h0;
      accessDataValid_pipe_pipe_v_1 <= 1'h0;
      shifterReg_9_0_valid <= 1'h0;
      shifterReg_9_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_2 <= 1'h0;
      sinkVec_tokenCheck_counter_2 <= 3'h0;
      sinkVec_shifterReg_2_0_valid <= 1'h0;
      sinkVec_shifterReg_2_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_2_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_2_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_2_0_bits_data <= 32'h0;
      sinkVec_shifterReg_2_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_3 <= 1'h0;
      sinkVec_tokenCheck_counter_3 <= 3'h0;
      sinkVec_shifterReg_3_0_valid <= 1'h0;
      sinkVec_shifterReg_3_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_3_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_3_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_3_0_bits_data <= 32'h0;
      sinkVec_shifterReg_3_0_bits_last <= 1'h0;
      sinkVec_shifterReg_3_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_1 <= 1'h0;
      view__writeRelease_0_pipe_v <= 1'h0;
      pipe_v <= 1'h0;
      instructionFinishedPipe_pipe_v <= 1'h0;
      pipe_v_1 <= 1'h0;
      pipe_pipe_v <= 1'h0;
      view__laneMaskSelect_0_pipe_v <= 1'h0;
      view__laneMaskSelect_0_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_0_pipe_v <= 1'h0;
      view__laneMaskSewSelect_0_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v <= 1'h0;
      maskLastPipe_pipe_v <= 1'h0;
      pipe_v_2 <= 1'h0;
      sinkVec_releasePipe_pipe_v_4 <= 1'h0;
      sinkVec_tokenCheck_counter_4 <= 3'h0;
      sinkVec_shifterReg_4_0_valid <= 1'h0;
      sinkVec_shifterReg_4_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_4_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_4_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_4_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_5 <= 1'h0;
      sinkVec_tokenCheck_counter_5 <= 3'h0;
      sinkVec_shifterReg_5_0_valid <= 1'h0;
      sinkVec_shifterReg_5_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_5_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_5_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_5_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_2 <= 1'h0;
      accessDataValid_pipe_v_2 <= 1'h0;
      accessDataValid_pipe_pipe_v_2 <= 1'h0;
      shifterReg_10_0_valid <= 1'h0;
      shifterReg_10_0_bits <= 32'h0;
      accessDataValid_pipe_v_3 <= 1'h0;
      accessDataValid_pipe_pipe_v_3 <= 1'h0;
      shifterReg_11_0_valid <= 1'h0;
      shifterReg_11_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_6 <= 1'h0;
      sinkVec_tokenCheck_counter_6 <= 3'h0;
      sinkVec_shifterReg_6_0_valid <= 1'h0;
      sinkVec_shifterReg_6_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_6_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_6_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_6_0_bits_data <= 32'h0;
      sinkVec_shifterReg_6_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_7 <= 1'h0;
      sinkVec_tokenCheck_counter_7 <= 3'h0;
      sinkVec_shifterReg_7_0_valid <= 1'h0;
      sinkVec_shifterReg_7_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_7_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_7_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_7_0_bits_data <= 32'h0;
      sinkVec_shifterReg_7_0_bits_last <= 1'h0;
      sinkVec_shifterReg_7_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_3 <= 1'h0;
      view__writeRelease_1_pipe_v <= 1'h0;
      pipe_v_3 <= 1'h0;
      instructionFinishedPipe_pipe_v_1 <= 1'h0;
      pipe_v_4 <= 1'h0;
      pipe_pipe_v_1 <= 1'h0;
      view__laneMaskSelect_1_pipe_v <= 1'h0;
      view__laneMaskSelect_1_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_1_pipe_v <= 1'h0;
      view__laneMaskSewSelect_1_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v_1 <= 1'h0;
      maskLastPipe_pipe_v_1 <= 1'h0;
      pipe_v_5 <= 1'h0;
      sinkVec_releasePipe_pipe_v_8 <= 1'h0;
      sinkVec_tokenCheck_counter_8 <= 3'h0;
      sinkVec_shifterReg_8_0_valid <= 1'h0;
      sinkVec_shifterReg_8_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_8_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_8_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_8_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_9 <= 1'h0;
      sinkVec_tokenCheck_counter_9 <= 3'h0;
      sinkVec_shifterReg_9_0_valid <= 1'h0;
      sinkVec_shifterReg_9_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_9_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_9_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_9_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_4 <= 1'h0;
      accessDataValid_pipe_v_4 <= 1'h0;
      accessDataValid_pipe_pipe_v_4 <= 1'h0;
      shifterReg_12_0_valid <= 1'h0;
      shifterReg_12_0_bits <= 32'h0;
      accessDataValid_pipe_v_5 <= 1'h0;
      accessDataValid_pipe_pipe_v_5 <= 1'h0;
      shifterReg_13_0_valid <= 1'h0;
      shifterReg_13_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_10 <= 1'h0;
      sinkVec_tokenCheck_counter_10 <= 3'h0;
      sinkVec_shifterReg_10_0_valid <= 1'h0;
      sinkVec_shifterReg_10_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_10_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_10_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_10_0_bits_data <= 32'h0;
      sinkVec_shifterReg_10_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_11 <= 1'h0;
      sinkVec_tokenCheck_counter_11 <= 3'h0;
      sinkVec_shifterReg_11_0_valid <= 1'h0;
      sinkVec_shifterReg_11_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_11_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_11_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_11_0_bits_data <= 32'h0;
      sinkVec_shifterReg_11_0_bits_last <= 1'h0;
      sinkVec_shifterReg_11_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_5 <= 1'h0;
      view__writeRelease_2_pipe_v <= 1'h0;
      pipe_v_6 <= 1'h0;
      instructionFinishedPipe_pipe_v_2 <= 1'h0;
      pipe_v_7 <= 1'h0;
      pipe_pipe_v_2 <= 1'h0;
      view__laneMaskSelect_2_pipe_v <= 1'h0;
      view__laneMaskSelect_2_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_2_pipe_v <= 1'h0;
      view__laneMaskSewSelect_2_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v_2 <= 1'h0;
      maskLastPipe_pipe_v_2 <= 1'h0;
      pipe_v_8 <= 1'h0;
      sinkVec_releasePipe_pipe_v_12 <= 1'h0;
      sinkVec_tokenCheck_counter_12 <= 3'h0;
      sinkVec_shifterReg_12_0_valid <= 1'h0;
      sinkVec_shifterReg_12_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_12_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_12_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_12_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_13 <= 1'h0;
      sinkVec_tokenCheck_counter_13 <= 3'h0;
      sinkVec_shifterReg_13_0_valid <= 1'h0;
      sinkVec_shifterReg_13_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_13_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_13_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_13_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_6 <= 1'h0;
      accessDataValid_pipe_v_6 <= 1'h0;
      accessDataValid_pipe_pipe_v_6 <= 1'h0;
      shifterReg_14_0_valid <= 1'h0;
      shifterReg_14_0_bits <= 32'h0;
      accessDataValid_pipe_v_7 <= 1'h0;
      accessDataValid_pipe_pipe_v_7 <= 1'h0;
      shifterReg_15_0_valid <= 1'h0;
      shifterReg_15_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_14 <= 1'h0;
      sinkVec_tokenCheck_counter_14 <= 3'h0;
      sinkVec_shifterReg_14_0_valid <= 1'h0;
      sinkVec_shifterReg_14_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_14_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_14_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_14_0_bits_data <= 32'h0;
      sinkVec_shifterReg_14_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_15 <= 1'h0;
      sinkVec_tokenCheck_counter_15 <= 3'h0;
      sinkVec_shifterReg_15_0_valid <= 1'h0;
      sinkVec_shifterReg_15_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_15_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_15_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_15_0_bits_data <= 32'h0;
      sinkVec_shifterReg_15_0_bits_last <= 1'h0;
      sinkVec_shifterReg_15_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_7 <= 1'h0;
      view__writeRelease_3_pipe_v <= 1'h0;
      pipe_v_9 <= 1'h0;
      instructionFinishedPipe_pipe_v_3 <= 1'h0;
      pipe_v_10 <= 1'h0;
      pipe_pipe_v_3 <= 1'h0;
      view__laneMaskSelect_3_pipe_v <= 1'h0;
      view__laneMaskSelect_3_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_3_pipe_v <= 1'h0;
      view__laneMaskSewSelect_3_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v_3 <= 1'h0;
      maskLastPipe_pipe_v_3 <= 1'h0;
      pipe_v_11 <= 1'h0;
      sinkVec_releasePipe_pipe_v_16 <= 1'h0;
      sinkVec_tokenCheck_counter_16 <= 3'h0;
      sinkVec_shifterReg_16_0_valid <= 1'h0;
      sinkVec_shifterReg_16_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_16_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_16_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_16_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_17 <= 1'h0;
      sinkVec_tokenCheck_counter_17 <= 3'h0;
      sinkVec_shifterReg_17_0_valid <= 1'h0;
      sinkVec_shifterReg_17_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_17_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_17_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_17_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_8 <= 1'h0;
      accessDataValid_pipe_v_8 <= 1'h0;
      accessDataValid_pipe_pipe_v_8 <= 1'h0;
      shifterReg_16_0_valid <= 1'h0;
      shifterReg_16_0_bits <= 32'h0;
      accessDataValid_pipe_v_9 <= 1'h0;
      accessDataValid_pipe_pipe_v_9 <= 1'h0;
      shifterReg_17_0_valid <= 1'h0;
      shifterReg_17_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_18 <= 1'h0;
      sinkVec_tokenCheck_counter_18 <= 3'h0;
      sinkVec_shifterReg_18_0_valid <= 1'h0;
      sinkVec_shifterReg_18_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_18_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_18_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_18_0_bits_data <= 32'h0;
      sinkVec_shifterReg_18_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_19 <= 1'h0;
      sinkVec_tokenCheck_counter_19 <= 3'h0;
      sinkVec_shifterReg_19_0_valid <= 1'h0;
      sinkVec_shifterReg_19_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_19_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_19_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_19_0_bits_data <= 32'h0;
      sinkVec_shifterReg_19_0_bits_last <= 1'h0;
      sinkVec_shifterReg_19_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_9 <= 1'h0;
      view__writeRelease_4_pipe_v <= 1'h0;
      pipe_v_12 <= 1'h0;
      instructionFinishedPipe_pipe_v_4 <= 1'h0;
      pipe_v_13 <= 1'h0;
      pipe_pipe_v_4 <= 1'h0;
      view__laneMaskSelect_4_pipe_v <= 1'h0;
      view__laneMaskSelect_4_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_4_pipe_v <= 1'h0;
      view__laneMaskSewSelect_4_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v_4 <= 1'h0;
      maskLastPipe_pipe_v_4 <= 1'h0;
      pipe_v_14 <= 1'h0;
      sinkVec_releasePipe_pipe_v_20 <= 1'h0;
      sinkVec_tokenCheck_counter_20 <= 3'h0;
      sinkVec_shifterReg_20_0_valid <= 1'h0;
      sinkVec_shifterReg_20_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_20_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_20_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_20_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_21 <= 1'h0;
      sinkVec_tokenCheck_counter_21 <= 3'h0;
      sinkVec_shifterReg_21_0_valid <= 1'h0;
      sinkVec_shifterReg_21_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_21_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_21_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_21_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_10 <= 1'h0;
      accessDataValid_pipe_v_10 <= 1'h0;
      accessDataValid_pipe_pipe_v_10 <= 1'h0;
      shifterReg_18_0_valid <= 1'h0;
      shifterReg_18_0_bits <= 32'h0;
      accessDataValid_pipe_v_11 <= 1'h0;
      accessDataValid_pipe_pipe_v_11 <= 1'h0;
      shifterReg_19_0_valid <= 1'h0;
      shifterReg_19_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_22 <= 1'h0;
      sinkVec_tokenCheck_counter_22 <= 3'h0;
      sinkVec_shifterReg_22_0_valid <= 1'h0;
      sinkVec_shifterReg_22_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_22_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_22_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_22_0_bits_data <= 32'h0;
      sinkVec_shifterReg_22_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_23 <= 1'h0;
      sinkVec_tokenCheck_counter_23 <= 3'h0;
      sinkVec_shifterReg_23_0_valid <= 1'h0;
      sinkVec_shifterReg_23_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_23_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_23_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_23_0_bits_data <= 32'h0;
      sinkVec_shifterReg_23_0_bits_last <= 1'h0;
      sinkVec_shifterReg_23_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_11 <= 1'h0;
      view__writeRelease_5_pipe_v <= 1'h0;
      pipe_v_15 <= 1'h0;
      instructionFinishedPipe_pipe_v_5 <= 1'h0;
      pipe_v_16 <= 1'h0;
      pipe_pipe_v_5 <= 1'h0;
      view__laneMaskSelect_5_pipe_v <= 1'h0;
      view__laneMaskSelect_5_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_5_pipe_v <= 1'h0;
      view__laneMaskSewSelect_5_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v_5 <= 1'h0;
      maskLastPipe_pipe_v_5 <= 1'h0;
      pipe_v_17 <= 1'h0;
      sinkVec_releasePipe_pipe_v_24 <= 1'h0;
      sinkVec_tokenCheck_counter_24 <= 3'h0;
      sinkVec_shifterReg_24_0_valid <= 1'h0;
      sinkVec_shifterReg_24_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_24_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_24_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_24_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_25 <= 1'h0;
      sinkVec_tokenCheck_counter_25 <= 3'h0;
      sinkVec_shifterReg_25_0_valid <= 1'h0;
      sinkVec_shifterReg_25_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_25_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_25_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_25_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_12 <= 1'h0;
      accessDataValid_pipe_v_12 <= 1'h0;
      accessDataValid_pipe_pipe_v_12 <= 1'h0;
      shifterReg_20_0_valid <= 1'h0;
      shifterReg_20_0_bits <= 32'h0;
      accessDataValid_pipe_v_13 <= 1'h0;
      accessDataValid_pipe_pipe_v_13 <= 1'h0;
      shifterReg_21_0_valid <= 1'h0;
      shifterReg_21_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_26 <= 1'h0;
      sinkVec_tokenCheck_counter_26 <= 3'h0;
      sinkVec_shifterReg_26_0_valid <= 1'h0;
      sinkVec_shifterReg_26_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_26_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_26_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_26_0_bits_data <= 32'h0;
      sinkVec_shifterReg_26_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_27 <= 1'h0;
      sinkVec_tokenCheck_counter_27 <= 3'h0;
      sinkVec_shifterReg_27_0_valid <= 1'h0;
      sinkVec_shifterReg_27_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_27_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_27_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_27_0_bits_data <= 32'h0;
      sinkVec_shifterReg_27_0_bits_last <= 1'h0;
      sinkVec_shifterReg_27_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_13 <= 1'h0;
      view__writeRelease_6_pipe_v <= 1'h0;
      pipe_v_18 <= 1'h0;
      instructionFinishedPipe_pipe_v_6 <= 1'h0;
      pipe_v_19 <= 1'h0;
      pipe_pipe_v_6 <= 1'h0;
      view__laneMaskSelect_6_pipe_v <= 1'h0;
      view__laneMaskSelect_6_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_6_pipe_v <= 1'h0;
      view__laneMaskSewSelect_6_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v_6 <= 1'h0;
      maskLastPipe_pipe_v_6 <= 1'h0;
      pipe_v_20 <= 1'h0;
      sinkVec_releasePipe_pipe_v_28 <= 1'h0;
      sinkVec_tokenCheck_counter_28 <= 3'h0;
      sinkVec_shifterReg_28_0_valid <= 1'h0;
      sinkVec_shifterReg_28_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_28_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_28_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_28_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_29 <= 1'h0;
      sinkVec_tokenCheck_counter_29 <= 3'h0;
      sinkVec_shifterReg_29_0_valid <= 1'h0;
      sinkVec_shifterReg_29_0_bits_vs <= 5'h0;
      sinkVec_shifterReg_29_0_bits_readSource <= 2'h0;
      sinkVec_shifterReg_29_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_29_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_14 <= 1'h0;
      accessDataValid_pipe_v_14 <= 1'h0;
      accessDataValid_pipe_pipe_v_14 <= 1'h0;
      shifterReg_22_0_valid <= 1'h0;
      shifterReg_22_0_bits <= 32'h0;
      accessDataValid_pipe_v_15 <= 1'h0;
      accessDataValid_pipe_pipe_v_15 <= 1'h0;
      shifterReg_23_0_valid <= 1'h0;
      shifterReg_23_0_bits <= 32'h0;
      sinkVec_releasePipe_pipe_v_30 <= 1'h0;
      sinkVec_tokenCheck_counter_30 <= 3'h0;
      sinkVec_shifterReg_30_0_valid <= 1'h0;
      sinkVec_shifterReg_30_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_30_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_30_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_30_0_bits_data <= 32'h0;
      sinkVec_shifterReg_30_0_bits_instructionIndex <= 3'h0;
      sinkVec_releasePipe_pipe_v_31 <= 1'h0;
      sinkVec_tokenCheck_counter_31 <= 3'h0;
      sinkVec_shifterReg_31_0_valid <= 1'h0;
      sinkVec_shifterReg_31_0_bits_vd <= 5'h0;
      sinkVec_shifterReg_31_0_bits_offset <= 3'h0;
      sinkVec_shifterReg_31_0_bits_mask <= 4'h0;
      sinkVec_shifterReg_31_0_bits_data <= 32'h0;
      sinkVec_shifterReg_31_0_bits_last <= 1'h0;
      sinkVec_shifterReg_31_0_bits_instructionIndex <= 3'h0;
      maskUnitFirst_15 <= 1'h0;
      view__writeRelease_7_pipe_v <= 1'h0;
      pipe_v_21 <= 1'h0;
      instructionFinishedPipe_pipe_v_7 <= 1'h0;
      pipe_v_22 <= 1'h0;
      pipe_pipe_v_7 <= 1'h0;
      view__laneMaskSelect_7_pipe_v <= 1'h0;
      view__laneMaskSelect_7_pipe_pipe_v <= 1'h0;
      view__laneMaskSewSelect_7_pipe_v <= 1'h0;
      view__laneMaskSewSelect_7_pipe_pipe_v <= 1'h0;
      lsuLastPipe_pipe_v_7 <= 1'h0;
      maskLastPipe_pipe_v_7 <= 1'h0;
      pipe_v_23 <= 1'h0;
      pipe_v_24 <= 1'h0;
      shifterReg_24_0_valid <= 1'h0;
      shifterReg_24_0_bits_data <= 32'h0;
      pipe_v_25 <= 1'h0;
      shifterReg_25_0_valid <= 1'h0;
      shifterReg_25_0_bits_data <= 32'h0;
      shifterReg_25_0_bits_mask <= 2'h0;
      shifterReg_25_0_bits_instructionIndex <= 3'h0;
      shifterReg_25_0_bits_counter <= 7'h0;
      pipe_v_26 <= 1'h0;
      shifterReg_26_0_valid <= 1'h0;
      shifterReg_26_0_bits_data <= 32'h0;
      pipe_v_27 <= 1'h0;
      shifterReg_27_0_valid <= 1'h0;
      shifterReg_27_0_bits_data <= 32'h0;
      shifterReg_27_0_bits_mask <= 2'h0;
      shifterReg_27_0_bits_instructionIndex <= 3'h0;
      shifterReg_27_0_bits_counter <= 7'h0;
      pipe_v_28 <= 1'h0;
      shifterReg_28_0_valid <= 1'h0;
      shifterReg_28_0_bits_data <= 32'h0;
      pipe_v_29 <= 1'h0;
      shifterReg_29_0_valid <= 1'h0;
      shifterReg_29_0_bits_data <= 32'h0;
      shifterReg_29_0_bits_mask <= 2'h0;
      shifterReg_29_0_bits_instructionIndex <= 3'h0;
      shifterReg_29_0_bits_counter <= 7'h0;
      pipe_v_30 <= 1'h0;
      shifterReg_30_0_valid <= 1'h0;
      shifterReg_30_0_bits_data <= 32'h0;
      pipe_v_31 <= 1'h0;
      shifterReg_31_0_valid <= 1'h0;
      shifterReg_31_0_bits_data <= 32'h0;
      shifterReg_31_0_bits_mask <= 2'h0;
      shifterReg_31_0_bits_instructionIndex <= 3'h0;
      shifterReg_31_0_bits_counter <= 7'h0;
      pipe_v_32 <= 1'h0;
      shifterReg_32_0_valid <= 1'h0;
      shifterReg_32_0_bits_data <= 32'h0;
      pipe_v_33 <= 1'h0;
      shifterReg_33_0_valid <= 1'h0;
      shifterReg_33_0_bits_data <= 32'h0;
      shifterReg_33_0_bits_mask <= 2'h0;
      shifterReg_33_0_bits_instructionIndex <= 3'h0;
      shifterReg_33_0_bits_counter <= 7'h0;
      pipe_v_34 <= 1'h0;
      shifterReg_34_0_valid <= 1'h0;
      shifterReg_34_0_bits_data <= 32'h0;
      pipe_v_35 <= 1'h0;
      shifterReg_35_0_valid <= 1'h0;
      shifterReg_35_0_bits_data <= 32'h0;
      shifterReg_35_0_bits_mask <= 2'h0;
      shifterReg_35_0_bits_instructionIndex <= 3'h0;
      shifterReg_35_0_bits_counter <= 7'h0;
      pipe_v_36 <= 1'h0;
      shifterReg_36_0_valid <= 1'h0;
      shifterReg_36_0_bits_data <= 32'h0;
      pipe_v_37 <= 1'h0;
      shifterReg_37_0_valid <= 1'h0;
      shifterReg_37_0_bits_data <= 32'h0;
      shifterReg_37_0_bits_mask <= 2'h0;
      shifterReg_37_0_bits_instructionIndex <= 3'h0;
      shifterReg_37_0_bits_counter <= 7'h0;
      pipe_v_38 <= 1'h0;
      shifterReg_38_0_valid <= 1'h0;
      shifterReg_38_0_bits_data <= 32'h0;
      pipe_v_39 <= 1'h0;
      shifterReg_39_0_valid <= 1'h0;
      shifterReg_39_0_bits_data <= 32'h0;
      shifterReg_39_0_bits_mask <= 2'h0;
      shifterReg_39_0_bits_instructionIndex <= 3'h0;
      shifterReg_39_0_bits_counter <= 7'h0;
      pipe_v_40 <= 1'h0;
      shifterReg_40_0_valid <= 1'h0;
      shifterReg_40_0_bits_data <= 32'h0;
      pipe_v_41 <= 1'h0;
      shifterReg_41_0_valid <= 1'h0;
      shifterReg_41_0_bits_data <= 32'h0;
      shifterReg_41_0_bits_mask <= 2'h0;
      shifterReg_41_0_bits_instructionIndex <= 3'h0;
      shifterReg_41_0_bits_counter <= 7'h0;
      pipe_v_42 <= 1'h0;
      shifterReg_42_0_valid <= 1'h0;
      shifterReg_42_0_bits_data <= 32'h0;
      pipe_v_43 <= 1'h0;
      shifterReg_43_0_valid <= 1'h0;
      shifterReg_43_0_bits_data <= 32'h0;
      shifterReg_43_0_bits_mask <= 2'h0;
      shifterReg_43_0_bits_instructionIndex <= 3'h0;
      shifterReg_43_0_bits_counter <= 7'h0;
      pipe_v_44 <= 1'h0;
      shifterReg_44_0_valid <= 1'h0;
      shifterReg_44_0_bits_data <= 32'h0;
      pipe_v_45 <= 1'h0;
      shifterReg_45_0_valid <= 1'h0;
      shifterReg_45_0_bits_data <= 32'h0;
      shifterReg_45_0_bits_mask <= 2'h0;
      shifterReg_45_0_bits_instructionIndex <= 3'h0;
      shifterReg_45_0_bits_counter <= 7'h0;
      pipe_v_46 <= 1'h0;
      shifterReg_46_0_valid <= 1'h0;
      shifterReg_46_0_bits_data <= 32'h0;
      pipe_v_47 <= 1'h0;
      shifterReg_47_0_valid <= 1'h0;
      shifterReg_47_0_bits_data <= 32'h0;
      shifterReg_47_0_bits_mask <= 2'h0;
      shifterReg_47_0_bits_instructionIndex <= 3'h0;
      shifterReg_47_0_bits_counter <= 7'h0;
      pipe_v_48 <= 1'h0;
      shifterReg_48_0_valid <= 1'h0;
      shifterReg_48_0_bits_data <= 32'h0;
      pipe_v_49 <= 1'h0;
      shifterReg_49_0_valid <= 1'h0;
      shifterReg_49_0_bits_data <= 32'h0;
      shifterReg_49_0_bits_mask <= 2'h0;
      shifterReg_49_0_bits_instructionIndex <= 3'h0;
      shifterReg_49_0_bits_counter <= 7'h0;
      pipe_v_50 <= 1'h0;
      shifterReg_50_0_valid <= 1'h0;
      shifterReg_50_0_bits_data <= 32'h0;
      pipe_v_51 <= 1'h0;
      shifterReg_51_0_valid <= 1'h0;
      shifterReg_51_0_bits_data <= 32'h0;
      shifterReg_51_0_bits_mask <= 2'h0;
      shifterReg_51_0_bits_instructionIndex <= 3'h0;
      shifterReg_51_0_bits_counter <= 7'h0;
      pipe_v_52 <= 1'h0;
      shifterReg_52_0_valid <= 1'h0;
      shifterReg_52_0_bits_data <= 32'h0;
      pipe_v_53 <= 1'h0;
      shifterReg_53_0_valid <= 1'h0;
      shifterReg_53_0_bits_data <= 32'h0;
      shifterReg_53_0_bits_mask <= 2'h0;
      shifterReg_53_0_bits_instructionIndex <= 3'h0;
      shifterReg_53_0_bits_counter <= 7'h0;
      pipe_v_54 <= 1'h0;
      shifterReg_54_0_valid <= 1'h0;
      shifterReg_54_0_bits_data <= 32'h0;
      pipe_v_55 <= 1'h0;
      shifterReg_55_0_valid <= 1'h0;
      shifterReg_55_0_bits_data <= 32'h0;
      shifterReg_55_0_bits_mask <= 2'h0;
      shifterReg_55_0_bits_instructionIndex <= 3'h0;
      shifterReg_55_0_bits_counter <= 7'h0;
    end
    else begin
      if (_probeWire_issue_valid_T) begin
        automatic logic [38:0] _requestReg_bits_writeByte_T_8 = {7'h0, issue_bits_vl_0} << issue_bits_vtype_0[5:3] + {2'h0, _decode_decodeResult_crossWrite};
        instructionCounter <= nextInstructionCounter;
        requestReg_bits_issue_instruction <= issue_bits_instruction_0;
        requestReg_bits_issue_rs1Data <= issue_bits_rs1Data_0;
        requestReg_bits_issue_rs2Data <= issue_bits_rs2Data_0;
        requestReg_bits_issue_vtype <= issue_bits_vtype_0;
        requestReg_bits_issue_vl <= issue_bits_vl_0;
        requestReg_bits_issue_vstart <= issue_bits_vstart_0;
        requestReg_bits_issue_vcsr <= issue_bits_vcsr_0;
        requestReg_bits_decodeResult_specialSlot <= _decode_decodeResult_specialSlot;
        requestReg_bits_decodeResult_topUop <= _decode_decodeResult_topUop;
        requestReg_bits_decodeResult_popCount <= _decode_decodeResult_popCount;
        requestReg_bits_decodeResult_ffo <= _decode_decodeResult_ffo;
        requestReg_bits_decodeResult_average <= _decode_decodeResult_average;
        requestReg_bits_decodeResult_reverse <= _decode_decodeResult_reverse;
        requestReg_bits_decodeResult_dontNeedExecuteInLane <= _decode_decodeResult_dontNeedExecuteInLane;
        requestReg_bits_decodeResult_scheduler <= _decode_decodeResult_scheduler;
        requestReg_bits_decodeResult_sReadVD <= _decode_decodeResult_sReadVD;
        requestReg_bits_decodeResult_vtype <= _decode_decodeResult_vtype;
        requestReg_bits_decodeResult_sWrite <= _decode_decodeResult_sWrite;
        requestReg_bits_decodeResult_crossRead <= _decode_decodeResult_crossRead;
        requestReg_bits_decodeResult_crossWrite <= _decode_decodeResult_crossWrite;
        requestReg_bits_decodeResult_maskUnit <= _decode_decodeResult_maskUnit;
        requestReg_bits_decodeResult_special <= _decode_decodeResult_special;
        requestReg_bits_decodeResult_saturate <= _decode_decodeResult_saturate;
        requestReg_bits_decodeResult_vwmacc <= _decode_decodeResult_vwmacc;
        requestReg_bits_decodeResult_readOnly <= _decode_decodeResult_readOnly;
        requestReg_bits_decodeResult_maskSource <= _decode_decodeResult_maskSource;
        requestReg_bits_decodeResult_maskDestination <= _decode_decodeResult_maskDestination;
        requestReg_bits_decodeResult_maskLogic <= _decode_decodeResult_maskLogic;
        requestReg_bits_decodeResult_uop <= _decode_decodeResult_uop;
        requestReg_bits_decodeResult_iota <= _decode_decodeResult_iota;
        requestReg_bits_decodeResult_mv <= _decode_decodeResult_mv;
        requestReg_bits_decodeResult_extend <= _decode_decodeResult_extend;
        requestReg_bits_decodeResult_unOrderWrite <= _decode_decodeResult_unOrderWrite;
        requestReg_bits_decodeResult_compress <= _decode_decodeResult_compress;
        requestReg_bits_decodeResult_gather16 <= _decode_decodeResult_gather16;
        requestReg_bits_decodeResult_gather <= _decode_decodeResult_gather;
        requestReg_bits_decodeResult_slid <= _decode_decodeResult_slid;
        requestReg_bits_decodeResult_targetRd <= _decode_decodeResult_targetRd;
        requestReg_bits_decodeResult_widenReduce <= _decode_decodeResult_widenReduce;
        requestReg_bits_decodeResult_red <= _decode_decodeResult_red;
        requestReg_bits_decodeResult_nr <= _decode_decodeResult_nr;
        requestReg_bits_decodeResult_itype <= _decode_decodeResult_itype;
        requestReg_bits_decodeResult_unsigned1 <= _decode_decodeResult_unsigned1;
        requestReg_bits_decodeResult_unsigned0 <= _decode_decodeResult_unsigned0;
        requestReg_bits_decodeResult_other <= _decode_decodeResult_other;
        requestReg_bits_decodeResult_multiCycle <= _decode_decodeResult_multiCycle;
        requestReg_bits_decodeResult_divider <= _decode_decodeResult_divider;
        requestReg_bits_decodeResult_multiplier <= _decode_decodeResult_multiplier;
        requestReg_bits_decodeResult_shift <= _decode_decodeResult_shift;
        requestReg_bits_decodeResult_adder <= _decode_decodeResult_adder;
        requestReg_bits_decodeResult_logic <= _decode_decodeResult_logic;
        requestReg_bits_instructionIndex <= instructionCounter;
        requestReg_bits_vdIsV0 <= issue_bits_instruction_0[11:7] == 5'h0 & (issue_bits_instruction_0[6] | ~(issue_bits_instruction_0[5]));
        requestReg_bits_writeByte <= _decode_decodeResult_red ? 12'h1 : _decode_decodeResult_maskDestination ? issue_bits_vl_0[14:3] + {11'h0, |(issue_bits_vl_0[2:0])} : _requestReg_bits_writeByte_T_8[11:0];
      end
      if (retire_1)
        responseCounter <= nextResponseCounter;
      if (_probeWire_issue_valid_T ^ maskUnit_gatherData_ready)
        requestReg_valid <= _probeWire_issue_valid_T;
      if (instructionToSlotOH[0]) begin
        slots_0_record_instructionIndex <= requestReg_bits_instructionIndex;
        slots_0_record_isLoadStore <= isLoadStoreType;
        slots_0_record_maskType <= maskType;
      end
      slots_0_state_wLast <= ~(instructionToSlotOH[0]) & (slots_laneAndLSUFinish & slots_v0WriteFinish | slots_0_state_wLast);
      slots_0_state_idle <= ~(instructionToSlotOH[0]) & (slots_0_state_sCommit & slots_0_state_wVRFWrite & slots_0_state_wMaskUnitLast | slots_0_state_idle);
      slots_0_state_wMaskUnitLast <= instructionToSlotOH[0] ? ~requestReg_bits_decodeResult_maskUnit : (|_maskUnit_lastReport) | slots_0_state_wMaskUnitLast;
      slots_0_state_wVRFWrite <= instructionToSlotOH[0] ? ~requestReg_bits_decodeResult_maskUnit : slots_0_state_wLast & slots_0_state_wMaskUnitLast & ~slots_dataInWritePipeCheck | slots_0_state_wVRFWrite;
      slots_0_state_sCommit <= ~(instructionToSlotOH[0]) & (responseCounter == slots_0_record_instructionIndex & retire_1 | slots_0_state_sCommit);
      slots_0_endTag_0 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_0 | instructionFinished_0_0;
      slots_0_endTag_1 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_1 | instructionFinished_1_0;
      slots_0_endTag_2 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_2 | instructionFinished_2_0;
      slots_0_endTag_3 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_3 | instructionFinished_3_0;
      slots_0_endTag_4 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_4 | instructionFinished_4_0;
      slots_0_endTag_5 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_5 | instructionFinished_5_0;
      slots_0_endTag_6 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_6 | instructionFinished_6_0;
      slots_0_endTag_7 <= instructionToSlotOH[0] ? skipLastFromLane : slots_0_endTag_7 | instructionFinished_7_0;
      slots_0_endTag_8 <= instructionToSlotOH[0] ? ~isLoadStoreType : slots_0_endTag_8 | slots_lsuFinished;
      slots_0_vxsat <= ~(instructionToSlotOH[0]) & (slots_vxsatUpdate | slots_0_vxsat);
      if (instructionToSlotOH[1]) begin
        slots_1_record_instructionIndex <= requestReg_bits_instructionIndex;
        slots_1_record_isLoadStore <= isLoadStoreType;
        slots_1_record_maskType <= maskType;
      end
      slots_1_state_wLast <= ~(instructionToSlotOH[1]) & (slots_laneAndLSUFinish_1 & slots_v0WriteFinish_1 | slots_1_state_wLast);
      slots_1_state_idle <= ~(instructionToSlotOH[1]) & (slots_1_state_sCommit & slots_1_state_wVRFWrite & slots_1_state_wMaskUnitLast | slots_1_state_idle);
      slots_1_state_wMaskUnitLast <= instructionToSlotOH[1] ? ~requestReg_bits_decodeResult_maskUnit : (|_maskUnit_lastReport) | slots_1_state_wMaskUnitLast;
      slots_1_state_wVRFWrite <= instructionToSlotOH[1] ? ~requestReg_bits_decodeResult_maskUnit : slots_1_state_wLast & slots_1_state_wMaskUnitLast & ~slots_dataInWritePipeCheck_1 | slots_1_state_wVRFWrite;
      slots_1_state_sCommit <= ~(instructionToSlotOH[1]) & (responseCounter == slots_1_record_instructionIndex & retire_1 | slots_1_state_sCommit);
      slots_1_endTag_0 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_0 | instructionFinished_0_1;
      slots_1_endTag_1 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_1 | instructionFinished_1_1;
      slots_1_endTag_2 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_2 | instructionFinished_2_1;
      slots_1_endTag_3 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_3 | instructionFinished_3_1;
      slots_1_endTag_4 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_4 | instructionFinished_4_1;
      slots_1_endTag_5 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_5 | instructionFinished_5_1;
      slots_1_endTag_6 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_6 | instructionFinished_6_1;
      slots_1_endTag_7 <= instructionToSlotOH[1] ? skipLastFromLane : slots_1_endTag_7 | instructionFinished_7_1;
      slots_1_endTag_8 <= instructionToSlotOH[1] ? ~isLoadStoreType : slots_1_endTag_8 | slots_lsuFinished_1;
      slots_1_vxsat <= ~(instructionToSlotOH[1]) & (slots_vxsatUpdate_1 | slots_1_vxsat);
      if (instructionToSlotOH[2]) begin
        slots_2_record_instructionIndex <= requestReg_bits_instructionIndex;
        slots_2_record_isLoadStore <= isLoadStoreType;
        slots_2_record_maskType <= maskType;
      end
      slots_2_state_wLast <= ~(instructionToSlotOH[2]) & (slots_laneAndLSUFinish_2 & slots_v0WriteFinish_2 | slots_2_state_wLast);
      slots_2_state_idle <= ~(instructionToSlotOH[2]) & (slots_2_state_sCommit & slots_2_state_wVRFWrite & slots_2_state_wMaskUnitLast | slots_2_state_idle);
      slots_2_state_wMaskUnitLast <= instructionToSlotOH[2] ? ~requestReg_bits_decodeResult_maskUnit : (|_maskUnit_lastReport) | slots_2_state_wMaskUnitLast;
      slots_2_state_wVRFWrite <= instructionToSlotOH[2] ? ~requestReg_bits_decodeResult_maskUnit : slots_2_state_wLast & slots_2_state_wMaskUnitLast & ~slots_dataInWritePipeCheck_2 | slots_2_state_wVRFWrite;
      slots_2_state_sCommit <= ~(instructionToSlotOH[2]) & (responseCounter == slots_2_record_instructionIndex & retire_1 | slots_2_state_sCommit);
      slots_2_endTag_0 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_0 | instructionFinished_0_2;
      slots_2_endTag_1 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_1 | instructionFinished_1_2;
      slots_2_endTag_2 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_2 | instructionFinished_2_2;
      slots_2_endTag_3 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_3 | instructionFinished_3_2;
      slots_2_endTag_4 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_4 | instructionFinished_4_2;
      slots_2_endTag_5 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_5 | instructionFinished_5_2;
      slots_2_endTag_6 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_6 | instructionFinished_6_2;
      slots_2_endTag_7 <= instructionToSlotOH[2] ? skipLastFromLane : slots_2_endTag_7 | instructionFinished_7_2;
      slots_2_endTag_8 <= instructionToSlotOH[2] ? ~isLoadStoreType : slots_2_endTag_8 | slots_lsuFinished_2;
      slots_2_vxsat <= ~(instructionToSlotOH[2]) & (slots_vxsatUpdate_2 | slots_2_vxsat);
      if (instructionToSlotOH[3]) begin
        slots_3_record_instructionIndex <= requestReg_bits_instructionIndex;
        slots_3_record_isLoadStore <= isLoadStoreType;
        slots_3_record_maskType <= maskType;
        slots_writeRD <= requestReg_bits_decodeResult_targetRd;
        slots_vd <= requestRegDequeue_bits_instruction[11:7];
      end
      slots_3_state_wLast <= ~(instructionToSlotOH[3]) & (slots_laneAndLSUFinish_3 & slots_v0WriteFinish_3 | slots_3_state_wLast);
      slots_3_state_idle <= ~(instructionToSlotOH[3]) & (slots_3_state_sCommit & slots_3_state_wVRFWrite & slots_3_state_wMaskUnitLast | slots_3_state_idle);
      slots_3_state_wMaskUnitLast <= instructionToSlotOH[3] ? ~requestReg_bits_decodeResult_maskUnit : (|_maskUnit_lastReport) | slots_3_state_wMaskUnitLast;
      slots_3_state_wVRFWrite <= instructionToSlotOH[3] ? ~requestReg_bits_decodeResult_maskUnit : slots_3_state_wLast & slots_3_state_wMaskUnitLast & ~slots_dataInWritePipeCheck_3 | slots_3_state_wVRFWrite;
      slots_3_state_sCommit <= ~(instructionToSlotOH[3]) & (responseCounter == slots_3_record_instructionIndex & retire_1 | slots_3_state_sCommit);
      slots_3_endTag_0 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_0 | instructionFinished_0_3;
      slots_3_endTag_1 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_1 | instructionFinished_1_3;
      slots_3_endTag_2 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_2 | instructionFinished_2_3;
      slots_3_endTag_3 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_3 | instructionFinished_3_3;
      slots_3_endTag_4 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_4 | instructionFinished_4_3;
      slots_3_endTag_5 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_5 | instructionFinished_5_3;
      slots_3_endTag_6 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_6 | instructionFinished_6_3;
      slots_3_endTag_7 <= instructionToSlotOH[3] ? skipLastFromLane : slots_3_endTag_7 | instructionFinished_7_3;
      slots_3_endTag_8 <= instructionToSlotOH[3] ? ~isLoadStoreType : slots_3_endTag_8 | slots_lsuFinished_3;
      slots_3_vxsat <= ~(instructionToSlotOH[3]) & (slots_vxsatUpdate_3 | slots_3_vxsat);
      releasePipe_pipe_v <= laneVec_0_laneRequest_bits_issueInst;
      if (validSource_valid ^ releasePipe_pipe_out_valid)
        tokenCheck_counter <= tokenCheck_counter + tokenCheck_counterChange;
      if (shifterValid) begin
        shifterReg_0_valid <= validSource_valid;
        shifterReg_0_bits_instructionIndex <= validSource_bits_instructionIndex;
        shifterReg_0_bits_decodeResult_specialSlot <= validSource_bits_decodeResult_specialSlot;
        shifterReg_0_bits_decodeResult_topUop <= validSource_bits_decodeResult_topUop;
        shifterReg_0_bits_decodeResult_popCount <= validSource_bits_decodeResult_popCount;
        shifterReg_0_bits_decodeResult_ffo <= validSource_bits_decodeResult_ffo;
        shifterReg_0_bits_decodeResult_average <= validSource_bits_decodeResult_average;
        shifterReg_0_bits_decodeResult_reverse <= validSource_bits_decodeResult_reverse;
        shifterReg_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_0_bits_decodeResult_scheduler <= validSource_bits_decodeResult_scheduler;
        shifterReg_0_bits_decodeResult_sReadVD <= validSource_bits_decodeResult_sReadVD;
        shifterReg_0_bits_decodeResult_vtype <= validSource_bits_decodeResult_vtype;
        shifterReg_0_bits_decodeResult_sWrite <= validSource_bits_decodeResult_sWrite;
        shifterReg_0_bits_decodeResult_crossRead <= validSource_bits_decodeResult_crossRead;
        shifterReg_0_bits_decodeResult_crossWrite <= validSource_bits_decodeResult_crossWrite;
        shifterReg_0_bits_decodeResult_maskUnit <= validSource_bits_decodeResult_maskUnit;
        shifterReg_0_bits_decodeResult_special <= validSource_bits_decodeResult_special;
        shifterReg_0_bits_decodeResult_saturate <= validSource_bits_decodeResult_saturate;
        shifterReg_0_bits_decodeResult_vwmacc <= validSource_bits_decodeResult_vwmacc;
        shifterReg_0_bits_decodeResult_readOnly <= validSource_bits_decodeResult_readOnly;
        shifterReg_0_bits_decodeResult_maskSource <= validSource_bits_decodeResult_maskSource;
        shifterReg_0_bits_decodeResult_maskDestination <= validSource_bits_decodeResult_maskDestination;
        shifterReg_0_bits_decodeResult_maskLogic <= validSource_bits_decodeResult_maskLogic;
        shifterReg_0_bits_decodeResult_uop <= validSource_bits_decodeResult_uop;
        shifterReg_0_bits_decodeResult_iota <= validSource_bits_decodeResult_iota;
        shifterReg_0_bits_decodeResult_mv <= validSource_bits_decodeResult_mv;
        shifterReg_0_bits_decodeResult_extend <= validSource_bits_decodeResult_extend;
        shifterReg_0_bits_decodeResult_unOrderWrite <= validSource_bits_decodeResult_unOrderWrite;
        shifterReg_0_bits_decodeResult_compress <= validSource_bits_decodeResult_compress;
        shifterReg_0_bits_decodeResult_gather16 <= validSource_bits_decodeResult_gather16;
        shifterReg_0_bits_decodeResult_gather <= validSource_bits_decodeResult_gather;
        shifterReg_0_bits_decodeResult_slid <= validSource_bits_decodeResult_slid;
        shifterReg_0_bits_decodeResult_targetRd <= validSource_bits_decodeResult_targetRd;
        shifterReg_0_bits_decodeResult_widenReduce <= validSource_bits_decodeResult_widenReduce;
        shifterReg_0_bits_decodeResult_red <= validSource_bits_decodeResult_red;
        shifterReg_0_bits_decodeResult_nr <= validSource_bits_decodeResult_nr;
        shifterReg_0_bits_decodeResult_itype <= validSource_bits_decodeResult_itype;
        shifterReg_0_bits_decodeResult_unsigned1 <= validSource_bits_decodeResult_unsigned1;
        shifterReg_0_bits_decodeResult_unsigned0 <= validSource_bits_decodeResult_unsigned0;
        shifterReg_0_bits_decodeResult_other <= validSource_bits_decodeResult_other;
        shifterReg_0_bits_decodeResult_multiCycle <= validSource_bits_decodeResult_multiCycle;
        shifterReg_0_bits_decodeResult_divider <= validSource_bits_decodeResult_divider;
        shifterReg_0_bits_decodeResult_multiplier <= validSource_bits_decodeResult_multiplier;
        shifterReg_0_bits_decodeResult_shift <= validSource_bits_decodeResult_shift;
        shifterReg_0_bits_decodeResult_adder <= validSource_bits_decodeResult_adder;
        shifterReg_0_bits_decodeResult_logic <= validSource_bits_decodeResult_logic;
        shifterReg_0_bits_loadStore <= validSource_bits_loadStore;
        shifterReg_0_bits_issueInst <= validSource_bits_issueInst;
        shifterReg_0_bits_store <= validSource_bits_store;
        shifterReg_0_bits_special <= validSource_bits_special;
        shifterReg_0_bits_lsWholeReg <= validSource_bits_lsWholeReg;
        shifterReg_0_bits_vs1 <= validSource_bits_vs1;
        shifterReg_0_bits_vs2 <= validSource_bits_vs2;
        shifterReg_0_bits_vd <= validSource_bits_vd;
        shifterReg_0_bits_loadStoreEEW <= validSource_bits_loadStoreEEW;
        shifterReg_0_bits_mask <= validSource_bits_mask;
        shifterReg_0_bits_segment <= validSource_bits_segment;
        shifterReg_0_bits_readFromScalar <= validSource_bits_readFromScalar;
        shifterReg_0_bits_csrInterface_vl <= validSource_bits_csrInterface_vl;
        shifterReg_0_bits_csrInterface_vStart <= validSource_bits_csrInterface_vStart;
        shifterReg_0_bits_csrInterface_vlmul <= validSource_bits_csrInterface_vlmul;
        shifterReg_0_bits_csrInterface_vSew <= validSource_bits_csrInterface_vSew;
        shifterReg_0_bits_csrInterface_vxrm <= validSource_bits_csrInterface_vxrm;
        shifterReg_0_bits_csrInterface_vta <= validSource_bits_csrInterface_vta;
        shifterReg_0_bits_csrInterface_vma <= validSource_bits_csrInterface_vma;
      end
      releasePipe_pipe_v_1 <= laneVec_1_laneRequest_bits_issueInst;
      if (validSource_1_valid ^ releasePipe_pipe_out_1_valid)
        tokenCheck_counter_1 <= tokenCheck_counter_1 + tokenCheck_counterChange_1;
      if (shifterValid_1) begin
        shifterReg_1_0_valid <= validSource_1_valid;
        shifterReg_1_0_bits_instructionIndex <= validSource_1_bits_instructionIndex;
        shifterReg_1_0_bits_decodeResult_specialSlot <= validSource_1_bits_decodeResult_specialSlot;
        shifterReg_1_0_bits_decodeResult_topUop <= validSource_1_bits_decodeResult_topUop;
        shifterReg_1_0_bits_decodeResult_popCount <= validSource_1_bits_decodeResult_popCount;
        shifterReg_1_0_bits_decodeResult_ffo <= validSource_1_bits_decodeResult_ffo;
        shifterReg_1_0_bits_decodeResult_average <= validSource_1_bits_decodeResult_average;
        shifterReg_1_0_bits_decodeResult_reverse <= validSource_1_bits_decodeResult_reverse;
        shifterReg_1_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_1_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_1_0_bits_decodeResult_scheduler <= validSource_1_bits_decodeResult_scheduler;
        shifterReg_1_0_bits_decodeResult_sReadVD <= validSource_1_bits_decodeResult_sReadVD;
        shifterReg_1_0_bits_decodeResult_vtype <= validSource_1_bits_decodeResult_vtype;
        shifterReg_1_0_bits_decodeResult_sWrite <= validSource_1_bits_decodeResult_sWrite;
        shifterReg_1_0_bits_decodeResult_crossRead <= validSource_1_bits_decodeResult_crossRead;
        shifterReg_1_0_bits_decodeResult_crossWrite <= validSource_1_bits_decodeResult_crossWrite;
        shifterReg_1_0_bits_decodeResult_maskUnit <= validSource_1_bits_decodeResult_maskUnit;
        shifterReg_1_0_bits_decodeResult_special <= validSource_1_bits_decodeResult_special;
        shifterReg_1_0_bits_decodeResult_saturate <= validSource_1_bits_decodeResult_saturate;
        shifterReg_1_0_bits_decodeResult_vwmacc <= validSource_1_bits_decodeResult_vwmacc;
        shifterReg_1_0_bits_decodeResult_readOnly <= validSource_1_bits_decodeResult_readOnly;
        shifterReg_1_0_bits_decodeResult_maskSource <= validSource_1_bits_decodeResult_maskSource;
        shifterReg_1_0_bits_decodeResult_maskDestination <= validSource_1_bits_decodeResult_maskDestination;
        shifterReg_1_0_bits_decodeResult_maskLogic <= validSource_1_bits_decodeResult_maskLogic;
        shifterReg_1_0_bits_decodeResult_uop <= validSource_1_bits_decodeResult_uop;
        shifterReg_1_0_bits_decodeResult_iota <= validSource_1_bits_decodeResult_iota;
        shifterReg_1_0_bits_decodeResult_mv <= validSource_1_bits_decodeResult_mv;
        shifterReg_1_0_bits_decodeResult_extend <= validSource_1_bits_decodeResult_extend;
        shifterReg_1_0_bits_decodeResult_unOrderWrite <= validSource_1_bits_decodeResult_unOrderWrite;
        shifterReg_1_0_bits_decodeResult_compress <= validSource_1_bits_decodeResult_compress;
        shifterReg_1_0_bits_decodeResult_gather16 <= validSource_1_bits_decodeResult_gather16;
        shifterReg_1_0_bits_decodeResult_gather <= validSource_1_bits_decodeResult_gather;
        shifterReg_1_0_bits_decodeResult_slid <= validSource_1_bits_decodeResult_slid;
        shifterReg_1_0_bits_decodeResult_targetRd <= validSource_1_bits_decodeResult_targetRd;
        shifterReg_1_0_bits_decodeResult_widenReduce <= validSource_1_bits_decodeResult_widenReduce;
        shifterReg_1_0_bits_decodeResult_red <= validSource_1_bits_decodeResult_red;
        shifterReg_1_0_bits_decodeResult_nr <= validSource_1_bits_decodeResult_nr;
        shifterReg_1_0_bits_decodeResult_itype <= validSource_1_bits_decodeResult_itype;
        shifterReg_1_0_bits_decodeResult_unsigned1 <= validSource_1_bits_decodeResult_unsigned1;
        shifterReg_1_0_bits_decodeResult_unsigned0 <= validSource_1_bits_decodeResult_unsigned0;
        shifterReg_1_0_bits_decodeResult_other <= validSource_1_bits_decodeResult_other;
        shifterReg_1_0_bits_decodeResult_multiCycle <= validSource_1_bits_decodeResult_multiCycle;
        shifterReg_1_0_bits_decodeResult_divider <= validSource_1_bits_decodeResult_divider;
        shifterReg_1_0_bits_decodeResult_multiplier <= validSource_1_bits_decodeResult_multiplier;
        shifterReg_1_0_bits_decodeResult_shift <= validSource_1_bits_decodeResult_shift;
        shifterReg_1_0_bits_decodeResult_adder <= validSource_1_bits_decodeResult_adder;
        shifterReg_1_0_bits_decodeResult_logic <= validSource_1_bits_decodeResult_logic;
        shifterReg_1_0_bits_loadStore <= validSource_1_bits_loadStore;
        shifterReg_1_0_bits_issueInst <= validSource_1_bits_issueInst;
        shifterReg_1_0_bits_store <= validSource_1_bits_store;
        shifterReg_1_0_bits_special <= validSource_1_bits_special;
        shifterReg_1_0_bits_lsWholeReg <= validSource_1_bits_lsWholeReg;
        shifterReg_1_0_bits_vs1 <= validSource_1_bits_vs1;
        shifterReg_1_0_bits_vs2 <= validSource_1_bits_vs2;
        shifterReg_1_0_bits_vd <= validSource_1_bits_vd;
        shifterReg_1_0_bits_loadStoreEEW <= validSource_1_bits_loadStoreEEW;
        shifterReg_1_0_bits_mask <= validSource_1_bits_mask;
        shifterReg_1_0_bits_segment <= validSource_1_bits_segment;
        shifterReg_1_0_bits_readFromScalar <= validSource_1_bits_readFromScalar;
        shifterReg_1_0_bits_csrInterface_vl <= validSource_1_bits_csrInterface_vl;
        shifterReg_1_0_bits_csrInterface_vStart <= validSource_1_bits_csrInterface_vStart;
        shifterReg_1_0_bits_csrInterface_vlmul <= validSource_1_bits_csrInterface_vlmul;
        shifterReg_1_0_bits_csrInterface_vSew <= validSource_1_bits_csrInterface_vSew;
        shifterReg_1_0_bits_csrInterface_vxrm <= validSource_1_bits_csrInterface_vxrm;
        shifterReg_1_0_bits_csrInterface_vta <= validSource_1_bits_csrInterface_vta;
        shifterReg_1_0_bits_csrInterface_vma <= validSource_1_bits_csrInterface_vma;
      end
      releasePipe_pipe_v_2 <= laneVec_2_laneRequest_bits_issueInst;
      if (validSource_2_valid ^ releasePipe_pipe_out_2_valid)
        tokenCheck_counter_2 <= tokenCheck_counter_2 + tokenCheck_counterChange_2;
      if (shifterValid_2) begin
        shifterReg_2_0_valid <= validSource_2_valid;
        shifterReg_2_0_bits_instructionIndex <= validSource_2_bits_instructionIndex;
        shifterReg_2_0_bits_decodeResult_specialSlot <= validSource_2_bits_decodeResult_specialSlot;
        shifterReg_2_0_bits_decodeResult_topUop <= validSource_2_bits_decodeResult_topUop;
        shifterReg_2_0_bits_decodeResult_popCount <= validSource_2_bits_decodeResult_popCount;
        shifterReg_2_0_bits_decodeResult_ffo <= validSource_2_bits_decodeResult_ffo;
        shifterReg_2_0_bits_decodeResult_average <= validSource_2_bits_decodeResult_average;
        shifterReg_2_0_bits_decodeResult_reverse <= validSource_2_bits_decodeResult_reverse;
        shifterReg_2_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_2_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_2_0_bits_decodeResult_scheduler <= validSource_2_bits_decodeResult_scheduler;
        shifterReg_2_0_bits_decodeResult_sReadVD <= validSource_2_bits_decodeResult_sReadVD;
        shifterReg_2_0_bits_decodeResult_vtype <= validSource_2_bits_decodeResult_vtype;
        shifterReg_2_0_bits_decodeResult_sWrite <= validSource_2_bits_decodeResult_sWrite;
        shifterReg_2_0_bits_decodeResult_crossRead <= validSource_2_bits_decodeResult_crossRead;
        shifterReg_2_0_bits_decodeResult_crossWrite <= validSource_2_bits_decodeResult_crossWrite;
        shifterReg_2_0_bits_decodeResult_maskUnit <= validSource_2_bits_decodeResult_maskUnit;
        shifterReg_2_0_bits_decodeResult_special <= validSource_2_bits_decodeResult_special;
        shifterReg_2_0_bits_decodeResult_saturate <= validSource_2_bits_decodeResult_saturate;
        shifterReg_2_0_bits_decodeResult_vwmacc <= validSource_2_bits_decodeResult_vwmacc;
        shifterReg_2_0_bits_decodeResult_readOnly <= validSource_2_bits_decodeResult_readOnly;
        shifterReg_2_0_bits_decodeResult_maskSource <= validSource_2_bits_decodeResult_maskSource;
        shifterReg_2_0_bits_decodeResult_maskDestination <= validSource_2_bits_decodeResult_maskDestination;
        shifterReg_2_0_bits_decodeResult_maskLogic <= validSource_2_bits_decodeResult_maskLogic;
        shifterReg_2_0_bits_decodeResult_uop <= validSource_2_bits_decodeResult_uop;
        shifterReg_2_0_bits_decodeResult_iota <= validSource_2_bits_decodeResult_iota;
        shifterReg_2_0_bits_decodeResult_mv <= validSource_2_bits_decodeResult_mv;
        shifterReg_2_0_bits_decodeResult_extend <= validSource_2_bits_decodeResult_extend;
        shifterReg_2_0_bits_decodeResult_unOrderWrite <= validSource_2_bits_decodeResult_unOrderWrite;
        shifterReg_2_0_bits_decodeResult_compress <= validSource_2_bits_decodeResult_compress;
        shifterReg_2_0_bits_decodeResult_gather16 <= validSource_2_bits_decodeResult_gather16;
        shifterReg_2_0_bits_decodeResult_gather <= validSource_2_bits_decodeResult_gather;
        shifterReg_2_0_bits_decodeResult_slid <= validSource_2_bits_decodeResult_slid;
        shifterReg_2_0_bits_decodeResult_targetRd <= validSource_2_bits_decodeResult_targetRd;
        shifterReg_2_0_bits_decodeResult_widenReduce <= validSource_2_bits_decodeResult_widenReduce;
        shifterReg_2_0_bits_decodeResult_red <= validSource_2_bits_decodeResult_red;
        shifterReg_2_0_bits_decodeResult_nr <= validSource_2_bits_decodeResult_nr;
        shifterReg_2_0_bits_decodeResult_itype <= validSource_2_bits_decodeResult_itype;
        shifterReg_2_0_bits_decodeResult_unsigned1 <= validSource_2_bits_decodeResult_unsigned1;
        shifterReg_2_0_bits_decodeResult_unsigned0 <= validSource_2_bits_decodeResult_unsigned0;
        shifterReg_2_0_bits_decodeResult_other <= validSource_2_bits_decodeResult_other;
        shifterReg_2_0_bits_decodeResult_multiCycle <= validSource_2_bits_decodeResult_multiCycle;
        shifterReg_2_0_bits_decodeResult_divider <= validSource_2_bits_decodeResult_divider;
        shifterReg_2_0_bits_decodeResult_multiplier <= validSource_2_bits_decodeResult_multiplier;
        shifterReg_2_0_bits_decodeResult_shift <= validSource_2_bits_decodeResult_shift;
        shifterReg_2_0_bits_decodeResult_adder <= validSource_2_bits_decodeResult_adder;
        shifterReg_2_0_bits_decodeResult_logic <= validSource_2_bits_decodeResult_logic;
        shifterReg_2_0_bits_loadStore <= validSource_2_bits_loadStore;
        shifterReg_2_0_bits_issueInst <= validSource_2_bits_issueInst;
        shifterReg_2_0_bits_store <= validSource_2_bits_store;
        shifterReg_2_0_bits_special <= validSource_2_bits_special;
        shifterReg_2_0_bits_lsWholeReg <= validSource_2_bits_lsWholeReg;
        shifterReg_2_0_bits_vs1 <= validSource_2_bits_vs1;
        shifterReg_2_0_bits_vs2 <= validSource_2_bits_vs2;
        shifterReg_2_0_bits_vd <= validSource_2_bits_vd;
        shifterReg_2_0_bits_loadStoreEEW <= validSource_2_bits_loadStoreEEW;
        shifterReg_2_0_bits_mask <= validSource_2_bits_mask;
        shifterReg_2_0_bits_segment <= validSource_2_bits_segment;
        shifterReg_2_0_bits_readFromScalar <= validSource_2_bits_readFromScalar;
        shifterReg_2_0_bits_csrInterface_vl <= validSource_2_bits_csrInterface_vl;
        shifterReg_2_0_bits_csrInterface_vStart <= validSource_2_bits_csrInterface_vStart;
        shifterReg_2_0_bits_csrInterface_vlmul <= validSource_2_bits_csrInterface_vlmul;
        shifterReg_2_0_bits_csrInterface_vSew <= validSource_2_bits_csrInterface_vSew;
        shifterReg_2_0_bits_csrInterface_vxrm <= validSource_2_bits_csrInterface_vxrm;
        shifterReg_2_0_bits_csrInterface_vta <= validSource_2_bits_csrInterface_vta;
        shifterReg_2_0_bits_csrInterface_vma <= validSource_2_bits_csrInterface_vma;
      end
      releasePipe_pipe_v_3 <= laneVec_3_laneRequest_bits_issueInst;
      if (validSource_3_valid ^ releasePipe_pipe_out_3_valid)
        tokenCheck_counter_3 <= tokenCheck_counter_3 + tokenCheck_counterChange_3;
      if (shifterValid_3) begin
        shifterReg_3_0_valid <= validSource_3_valid;
        shifterReg_3_0_bits_instructionIndex <= validSource_3_bits_instructionIndex;
        shifterReg_3_0_bits_decodeResult_specialSlot <= validSource_3_bits_decodeResult_specialSlot;
        shifterReg_3_0_bits_decodeResult_topUop <= validSource_3_bits_decodeResult_topUop;
        shifterReg_3_0_bits_decodeResult_popCount <= validSource_3_bits_decodeResult_popCount;
        shifterReg_3_0_bits_decodeResult_ffo <= validSource_3_bits_decodeResult_ffo;
        shifterReg_3_0_bits_decodeResult_average <= validSource_3_bits_decodeResult_average;
        shifterReg_3_0_bits_decodeResult_reverse <= validSource_3_bits_decodeResult_reverse;
        shifterReg_3_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_3_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_3_0_bits_decodeResult_scheduler <= validSource_3_bits_decodeResult_scheduler;
        shifterReg_3_0_bits_decodeResult_sReadVD <= validSource_3_bits_decodeResult_sReadVD;
        shifterReg_3_0_bits_decodeResult_vtype <= validSource_3_bits_decodeResult_vtype;
        shifterReg_3_0_bits_decodeResult_sWrite <= validSource_3_bits_decodeResult_sWrite;
        shifterReg_3_0_bits_decodeResult_crossRead <= validSource_3_bits_decodeResult_crossRead;
        shifterReg_3_0_bits_decodeResult_crossWrite <= validSource_3_bits_decodeResult_crossWrite;
        shifterReg_3_0_bits_decodeResult_maskUnit <= validSource_3_bits_decodeResult_maskUnit;
        shifterReg_3_0_bits_decodeResult_special <= validSource_3_bits_decodeResult_special;
        shifterReg_3_0_bits_decodeResult_saturate <= validSource_3_bits_decodeResult_saturate;
        shifterReg_3_0_bits_decodeResult_vwmacc <= validSource_3_bits_decodeResult_vwmacc;
        shifterReg_3_0_bits_decodeResult_readOnly <= validSource_3_bits_decodeResult_readOnly;
        shifterReg_3_0_bits_decodeResult_maskSource <= validSource_3_bits_decodeResult_maskSource;
        shifterReg_3_0_bits_decodeResult_maskDestination <= validSource_3_bits_decodeResult_maskDestination;
        shifterReg_3_0_bits_decodeResult_maskLogic <= validSource_3_bits_decodeResult_maskLogic;
        shifterReg_3_0_bits_decodeResult_uop <= validSource_3_bits_decodeResult_uop;
        shifterReg_3_0_bits_decodeResult_iota <= validSource_3_bits_decodeResult_iota;
        shifterReg_3_0_bits_decodeResult_mv <= validSource_3_bits_decodeResult_mv;
        shifterReg_3_0_bits_decodeResult_extend <= validSource_3_bits_decodeResult_extend;
        shifterReg_3_0_bits_decodeResult_unOrderWrite <= validSource_3_bits_decodeResult_unOrderWrite;
        shifterReg_3_0_bits_decodeResult_compress <= validSource_3_bits_decodeResult_compress;
        shifterReg_3_0_bits_decodeResult_gather16 <= validSource_3_bits_decodeResult_gather16;
        shifterReg_3_0_bits_decodeResult_gather <= validSource_3_bits_decodeResult_gather;
        shifterReg_3_0_bits_decodeResult_slid <= validSource_3_bits_decodeResult_slid;
        shifterReg_3_0_bits_decodeResult_targetRd <= validSource_3_bits_decodeResult_targetRd;
        shifterReg_3_0_bits_decodeResult_widenReduce <= validSource_3_bits_decodeResult_widenReduce;
        shifterReg_3_0_bits_decodeResult_red <= validSource_3_bits_decodeResult_red;
        shifterReg_3_0_bits_decodeResult_nr <= validSource_3_bits_decodeResult_nr;
        shifterReg_3_0_bits_decodeResult_itype <= validSource_3_bits_decodeResult_itype;
        shifterReg_3_0_bits_decodeResult_unsigned1 <= validSource_3_bits_decodeResult_unsigned1;
        shifterReg_3_0_bits_decodeResult_unsigned0 <= validSource_3_bits_decodeResult_unsigned0;
        shifterReg_3_0_bits_decodeResult_other <= validSource_3_bits_decodeResult_other;
        shifterReg_3_0_bits_decodeResult_multiCycle <= validSource_3_bits_decodeResult_multiCycle;
        shifterReg_3_0_bits_decodeResult_divider <= validSource_3_bits_decodeResult_divider;
        shifterReg_3_0_bits_decodeResult_multiplier <= validSource_3_bits_decodeResult_multiplier;
        shifterReg_3_0_bits_decodeResult_shift <= validSource_3_bits_decodeResult_shift;
        shifterReg_3_0_bits_decodeResult_adder <= validSource_3_bits_decodeResult_adder;
        shifterReg_3_0_bits_decodeResult_logic <= validSource_3_bits_decodeResult_logic;
        shifterReg_3_0_bits_loadStore <= validSource_3_bits_loadStore;
        shifterReg_3_0_bits_issueInst <= validSource_3_bits_issueInst;
        shifterReg_3_0_bits_store <= validSource_3_bits_store;
        shifterReg_3_0_bits_special <= validSource_3_bits_special;
        shifterReg_3_0_bits_lsWholeReg <= validSource_3_bits_lsWholeReg;
        shifterReg_3_0_bits_vs1 <= validSource_3_bits_vs1;
        shifterReg_3_0_bits_vs2 <= validSource_3_bits_vs2;
        shifterReg_3_0_bits_vd <= validSource_3_bits_vd;
        shifterReg_3_0_bits_loadStoreEEW <= validSource_3_bits_loadStoreEEW;
        shifterReg_3_0_bits_mask <= validSource_3_bits_mask;
        shifterReg_3_0_bits_segment <= validSource_3_bits_segment;
        shifterReg_3_0_bits_readFromScalar <= validSource_3_bits_readFromScalar;
        shifterReg_3_0_bits_csrInterface_vl <= validSource_3_bits_csrInterface_vl;
        shifterReg_3_0_bits_csrInterface_vStart <= validSource_3_bits_csrInterface_vStart;
        shifterReg_3_0_bits_csrInterface_vlmul <= validSource_3_bits_csrInterface_vlmul;
        shifterReg_3_0_bits_csrInterface_vSew <= validSource_3_bits_csrInterface_vSew;
        shifterReg_3_0_bits_csrInterface_vxrm <= validSource_3_bits_csrInterface_vxrm;
        shifterReg_3_0_bits_csrInterface_vta <= validSource_3_bits_csrInterface_vta;
        shifterReg_3_0_bits_csrInterface_vma <= validSource_3_bits_csrInterface_vma;
      end
      releasePipe_pipe_v_4 <= laneVec_4_laneRequest_bits_issueInst;
      if (validSource_4_valid ^ releasePipe_pipe_out_4_valid)
        tokenCheck_counter_4 <= tokenCheck_counter_4 + tokenCheck_counterChange_4;
      if (shifterValid_4) begin
        shifterReg_4_0_valid <= validSource_4_valid;
        shifterReg_4_0_bits_instructionIndex <= validSource_4_bits_instructionIndex;
        shifterReg_4_0_bits_decodeResult_specialSlot <= validSource_4_bits_decodeResult_specialSlot;
        shifterReg_4_0_bits_decodeResult_topUop <= validSource_4_bits_decodeResult_topUop;
        shifterReg_4_0_bits_decodeResult_popCount <= validSource_4_bits_decodeResult_popCount;
        shifterReg_4_0_bits_decodeResult_ffo <= validSource_4_bits_decodeResult_ffo;
        shifterReg_4_0_bits_decodeResult_average <= validSource_4_bits_decodeResult_average;
        shifterReg_4_0_bits_decodeResult_reverse <= validSource_4_bits_decodeResult_reverse;
        shifterReg_4_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_4_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_4_0_bits_decodeResult_scheduler <= validSource_4_bits_decodeResult_scheduler;
        shifterReg_4_0_bits_decodeResult_sReadVD <= validSource_4_bits_decodeResult_sReadVD;
        shifterReg_4_0_bits_decodeResult_vtype <= validSource_4_bits_decodeResult_vtype;
        shifterReg_4_0_bits_decodeResult_sWrite <= validSource_4_bits_decodeResult_sWrite;
        shifterReg_4_0_bits_decodeResult_crossRead <= validSource_4_bits_decodeResult_crossRead;
        shifterReg_4_0_bits_decodeResult_crossWrite <= validSource_4_bits_decodeResult_crossWrite;
        shifterReg_4_0_bits_decodeResult_maskUnit <= validSource_4_bits_decodeResult_maskUnit;
        shifterReg_4_0_bits_decodeResult_special <= validSource_4_bits_decodeResult_special;
        shifterReg_4_0_bits_decodeResult_saturate <= validSource_4_bits_decodeResult_saturate;
        shifterReg_4_0_bits_decodeResult_vwmacc <= validSource_4_bits_decodeResult_vwmacc;
        shifterReg_4_0_bits_decodeResult_readOnly <= validSource_4_bits_decodeResult_readOnly;
        shifterReg_4_0_bits_decodeResult_maskSource <= validSource_4_bits_decodeResult_maskSource;
        shifterReg_4_0_bits_decodeResult_maskDestination <= validSource_4_bits_decodeResult_maskDestination;
        shifterReg_4_0_bits_decodeResult_maskLogic <= validSource_4_bits_decodeResult_maskLogic;
        shifterReg_4_0_bits_decodeResult_uop <= validSource_4_bits_decodeResult_uop;
        shifterReg_4_0_bits_decodeResult_iota <= validSource_4_bits_decodeResult_iota;
        shifterReg_4_0_bits_decodeResult_mv <= validSource_4_bits_decodeResult_mv;
        shifterReg_4_0_bits_decodeResult_extend <= validSource_4_bits_decodeResult_extend;
        shifterReg_4_0_bits_decodeResult_unOrderWrite <= validSource_4_bits_decodeResult_unOrderWrite;
        shifterReg_4_0_bits_decodeResult_compress <= validSource_4_bits_decodeResult_compress;
        shifterReg_4_0_bits_decodeResult_gather16 <= validSource_4_bits_decodeResult_gather16;
        shifterReg_4_0_bits_decodeResult_gather <= validSource_4_bits_decodeResult_gather;
        shifterReg_4_0_bits_decodeResult_slid <= validSource_4_bits_decodeResult_slid;
        shifterReg_4_0_bits_decodeResult_targetRd <= validSource_4_bits_decodeResult_targetRd;
        shifterReg_4_0_bits_decodeResult_widenReduce <= validSource_4_bits_decodeResult_widenReduce;
        shifterReg_4_0_bits_decodeResult_red <= validSource_4_bits_decodeResult_red;
        shifterReg_4_0_bits_decodeResult_nr <= validSource_4_bits_decodeResult_nr;
        shifterReg_4_0_bits_decodeResult_itype <= validSource_4_bits_decodeResult_itype;
        shifterReg_4_0_bits_decodeResult_unsigned1 <= validSource_4_bits_decodeResult_unsigned1;
        shifterReg_4_0_bits_decodeResult_unsigned0 <= validSource_4_bits_decodeResult_unsigned0;
        shifterReg_4_0_bits_decodeResult_other <= validSource_4_bits_decodeResult_other;
        shifterReg_4_0_bits_decodeResult_multiCycle <= validSource_4_bits_decodeResult_multiCycle;
        shifterReg_4_0_bits_decodeResult_divider <= validSource_4_bits_decodeResult_divider;
        shifterReg_4_0_bits_decodeResult_multiplier <= validSource_4_bits_decodeResult_multiplier;
        shifterReg_4_0_bits_decodeResult_shift <= validSource_4_bits_decodeResult_shift;
        shifterReg_4_0_bits_decodeResult_adder <= validSource_4_bits_decodeResult_adder;
        shifterReg_4_0_bits_decodeResult_logic <= validSource_4_bits_decodeResult_logic;
        shifterReg_4_0_bits_loadStore <= validSource_4_bits_loadStore;
        shifterReg_4_0_bits_issueInst <= validSource_4_bits_issueInst;
        shifterReg_4_0_bits_store <= validSource_4_bits_store;
        shifterReg_4_0_bits_special <= validSource_4_bits_special;
        shifterReg_4_0_bits_lsWholeReg <= validSource_4_bits_lsWholeReg;
        shifterReg_4_0_bits_vs1 <= validSource_4_bits_vs1;
        shifterReg_4_0_bits_vs2 <= validSource_4_bits_vs2;
        shifterReg_4_0_bits_vd <= validSource_4_bits_vd;
        shifterReg_4_0_bits_loadStoreEEW <= validSource_4_bits_loadStoreEEW;
        shifterReg_4_0_bits_mask <= validSource_4_bits_mask;
        shifterReg_4_0_bits_segment <= validSource_4_bits_segment;
        shifterReg_4_0_bits_readFromScalar <= validSource_4_bits_readFromScalar;
        shifterReg_4_0_bits_csrInterface_vl <= validSource_4_bits_csrInterface_vl;
        shifterReg_4_0_bits_csrInterface_vStart <= validSource_4_bits_csrInterface_vStart;
        shifterReg_4_0_bits_csrInterface_vlmul <= validSource_4_bits_csrInterface_vlmul;
        shifterReg_4_0_bits_csrInterface_vSew <= validSource_4_bits_csrInterface_vSew;
        shifterReg_4_0_bits_csrInterface_vxrm <= validSource_4_bits_csrInterface_vxrm;
        shifterReg_4_0_bits_csrInterface_vta <= validSource_4_bits_csrInterface_vta;
        shifterReg_4_0_bits_csrInterface_vma <= validSource_4_bits_csrInterface_vma;
      end
      releasePipe_pipe_v_5 <= laneVec_5_laneRequest_bits_issueInst;
      if (validSource_5_valid ^ releasePipe_pipe_out_5_valid)
        tokenCheck_counter_5 <= tokenCheck_counter_5 + tokenCheck_counterChange_5;
      if (shifterValid_5) begin
        shifterReg_5_0_valid <= validSource_5_valid;
        shifterReg_5_0_bits_instructionIndex <= validSource_5_bits_instructionIndex;
        shifterReg_5_0_bits_decodeResult_specialSlot <= validSource_5_bits_decodeResult_specialSlot;
        shifterReg_5_0_bits_decodeResult_topUop <= validSource_5_bits_decodeResult_topUop;
        shifterReg_5_0_bits_decodeResult_popCount <= validSource_5_bits_decodeResult_popCount;
        shifterReg_5_0_bits_decodeResult_ffo <= validSource_5_bits_decodeResult_ffo;
        shifterReg_5_0_bits_decodeResult_average <= validSource_5_bits_decodeResult_average;
        shifterReg_5_0_bits_decodeResult_reverse <= validSource_5_bits_decodeResult_reverse;
        shifterReg_5_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_5_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_5_0_bits_decodeResult_scheduler <= validSource_5_bits_decodeResult_scheduler;
        shifterReg_5_0_bits_decodeResult_sReadVD <= validSource_5_bits_decodeResult_sReadVD;
        shifterReg_5_0_bits_decodeResult_vtype <= validSource_5_bits_decodeResult_vtype;
        shifterReg_5_0_bits_decodeResult_sWrite <= validSource_5_bits_decodeResult_sWrite;
        shifterReg_5_0_bits_decodeResult_crossRead <= validSource_5_bits_decodeResult_crossRead;
        shifterReg_5_0_bits_decodeResult_crossWrite <= validSource_5_bits_decodeResult_crossWrite;
        shifterReg_5_0_bits_decodeResult_maskUnit <= validSource_5_bits_decodeResult_maskUnit;
        shifterReg_5_0_bits_decodeResult_special <= validSource_5_bits_decodeResult_special;
        shifterReg_5_0_bits_decodeResult_saturate <= validSource_5_bits_decodeResult_saturate;
        shifterReg_5_0_bits_decodeResult_vwmacc <= validSource_5_bits_decodeResult_vwmacc;
        shifterReg_5_0_bits_decodeResult_readOnly <= validSource_5_bits_decodeResult_readOnly;
        shifterReg_5_0_bits_decodeResult_maskSource <= validSource_5_bits_decodeResult_maskSource;
        shifterReg_5_0_bits_decodeResult_maskDestination <= validSource_5_bits_decodeResult_maskDestination;
        shifterReg_5_0_bits_decodeResult_maskLogic <= validSource_5_bits_decodeResult_maskLogic;
        shifterReg_5_0_bits_decodeResult_uop <= validSource_5_bits_decodeResult_uop;
        shifterReg_5_0_bits_decodeResult_iota <= validSource_5_bits_decodeResult_iota;
        shifterReg_5_0_bits_decodeResult_mv <= validSource_5_bits_decodeResult_mv;
        shifterReg_5_0_bits_decodeResult_extend <= validSource_5_bits_decodeResult_extend;
        shifterReg_5_0_bits_decodeResult_unOrderWrite <= validSource_5_bits_decodeResult_unOrderWrite;
        shifterReg_5_0_bits_decodeResult_compress <= validSource_5_bits_decodeResult_compress;
        shifterReg_5_0_bits_decodeResult_gather16 <= validSource_5_bits_decodeResult_gather16;
        shifterReg_5_0_bits_decodeResult_gather <= validSource_5_bits_decodeResult_gather;
        shifterReg_5_0_bits_decodeResult_slid <= validSource_5_bits_decodeResult_slid;
        shifterReg_5_0_bits_decodeResult_targetRd <= validSource_5_bits_decodeResult_targetRd;
        shifterReg_5_0_bits_decodeResult_widenReduce <= validSource_5_bits_decodeResult_widenReduce;
        shifterReg_5_0_bits_decodeResult_red <= validSource_5_bits_decodeResult_red;
        shifterReg_5_0_bits_decodeResult_nr <= validSource_5_bits_decodeResult_nr;
        shifterReg_5_0_bits_decodeResult_itype <= validSource_5_bits_decodeResult_itype;
        shifterReg_5_0_bits_decodeResult_unsigned1 <= validSource_5_bits_decodeResult_unsigned1;
        shifterReg_5_0_bits_decodeResult_unsigned0 <= validSource_5_bits_decodeResult_unsigned0;
        shifterReg_5_0_bits_decodeResult_other <= validSource_5_bits_decodeResult_other;
        shifterReg_5_0_bits_decodeResult_multiCycle <= validSource_5_bits_decodeResult_multiCycle;
        shifterReg_5_0_bits_decodeResult_divider <= validSource_5_bits_decodeResult_divider;
        shifterReg_5_0_bits_decodeResult_multiplier <= validSource_5_bits_decodeResult_multiplier;
        shifterReg_5_0_bits_decodeResult_shift <= validSource_5_bits_decodeResult_shift;
        shifterReg_5_0_bits_decodeResult_adder <= validSource_5_bits_decodeResult_adder;
        shifterReg_5_0_bits_decodeResult_logic <= validSource_5_bits_decodeResult_logic;
        shifterReg_5_0_bits_loadStore <= validSource_5_bits_loadStore;
        shifterReg_5_0_bits_issueInst <= validSource_5_bits_issueInst;
        shifterReg_5_0_bits_store <= validSource_5_bits_store;
        shifterReg_5_0_bits_special <= validSource_5_bits_special;
        shifterReg_5_0_bits_lsWholeReg <= validSource_5_bits_lsWholeReg;
        shifterReg_5_0_bits_vs1 <= validSource_5_bits_vs1;
        shifterReg_5_0_bits_vs2 <= validSource_5_bits_vs2;
        shifterReg_5_0_bits_vd <= validSource_5_bits_vd;
        shifterReg_5_0_bits_loadStoreEEW <= validSource_5_bits_loadStoreEEW;
        shifterReg_5_0_bits_mask <= validSource_5_bits_mask;
        shifterReg_5_0_bits_segment <= validSource_5_bits_segment;
        shifterReg_5_0_bits_readFromScalar <= validSource_5_bits_readFromScalar;
        shifterReg_5_0_bits_csrInterface_vl <= validSource_5_bits_csrInterface_vl;
        shifterReg_5_0_bits_csrInterface_vStart <= validSource_5_bits_csrInterface_vStart;
        shifterReg_5_0_bits_csrInterface_vlmul <= validSource_5_bits_csrInterface_vlmul;
        shifterReg_5_0_bits_csrInterface_vSew <= validSource_5_bits_csrInterface_vSew;
        shifterReg_5_0_bits_csrInterface_vxrm <= validSource_5_bits_csrInterface_vxrm;
        shifterReg_5_0_bits_csrInterface_vta <= validSource_5_bits_csrInterface_vta;
        shifterReg_5_0_bits_csrInterface_vma <= validSource_5_bits_csrInterface_vma;
      end
      releasePipe_pipe_v_6 <= laneVec_6_laneRequest_bits_issueInst;
      if (validSource_6_valid ^ releasePipe_pipe_out_6_valid)
        tokenCheck_counter_6 <= tokenCheck_counter_6 + tokenCheck_counterChange_6;
      if (shifterValid_6) begin
        shifterReg_6_0_valid <= validSource_6_valid;
        shifterReg_6_0_bits_instructionIndex <= validSource_6_bits_instructionIndex;
        shifterReg_6_0_bits_decodeResult_specialSlot <= validSource_6_bits_decodeResult_specialSlot;
        shifterReg_6_0_bits_decodeResult_topUop <= validSource_6_bits_decodeResult_topUop;
        shifterReg_6_0_bits_decodeResult_popCount <= validSource_6_bits_decodeResult_popCount;
        shifterReg_6_0_bits_decodeResult_ffo <= validSource_6_bits_decodeResult_ffo;
        shifterReg_6_0_bits_decodeResult_average <= validSource_6_bits_decodeResult_average;
        shifterReg_6_0_bits_decodeResult_reverse <= validSource_6_bits_decodeResult_reverse;
        shifterReg_6_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_6_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_6_0_bits_decodeResult_scheduler <= validSource_6_bits_decodeResult_scheduler;
        shifterReg_6_0_bits_decodeResult_sReadVD <= validSource_6_bits_decodeResult_sReadVD;
        shifterReg_6_0_bits_decodeResult_vtype <= validSource_6_bits_decodeResult_vtype;
        shifterReg_6_0_bits_decodeResult_sWrite <= validSource_6_bits_decodeResult_sWrite;
        shifterReg_6_0_bits_decodeResult_crossRead <= validSource_6_bits_decodeResult_crossRead;
        shifterReg_6_0_bits_decodeResult_crossWrite <= validSource_6_bits_decodeResult_crossWrite;
        shifterReg_6_0_bits_decodeResult_maskUnit <= validSource_6_bits_decodeResult_maskUnit;
        shifterReg_6_0_bits_decodeResult_special <= validSource_6_bits_decodeResult_special;
        shifterReg_6_0_bits_decodeResult_saturate <= validSource_6_bits_decodeResult_saturate;
        shifterReg_6_0_bits_decodeResult_vwmacc <= validSource_6_bits_decodeResult_vwmacc;
        shifterReg_6_0_bits_decodeResult_readOnly <= validSource_6_bits_decodeResult_readOnly;
        shifterReg_6_0_bits_decodeResult_maskSource <= validSource_6_bits_decodeResult_maskSource;
        shifterReg_6_0_bits_decodeResult_maskDestination <= validSource_6_bits_decodeResult_maskDestination;
        shifterReg_6_0_bits_decodeResult_maskLogic <= validSource_6_bits_decodeResult_maskLogic;
        shifterReg_6_0_bits_decodeResult_uop <= validSource_6_bits_decodeResult_uop;
        shifterReg_6_0_bits_decodeResult_iota <= validSource_6_bits_decodeResult_iota;
        shifterReg_6_0_bits_decodeResult_mv <= validSource_6_bits_decodeResult_mv;
        shifterReg_6_0_bits_decodeResult_extend <= validSource_6_bits_decodeResult_extend;
        shifterReg_6_0_bits_decodeResult_unOrderWrite <= validSource_6_bits_decodeResult_unOrderWrite;
        shifterReg_6_0_bits_decodeResult_compress <= validSource_6_bits_decodeResult_compress;
        shifterReg_6_0_bits_decodeResult_gather16 <= validSource_6_bits_decodeResult_gather16;
        shifterReg_6_0_bits_decodeResult_gather <= validSource_6_bits_decodeResult_gather;
        shifterReg_6_0_bits_decodeResult_slid <= validSource_6_bits_decodeResult_slid;
        shifterReg_6_0_bits_decodeResult_targetRd <= validSource_6_bits_decodeResult_targetRd;
        shifterReg_6_0_bits_decodeResult_widenReduce <= validSource_6_bits_decodeResult_widenReduce;
        shifterReg_6_0_bits_decodeResult_red <= validSource_6_bits_decodeResult_red;
        shifterReg_6_0_bits_decodeResult_nr <= validSource_6_bits_decodeResult_nr;
        shifterReg_6_0_bits_decodeResult_itype <= validSource_6_bits_decodeResult_itype;
        shifterReg_6_0_bits_decodeResult_unsigned1 <= validSource_6_bits_decodeResult_unsigned1;
        shifterReg_6_0_bits_decodeResult_unsigned0 <= validSource_6_bits_decodeResult_unsigned0;
        shifterReg_6_0_bits_decodeResult_other <= validSource_6_bits_decodeResult_other;
        shifterReg_6_0_bits_decodeResult_multiCycle <= validSource_6_bits_decodeResult_multiCycle;
        shifterReg_6_0_bits_decodeResult_divider <= validSource_6_bits_decodeResult_divider;
        shifterReg_6_0_bits_decodeResult_multiplier <= validSource_6_bits_decodeResult_multiplier;
        shifterReg_6_0_bits_decodeResult_shift <= validSource_6_bits_decodeResult_shift;
        shifterReg_6_0_bits_decodeResult_adder <= validSource_6_bits_decodeResult_adder;
        shifterReg_6_0_bits_decodeResult_logic <= validSource_6_bits_decodeResult_logic;
        shifterReg_6_0_bits_loadStore <= validSource_6_bits_loadStore;
        shifterReg_6_0_bits_issueInst <= validSource_6_bits_issueInst;
        shifterReg_6_0_bits_store <= validSource_6_bits_store;
        shifterReg_6_0_bits_special <= validSource_6_bits_special;
        shifterReg_6_0_bits_lsWholeReg <= validSource_6_bits_lsWholeReg;
        shifterReg_6_0_bits_vs1 <= validSource_6_bits_vs1;
        shifterReg_6_0_bits_vs2 <= validSource_6_bits_vs2;
        shifterReg_6_0_bits_vd <= validSource_6_bits_vd;
        shifterReg_6_0_bits_loadStoreEEW <= validSource_6_bits_loadStoreEEW;
        shifterReg_6_0_bits_mask <= validSource_6_bits_mask;
        shifterReg_6_0_bits_segment <= validSource_6_bits_segment;
        shifterReg_6_0_bits_readFromScalar <= validSource_6_bits_readFromScalar;
        shifterReg_6_0_bits_csrInterface_vl <= validSource_6_bits_csrInterface_vl;
        shifterReg_6_0_bits_csrInterface_vStart <= validSource_6_bits_csrInterface_vStart;
        shifterReg_6_0_bits_csrInterface_vlmul <= validSource_6_bits_csrInterface_vlmul;
        shifterReg_6_0_bits_csrInterface_vSew <= validSource_6_bits_csrInterface_vSew;
        shifterReg_6_0_bits_csrInterface_vxrm <= validSource_6_bits_csrInterface_vxrm;
        shifterReg_6_0_bits_csrInterface_vta <= validSource_6_bits_csrInterface_vta;
        shifterReg_6_0_bits_csrInterface_vma <= validSource_6_bits_csrInterface_vma;
      end
      releasePipe_pipe_v_7 <= laneVec_7_laneRequest_bits_issueInst;
      if (validSource_7_valid ^ releasePipe_pipe_out_7_valid)
        tokenCheck_counter_7 <= tokenCheck_counter_7 + tokenCheck_counterChange_7;
      if (shifterValid_7) begin
        shifterReg_7_0_valid <= validSource_7_valid;
        shifterReg_7_0_bits_instructionIndex <= validSource_7_bits_instructionIndex;
        shifterReg_7_0_bits_decodeResult_specialSlot <= validSource_7_bits_decodeResult_specialSlot;
        shifterReg_7_0_bits_decodeResult_topUop <= validSource_7_bits_decodeResult_topUop;
        shifterReg_7_0_bits_decodeResult_popCount <= validSource_7_bits_decodeResult_popCount;
        shifterReg_7_0_bits_decodeResult_ffo <= validSource_7_bits_decodeResult_ffo;
        shifterReg_7_0_bits_decodeResult_average <= validSource_7_bits_decodeResult_average;
        shifterReg_7_0_bits_decodeResult_reverse <= validSource_7_bits_decodeResult_reverse;
        shifterReg_7_0_bits_decodeResult_dontNeedExecuteInLane <= validSource_7_bits_decodeResult_dontNeedExecuteInLane;
        shifterReg_7_0_bits_decodeResult_scheduler <= validSource_7_bits_decodeResult_scheduler;
        shifterReg_7_0_bits_decodeResult_sReadVD <= validSource_7_bits_decodeResult_sReadVD;
        shifterReg_7_0_bits_decodeResult_vtype <= validSource_7_bits_decodeResult_vtype;
        shifterReg_7_0_bits_decodeResult_sWrite <= validSource_7_bits_decodeResult_sWrite;
        shifterReg_7_0_bits_decodeResult_crossRead <= validSource_7_bits_decodeResult_crossRead;
        shifterReg_7_0_bits_decodeResult_crossWrite <= validSource_7_bits_decodeResult_crossWrite;
        shifterReg_7_0_bits_decodeResult_maskUnit <= validSource_7_bits_decodeResult_maskUnit;
        shifterReg_7_0_bits_decodeResult_special <= validSource_7_bits_decodeResult_special;
        shifterReg_7_0_bits_decodeResult_saturate <= validSource_7_bits_decodeResult_saturate;
        shifterReg_7_0_bits_decodeResult_vwmacc <= validSource_7_bits_decodeResult_vwmacc;
        shifterReg_7_0_bits_decodeResult_readOnly <= validSource_7_bits_decodeResult_readOnly;
        shifterReg_7_0_bits_decodeResult_maskSource <= validSource_7_bits_decodeResult_maskSource;
        shifterReg_7_0_bits_decodeResult_maskDestination <= validSource_7_bits_decodeResult_maskDestination;
        shifterReg_7_0_bits_decodeResult_maskLogic <= validSource_7_bits_decodeResult_maskLogic;
        shifterReg_7_0_bits_decodeResult_uop <= validSource_7_bits_decodeResult_uop;
        shifterReg_7_0_bits_decodeResult_iota <= validSource_7_bits_decodeResult_iota;
        shifterReg_7_0_bits_decodeResult_mv <= validSource_7_bits_decodeResult_mv;
        shifterReg_7_0_bits_decodeResult_extend <= validSource_7_bits_decodeResult_extend;
        shifterReg_7_0_bits_decodeResult_unOrderWrite <= validSource_7_bits_decodeResult_unOrderWrite;
        shifterReg_7_0_bits_decodeResult_compress <= validSource_7_bits_decodeResult_compress;
        shifterReg_7_0_bits_decodeResult_gather16 <= validSource_7_bits_decodeResult_gather16;
        shifterReg_7_0_bits_decodeResult_gather <= validSource_7_bits_decodeResult_gather;
        shifterReg_7_0_bits_decodeResult_slid <= validSource_7_bits_decodeResult_slid;
        shifterReg_7_0_bits_decodeResult_targetRd <= validSource_7_bits_decodeResult_targetRd;
        shifterReg_7_0_bits_decodeResult_widenReduce <= validSource_7_bits_decodeResult_widenReduce;
        shifterReg_7_0_bits_decodeResult_red <= validSource_7_bits_decodeResult_red;
        shifterReg_7_0_bits_decodeResult_nr <= validSource_7_bits_decodeResult_nr;
        shifterReg_7_0_bits_decodeResult_itype <= validSource_7_bits_decodeResult_itype;
        shifterReg_7_0_bits_decodeResult_unsigned1 <= validSource_7_bits_decodeResult_unsigned1;
        shifterReg_7_0_bits_decodeResult_unsigned0 <= validSource_7_bits_decodeResult_unsigned0;
        shifterReg_7_0_bits_decodeResult_other <= validSource_7_bits_decodeResult_other;
        shifterReg_7_0_bits_decodeResult_multiCycle <= validSource_7_bits_decodeResult_multiCycle;
        shifterReg_7_0_bits_decodeResult_divider <= validSource_7_bits_decodeResult_divider;
        shifterReg_7_0_bits_decodeResult_multiplier <= validSource_7_bits_decodeResult_multiplier;
        shifterReg_7_0_bits_decodeResult_shift <= validSource_7_bits_decodeResult_shift;
        shifterReg_7_0_bits_decodeResult_adder <= validSource_7_bits_decodeResult_adder;
        shifterReg_7_0_bits_decodeResult_logic <= validSource_7_bits_decodeResult_logic;
        shifterReg_7_0_bits_loadStore <= validSource_7_bits_loadStore;
        shifterReg_7_0_bits_issueInst <= validSource_7_bits_issueInst;
        shifterReg_7_0_bits_store <= validSource_7_bits_store;
        shifterReg_7_0_bits_special <= validSource_7_bits_special;
        shifterReg_7_0_bits_lsWholeReg <= validSource_7_bits_lsWholeReg;
        shifterReg_7_0_bits_vs1 <= validSource_7_bits_vs1;
        shifterReg_7_0_bits_vs2 <= validSource_7_bits_vs2;
        shifterReg_7_0_bits_vd <= validSource_7_bits_vd;
        shifterReg_7_0_bits_loadStoreEEW <= validSource_7_bits_loadStoreEEW;
        shifterReg_7_0_bits_mask <= validSource_7_bits_mask;
        shifterReg_7_0_bits_segment <= validSource_7_bits_segment;
        shifterReg_7_0_bits_readFromScalar <= validSource_7_bits_readFromScalar;
        shifterReg_7_0_bits_csrInterface_vl <= validSource_7_bits_csrInterface_vl;
        shifterReg_7_0_bits_csrInterface_vStart <= validSource_7_bits_csrInterface_vStart;
        shifterReg_7_0_bits_csrInterface_vlmul <= validSource_7_bits_csrInterface_vlmul;
        shifterReg_7_0_bits_csrInterface_vSew <= validSource_7_bits_csrInterface_vSew;
        shifterReg_7_0_bits_csrInterface_vxrm <= validSource_7_bits_csrInterface_vxrm;
        shifterReg_7_0_bits_csrInterface_vta <= validSource_7_bits_csrInterface_vta;
        shifterReg_7_0_bits_csrInterface_vma <= validSource_7_bits_csrInterface_vma;
      end
      sinkVec_releasePipe_pipe_v <= sinkVec_sinkWire_ready & sinkVec_sinkWire_valid;
      if (sinkVec_validSource_valid ^ sinkVec_releasePipe_pipe_out_valid)
        sinkVec_tokenCheck_counter <= sinkVec_tokenCheck_counter + sinkVec_tokenCheck_counterChange;
      if (sinkVec_shifterValid) begin
        sinkVec_shifterReg_0_valid <= sinkVec_validSource_valid;
        sinkVec_shifterReg_0_bits_vs <= sinkVec_validSource_bits_vs;
        sinkVec_shifterReg_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_0_bits_offset <= sinkVec_validSource_bits_offset;
        sinkVec_shifterReg_0_bits_instructionIndex <= sinkVec_validSource_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_1 <= sinkVec_sinkWire_1_ready & sinkVec_sinkWire_1_valid;
      if (sinkVec_validSource_1_valid ^ sinkVec_releasePipe_pipe_out_1_valid)
        sinkVec_tokenCheck_counter_1 <= sinkVec_tokenCheck_counter_1 + sinkVec_tokenCheck_counterChange_1;
      if (sinkVec_shifterValid_1) begin
        sinkVec_shifterReg_1_0_valid <= sinkVec_validSource_1_valid;
        sinkVec_shifterReg_1_0_bits_vs <= sinkVec_validSource_1_bits_vs;
        sinkVec_shifterReg_1_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_1_0_bits_offset <= sinkVec_validSource_1_bits_offset;
        sinkVec_shifterReg_1_0_bits_instructionIndex <= sinkVec_validSource_1_bits_instructionIndex;
      end
      maskUnitFirst <= tryToRead & ~(sinkWire_ready & sinkWire_valid) ^ maskUnitFirst;
      accessDataValid_pipe_v <= sinkVec_0_ready & sinkVec_0_valid;
      accessDataValid_pipe_pipe_v <= accessDataValid_pipe_v;
      if (shifterValid_8) begin
        shifterReg_8_0_valid <= accessDataSource_valid;
        shifterReg_8_0_bits <= accessDataSource_bits;
      end
      accessDataValid_pipe_v_1 <= sinkVec_1_ready & sinkVec_1_valid;
      accessDataValid_pipe_pipe_v_1 <= accessDataValid_pipe_v_1;
      if (shifterValid_9) begin
        shifterReg_9_0_valid <= accessDataSource_1_valid;
        shifterReg_9_0_bits <= accessDataSource_1_bits;
      end
      sinkVec_releasePipe_pipe_v_2 <= sinkVec_sinkWire_2_ready & sinkVec_sinkWire_2_valid;
      if (sinkVec_validSource_2_valid ^ sinkVec_releasePipe_pipe_out_2_valid)
        sinkVec_tokenCheck_counter_2 <= sinkVec_tokenCheck_counter_2 + sinkVec_tokenCheck_counterChange_2;
      if (sinkVec_shifterValid_2) begin
        sinkVec_shifterReg_2_0_valid <= sinkVec_validSource_2_valid;
        sinkVec_shifterReg_2_0_bits_vd <= sinkVec_validSource_2_bits_vd;
        sinkVec_shifterReg_2_0_bits_offset <= sinkVec_validSource_2_bits_offset;
        sinkVec_shifterReg_2_0_bits_mask <= sinkVec_validSource_2_bits_mask;
        sinkVec_shifterReg_2_0_bits_data <= sinkVec_validSource_2_bits_data;
        sinkVec_shifterReg_2_0_bits_instructionIndex <= sinkVec_validSource_2_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_3 <= sinkVec_sinkWire_3_ready & sinkVec_sinkWire_3_valid;
      if (sinkVec_validSource_3_valid ^ sinkVec_releasePipe_pipe_out_3_valid)
        sinkVec_tokenCheck_counter_3 <= sinkVec_tokenCheck_counter_3 + sinkVec_tokenCheck_counterChange_3;
      if (sinkVec_shifterValid_3) begin
        sinkVec_shifterReg_3_0_valid <= sinkVec_validSource_3_valid;
        sinkVec_shifterReg_3_0_bits_vd <= sinkVec_validSource_3_bits_vd;
        sinkVec_shifterReg_3_0_bits_offset <= sinkVec_validSource_3_bits_offset;
        sinkVec_shifterReg_3_0_bits_mask <= sinkVec_validSource_3_bits_mask;
        sinkVec_shifterReg_3_0_bits_data <= sinkVec_validSource_3_bits_data;
        sinkVec_shifterReg_3_0_bits_last <= sinkVec_validSource_3_bits_last;
        sinkVec_shifterReg_3_0_bits_instructionIndex <= sinkVec_validSource_3_bits_instructionIndex;
      end
      maskUnitFirst_1 <= tryToRead_1 & ~(sinkWire_1_ready & sinkWire_1_valid) ^ maskUnitFirst_1;
      view__writeRelease_0_pipe_v <= sinkVec_1_0_ready & sinkVec_1_0_valid;
      pipe_v <= sinkVec_1_1_ready & sinkVec_1_1_valid;
      instructionFinishedPipe_pipe_v <= 1'h1;
      pipe_v_1 <= 1'h1;
      pipe_pipe_v <= pipe_v_1;
      view__laneMaskSelect_0_pipe_v <= 1'h1;
      view__laneMaskSelect_0_pipe_pipe_v <= view__laneMaskSelect_0_pipe_v;
      view__laneMaskSewSelect_0_pipe_v <= 1'h1;
      view__laneMaskSewSelect_0_pipe_pipe_v <= view__laneMaskSewSelect_0_pipe_v;
      lsuLastPipe_pipe_v <= 1'h1;
      maskLastPipe_pipe_v <= 1'h1;
      pipe_v_2 <= 1'h1;
      sinkVec_releasePipe_pipe_v_4 <= sinkVec_sinkWire_4_ready & sinkVec_sinkWire_4_valid;
      if (sinkVec_validSource_4_valid ^ sinkVec_releasePipe_pipe_out_4_valid)
        sinkVec_tokenCheck_counter_4 <= sinkVec_tokenCheck_counter_4 + sinkVec_tokenCheck_counterChange_4;
      if (sinkVec_shifterValid_4) begin
        sinkVec_shifterReg_4_0_valid <= sinkVec_validSource_4_valid;
        sinkVec_shifterReg_4_0_bits_vs <= sinkVec_validSource_4_bits_vs;
        sinkVec_shifterReg_4_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_4_0_bits_offset <= sinkVec_validSource_4_bits_offset;
        sinkVec_shifterReg_4_0_bits_instructionIndex <= sinkVec_validSource_4_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_5 <= sinkVec_sinkWire_5_ready & sinkVec_sinkWire_5_valid;
      if (sinkVec_validSource_5_valid ^ sinkVec_releasePipe_pipe_out_5_valid)
        sinkVec_tokenCheck_counter_5 <= sinkVec_tokenCheck_counter_5 + sinkVec_tokenCheck_counterChange_5;
      if (sinkVec_shifterValid_5) begin
        sinkVec_shifterReg_5_0_valid <= sinkVec_validSource_5_valid;
        sinkVec_shifterReg_5_0_bits_vs <= sinkVec_validSource_5_bits_vs;
        sinkVec_shifterReg_5_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_5_0_bits_offset <= sinkVec_validSource_5_bits_offset;
        sinkVec_shifterReg_5_0_bits_instructionIndex <= sinkVec_validSource_5_bits_instructionIndex;
      end
      maskUnitFirst_2 <= tryToRead_2 & ~(sinkWire_2_ready & sinkWire_2_valid) ^ maskUnitFirst_2;
      accessDataValid_pipe_v_2 <= sinkVec_2_0_ready & sinkVec_2_0_valid;
      accessDataValid_pipe_pipe_v_2 <= accessDataValid_pipe_v_2;
      if (shifterValid_10) begin
        shifterReg_10_0_valid <= accessDataSource_2_valid;
        shifterReg_10_0_bits <= accessDataSource_2_bits;
      end
      accessDataValid_pipe_v_3 <= sinkVec_2_1_ready & sinkVec_2_1_valid;
      accessDataValid_pipe_pipe_v_3 <= accessDataValid_pipe_v_3;
      if (shifterValid_11) begin
        shifterReg_11_0_valid <= accessDataSource_3_valid;
        shifterReg_11_0_bits <= accessDataSource_3_bits;
      end
      sinkVec_releasePipe_pipe_v_6 <= sinkVec_sinkWire_6_ready & sinkVec_sinkWire_6_valid;
      if (sinkVec_validSource_6_valid ^ sinkVec_releasePipe_pipe_out_6_valid)
        sinkVec_tokenCheck_counter_6 <= sinkVec_tokenCheck_counter_6 + sinkVec_tokenCheck_counterChange_6;
      if (sinkVec_shifterValid_6) begin
        sinkVec_shifterReg_6_0_valid <= sinkVec_validSource_6_valid;
        sinkVec_shifterReg_6_0_bits_vd <= sinkVec_validSource_6_bits_vd;
        sinkVec_shifterReg_6_0_bits_offset <= sinkVec_validSource_6_bits_offset;
        sinkVec_shifterReg_6_0_bits_mask <= sinkVec_validSource_6_bits_mask;
        sinkVec_shifterReg_6_0_bits_data <= sinkVec_validSource_6_bits_data;
        sinkVec_shifterReg_6_0_bits_instructionIndex <= sinkVec_validSource_6_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_7 <= sinkVec_sinkWire_7_ready & sinkVec_sinkWire_7_valid;
      if (sinkVec_validSource_7_valid ^ sinkVec_releasePipe_pipe_out_7_valid)
        sinkVec_tokenCheck_counter_7 <= sinkVec_tokenCheck_counter_7 + sinkVec_tokenCheck_counterChange_7;
      if (sinkVec_shifterValid_7) begin
        sinkVec_shifterReg_7_0_valid <= sinkVec_validSource_7_valid;
        sinkVec_shifterReg_7_0_bits_vd <= sinkVec_validSource_7_bits_vd;
        sinkVec_shifterReg_7_0_bits_offset <= sinkVec_validSource_7_bits_offset;
        sinkVec_shifterReg_7_0_bits_mask <= sinkVec_validSource_7_bits_mask;
        sinkVec_shifterReg_7_0_bits_data <= sinkVec_validSource_7_bits_data;
        sinkVec_shifterReg_7_0_bits_last <= sinkVec_validSource_7_bits_last;
        sinkVec_shifterReg_7_0_bits_instructionIndex <= sinkVec_validSource_7_bits_instructionIndex;
      end
      maskUnitFirst_3 <= tryToRead_3 & ~(sinkWire_3_ready & sinkWire_3_valid) ^ maskUnitFirst_3;
      view__writeRelease_1_pipe_v <= sinkVec_3_0_ready & sinkVec_3_0_valid;
      pipe_v_3 <= sinkVec_3_1_ready & sinkVec_3_1_valid;
      instructionFinishedPipe_pipe_v_1 <= 1'h1;
      pipe_v_4 <= 1'h1;
      pipe_pipe_v_1 <= pipe_v_4;
      view__laneMaskSelect_1_pipe_v <= 1'h1;
      view__laneMaskSelect_1_pipe_pipe_v <= view__laneMaskSelect_1_pipe_v;
      view__laneMaskSewSelect_1_pipe_v <= 1'h1;
      view__laneMaskSewSelect_1_pipe_pipe_v <= view__laneMaskSewSelect_1_pipe_v;
      lsuLastPipe_pipe_v_1 <= 1'h1;
      maskLastPipe_pipe_v_1 <= 1'h1;
      pipe_v_5 <= 1'h1;
      sinkVec_releasePipe_pipe_v_8 <= sinkVec_sinkWire_8_ready & sinkVec_sinkWire_8_valid;
      if (sinkVec_validSource_8_valid ^ sinkVec_releasePipe_pipe_out_8_valid)
        sinkVec_tokenCheck_counter_8 <= sinkVec_tokenCheck_counter_8 + sinkVec_tokenCheck_counterChange_8;
      if (sinkVec_shifterValid_8) begin
        sinkVec_shifterReg_8_0_valid <= sinkVec_validSource_8_valid;
        sinkVec_shifterReg_8_0_bits_vs <= sinkVec_validSource_8_bits_vs;
        sinkVec_shifterReg_8_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_8_0_bits_offset <= sinkVec_validSource_8_bits_offset;
        sinkVec_shifterReg_8_0_bits_instructionIndex <= sinkVec_validSource_8_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_9 <= sinkVec_sinkWire_9_ready & sinkVec_sinkWire_9_valid;
      if (sinkVec_validSource_9_valid ^ sinkVec_releasePipe_pipe_out_9_valid)
        sinkVec_tokenCheck_counter_9 <= sinkVec_tokenCheck_counter_9 + sinkVec_tokenCheck_counterChange_9;
      if (sinkVec_shifterValid_9) begin
        sinkVec_shifterReg_9_0_valid <= sinkVec_validSource_9_valid;
        sinkVec_shifterReg_9_0_bits_vs <= sinkVec_validSource_9_bits_vs;
        sinkVec_shifterReg_9_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_9_0_bits_offset <= sinkVec_validSource_9_bits_offset;
        sinkVec_shifterReg_9_0_bits_instructionIndex <= sinkVec_validSource_9_bits_instructionIndex;
      end
      maskUnitFirst_4 <= tryToRead_4 & ~(sinkWire_4_ready & sinkWire_4_valid) ^ maskUnitFirst_4;
      accessDataValid_pipe_v_4 <= sinkVec_4_0_ready & sinkVec_4_0_valid;
      accessDataValid_pipe_pipe_v_4 <= accessDataValid_pipe_v_4;
      if (shifterValid_12) begin
        shifterReg_12_0_valid <= accessDataSource_4_valid;
        shifterReg_12_0_bits <= accessDataSource_4_bits;
      end
      accessDataValid_pipe_v_5 <= sinkVec_4_1_ready & sinkVec_4_1_valid;
      accessDataValid_pipe_pipe_v_5 <= accessDataValid_pipe_v_5;
      if (shifterValid_13) begin
        shifterReg_13_0_valid <= accessDataSource_5_valid;
        shifterReg_13_0_bits <= accessDataSource_5_bits;
      end
      sinkVec_releasePipe_pipe_v_10 <= sinkVec_sinkWire_10_ready & sinkVec_sinkWire_10_valid;
      if (sinkVec_validSource_10_valid ^ sinkVec_releasePipe_pipe_out_10_valid)
        sinkVec_tokenCheck_counter_10 <= sinkVec_tokenCheck_counter_10 + sinkVec_tokenCheck_counterChange_10;
      if (sinkVec_shifterValid_10) begin
        sinkVec_shifterReg_10_0_valid <= sinkVec_validSource_10_valid;
        sinkVec_shifterReg_10_0_bits_vd <= sinkVec_validSource_10_bits_vd;
        sinkVec_shifterReg_10_0_bits_offset <= sinkVec_validSource_10_bits_offset;
        sinkVec_shifterReg_10_0_bits_mask <= sinkVec_validSource_10_bits_mask;
        sinkVec_shifterReg_10_0_bits_data <= sinkVec_validSource_10_bits_data;
        sinkVec_shifterReg_10_0_bits_instructionIndex <= sinkVec_validSource_10_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_11 <= sinkVec_sinkWire_11_ready & sinkVec_sinkWire_11_valid;
      if (sinkVec_validSource_11_valid ^ sinkVec_releasePipe_pipe_out_11_valid)
        sinkVec_tokenCheck_counter_11 <= sinkVec_tokenCheck_counter_11 + sinkVec_tokenCheck_counterChange_11;
      if (sinkVec_shifterValid_11) begin
        sinkVec_shifterReg_11_0_valid <= sinkVec_validSource_11_valid;
        sinkVec_shifterReg_11_0_bits_vd <= sinkVec_validSource_11_bits_vd;
        sinkVec_shifterReg_11_0_bits_offset <= sinkVec_validSource_11_bits_offset;
        sinkVec_shifterReg_11_0_bits_mask <= sinkVec_validSource_11_bits_mask;
        sinkVec_shifterReg_11_0_bits_data <= sinkVec_validSource_11_bits_data;
        sinkVec_shifterReg_11_0_bits_last <= sinkVec_validSource_11_bits_last;
        sinkVec_shifterReg_11_0_bits_instructionIndex <= sinkVec_validSource_11_bits_instructionIndex;
      end
      maskUnitFirst_5 <= tryToRead_5 & ~(sinkWire_5_ready & sinkWire_5_valid) ^ maskUnitFirst_5;
      view__writeRelease_2_pipe_v <= sinkVec_5_0_ready & sinkVec_5_0_valid;
      pipe_v_6 <= sinkVec_5_1_ready & sinkVec_5_1_valid;
      instructionFinishedPipe_pipe_v_2 <= 1'h1;
      pipe_v_7 <= 1'h1;
      pipe_pipe_v_2 <= pipe_v_7;
      view__laneMaskSelect_2_pipe_v <= 1'h1;
      view__laneMaskSelect_2_pipe_pipe_v <= view__laneMaskSelect_2_pipe_v;
      view__laneMaskSewSelect_2_pipe_v <= 1'h1;
      view__laneMaskSewSelect_2_pipe_pipe_v <= view__laneMaskSewSelect_2_pipe_v;
      lsuLastPipe_pipe_v_2 <= 1'h1;
      maskLastPipe_pipe_v_2 <= 1'h1;
      pipe_v_8 <= 1'h1;
      sinkVec_releasePipe_pipe_v_12 <= sinkVec_sinkWire_12_ready & sinkVec_sinkWire_12_valid;
      if (sinkVec_validSource_12_valid ^ sinkVec_releasePipe_pipe_out_12_valid)
        sinkVec_tokenCheck_counter_12 <= sinkVec_tokenCheck_counter_12 + sinkVec_tokenCheck_counterChange_12;
      if (sinkVec_shifterValid_12) begin
        sinkVec_shifterReg_12_0_valid <= sinkVec_validSource_12_valid;
        sinkVec_shifterReg_12_0_bits_vs <= sinkVec_validSource_12_bits_vs;
        sinkVec_shifterReg_12_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_12_0_bits_offset <= sinkVec_validSource_12_bits_offset;
        sinkVec_shifterReg_12_0_bits_instructionIndex <= sinkVec_validSource_12_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_13 <= sinkVec_sinkWire_13_ready & sinkVec_sinkWire_13_valid;
      if (sinkVec_validSource_13_valid ^ sinkVec_releasePipe_pipe_out_13_valid)
        sinkVec_tokenCheck_counter_13 <= sinkVec_tokenCheck_counter_13 + sinkVec_tokenCheck_counterChange_13;
      if (sinkVec_shifterValid_13) begin
        sinkVec_shifterReg_13_0_valid <= sinkVec_validSource_13_valid;
        sinkVec_shifterReg_13_0_bits_vs <= sinkVec_validSource_13_bits_vs;
        sinkVec_shifterReg_13_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_13_0_bits_offset <= sinkVec_validSource_13_bits_offset;
        sinkVec_shifterReg_13_0_bits_instructionIndex <= sinkVec_validSource_13_bits_instructionIndex;
      end
      maskUnitFirst_6 <= tryToRead_6 & ~(sinkWire_6_ready & sinkWire_6_valid) ^ maskUnitFirst_6;
      accessDataValid_pipe_v_6 <= sinkVec_6_0_ready & sinkVec_6_0_valid;
      accessDataValid_pipe_pipe_v_6 <= accessDataValid_pipe_v_6;
      if (shifterValid_14) begin
        shifterReg_14_0_valid <= accessDataSource_6_valid;
        shifterReg_14_0_bits <= accessDataSource_6_bits;
      end
      accessDataValid_pipe_v_7 <= sinkVec_6_1_ready & sinkVec_6_1_valid;
      accessDataValid_pipe_pipe_v_7 <= accessDataValid_pipe_v_7;
      if (shifterValid_15) begin
        shifterReg_15_0_valid <= accessDataSource_7_valid;
        shifterReg_15_0_bits <= accessDataSource_7_bits;
      end
      sinkVec_releasePipe_pipe_v_14 <= sinkVec_sinkWire_14_ready & sinkVec_sinkWire_14_valid;
      if (sinkVec_validSource_14_valid ^ sinkVec_releasePipe_pipe_out_14_valid)
        sinkVec_tokenCheck_counter_14 <= sinkVec_tokenCheck_counter_14 + sinkVec_tokenCheck_counterChange_14;
      if (sinkVec_shifterValid_14) begin
        sinkVec_shifterReg_14_0_valid <= sinkVec_validSource_14_valid;
        sinkVec_shifterReg_14_0_bits_vd <= sinkVec_validSource_14_bits_vd;
        sinkVec_shifterReg_14_0_bits_offset <= sinkVec_validSource_14_bits_offset;
        sinkVec_shifterReg_14_0_bits_mask <= sinkVec_validSource_14_bits_mask;
        sinkVec_shifterReg_14_0_bits_data <= sinkVec_validSource_14_bits_data;
        sinkVec_shifterReg_14_0_bits_instructionIndex <= sinkVec_validSource_14_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_15 <= sinkVec_sinkWire_15_ready & sinkVec_sinkWire_15_valid;
      if (sinkVec_validSource_15_valid ^ sinkVec_releasePipe_pipe_out_15_valid)
        sinkVec_tokenCheck_counter_15 <= sinkVec_tokenCheck_counter_15 + sinkVec_tokenCheck_counterChange_15;
      if (sinkVec_shifterValid_15) begin
        sinkVec_shifterReg_15_0_valid <= sinkVec_validSource_15_valid;
        sinkVec_shifterReg_15_0_bits_vd <= sinkVec_validSource_15_bits_vd;
        sinkVec_shifterReg_15_0_bits_offset <= sinkVec_validSource_15_bits_offset;
        sinkVec_shifterReg_15_0_bits_mask <= sinkVec_validSource_15_bits_mask;
        sinkVec_shifterReg_15_0_bits_data <= sinkVec_validSource_15_bits_data;
        sinkVec_shifterReg_15_0_bits_last <= sinkVec_validSource_15_bits_last;
        sinkVec_shifterReg_15_0_bits_instructionIndex <= sinkVec_validSource_15_bits_instructionIndex;
      end
      maskUnitFirst_7 <= tryToRead_7 & ~(sinkWire_7_ready & sinkWire_7_valid) ^ maskUnitFirst_7;
      view__writeRelease_3_pipe_v <= sinkVec_7_0_ready & sinkVec_7_0_valid;
      pipe_v_9 <= sinkVec_7_1_ready & sinkVec_7_1_valid;
      instructionFinishedPipe_pipe_v_3 <= 1'h1;
      pipe_v_10 <= 1'h1;
      pipe_pipe_v_3 <= pipe_v_10;
      view__laneMaskSelect_3_pipe_v <= 1'h1;
      view__laneMaskSelect_3_pipe_pipe_v <= view__laneMaskSelect_3_pipe_v;
      view__laneMaskSewSelect_3_pipe_v <= 1'h1;
      view__laneMaskSewSelect_3_pipe_pipe_v <= view__laneMaskSewSelect_3_pipe_v;
      lsuLastPipe_pipe_v_3 <= 1'h1;
      maskLastPipe_pipe_v_3 <= 1'h1;
      pipe_v_11 <= 1'h1;
      sinkVec_releasePipe_pipe_v_16 <= sinkVec_sinkWire_16_ready & sinkVec_sinkWire_16_valid;
      if (sinkVec_validSource_16_valid ^ sinkVec_releasePipe_pipe_out_16_valid)
        sinkVec_tokenCheck_counter_16 <= sinkVec_tokenCheck_counter_16 + sinkVec_tokenCheck_counterChange_16;
      if (sinkVec_shifterValid_16) begin
        sinkVec_shifterReg_16_0_valid <= sinkVec_validSource_16_valid;
        sinkVec_shifterReg_16_0_bits_vs <= sinkVec_validSource_16_bits_vs;
        sinkVec_shifterReg_16_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_16_0_bits_offset <= sinkVec_validSource_16_bits_offset;
        sinkVec_shifterReg_16_0_bits_instructionIndex <= sinkVec_validSource_16_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_17 <= sinkVec_sinkWire_17_ready & sinkVec_sinkWire_17_valid;
      if (sinkVec_validSource_17_valid ^ sinkVec_releasePipe_pipe_out_17_valid)
        sinkVec_tokenCheck_counter_17 <= sinkVec_tokenCheck_counter_17 + sinkVec_tokenCheck_counterChange_17;
      if (sinkVec_shifterValid_17) begin
        sinkVec_shifterReg_17_0_valid <= sinkVec_validSource_17_valid;
        sinkVec_shifterReg_17_0_bits_vs <= sinkVec_validSource_17_bits_vs;
        sinkVec_shifterReg_17_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_17_0_bits_offset <= sinkVec_validSource_17_bits_offset;
        sinkVec_shifterReg_17_0_bits_instructionIndex <= sinkVec_validSource_17_bits_instructionIndex;
      end
      maskUnitFirst_8 <= tryToRead_8 & ~(sinkWire_8_ready & sinkWire_8_valid) ^ maskUnitFirst_8;
      accessDataValid_pipe_v_8 <= sinkVec_8_0_ready & sinkVec_8_0_valid;
      accessDataValid_pipe_pipe_v_8 <= accessDataValid_pipe_v_8;
      if (shifterValid_16) begin
        shifterReg_16_0_valid <= accessDataSource_8_valid;
        shifterReg_16_0_bits <= accessDataSource_8_bits;
      end
      accessDataValid_pipe_v_9 <= sinkVec_8_1_ready & sinkVec_8_1_valid;
      accessDataValid_pipe_pipe_v_9 <= accessDataValid_pipe_v_9;
      if (shifterValid_17) begin
        shifterReg_17_0_valid <= accessDataSource_9_valid;
        shifterReg_17_0_bits <= accessDataSource_9_bits;
      end
      sinkVec_releasePipe_pipe_v_18 <= sinkVec_sinkWire_18_ready & sinkVec_sinkWire_18_valid;
      if (sinkVec_validSource_18_valid ^ sinkVec_releasePipe_pipe_out_18_valid)
        sinkVec_tokenCheck_counter_18 <= sinkVec_tokenCheck_counter_18 + sinkVec_tokenCheck_counterChange_18;
      if (sinkVec_shifterValid_18) begin
        sinkVec_shifterReg_18_0_valid <= sinkVec_validSource_18_valid;
        sinkVec_shifterReg_18_0_bits_vd <= sinkVec_validSource_18_bits_vd;
        sinkVec_shifterReg_18_0_bits_offset <= sinkVec_validSource_18_bits_offset;
        sinkVec_shifterReg_18_0_bits_mask <= sinkVec_validSource_18_bits_mask;
        sinkVec_shifterReg_18_0_bits_data <= sinkVec_validSource_18_bits_data;
        sinkVec_shifterReg_18_0_bits_instructionIndex <= sinkVec_validSource_18_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_19 <= sinkVec_sinkWire_19_ready & sinkVec_sinkWire_19_valid;
      if (sinkVec_validSource_19_valid ^ sinkVec_releasePipe_pipe_out_19_valid)
        sinkVec_tokenCheck_counter_19 <= sinkVec_tokenCheck_counter_19 + sinkVec_tokenCheck_counterChange_19;
      if (sinkVec_shifterValid_19) begin
        sinkVec_shifterReg_19_0_valid <= sinkVec_validSource_19_valid;
        sinkVec_shifterReg_19_0_bits_vd <= sinkVec_validSource_19_bits_vd;
        sinkVec_shifterReg_19_0_bits_offset <= sinkVec_validSource_19_bits_offset;
        sinkVec_shifterReg_19_0_bits_mask <= sinkVec_validSource_19_bits_mask;
        sinkVec_shifterReg_19_0_bits_data <= sinkVec_validSource_19_bits_data;
        sinkVec_shifterReg_19_0_bits_last <= sinkVec_validSource_19_bits_last;
        sinkVec_shifterReg_19_0_bits_instructionIndex <= sinkVec_validSource_19_bits_instructionIndex;
      end
      maskUnitFirst_9 <= tryToRead_9 & ~(sinkWire_9_ready & sinkWire_9_valid) ^ maskUnitFirst_9;
      view__writeRelease_4_pipe_v <= sinkVec_9_0_ready & sinkVec_9_0_valid;
      pipe_v_12 <= sinkVec_9_1_ready & sinkVec_9_1_valid;
      instructionFinishedPipe_pipe_v_4 <= 1'h1;
      pipe_v_13 <= 1'h1;
      pipe_pipe_v_4 <= pipe_v_13;
      view__laneMaskSelect_4_pipe_v <= 1'h1;
      view__laneMaskSelect_4_pipe_pipe_v <= view__laneMaskSelect_4_pipe_v;
      view__laneMaskSewSelect_4_pipe_v <= 1'h1;
      view__laneMaskSewSelect_4_pipe_pipe_v <= view__laneMaskSewSelect_4_pipe_v;
      lsuLastPipe_pipe_v_4 <= 1'h1;
      maskLastPipe_pipe_v_4 <= 1'h1;
      pipe_v_14 <= 1'h1;
      sinkVec_releasePipe_pipe_v_20 <= sinkVec_sinkWire_20_ready & sinkVec_sinkWire_20_valid;
      if (sinkVec_validSource_20_valid ^ sinkVec_releasePipe_pipe_out_20_valid)
        sinkVec_tokenCheck_counter_20 <= sinkVec_tokenCheck_counter_20 + sinkVec_tokenCheck_counterChange_20;
      if (sinkVec_shifterValid_20) begin
        sinkVec_shifterReg_20_0_valid <= sinkVec_validSource_20_valid;
        sinkVec_shifterReg_20_0_bits_vs <= sinkVec_validSource_20_bits_vs;
        sinkVec_shifterReg_20_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_20_0_bits_offset <= sinkVec_validSource_20_bits_offset;
        sinkVec_shifterReg_20_0_bits_instructionIndex <= sinkVec_validSource_20_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_21 <= sinkVec_sinkWire_21_ready & sinkVec_sinkWire_21_valid;
      if (sinkVec_validSource_21_valid ^ sinkVec_releasePipe_pipe_out_21_valid)
        sinkVec_tokenCheck_counter_21 <= sinkVec_tokenCheck_counter_21 + sinkVec_tokenCheck_counterChange_21;
      if (sinkVec_shifterValid_21) begin
        sinkVec_shifterReg_21_0_valid <= sinkVec_validSource_21_valid;
        sinkVec_shifterReg_21_0_bits_vs <= sinkVec_validSource_21_bits_vs;
        sinkVec_shifterReg_21_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_21_0_bits_offset <= sinkVec_validSource_21_bits_offset;
        sinkVec_shifterReg_21_0_bits_instructionIndex <= sinkVec_validSource_21_bits_instructionIndex;
      end
      maskUnitFirst_10 <= tryToRead_10 & ~(sinkWire_10_ready & sinkWire_10_valid) ^ maskUnitFirst_10;
      accessDataValid_pipe_v_10 <= sinkVec_10_0_ready & sinkVec_10_0_valid;
      accessDataValid_pipe_pipe_v_10 <= accessDataValid_pipe_v_10;
      if (shifterValid_18) begin
        shifterReg_18_0_valid <= accessDataSource_10_valid;
        shifterReg_18_0_bits <= accessDataSource_10_bits;
      end
      accessDataValid_pipe_v_11 <= sinkVec_10_1_ready & sinkVec_10_1_valid;
      accessDataValid_pipe_pipe_v_11 <= accessDataValid_pipe_v_11;
      if (shifterValid_19) begin
        shifterReg_19_0_valid <= accessDataSource_11_valid;
        shifterReg_19_0_bits <= accessDataSource_11_bits;
      end
      sinkVec_releasePipe_pipe_v_22 <= sinkVec_sinkWire_22_ready & sinkVec_sinkWire_22_valid;
      if (sinkVec_validSource_22_valid ^ sinkVec_releasePipe_pipe_out_22_valid)
        sinkVec_tokenCheck_counter_22 <= sinkVec_tokenCheck_counter_22 + sinkVec_tokenCheck_counterChange_22;
      if (sinkVec_shifterValid_22) begin
        sinkVec_shifterReg_22_0_valid <= sinkVec_validSource_22_valid;
        sinkVec_shifterReg_22_0_bits_vd <= sinkVec_validSource_22_bits_vd;
        sinkVec_shifterReg_22_0_bits_offset <= sinkVec_validSource_22_bits_offset;
        sinkVec_shifterReg_22_0_bits_mask <= sinkVec_validSource_22_bits_mask;
        sinkVec_shifterReg_22_0_bits_data <= sinkVec_validSource_22_bits_data;
        sinkVec_shifterReg_22_0_bits_instructionIndex <= sinkVec_validSource_22_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_23 <= sinkVec_sinkWire_23_ready & sinkVec_sinkWire_23_valid;
      if (sinkVec_validSource_23_valid ^ sinkVec_releasePipe_pipe_out_23_valid)
        sinkVec_tokenCheck_counter_23 <= sinkVec_tokenCheck_counter_23 + sinkVec_tokenCheck_counterChange_23;
      if (sinkVec_shifterValid_23) begin
        sinkVec_shifterReg_23_0_valid <= sinkVec_validSource_23_valid;
        sinkVec_shifterReg_23_0_bits_vd <= sinkVec_validSource_23_bits_vd;
        sinkVec_shifterReg_23_0_bits_offset <= sinkVec_validSource_23_bits_offset;
        sinkVec_shifterReg_23_0_bits_mask <= sinkVec_validSource_23_bits_mask;
        sinkVec_shifterReg_23_0_bits_data <= sinkVec_validSource_23_bits_data;
        sinkVec_shifterReg_23_0_bits_last <= sinkVec_validSource_23_bits_last;
        sinkVec_shifterReg_23_0_bits_instructionIndex <= sinkVec_validSource_23_bits_instructionIndex;
      end
      maskUnitFirst_11 <= tryToRead_11 & ~(sinkWire_11_ready & sinkWire_11_valid) ^ maskUnitFirst_11;
      view__writeRelease_5_pipe_v <= sinkVec_11_0_ready & sinkVec_11_0_valid;
      pipe_v_15 <= sinkVec_11_1_ready & sinkVec_11_1_valid;
      instructionFinishedPipe_pipe_v_5 <= 1'h1;
      pipe_v_16 <= 1'h1;
      pipe_pipe_v_5 <= pipe_v_16;
      view__laneMaskSelect_5_pipe_v <= 1'h1;
      view__laneMaskSelect_5_pipe_pipe_v <= view__laneMaskSelect_5_pipe_v;
      view__laneMaskSewSelect_5_pipe_v <= 1'h1;
      view__laneMaskSewSelect_5_pipe_pipe_v <= view__laneMaskSewSelect_5_pipe_v;
      lsuLastPipe_pipe_v_5 <= 1'h1;
      maskLastPipe_pipe_v_5 <= 1'h1;
      pipe_v_17 <= 1'h1;
      sinkVec_releasePipe_pipe_v_24 <= sinkVec_sinkWire_24_ready & sinkVec_sinkWire_24_valid;
      if (sinkVec_validSource_24_valid ^ sinkVec_releasePipe_pipe_out_24_valid)
        sinkVec_tokenCheck_counter_24 <= sinkVec_tokenCheck_counter_24 + sinkVec_tokenCheck_counterChange_24;
      if (sinkVec_shifterValid_24) begin
        sinkVec_shifterReg_24_0_valid <= sinkVec_validSource_24_valid;
        sinkVec_shifterReg_24_0_bits_vs <= sinkVec_validSource_24_bits_vs;
        sinkVec_shifterReg_24_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_24_0_bits_offset <= sinkVec_validSource_24_bits_offset;
        sinkVec_shifterReg_24_0_bits_instructionIndex <= sinkVec_validSource_24_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_25 <= sinkVec_sinkWire_25_ready & sinkVec_sinkWire_25_valid;
      if (sinkVec_validSource_25_valid ^ sinkVec_releasePipe_pipe_out_25_valid)
        sinkVec_tokenCheck_counter_25 <= sinkVec_tokenCheck_counter_25 + sinkVec_tokenCheck_counterChange_25;
      if (sinkVec_shifterValid_25) begin
        sinkVec_shifterReg_25_0_valid <= sinkVec_validSource_25_valid;
        sinkVec_shifterReg_25_0_bits_vs <= sinkVec_validSource_25_bits_vs;
        sinkVec_shifterReg_25_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_25_0_bits_offset <= sinkVec_validSource_25_bits_offset;
        sinkVec_shifterReg_25_0_bits_instructionIndex <= sinkVec_validSource_25_bits_instructionIndex;
      end
      maskUnitFirst_12 <= tryToRead_12 & ~(sinkWire_12_ready & sinkWire_12_valid) ^ maskUnitFirst_12;
      accessDataValid_pipe_v_12 <= sinkVec_12_0_ready & sinkVec_12_0_valid;
      accessDataValid_pipe_pipe_v_12 <= accessDataValid_pipe_v_12;
      if (shifterValid_20) begin
        shifterReg_20_0_valid <= accessDataSource_12_valid;
        shifterReg_20_0_bits <= accessDataSource_12_bits;
      end
      accessDataValid_pipe_v_13 <= sinkVec_12_1_ready & sinkVec_12_1_valid;
      accessDataValid_pipe_pipe_v_13 <= accessDataValid_pipe_v_13;
      if (shifterValid_21) begin
        shifterReg_21_0_valid <= accessDataSource_13_valid;
        shifterReg_21_0_bits <= accessDataSource_13_bits;
      end
      sinkVec_releasePipe_pipe_v_26 <= sinkVec_sinkWire_26_ready & sinkVec_sinkWire_26_valid;
      if (sinkVec_validSource_26_valid ^ sinkVec_releasePipe_pipe_out_26_valid)
        sinkVec_tokenCheck_counter_26 <= sinkVec_tokenCheck_counter_26 + sinkVec_tokenCheck_counterChange_26;
      if (sinkVec_shifterValid_26) begin
        sinkVec_shifterReg_26_0_valid <= sinkVec_validSource_26_valid;
        sinkVec_shifterReg_26_0_bits_vd <= sinkVec_validSource_26_bits_vd;
        sinkVec_shifterReg_26_0_bits_offset <= sinkVec_validSource_26_bits_offset;
        sinkVec_shifterReg_26_0_bits_mask <= sinkVec_validSource_26_bits_mask;
        sinkVec_shifterReg_26_0_bits_data <= sinkVec_validSource_26_bits_data;
        sinkVec_shifterReg_26_0_bits_instructionIndex <= sinkVec_validSource_26_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_27 <= sinkVec_sinkWire_27_ready & sinkVec_sinkWire_27_valid;
      if (sinkVec_validSource_27_valid ^ sinkVec_releasePipe_pipe_out_27_valid)
        sinkVec_tokenCheck_counter_27 <= sinkVec_tokenCheck_counter_27 + sinkVec_tokenCheck_counterChange_27;
      if (sinkVec_shifterValid_27) begin
        sinkVec_shifterReg_27_0_valid <= sinkVec_validSource_27_valid;
        sinkVec_shifterReg_27_0_bits_vd <= sinkVec_validSource_27_bits_vd;
        sinkVec_shifterReg_27_0_bits_offset <= sinkVec_validSource_27_bits_offset;
        sinkVec_shifterReg_27_0_bits_mask <= sinkVec_validSource_27_bits_mask;
        sinkVec_shifterReg_27_0_bits_data <= sinkVec_validSource_27_bits_data;
        sinkVec_shifterReg_27_0_bits_last <= sinkVec_validSource_27_bits_last;
        sinkVec_shifterReg_27_0_bits_instructionIndex <= sinkVec_validSource_27_bits_instructionIndex;
      end
      maskUnitFirst_13 <= tryToRead_13 & ~(sinkWire_13_ready & sinkWire_13_valid) ^ maskUnitFirst_13;
      view__writeRelease_6_pipe_v <= sinkVec_13_0_ready & sinkVec_13_0_valid;
      pipe_v_18 <= sinkVec_13_1_ready & sinkVec_13_1_valid;
      instructionFinishedPipe_pipe_v_6 <= 1'h1;
      pipe_v_19 <= 1'h1;
      pipe_pipe_v_6 <= pipe_v_19;
      view__laneMaskSelect_6_pipe_v <= 1'h1;
      view__laneMaskSelect_6_pipe_pipe_v <= view__laneMaskSelect_6_pipe_v;
      view__laneMaskSewSelect_6_pipe_v <= 1'h1;
      view__laneMaskSewSelect_6_pipe_pipe_v <= view__laneMaskSewSelect_6_pipe_v;
      lsuLastPipe_pipe_v_6 <= 1'h1;
      maskLastPipe_pipe_v_6 <= 1'h1;
      pipe_v_20 <= 1'h1;
      sinkVec_releasePipe_pipe_v_28 <= sinkVec_sinkWire_28_ready & sinkVec_sinkWire_28_valid;
      if (sinkVec_validSource_28_valid ^ sinkVec_releasePipe_pipe_out_28_valid)
        sinkVec_tokenCheck_counter_28 <= sinkVec_tokenCheck_counter_28 + sinkVec_tokenCheck_counterChange_28;
      if (sinkVec_shifterValid_28) begin
        sinkVec_shifterReg_28_0_valid <= sinkVec_validSource_28_valid;
        sinkVec_shifterReg_28_0_bits_vs <= sinkVec_validSource_28_bits_vs;
        sinkVec_shifterReg_28_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_28_0_bits_offset <= sinkVec_validSource_28_bits_offset;
        sinkVec_shifterReg_28_0_bits_instructionIndex <= sinkVec_validSource_28_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_29 <= sinkVec_sinkWire_29_ready & sinkVec_sinkWire_29_valid;
      if (sinkVec_validSource_29_valid ^ sinkVec_releasePipe_pipe_out_29_valid)
        sinkVec_tokenCheck_counter_29 <= sinkVec_tokenCheck_counter_29 + sinkVec_tokenCheck_counterChange_29;
      if (sinkVec_shifterValid_29) begin
        sinkVec_shifterReg_29_0_valid <= sinkVec_validSource_29_valid;
        sinkVec_shifterReg_29_0_bits_vs <= sinkVec_validSource_29_bits_vs;
        sinkVec_shifterReg_29_0_bits_readSource <= 2'h2;
        sinkVec_shifterReg_29_0_bits_offset <= sinkVec_validSource_29_bits_offset;
        sinkVec_shifterReg_29_0_bits_instructionIndex <= sinkVec_validSource_29_bits_instructionIndex;
      end
      maskUnitFirst_14 <= tryToRead_14 & ~(sinkWire_14_ready & sinkWire_14_valid) ^ maskUnitFirst_14;
      accessDataValid_pipe_v_14 <= sinkVec_14_0_ready & sinkVec_14_0_valid;
      accessDataValid_pipe_pipe_v_14 <= accessDataValid_pipe_v_14;
      if (shifterValid_22) begin
        shifterReg_22_0_valid <= accessDataSource_14_valid;
        shifterReg_22_0_bits <= accessDataSource_14_bits;
      end
      accessDataValid_pipe_v_15 <= sinkVec_14_1_ready & sinkVec_14_1_valid;
      accessDataValid_pipe_pipe_v_15 <= accessDataValid_pipe_v_15;
      if (shifterValid_23) begin
        shifterReg_23_0_valid <= accessDataSource_15_valid;
        shifterReg_23_0_bits <= accessDataSource_15_bits;
      end
      sinkVec_releasePipe_pipe_v_30 <= sinkVec_sinkWire_30_ready & sinkVec_sinkWire_30_valid;
      if (sinkVec_validSource_30_valid ^ sinkVec_releasePipe_pipe_out_30_valid)
        sinkVec_tokenCheck_counter_30 <= sinkVec_tokenCheck_counter_30 + sinkVec_tokenCheck_counterChange_30;
      if (sinkVec_shifterValid_30) begin
        sinkVec_shifterReg_30_0_valid <= sinkVec_validSource_30_valid;
        sinkVec_shifterReg_30_0_bits_vd <= sinkVec_validSource_30_bits_vd;
        sinkVec_shifterReg_30_0_bits_offset <= sinkVec_validSource_30_bits_offset;
        sinkVec_shifterReg_30_0_bits_mask <= sinkVec_validSource_30_bits_mask;
        sinkVec_shifterReg_30_0_bits_data <= sinkVec_validSource_30_bits_data;
        sinkVec_shifterReg_30_0_bits_instructionIndex <= sinkVec_validSource_30_bits_instructionIndex;
      end
      sinkVec_releasePipe_pipe_v_31 <= sinkVec_sinkWire_31_ready & sinkVec_sinkWire_31_valid;
      if (sinkVec_validSource_31_valid ^ sinkVec_releasePipe_pipe_out_31_valid)
        sinkVec_tokenCheck_counter_31 <= sinkVec_tokenCheck_counter_31 + sinkVec_tokenCheck_counterChange_31;
      if (sinkVec_shifterValid_31) begin
        sinkVec_shifterReg_31_0_valid <= sinkVec_validSource_31_valid;
        sinkVec_shifterReg_31_0_bits_vd <= sinkVec_validSource_31_bits_vd;
        sinkVec_shifterReg_31_0_bits_offset <= sinkVec_validSource_31_bits_offset;
        sinkVec_shifterReg_31_0_bits_mask <= sinkVec_validSource_31_bits_mask;
        sinkVec_shifterReg_31_0_bits_data <= sinkVec_validSource_31_bits_data;
        sinkVec_shifterReg_31_0_bits_last <= sinkVec_validSource_31_bits_last;
        sinkVec_shifterReg_31_0_bits_instructionIndex <= sinkVec_validSource_31_bits_instructionIndex;
      end
      maskUnitFirst_15 <= tryToRead_15 & ~(sinkWire_15_ready & sinkWire_15_valid) ^ maskUnitFirst_15;
      view__writeRelease_7_pipe_v <= sinkVec_15_0_ready & sinkVec_15_0_valid;
      pipe_v_21 <= sinkVec_15_1_ready & sinkVec_15_1_valid;
      instructionFinishedPipe_pipe_v_7 <= 1'h1;
      pipe_v_22 <= 1'h1;
      pipe_pipe_v_7 <= pipe_v_22;
      view__laneMaskSelect_7_pipe_v <= 1'h1;
      view__laneMaskSelect_7_pipe_pipe_v <= view__laneMaskSelect_7_pipe_v;
      view__laneMaskSewSelect_7_pipe_v <= 1'h1;
      view__laneMaskSewSelect_7_pipe_pipe_v <= view__laneMaskSewSelect_7_pipe_v;
      lsuLastPipe_pipe_v_7 <= 1'h1;
      maskLastPipe_pipe_v_7 <= 1'h1;
      pipe_v_23 <= 1'h1;
      pipe_v_24 <= _laneVec_0_readBusPort_0_enqRelease;
      if (shifterValid_24) begin
        shifterReg_24_0_valid <= _laneVec_0_readBusPort_0_deq_valid;
        shifterReg_24_0_bits_data <= _laneVec_0_readBusPort_0_deq_bits_data;
      end
      pipe_v_25 <= _laneVec_0_writeBusPort_0_enqRelease;
      if (shifterValid_25) begin
        shifterReg_25_0_valid <= _laneVec_0_writeBusPort_0_deq_valid;
        shifterReg_25_0_bits_data <= _laneVec_0_writeBusPort_0_deq_bits_data;
        shifterReg_25_0_bits_mask <= _laneVec_0_writeBusPort_0_deq_bits_mask;
        shifterReg_25_0_bits_instructionIndex <= _laneVec_0_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_25_0_bits_counter <= _laneVec_0_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_26 <= _laneVec_0_readBusPort_1_enqRelease;
      if (shifterValid_26) begin
        shifterReg_26_0_valid <= _laneVec_1_readBusPort_0_deq_valid;
        shifterReg_26_0_bits_data <= _laneVec_1_readBusPort_0_deq_bits_data;
      end
      pipe_v_27 <= _laneVec_1_writeBusPort_0_enqRelease;
      if (shifterValid_27) begin
        shifterReg_27_0_valid <= _laneVec_0_writeBusPort_1_deq_valid;
        shifterReg_27_0_bits_data <= _laneVec_0_writeBusPort_1_deq_bits_data;
        shifterReg_27_0_bits_mask <= _laneVec_0_writeBusPort_1_deq_bits_mask;
        shifterReg_27_0_bits_instructionIndex <= _laneVec_0_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_27_0_bits_counter <= _laneVec_0_writeBusPort_1_deq_bits_counter;
      end
      pipe_v_28 <= _laneVec_1_readBusPort_0_enqRelease;
      if (shifterValid_28) begin
        shifterReg_28_0_valid <= _laneVec_2_readBusPort_0_deq_valid;
        shifterReg_28_0_bits_data <= _laneVec_2_readBusPort_0_deq_bits_data;
      end
      pipe_v_29 <= _laneVec_2_writeBusPort_0_enqRelease;
      if (shifterValid_29) begin
        shifterReg_29_0_valid <= _laneVec_1_writeBusPort_0_deq_valid;
        shifterReg_29_0_bits_data <= _laneVec_1_writeBusPort_0_deq_bits_data;
        shifterReg_29_0_bits_mask <= _laneVec_1_writeBusPort_0_deq_bits_mask;
        shifterReg_29_0_bits_instructionIndex <= _laneVec_1_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_29_0_bits_counter <= _laneVec_1_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_30 <= _laneVec_1_readBusPort_1_enqRelease;
      if (shifterValid_30) begin
        shifterReg_30_0_valid <= _laneVec_3_readBusPort_0_deq_valid;
        shifterReg_30_0_bits_data <= _laneVec_3_readBusPort_0_deq_bits_data;
      end
      pipe_v_31 <= _laneVec_3_writeBusPort_0_enqRelease;
      if (shifterValid_31) begin
        shifterReg_31_0_valid <= _laneVec_1_writeBusPort_1_deq_valid;
        shifterReg_31_0_bits_data <= _laneVec_1_writeBusPort_1_deq_bits_data;
        shifterReg_31_0_bits_mask <= _laneVec_1_writeBusPort_1_deq_bits_mask;
        shifterReg_31_0_bits_instructionIndex <= _laneVec_1_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_31_0_bits_counter <= _laneVec_1_writeBusPort_1_deq_bits_counter;
      end
      pipe_v_32 <= _laneVec_2_readBusPort_0_enqRelease;
      if (shifterValid_32) begin
        shifterReg_32_0_valid <= _laneVec_4_readBusPort_0_deq_valid;
        shifterReg_32_0_bits_data <= _laneVec_4_readBusPort_0_deq_bits_data;
      end
      pipe_v_33 <= _laneVec_4_writeBusPort_0_enqRelease;
      if (shifterValid_33) begin
        shifterReg_33_0_valid <= _laneVec_2_writeBusPort_0_deq_valid;
        shifterReg_33_0_bits_data <= _laneVec_2_writeBusPort_0_deq_bits_data;
        shifterReg_33_0_bits_mask <= _laneVec_2_writeBusPort_0_deq_bits_mask;
        shifterReg_33_0_bits_instructionIndex <= _laneVec_2_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_33_0_bits_counter <= _laneVec_2_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_34 <= _laneVec_2_readBusPort_1_enqRelease;
      if (shifterValid_34) begin
        shifterReg_34_0_valid <= _laneVec_5_readBusPort_0_deq_valid;
        shifterReg_34_0_bits_data <= _laneVec_5_readBusPort_0_deq_bits_data;
      end
      pipe_v_35 <= _laneVec_5_writeBusPort_0_enqRelease;
      if (shifterValid_35) begin
        shifterReg_35_0_valid <= _laneVec_2_writeBusPort_1_deq_valid;
        shifterReg_35_0_bits_data <= _laneVec_2_writeBusPort_1_deq_bits_data;
        shifterReg_35_0_bits_mask <= _laneVec_2_writeBusPort_1_deq_bits_mask;
        shifterReg_35_0_bits_instructionIndex <= _laneVec_2_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_35_0_bits_counter <= _laneVec_2_writeBusPort_1_deq_bits_counter;
      end
      pipe_v_36 <= _laneVec_3_readBusPort_0_enqRelease;
      if (shifterValid_36) begin
        shifterReg_36_0_valid <= _laneVec_6_readBusPort_0_deq_valid;
        shifterReg_36_0_bits_data <= _laneVec_6_readBusPort_0_deq_bits_data;
      end
      pipe_v_37 <= _laneVec_6_writeBusPort_0_enqRelease;
      if (shifterValid_37) begin
        shifterReg_37_0_valid <= _laneVec_3_writeBusPort_0_deq_valid;
        shifterReg_37_0_bits_data <= _laneVec_3_writeBusPort_0_deq_bits_data;
        shifterReg_37_0_bits_mask <= _laneVec_3_writeBusPort_0_deq_bits_mask;
        shifterReg_37_0_bits_instructionIndex <= _laneVec_3_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_37_0_bits_counter <= _laneVec_3_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_38 <= _laneVec_3_readBusPort_1_enqRelease;
      if (shifterValid_38) begin
        shifterReg_38_0_valid <= _laneVec_7_readBusPort_0_deq_valid;
        shifterReg_38_0_bits_data <= _laneVec_7_readBusPort_0_deq_bits_data;
      end
      pipe_v_39 <= _laneVec_7_writeBusPort_0_enqRelease;
      if (shifterValid_39) begin
        shifterReg_39_0_valid <= _laneVec_3_writeBusPort_1_deq_valid;
        shifterReg_39_0_bits_data <= _laneVec_3_writeBusPort_1_deq_bits_data;
        shifterReg_39_0_bits_mask <= _laneVec_3_writeBusPort_1_deq_bits_mask;
        shifterReg_39_0_bits_instructionIndex <= _laneVec_3_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_39_0_bits_counter <= _laneVec_3_writeBusPort_1_deq_bits_counter;
      end
      pipe_v_40 <= _laneVec_4_readBusPort_0_enqRelease;
      if (shifterValid_40) begin
        shifterReg_40_0_valid <= _laneVec_0_readBusPort_1_deq_valid;
        shifterReg_40_0_bits_data <= _laneVec_0_readBusPort_1_deq_bits_data;
      end
      pipe_v_41 <= _laneVec_0_writeBusPort_1_enqRelease;
      if (shifterValid_41) begin
        shifterReg_41_0_valid <= _laneVec_4_writeBusPort_0_deq_valid;
        shifterReg_41_0_bits_data <= _laneVec_4_writeBusPort_0_deq_bits_data;
        shifterReg_41_0_bits_mask <= _laneVec_4_writeBusPort_0_deq_bits_mask;
        shifterReg_41_0_bits_instructionIndex <= _laneVec_4_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_41_0_bits_counter <= _laneVec_4_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_42 <= _laneVec_4_readBusPort_1_enqRelease;
      if (shifterValid_42) begin
        shifterReg_42_0_valid <= _laneVec_1_readBusPort_1_deq_valid;
        shifterReg_42_0_bits_data <= _laneVec_1_readBusPort_1_deq_bits_data;
      end
      pipe_v_43 <= _laneVec_1_writeBusPort_1_enqRelease;
      if (shifterValid_43) begin
        shifterReg_43_0_valid <= _laneVec_4_writeBusPort_1_deq_valid;
        shifterReg_43_0_bits_data <= _laneVec_4_writeBusPort_1_deq_bits_data;
        shifterReg_43_0_bits_mask <= _laneVec_4_writeBusPort_1_deq_bits_mask;
        shifterReg_43_0_bits_instructionIndex <= _laneVec_4_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_43_0_bits_counter <= _laneVec_4_writeBusPort_1_deq_bits_counter;
      end
      pipe_v_44 <= _laneVec_5_readBusPort_0_enqRelease;
      if (shifterValid_44) begin
        shifterReg_44_0_valid <= _laneVec_2_readBusPort_1_deq_valid;
        shifterReg_44_0_bits_data <= _laneVec_2_readBusPort_1_deq_bits_data;
      end
      pipe_v_45 <= _laneVec_2_writeBusPort_1_enqRelease;
      if (shifterValid_45) begin
        shifterReg_45_0_valid <= _laneVec_5_writeBusPort_0_deq_valid;
        shifterReg_45_0_bits_data <= _laneVec_5_writeBusPort_0_deq_bits_data;
        shifterReg_45_0_bits_mask <= _laneVec_5_writeBusPort_0_deq_bits_mask;
        shifterReg_45_0_bits_instructionIndex <= _laneVec_5_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_45_0_bits_counter <= _laneVec_5_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_46 <= _laneVec_5_readBusPort_1_enqRelease;
      if (shifterValid_46) begin
        shifterReg_46_0_valid <= _laneVec_3_readBusPort_1_deq_valid;
        shifterReg_46_0_bits_data <= _laneVec_3_readBusPort_1_deq_bits_data;
      end
      pipe_v_47 <= _laneVec_3_writeBusPort_1_enqRelease;
      if (shifterValid_47) begin
        shifterReg_47_0_valid <= _laneVec_5_writeBusPort_1_deq_valid;
        shifterReg_47_0_bits_data <= _laneVec_5_writeBusPort_1_deq_bits_data;
        shifterReg_47_0_bits_mask <= _laneVec_5_writeBusPort_1_deq_bits_mask;
        shifterReg_47_0_bits_instructionIndex <= _laneVec_5_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_47_0_bits_counter <= _laneVec_5_writeBusPort_1_deq_bits_counter;
      end
      pipe_v_48 <= _laneVec_6_readBusPort_0_enqRelease;
      if (shifterValid_48) begin
        shifterReg_48_0_valid <= _laneVec_4_readBusPort_1_deq_valid;
        shifterReg_48_0_bits_data <= _laneVec_4_readBusPort_1_deq_bits_data;
      end
      pipe_v_49 <= _laneVec_4_writeBusPort_1_enqRelease;
      if (shifterValid_49) begin
        shifterReg_49_0_valid <= _laneVec_6_writeBusPort_0_deq_valid;
        shifterReg_49_0_bits_data <= _laneVec_6_writeBusPort_0_deq_bits_data;
        shifterReg_49_0_bits_mask <= _laneVec_6_writeBusPort_0_deq_bits_mask;
        shifterReg_49_0_bits_instructionIndex <= _laneVec_6_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_49_0_bits_counter <= _laneVec_6_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_50 <= _laneVec_6_readBusPort_1_enqRelease;
      if (shifterValid_50) begin
        shifterReg_50_0_valid <= _laneVec_5_readBusPort_1_deq_valid;
        shifterReg_50_0_bits_data <= _laneVec_5_readBusPort_1_deq_bits_data;
      end
      pipe_v_51 <= _laneVec_5_writeBusPort_1_enqRelease;
      if (shifterValid_51) begin
        shifterReg_51_0_valid <= _laneVec_6_writeBusPort_1_deq_valid;
        shifterReg_51_0_bits_data <= _laneVec_6_writeBusPort_1_deq_bits_data;
        shifterReg_51_0_bits_mask <= _laneVec_6_writeBusPort_1_deq_bits_mask;
        shifterReg_51_0_bits_instructionIndex <= _laneVec_6_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_51_0_bits_counter <= _laneVec_6_writeBusPort_1_deq_bits_counter;
      end
      pipe_v_52 <= _laneVec_7_readBusPort_0_enqRelease;
      if (shifterValid_52) begin
        shifterReg_52_0_valid <= _laneVec_6_readBusPort_1_deq_valid;
        shifterReg_52_0_bits_data <= _laneVec_6_readBusPort_1_deq_bits_data;
      end
      pipe_v_53 <= _laneVec_6_writeBusPort_1_enqRelease;
      if (shifterValid_53) begin
        shifterReg_53_0_valid <= _laneVec_7_writeBusPort_0_deq_valid;
        shifterReg_53_0_bits_data <= _laneVec_7_writeBusPort_0_deq_bits_data;
        shifterReg_53_0_bits_mask <= _laneVec_7_writeBusPort_0_deq_bits_mask;
        shifterReg_53_0_bits_instructionIndex <= _laneVec_7_writeBusPort_0_deq_bits_instructionIndex;
        shifterReg_53_0_bits_counter <= _laneVec_7_writeBusPort_0_deq_bits_counter;
      end
      pipe_v_54 <= _laneVec_7_readBusPort_1_enqRelease;
      if (shifterValid_54) begin
        shifterReg_54_0_valid <= _laneVec_7_readBusPort_1_deq_valid;
        shifterReg_54_0_bits_data <= _laneVec_7_readBusPort_1_deq_bits_data;
      end
      pipe_v_55 <= _laneVec_7_writeBusPort_1_enqRelease;
      if (shifterValid_55) begin
        shifterReg_55_0_valid <= _laneVec_7_writeBusPort_1_deq_valid;
        shifterReg_55_0_bits_data <= _laneVec_7_writeBusPort_1_deq_bits_data;
        shifterReg_55_0_bits_mask <= _laneVec_7_writeBusPort_1_deq_bits_mask;
        shifterReg_55_0_bits_instructionIndex <= _laneVec_7_writeBusPort_1_deq_bits_instructionIndex;
        shifterReg_55_0_bits_counter <= _laneVec_7_writeBusPort_1_deq_bits_counter;
      end
    end
    instructionFinishedPipe_pipe_b <= _laneVec_0_instructionFinished;
    pipe_b_1 <= _maskUnit_laneMaskInput_0;
    if (pipe_v_1)
      pipe_pipe_b <= pipe_b_1;
    view__laneMaskSelect_0_pipe_b <= _laneVec_0_maskSelect;
    if (view__laneMaskSelect_0_pipe_v)
      view__laneMaskSelect_0_pipe_pipe_b <= view__laneMaskSelect_0_pipe_b;
    view__laneMaskSewSelect_0_pipe_b <= _laneVec_0_maskSelectSew;
    if (view__laneMaskSewSelect_0_pipe_v)
      view__laneMaskSewSelect_0_pipe_pipe_b <= view__laneMaskSewSelect_0_pipe_b;
    lsuLastPipe_pipe_b <= _lsu_lastReport;
    maskLastPipe_pipe_b <= _maskUnit_lastReport;
    pipe_b_2 <= writeCounter;
    instructionFinishedPipe_pipe_b_1 <= _laneVec_1_instructionFinished;
    pipe_b_4 <= _maskUnit_laneMaskInput_1;
    if (pipe_v_4)
      pipe_pipe_b_1 <= pipe_b_4;
    view__laneMaskSelect_1_pipe_b <= _laneVec_1_maskSelect;
    if (view__laneMaskSelect_1_pipe_v)
      view__laneMaskSelect_1_pipe_pipe_b <= view__laneMaskSelect_1_pipe_b;
    view__laneMaskSewSelect_1_pipe_b <= _laneVec_1_maskSelectSew;
    if (view__laneMaskSewSelect_1_pipe_v)
      view__laneMaskSewSelect_1_pipe_pipe_b <= view__laneMaskSewSelect_1_pipe_b;
    lsuLastPipe_pipe_b_1 <= _lsu_lastReport;
    maskLastPipe_pipe_b_1 <= _maskUnit_lastReport;
    pipe_b_5 <= writeCounter_1;
    instructionFinishedPipe_pipe_b_2 <= _laneVec_2_instructionFinished;
    pipe_b_7 <= _maskUnit_laneMaskInput_2;
    if (pipe_v_7)
      pipe_pipe_b_2 <= pipe_b_7;
    view__laneMaskSelect_2_pipe_b <= _laneVec_2_maskSelect;
    if (view__laneMaskSelect_2_pipe_v)
      view__laneMaskSelect_2_pipe_pipe_b <= view__laneMaskSelect_2_pipe_b;
    view__laneMaskSewSelect_2_pipe_b <= _laneVec_2_maskSelectSew;
    if (view__laneMaskSewSelect_2_pipe_v)
      view__laneMaskSewSelect_2_pipe_pipe_b <= view__laneMaskSewSelect_2_pipe_b;
    lsuLastPipe_pipe_b_2 <= _lsu_lastReport;
    maskLastPipe_pipe_b_2 <= _maskUnit_lastReport;
    pipe_b_8 <= writeCounter_2;
    instructionFinishedPipe_pipe_b_3 <= _laneVec_3_instructionFinished;
    pipe_b_10 <= _maskUnit_laneMaskInput_3;
    if (pipe_v_10)
      pipe_pipe_b_3 <= pipe_b_10;
    view__laneMaskSelect_3_pipe_b <= _laneVec_3_maskSelect;
    if (view__laneMaskSelect_3_pipe_v)
      view__laneMaskSelect_3_pipe_pipe_b <= view__laneMaskSelect_3_pipe_b;
    view__laneMaskSewSelect_3_pipe_b <= _laneVec_3_maskSelectSew;
    if (view__laneMaskSewSelect_3_pipe_v)
      view__laneMaskSewSelect_3_pipe_pipe_b <= view__laneMaskSewSelect_3_pipe_b;
    lsuLastPipe_pipe_b_3 <= _lsu_lastReport;
    maskLastPipe_pipe_b_3 <= _maskUnit_lastReport;
    pipe_b_11 <= writeCounter_3;
    instructionFinishedPipe_pipe_b_4 <= _laneVec_4_instructionFinished;
    pipe_b_13 <= _maskUnit_laneMaskInput_4;
    if (pipe_v_13)
      pipe_pipe_b_4 <= pipe_b_13;
    view__laneMaskSelect_4_pipe_b <= _laneVec_4_maskSelect;
    if (view__laneMaskSelect_4_pipe_v)
      view__laneMaskSelect_4_pipe_pipe_b <= view__laneMaskSelect_4_pipe_b;
    view__laneMaskSewSelect_4_pipe_b <= _laneVec_4_maskSelectSew;
    if (view__laneMaskSewSelect_4_pipe_v)
      view__laneMaskSewSelect_4_pipe_pipe_b <= view__laneMaskSewSelect_4_pipe_b;
    lsuLastPipe_pipe_b_4 <= _lsu_lastReport;
    maskLastPipe_pipe_b_4 <= _maskUnit_lastReport;
    pipe_b_14 <= writeCounter_4;
    instructionFinishedPipe_pipe_b_5 <= _laneVec_5_instructionFinished;
    pipe_b_16 <= _maskUnit_laneMaskInput_5;
    if (pipe_v_16)
      pipe_pipe_b_5 <= pipe_b_16;
    view__laneMaskSelect_5_pipe_b <= _laneVec_5_maskSelect;
    if (view__laneMaskSelect_5_pipe_v)
      view__laneMaskSelect_5_pipe_pipe_b <= view__laneMaskSelect_5_pipe_b;
    view__laneMaskSewSelect_5_pipe_b <= _laneVec_5_maskSelectSew;
    if (view__laneMaskSewSelect_5_pipe_v)
      view__laneMaskSewSelect_5_pipe_pipe_b <= view__laneMaskSewSelect_5_pipe_b;
    lsuLastPipe_pipe_b_5 <= _lsu_lastReport;
    maskLastPipe_pipe_b_5 <= _maskUnit_lastReport;
    pipe_b_17 <= writeCounter_5;
    instructionFinishedPipe_pipe_b_6 <= _laneVec_6_instructionFinished;
    pipe_b_19 <= _maskUnit_laneMaskInput_6;
    if (pipe_v_19)
      pipe_pipe_b_6 <= pipe_b_19;
    view__laneMaskSelect_6_pipe_b <= _laneVec_6_maskSelect;
    if (view__laneMaskSelect_6_pipe_v)
      view__laneMaskSelect_6_pipe_pipe_b <= view__laneMaskSelect_6_pipe_b;
    view__laneMaskSewSelect_6_pipe_b <= _laneVec_6_maskSelectSew;
    if (view__laneMaskSewSelect_6_pipe_v)
      view__laneMaskSewSelect_6_pipe_pipe_b <= view__laneMaskSewSelect_6_pipe_b;
    lsuLastPipe_pipe_b_6 <= _lsu_lastReport;
    maskLastPipe_pipe_b_6 <= _maskUnit_lastReport;
    pipe_b_20 <= writeCounter_6;
    instructionFinishedPipe_pipe_b_7 <= _laneVec_7_instructionFinished;
    pipe_b_22 <= _maskUnit_laneMaskInput_7;
    if (pipe_v_22)
      pipe_pipe_b_7 <= pipe_b_22;
    view__laneMaskSelect_7_pipe_b <= _laneVec_7_maskSelect;
    if (view__laneMaskSelect_7_pipe_v)
      view__laneMaskSelect_7_pipe_pipe_b <= view__laneMaskSelect_7_pipe_b;
    view__laneMaskSewSelect_7_pipe_b <= _laneVec_7_maskSelectSew;
    if (view__laneMaskSewSelect_7_pipe_v)
      view__laneMaskSewSelect_7_pipe_pipe_b <= view__laneMaskSewSelect_7_pipe_b;
    lsuLastPipe_pipe_b_7 <= _lsu_lastReport;
    maskLastPipe_pipe_b_7 <= _maskUnit_lastReport;
    pipe_b_23 <= writeCounter_7;
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:174];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [7:0] i = 8'h0; i < 8'hAF; i += 8'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        instructionCounter = _RANDOM[8'h0][2:0];
        responseCounter = _RANDOM[8'h0][5:3];
        requestReg_valid = _RANDOM[8'h0][6];
        requestReg_bits_issue_instruction = {_RANDOM[8'h0][31:7], _RANDOM[8'h1][6:0]};
        requestReg_bits_issue_rs1Data = {_RANDOM[8'h1][31:7], _RANDOM[8'h2][6:0]};
        requestReg_bits_issue_rs2Data = {_RANDOM[8'h2][31:7], _RANDOM[8'h3][6:0]};
        requestReg_bits_issue_vtype = {_RANDOM[8'h3][31:7], _RANDOM[8'h4][6:0]};
        requestReg_bits_issue_vl = {_RANDOM[8'h4][31:7], _RANDOM[8'h5][6:0]};
        requestReg_bits_issue_vstart = {_RANDOM[8'h5][31:7], _RANDOM[8'h6][6:0]};
        requestReg_bits_issue_vcsr = {_RANDOM[8'h6][31:7], _RANDOM[8'h7][6:0]};
        requestReg_bits_decodeResult_specialSlot = _RANDOM[8'h7][7];
        requestReg_bits_decodeResult_topUop = _RANDOM[8'h7][12:8];
        requestReg_bits_decodeResult_popCount = _RANDOM[8'h7][13];
        requestReg_bits_decodeResult_ffo = _RANDOM[8'h7][14];
        requestReg_bits_decodeResult_average = _RANDOM[8'h7][15];
        requestReg_bits_decodeResult_reverse = _RANDOM[8'h7][16];
        requestReg_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[8'h7][17];
        requestReg_bits_decodeResult_scheduler = _RANDOM[8'h7][18];
        requestReg_bits_decodeResult_sReadVD = _RANDOM[8'h7][19];
        requestReg_bits_decodeResult_vtype = _RANDOM[8'h7][20];
        requestReg_bits_decodeResult_sWrite = _RANDOM[8'h7][21];
        requestReg_bits_decodeResult_crossRead = _RANDOM[8'h7][22];
        requestReg_bits_decodeResult_crossWrite = _RANDOM[8'h7][23];
        requestReg_bits_decodeResult_maskUnit = _RANDOM[8'h7][24];
        requestReg_bits_decodeResult_special = _RANDOM[8'h7][25];
        requestReg_bits_decodeResult_saturate = _RANDOM[8'h7][26];
        requestReg_bits_decodeResult_vwmacc = _RANDOM[8'h7][27];
        requestReg_bits_decodeResult_readOnly = _RANDOM[8'h7][28];
        requestReg_bits_decodeResult_maskSource = _RANDOM[8'h7][29];
        requestReg_bits_decodeResult_maskDestination = _RANDOM[8'h7][30];
        requestReg_bits_decodeResult_maskLogic = _RANDOM[8'h7][31];
        requestReg_bits_decodeResult_uop = _RANDOM[8'h8][3:0];
        requestReg_bits_decodeResult_iota = _RANDOM[8'h8][4];
        requestReg_bits_decodeResult_mv = _RANDOM[8'h8][5];
        requestReg_bits_decodeResult_extend = _RANDOM[8'h8][6];
        requestReg_bits_decodeResult_unOrderWrite = _RANDOM[8'h8][7];
        requestReg_bits_decodeResult_compress = _RANDOM[8'h8][8];
        requestReg_bits_decodeResult_gather16 = _RANDOM[8'h8][9];
        requestReg_bits_decodeResult_gather = _RANDOM[8'h8][10];
        requestReg_bits_decodeResult_slid = _RANDOM[8'h8][11];
        requestReg_bits_decodeResult_targetRd = _RANDOM[8'h8][12];
        requestReg_bits_decodeResult_widenReduce = _RANDOM[8'h8][13];
        requestReg_bits_decodeResult_red = _RANDOM[8'h8][14];
        requestReg_bits_decodeResult_nr = _RANDOM[8'h8][15];
        requestReg_bits_decodeResult_itype = _RANDOM[8'h8][16];
        requestReg_bits_decodeResult_unsigned1 = _RANDOM[8'h8][17];
        requestReg_bits_decodeResult_unsigned0 = _RANDOM[8'h8][18];
        requestReg_bits_decodeResult_other = _RANDOM[8'h8][19];
        requestReg_bits_decodeResult_multiCycle = _RANDOM[8'h8][20];
        requestReg_bits_decodeResult_divider = _RANDOM[8'h8][21];
        requestReg_bits_decodeResult_multiplier = _RANDOM[8'h8][22];
        requestReg_bits_decodeResult_shift = _RANDOM[8'h8][23];
        requestReg_bits_decodeResult_adder = _RANDOM[8'h8][24];
        requestReg_bits_decodeResult_logic = _RANDOM[8'h8][25];
        requestReg_bits_instructionIndex = _RANDOM[8'h8][28:26];
        requestReg_bits_vdIsV0 = _RANDOM[8'h8][29];
        requestReg_bits_writeByte = {_RANDOM[8'h8][31:30], _RANDOM[8'h9][9:0]};
        slots_0_record_instructionIndex = _RANDOM[8'hA][13:11];
        slots_0_record_isLoadStore = _RANDOM[8'hA][14];
        slots_0_record_maskType = _RANDOM[8'hA][15];
        slots_0_state_wLast = _RANDOM[8'hA][16];
        slots_0_state_idle = _RANDOM[8'hA][17];
        slots_0_state_wMaskUnitLast = _RANDOM[8'hA][18];
        slots_0_state_wVRFWrite = _RANDOM[8'hA][19];
        slots_0_state_sCommit = _RANDOM[8'hA][20];
        slots_0_endTag_0 = _RANDOM[8'hA][21];
        slots_0_endTag_1 = _RANDOM[8'hA][22];
        slots_0_endTag_2 = _RANDOM[8'hA][23];
        slots_0_endTag_3 = _RANDOM[8'hA][24];
        slots_0_endTag_4 = _RANDOM[8'hA][25];
        slots_0_endTag_5 = _RANDOM[8'hA][26];
        slots_0_endTag_6 = _RANDOM[8'hA][27];
        slots_0_endTag_7 = _RANDOM[8'hA][28];
        slots_0_endTag_8 = _RANDOM[8'hA][29];
        slots_0_vxsat = _RANDOM[8'hA][30];
        slots_1_record_instructionIndex = {_RANDOM[8'hA][31], _RANDOM[8'hB][1:0]};
        slots_1_record_isLoadStore = _RANDOM[8'hB][2];
        slots_1_record_maskType = _RANDOM[8'hB][3];
        slots_1_state_wLast = _RANDOM[8'hB][4];
        slots_1_state_idle = _RANDOM[8'hB][5];
        slots_1_state_wMaskUnitLast = _RANDOM[8'hB][6];
        slots_1_state_wVRFWrite = _RANDOM[8'hB][7];
        slots_1_state_sCommit = _RANDOM[8'hB][8];
        slots_1_endTag_0 = _RANDOM[8'hB][9];
        slots_1_endTag_1 = _RANDOM[8'hB][10];
        slots_1_endTag_2 = _RANDOM[8'hB][11];
        slots_1_endTag_3 = _RANDOM[8'hB][12];
        slots_1_endTag_4 = _RANDOM[8'hB][13];
        slots_1_endTag_5 = _RANDOM[8'hB][14];
        slots_1_endTag_6 = _RANDOM[8'hB][15];
        slots_1_endTag_7 = _RANDOM[8'hB][16];
        slots_1_endTag_8 = _RANDOM[8'hB][17];
        slots_1_vxsat = _RANDOM[8'hB][18];
        slots_2_record_instructionIndex = _RANDOM[8'hB][21:19];
        slots_2_record_isLoadStore = _RANDOM[8'hB][22];
        slots_2_record_maskType = _RANDOM[8'hB][23];
        slots_2_state_wLast = _RANDOM[8'hB][24];
        slots_2_state_idle = _RANDOM[8'hB][25];
        slots_2_state_wMaskUnitLast = _RANDOM[8'hB][26];
        slots_2_state_wVRFWrite = _RANDOM[8'hB][27];
        slots_2_state_sCommit = _RANDOM[8'hB][28];
        slots_2_endTag_0 = _RANDOM[8'hB][29];
        slots_2_endTag_1 = _RANDOM[8'hB][30];
        slots_2_endTag_2 = _RANDOM[8'hB][31];
        slots_2_endTag_3 = _RANDOM[8'hC][0];
        slots_2_endTag_4 = _RANDOM[8'hC][1];
        slots_2_endTag_5 = _RANDOM[8'hC][2];
        slots_2_endTag_6 = _RANDOM[8'hC][3];
        slots_2_endTag_7 = _RANDOM[8'hC][4];
        slots_2_endTag_8 = _RANDOM[8'hC][5];
        slots_2_vxsat = _RANDOM[8'hC][6];
        slots_3_record_instructionIndex = _RANDOM[8'hC][9:7];
        slots_3_record_isLoadStore = _RANDOM[8'hC][10];
        slots_3_record_maskType = _RANDOM[8'hC][11];
        slots_3_state_wLast = _RANDOM[8'hC][12];
        slots_3_state_idle = _RANDOM[8'hC][13];
        slots_3_state_wMaskUnitLast = _RANDOM[8'hC][14];
        slots_3_state_wVRFWrite = _RANDOM[8'hC][15];
        slots_3_state_sCommit = _RANDOM[8'hC][16];
        slots_3_endTag_0 = _RANDOM[8'hC][17];
        slots_3_endTag_1 = _RANDOM[8'hC][18];
        slots_3_endTag_2 = _RANDOM[8'hC][19];
        slots_3_endTag_3 = _RANDOM[8'hC][20];
        slots_3_endTag_4 = _RANDOM[8'hC][21];
        slots_3_endTag_5 = _RANDOM[8'hC][22];
        slots_3_endTag_6 = _RANDOM[8'hC][23];
        slots_3_endTag_7 = _RANDOM[8'hC][24];
        slots_3_endTag_8 = _RANDOM[8'hC][25];
        slots_3_vxsat = _RANDOM[8'hC][26];
        slots_writeRD = _RANDOM[8'hC][27];
        slots_vd = {_RANDOM[8'hC][31:28], _RANDOM[8'hD][0]};
        releasePipe_pipe_v = _RANDOM[8'hD][1];
        tokenCheck_counter = _RANDOM[8'hD][4:2];
        shifterReg_0_valid = _RANDOM[8'hD][5];
        shifterReg_0_bits_instructionIndex = _RANDOM[8'hD][8:6];
        shifterReg_0_bits_decodeResult_specialSlot = _RANDOM[8'hD][9];
        shifterReg_0_bits_decodeResult_topUop = _RANDOM[8'hD][14:10];
        shifterReg_0_bits_decodeResult_popCount = _RANDOM[8'hD][15];
        shifterReg_0_bits_decodeResult_ffo = _RANDOM[8'hD][16];
        shifterReg_0_bits_decodeResult_average = _RANDOM[8'hD][17];
        shifterReg_0_bits_decodeResult_reverse = _RANDOM[8'hD][18];
        shifterReg_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[8'hD][19];
        shifterReg_0_bits_decodeResult_scheduler = _RANDOM[8'hD][20];
        shifterReg_0_bits_decodeResult_sReadVD = _RANDOM[8'hD][21];
        shifterReg_0_bits_decodeResult_vtype = _RANDOM[8'hD][22];
        shifterReg_0_bits_decodeResult_sWrite = _RANDOM[8'hD][23];
        shifterReg_0_bits_decodeResult_crossRead = _RANDOM[8'hD][24];
        shifterReg_0_bits_decodeResult_crossWrite = _RANDOM[8'hD][25];
        shifterReg_0_bits_decodeResult_maskUnit = _RANDOM[8'hD][26];
        shifterReg_0_bits_decodeResult_special = _RANDOM[8'hD][27];
        shifterReg_0_bits_decodeResult_saturate = _RANDOM[8'hD][28];
        shifterReg_0_bits_decodeResult_vwmacc = _RANDOM[8'hD][29];
        shifterReg_0_bits_decodeResult_readOnly = _RANDOM[8'hD][30];
        shifterReg_0_bits_decodeResult_maskSource = _RANDOM[8'hD][31];
        shifterReg_0_bits_decodeResult_maskDestination = _RANDOM[8'hE][0];
        shifterReg_0_bits_decodeResult_maskLogic = _RANDOM[8'hE][1];
        shifterReg_0_bits_decodeResult_uop = _RANDOM[8'hE][5:2];
        shifterReg_0_bits_decodeResult_iota = _RANDOM[8'hE][6];
        shifterReg_0_bits_decodeResult_mv = _RANDOM[8'hE][7];
        shifterReg_0_bits_decodeResult_extend = _RANDOM[8'hE][8];
        shifterReg_0_bits_decodeResult_unOrderWrite = _RANDOM[8'hE][9];
        shifterReg_0_bits_decodeResult_compress = _RANDOM[8'hE][10];
        shifterReg_0_bits_decodeResult_gather16 = _RANDOM[8'hE][11];
        shifterReg_0_bits_decodeResult_gather = _RANDOM[8'hE][12];
        shifterReg_0_bits_decodeResult_slid = _RANDOM[8'hE][13];
        shifterReg_0_bits_decodeResult_targetRd = _RANDOM[8'hE][14];
        shifterReg_0_bits_decodeResult_widenReduce = _RANDOM[8'hE][15];
        shifterReg_0_bits_decodeResult_red = _RANDOM[8'hE][16];
        shifterReg_0_bits_decodeResult_nr = _RANDOM[8'hE][17];
        shifterReg_0_bits_decodeResult_itype = _RANDOM[8'hE][18];
        shifterReg_0_bits_decodeResult_unsigned1 = _RANDOM[8'hE][19];
        shifterReg_0_bits_decodeResult_unsigned0 = _RANDOM[8'hE][20];
        shifterReg_0_bits_decodeResult_other = _RANDOM[8'hE][21];
        shifterReg_0_bits_decodeResult_multiCycle = _RANDOM[8'hE][22];
        shifterReg_0_bits_decodeResult_divider = _RANDOM[8'hE][23];
        shifterReg_0_bits_decodeResult_multiplier = _RANDOM[8'hE][24];
        shifterReg_0_bits_decodeResult_shift = _RANDOM[8'hE][25];
        shifterReg_0_bits_decodeResult_adder = _RANDOM[8'hE][26];
        shifterReg_0_bits_decodeResult_logic = _RANDOM[8'hE][27];
        shifterReg_0_bits_loadStore = _RANDOM[8'hE][28];
        shifterReg_0_bits_issueInst = _RANDOM[8'hE][29];
        shifterReg_0_bits_store = _RANDOM[8'hE][30];
        shifterReg_0_bits_special = _RANDOM[8'hE][31];
        shifterReg_0_bits_lsWholeReg = _RANDOM[8'hF][0];
        shifterReg_0_bits_vs1 = _RANDOM[8'hF][5:1];
        shifterReg_0_bits_vs2 = _RANDOM[8'hF][10:6];
        shifterReg_0_bits_vd = _RANDOM[8'hF][15:11];
        shifterReg_0_bits_loadStoreEEW = _RANDOM[8'hF][17:16];
        shifterReg_0_bits_mask = _RANDOM[8'hF][18];
        shifterReg_0_bits_segment = _RANDOM[8'hF][21:19];
        shifterReg_0_bits_readFromScalar = {_RANDOM[8'hF][31:22], _RANDOM[8'h10][21:0]};
        shifterReg_0_bits_csrInterface_vl = {_RANDOM[8'h10][31:22], _RANDOM[8'h11][1:0]};
        shifterReg_0_bits_csrInterface_vStart = _RANDOM[8'h11][13:2];
        shifterReg_0_bits_csrInterface_vlmul = _RANDOM[8'h11][16:14];
        shifterReg_0_bits_csrInterface_vSew = _RANDOM[8'h11][18:17];
        shifterReg_0_bits_csrInterface_vxrm = _RANDOM[8'h11][20:19];
        shifterReg_0_bits_csrInterface_vta = _RANDOM[8'h11][21];
        shifterReg_0_bits_csrInterface_vma = _RANDOM[8'h11][22];
        releasePipe_pipe_v_1 = _RANDOM[8'h11][23];
        tokenCheck_counter_1 = _RANDOM[8'h11][26:24];
        shifterReg_1_0_valid = _RANDOM[8'h11][27];
        shifterReg_1_0_bits_instructionIndex = _RANDOM[8'h11][30:28];
        shifterReg_1_0_bits_decodeResult_specialSlot = _RANDOM[8'h11][31];
        shifterReg_1_0_bits_decodeResult_topUop = _RANDOM[8'h12][4:0];
        shifterReg_1_0_bits_decodeResult_popCount = _RANDOM[8'h12][5];
        shifterReg_1_0_bits_decodeResult_ffo = _RANDOM[8'h12][6];
        shifterReg_1_0_bits_decodeResult_average = _RANDOM[8'h12][7];
        shifterReg_1_0_bits_decodeResult_reverse = _RANDOM[8'h12][8];
        shifterReg_1_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[8'h12][9];
        shifterReg_1_0_bits_decodeResult_scheduler = _RANDOM[8'h12][10];
        shifterReg_1_0_bits_decodeResult_sReadVD = _RANDOM[8'h12][11];
        shifterReg_1_0_bits_decodeResult_vtype = _RANDOM[8'h12][12];
        shifterReg_1_0_bits_decodeResult_sWrite = _RANDOM[8'h12][13];
        shifterReg_1_0_bits_decodeResult_crossRead = _RANDOM[8'h12][14];
        shifterReg_1_0_bits_decodeResult_crossWrite = _RANDOM[8'h12][15];
        shifterReg_1_0_bits_decodeResult_maskUnit = _RANDOM[8'h12][16];
        shifterReg_1_0_bits_decodeResult_special = _RANDOM[8'h12][17];
        shifterReg_1_0_bits_decodeResult_saturate = _RANDOM[8'h12][18];
        shifterReg_1_0_bits_decodeResult_vwmacc = _RANDOM[8'h12][19];
        shifterReg_1_0_bits_decodeResult_readOnly = _RANDOM[8'h12][20];
        shifterReg_1_0_bits_decodeResult_maskSource = _RANDOM[8'h12][21];
        shifterReg_1_0_bits_decodeResult_maskDestination = _RANDOM[8'h12][22];
        shifterReg_1_0_bits_decodeResult_maskLogic = _RANDOM[8'h12][23];
        shifterReg_1_0_bits_decodeResult_uop = _RANDOM[8'h12][27:24];
        shifterReg_1_0_bits_decodeResult_iota = _RANDOM[8'h12][28];
        shifterReg_1_0_bits_decodeResult_mv = _RANDOM[8'h12][29];
        shifterReg_1_0_bits_decodeResult_extend = _RANDOM[8'h12][30];
        shifterReg_1_0_bits_decodeResult_unOrderWrite = _RANDOM[8'h12][31];
        shifterReg_1_0_bits_decodeResult_compress = _RANDOM[8'h13][0];
        shifterReg_1_0_bits_decodeResult_gather16 = _RANDOM[8'h13][1];
        shifterReg_1_0_bits_decodeResult_gather = _RANDOM[8'h13][2];
        shifterReg_1_0_bits_decodeResult_slid = _RANDOM[8'h13][3];
        shifterReg_1_0_bits_decodeResult_targetRd = _RANDOM[8'h13][4];
        shifterReg_1_0_bits_decodeResult_widenReduce = _RANDOM[8'h13][5];
        shifterReg_1_0_bits_decodeResult_red = _RANDOM[8'h13][6];
        shifterReg_1_0_bits_decodeResult_nr = _RANDOM[8'h13][7];
        shifterReg_1_0_bits_decodeResult_itype = _RANDOM[8'h13][8];
        shifterReg_1_0_bits_decodeResult_unsigned1 = _RANDOM[8'h13][9];
        shifterReg_1_0_bits_decodeResult_unsigned0 = _RANDOM[8'h13][10];
        shifterReg_1_0_bits_decodeResult_other = _RANDOM[8'h13][11];
        shifterReg_1_0_bits_decodeResult_multiCycle = _RANDOM[8'h13][12];
        shifterReg_1_0_bits_decodeResult_divider = _RANDOM[8'h13][13];
        shifterReg_1_0_bits_decodeResult_multiplier = _RANDOM[8'h13][14];
        shifterReg_1_0_bits_decodeResult_shift = _RANDOM[8'h13][15];
        shifterReg_1_0_bits_decodeResult_adder = _RANDOM[8'h13][16];
        shifterReg_1_0_bits_decodeResult_logic = _RANDOM[8'h13][17];
        shifterReg_1_0_bits_loadStore = _RANDOM[8'h13][18];
        shifterReg_1_0_bits_issueInst = _RANDOM[8'h13][19];
        shifterReg_1_0_bits_store = _RANDOM[8'h13][20];
        shifterReg_1_0_bits_special = _RANDOM[8'h13][21];
        shifterReg_1_0_bits_lsWholeReg = _RANDOM[8'h13][22];
        shifterReg_1_0_bits_vs1 = _RANDOM[8'h13][27:23];
        shifterReg_1_0_bits_vs2 = {_RANDOM[8'h13][31:28], _RANDOM[8'h14][0]};
        shifterReg_1_0_bits_vd = _RANDOM[8'h14][5:1];
        shifterReg_1_0_bits_loadStoreEEW = _RANDOM[8'h14][7:6];
        shifterReg_1_0_bits_mask = _RANDOM[8'h14][8];
        shifterReg_1_0_bits_segment = _RANDOM[8'h14][11:9];
        shifterReg_1_0_bits_readFromScalar = {_RANDOM[8'h14][31:12], _RANDOM[8'h15][11:0]};
        shifterReg_1_0_bits_csrInterface_vl = _RANDOM[8'h15][23:12];
        shifterReg_1_0_bits_csrInterface_vStart = {_RANDOM[8'h15][31:24], _RANDOM[8'h16][3:0]};
        shifterReg_1_0_bits_csrInterface_vlmul = _RANDOM[8'h16][6:4];
        shifterReg_1_0_bits_csrInterface_vSew = _RANDOM[8'h16][8:7];
        shifterReg_1_0_bits_csrInterface_vxrm = _RANDOM[8'h16][10:9];
        shifterReg_1_0_bits_csrInterface_vta = _RANDOM[8'h16][11];
        shifterReg_1_0_bits_csrInterface_vma = _RANDOM[8'h16][12];
        releasePipe_pipe_v_2 = _RANDOM[8'h16][13];
        tokenCheck_counter_2 = _RANDOM[8'h16][16:14];
        shifterReg_2_0_valid = _RANDOM[8'h16][17];
        shifterReg_2_0_bits_instructionIndex = _RANDOM[8'h16][20:18];
        shifterReg_2_0_bits_decodeResult_specialSlot = _RANDOM[8'h16][21];
        shifterReg_2_0_bits_decodeResult_topUop = _RANDOM[8'h16][26:22];
        shifterReg_2_0_bits_decodeResult_popCount = _RANDOM[8'h16][27];
        shifterReg_2_0_bits_decodeResult_ffo = _RANDOM[8'h16][28];
        shifterReg_2_0_bits_decodeResult_average = _RANDOM[8'h16][29];
        shifterReg_2_0_bits_decodeResult_reverse = _RANDOM[8'h16][30];
        shifterReg_2_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[8'h16][31];
        shifterReg_2_0_bits_decodeResult_scheduler = _RANDOM[8'h17][0];
        shifterReg_2_0_bits_decodeResult_sReadVD = _RANDOM[8'h17][1];
        shifterReg_2_0_bits_decodeResult_vtype = _RANDOM[8'h17][2];
        shifterReg_2_0_bits_decodeResult_sWrite = _RANDOM[8'h17][3];
        shifterReg_2_0_bits_decodeResult_crossRead = _RANDOM[8'h17][4];
        shifterReg_2_0_bits_decodeResult_crossWrite = _RANDOM[8'h17][5];
        shifterReg_2_0_bits_decodeResult_maskUnit = _RANDOM[8'h17][6];
        shifterReg_2_0_bits_decodeResult_special = _RANDOM[8'h17][7];
        shifterReg_2_0_bits_decodeResult_saturate = _RANDOM[8'h17][8];
        shifterReg_2_0_bits_decodeResult_vwmacc = _RANDOM[8'h17][9];
        shifterReg_2_0_bits_decodeResult_readOnly = _RANDOM[8'h17][10];
        shifterReg_2_0_bits_decodeResult_maskSource = _RANDOM[8'h17][11];
        shifterReg_2_0_bits_decodeResult_maskDestination = _RANDOM[8'h17][12];
        shifterReg_2_0_bits_decodeResult_maskLogic = _RANDOM[8'h17][13];
        shifterReg_2_0_bits_decodeResult_uop = _RANDOM[8'h17][17:14];
        shifterReg_2_0_bits_decodeResult_iota = _RANDOM[8'h17][18];
        shifterReg_2_0_bits_decodeResult_mv = _RANDOM[8'h17][19];
        shifterReg_2_0_bits_decodeResult_extend = _RANDOM[8'h17][20];
        shifterReg_2_0_bits_decodeResult_unOrderWrite = _RANDOM[8'h17][21];
        shifterReg_2_0_bits_decodeResult_compress = _RANDOM[8'h17][22];
        shifterReg_2_0_bits_decodeResult_gather16 = _RANDOM[8'h17][23];
        shifterReg_2_0_bits_decodeResult_gather = _RANDOM[8'h17][24];
        shifterReg_2_0_bits_decodeResult_slid = _RANDOM[8'h17][25];
        shifterReg_2_0_bits_decodeResult_targetRd = _RANDOM[8'h17][26];
        shifterReg_2_0_bits_decodeResult_widenReduce = _RANDOM[8'h17][27];
        shifterReg_2_0_bits_decodeResult_red = _RANDOM[8'h17][28];
        shifterReg_2_0_bits_decodeResult_nr = _RANDOM[8'h17][29];
        shifterReg_2_0_bits_decodeResult_itype = _RANDOM[8'h17][30];
        shifterReg_2_0_bits_decodeResult_unsigned1 = _RANDOM[8'h17][31];
        shifterReg_2_0_bits_decodeResult_unsigned0 = _RANDOM[8'h18][0];
        shifterReg_2_0_bits_decodeResult_other = _RANDOM[8'h18][1];
        shifterReg_2_0_bits_decodeResult_multiCycle = _RANDOM[8'h18][2];
        shifterReg_2_0_bits_decodeResult_divider = _RANDOM[8'h18][3];
        shifterReg_2_0_bits_decodeResult_multiplier = _RANDOM[8'h18][4];
        shifterReg_2_0_bits_decodeResult_shift = _RANDOM[8'h18][5];
        shifterReg_2_0_bits_decodeResult_adder = _RANDOM[8'h18][6];
        shifterReg_2_0_bits_decodeResult_logic = _RANDOM[8'h18][7];
        shifterReg_2_0_bits_loadStore = _RANDOM[8'h18][8];
        shifterReg_2_0_bits_issueInst = _RANDOM[8'h18][9];
        shifterReg_2_0_bits_store = _RANDOM[8'h18][10];
        shifterReg_2_0_bits_special = _RANDOM[8'h18][11];
        shifterReg_2_0_bits_lsWholeReg = _RANDOM[8'h18][12];
        shifterReg_2_0_bits_vs1 = _RANDOM[8'h18][17:13];
        shifterReg_2_0_bits_vs2 = _RANDOM[8'h18][22:18];
        shifterReg_2_0_bits_vd = _RANDOM[8'h18][27:23];
        shifterReg_2_0_bits_loadStoreEEW = _RANDOM[8'h18][29:28];
        shifterReg_2_0_bits_mask = _RANDOM[8'h18][30];
        shifterReg_2_0_bits_segment = {_RANDOM[8'h18][31], _RANDOM[8'h19][1:0]};
        shifterReg_2_0_bits_readFromScalar = {_RANDOM[8'h19][31:2], _RANDOM[8'h1A][1:0]};
        shifterReg_2_0_bits_csrInterface_vl = _RANDOM[8'h1A][13:2];
        shifterReg_2_0_bits_csrInterface_vStart = _RANDOM[8'h1A][25:14];
        shifterReg_2_0_bits_csrInterface_vlmul = _RANDOM[8'h1A][28:26];
        shifterReg_2_0_bits_csrInterface_vSew = _RANDOM[8'h1A][30:29];
        shifterReg_2_0_bits_csrInterface_vxrm = {_RANDOM[8'h1A][31], _RANDOM[8'h1B][0]};
        shifterReg_2_0_bits_csrInterface_vta = _RANDOM[8'h1B][1];
        shifterReg_2_0_bits_csrInterface_vma = _RANDOM[8'h1B][2];
        releasePipe_pipe_v_3 = _RANDOM[8'h1B][3];
        tokenCheck_counter_3 = _RANDOM[8'h1B][6:4];
        shifterReg_3_0_valid = _RANDOM[8'h1B][7];
        shifterReg_3_0_bits_instructionIndex = _RANDOM[8'h1B][10:8];
        shifterReg_3_0_bits_decodeResult_specialSlot = _RANDOM[8'h1B][11];
        shifterReg_3_0_bits_decodeResult_topUop = _RANDOM[8'h1B][16:12];
        shifterReg_3_0_bits_decodeResult_popCount = _RANDOM[8'h1B][17];
        shifterReg_3_0_bits_decodeResult_ffo = _RANDOM[8'h1B][18];
        shifterReg_3_0_bits_decodeResult_average = _RANDOM[8'h1B][19];
        shifterReg_3_0_bits_decodeResult_reverse = _RANDOM[8'h1B][20];
        shifterReg_3_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[8'h1B][21];
        shifterReg_3_0_bits_decodeResult_scheduler = _RANDOM[8'h1B][22];
        shifterReg_3_0_bits_decodeResult_sReadVD = _RANDOM[8'h1B][23];
        shifterReg_3_0_bits_decodeResult_vtype = _RANDOM[8'h1B][24];
        shifterReg_3_0_bits_decodeResult_sWrite = _RANDOM[8'h1B][25];
        shifterReg_3_0_bits_decodeResult_crossRead = _RANDOM[8'h1B][26];
        shifterReg_3_0_bits_decodeResult_crossWrite = _RANDOM[8'h1B][27];
        shifterReg_3_0_bits_decodeResult_maskUnit = _RANDOM[8'h1B][28];
        shifterReg_3_0_bits_decodeResult_special = _RANDOM[8'h1B][29];
        shifterReg_3_0_bits_decodeResult_saturate = _RANDOM[8'h1B][30];
        shifterReg_3_0_bits_decodeResult_vwmacc = _RANDOM[8'h1B][31];
        shifterReg_3_0_bits_decodeResult_readOnly = _RANDOM[8'h1C][0];
        shifterReg_3_0_bits_decodeResult_maskSource = _RANDOM[8'h1C][1];
        shifterReg_3_0_bits_decodeResult_maskDestination = _RANDOM[8'h1C][2];
        shifterReg_3_0_bits_decodeResult_maskLogic = _RANDOM[8'h1C][3];
        shifterReg_3_0_bits_decodeResult_uop = _RANDOM[8'h1C][7:4];
        shifterReg_3_0_bits_decodeResult_iota = _RANDOM[8'h1C][8];
        shifterReg_3_0_bits_decodeResult_mv = _RANDOM[8'h1C][9];
        shifterReg_3_0_bits_decodeResult_extend = _RANDOM[8'h1C][10];
        shifterReg_3_0_bits_decodeResult_unOrderWrite = _RANDOM[8'h1C][11];
        shifterReg_3_0_bits_decodeResult_compress = _RANDOM[8'h1C][12];
        shifterReg_3_0_bits_decodeResult_gather16 = _RANDOM[8'h1C][13];
        shifterReg_3_0_bits_decodeResult_gather = _RANDOM[8'h1C][14];
        shifterReg_3_0_bits_decodeResult_slid = _RANDOM[8'h1C][15];
        shifterReg_3_0_bits_decodeResult_targetRd = _RANDOM[8'h1C][16];
        shifterReg_3_0_bits_decodeResult_widenReduce = _RANDOM[8'h1C][17];
        shifterReg_3_0_bits_decodeResult_red = _RANDOM[8'h1C][18];
        shifterReg_3_0_bits_decodeResult_nr = _RANDOM[8'h1C][19];
        shifterReg_3_0_bits_decodeResult_itype = _RANDOM[8'h1C][20];
        shifterReg_3_0_bits_decodeResult_unsigned1 = _RANDOM[8'h1C][21];
        shifterReg_3_0_bits_decodeResult_unsigned0 = _RANDOM[8'h1C][22];
        shifterReg_3_0_bits_decodeResult_other = _RANDOM[8'h1C][23];
        shifterReg_3_0_bits_decodeResult_multiCycle = _RANDOM[8'h1C][24];
        shifterReg_3_0_bits_decodeResult_divider = _RANDOM[8'h1C][25];
        shifterReg_3_0_bits_decodeResult_multiplier = _RANDOM[8'h1C][26];
        shifterReg_3_0_bits_decodeResult_shift = _RANDOM[8'h1C][27];
        shifterReg_3_0_bits_decodeResult_adder = _RANDOM[8'h1C][28];
        shifterReg_3_0_bits_decodeResult_logic = _RANDOM[8'h1C][29];
        shifterReg_3_0_bits_loadStore = _RANDOM[8'h1C][30];
        shifterReg_3_0_bits_issueInst = _RANDOM[8'h1C][31];
        shifterReg_3_0_bits_store = _RANDOM[8'h1D][0];
        shifterReg_3_0_bits_special = _RANDOM[8'h1D][1];
        shifterReg_3_0_bits_lsWholeReg = _RANDOM[8'h1D][2];
        shifterReg_3_0_bits_vs1 = _RANDOM[8'h1D][7:3];
        shifterReg_3_0_bits_vs2 = _RANDOM[8'h1D][12:8];
        shifterReg_3_0_bits_vd = _RANDOM[8'h1D][17:13];
        shifterReg_3_0_bits_loadStoreEEW = _RANDOM[8'h1D][19:18];
        shifterReg_3_0_bits_mask = _RANDOM[8'h1D][20];
        shifterReg_3_0_bits_segment = _RANDOM[8'h1D][23:21];
        shifterReg_3_0_bits_readFromScalar = {_RANDOM[8'h1D][31:24], _RANDOM[8'h1E][23:0]};
        shifterReg_3_0_bits_csrInterface_vl = {_RANDOM[8'h1E][31:24], _RANDOM[8'h1F][3:0]};
        shifterReg_3_0_bits_csrInterface_vStart = _RANDOM[8'h1F][15:4];
        shifterReg_3_0_bits_csrInterface_vlmul = _RANDOM[8'h1F][18:16];
        shifterReg_3_0_bits_csrInterface_vSew = _RANDOM[8'h1F][20:19];
        shifterReg_3_0_bits_csrInterface_vxrm = _RANDOM[8'h1F][22:21];
        shifterReg_3_0_bits_csrInterface_vta = _RANDOM[8'h1F][23];
        shifterReg_3_0_bits_csrInterface_vma = _RANDOM[8'h1F][24];
        releasePipe_pipe_v_4 = _RANDOM[8'h1F][25];
        tokenCheck_counter_4 = _RANDOM[8'h1F][28:26];
        shifterReg_4_0_valid = _RANDOM[8'h1F][29];
        shifterReg_4_0_bits_instructionIndex = {_RANDOM[8'h1F][31:30], _RANDOM[8'h20][0]};
        shifterReg_4_0_bits_decodeResult_specialSlot = _RANDOM[8'h20][1];
        shifterReg_4_0_bits_decodeResult_topUop = _RANDOM[8'h20][6:2];
        shifterReg_4_0_bits_decodeResult_popCount = _RANDOM[8'h20][7];
        shifterReg_4_0_bits_decodeResult_ffo = _RANDOM[8'h20][8];
        shifterReg_4_0_bits_decodeResult_average = _RANDOM[8'h20][9];
        shifterReg_4_0_bits_decodeResult_reverse = _RANDOM[8'h20][10];
        shifterReg_4_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[8'h20][11];
        shifterReg_4_0_bits_decodeResult_scheduler = _RANDOM[8'h20][12];
        shifterReg_4_0_bits_decodeResult_sReadVD = _RANDOM[8'h20][13];
        shifterReg_4_0_bits_decodeResult_vtype = _RANDOM[8'h20][14];
        shifterReg_4_0_bits_decodeResult_sWrite = _RANDOM[8'h20][15];
        shifterReg_4_0_bits_decodeResult_crossRead = _RANDOM[8'h20][16];
        shifterReg_4_0_bits_decodeResult_crossWrite = _RANDOM[8'h20][17];
        shifterReg_4_0_bits_decodeResult_maskUnit = _RANDOM[8'h20][18];
        shifterReg_4_0_bits_decodeResult_special = _RANDOM[8'h20][19];
        shifterReg_4_0_bits_decodeResult_saturate = _RANDOM[8'h20][20];
        shifterReg_4_0_bits_decodeResult_vwmacc = _RANDOM[8'h20][21];
        shifterReg_4_0_bits_decodeResult_readOnly = _RANDOM[8'h20][22];
        shifterReg_4_0_bits_decodeResult_maskSource = _RANDOM[8'h20][23];
        shifterReg_4_0_bits_decodeResult_maskDestination = _RANDOM[8'h20][24];
        shifterReg_4_0_bits_decodeResult_maskLogic = _RANDOM[8'h20][25];
        shifterReg_4_0_bits_decodeResult_uop = _RANDOM[8'h20][29:26];
        shifterReg_4_0_bits_decodeResult_iota = _RANDOM[8'h20][30];
        shifterReg_4_0_bits_decodeResult_mv = _RANDOM[8'h20][31];
        shifterReg_4_0_bits_decodeResult_extend = _RANDOM[8'h21][0];
        shifterReg_4_0_bits_decodeResult_unOrderWrite = _RANDOM[8'h21][1];
        shifterReg_4_0_bits_decodeResult_compress = _RANDOM[8'h21][2];
        shifterReg_4_0_bits_decodeResult_gather16 = _RANDOM[8'h21][3];
        shifterReg_4_0_bits_decodeResult_gather = _RANDOM[8'h21][4];
        shifterReg_4_0_bits_decodeResult_slid = _RANDOM[8'h21][5];
        shifterReg_4_0_bits_decodeResult_targetRd = _RANDOM[8'h21][6];
        shifterReg_4_0_bits_decodeResult_widenReduce = _RANDOM[8'h21][7];
        shifterReg_4_0_bits_decodeResult_red = _RANDOM[8'h21][8];
        shifterReg_4_0_bits_decodeResult_nr = _RANDOM[8'h21][9];
        shifterReg_4_0_bits_decodeResult_itype = _RANDOM[8'h21][10];
        shifterReg_4_0_bits_decodeResult_unsigned1 = _RANDOM[8'h21][11];
        shifterReg_4_0_bits_decodeResult_unsigned0 = _RANDOM[8'h21][12];
        shifterReg_4_0_bits_decodeResult_other = _RANDOM[8'h21][13];
        shifterReg_4_0_bits_decodeResult_multiCycle = _RANDOM[8'h21][14];
        shifterReg_4_0_bits_decodeResult_divider = _RANDOM[8'h21][15];
        shifterReg_4_0_bits_decodeResult_multiplier = _RANDOM[8'h21][16];
        shifterReg_4_0_bits_decodeResult_shift = _RANDOM[8'h21][17];
        shifterReg_4_0_bits_decodeResult_adder = _RANDOM[8'h21][18];
        shifterReg_4_0_bits_decodeResult_logic = _RANDOM[8'h21][19];
        shifterReg_4_0_bits_loadStore = _RANDOM[8'h21][20];
        shifterReg_4_0_bits_issueInst = _RANDOM[8'h21][21];
        shifterReg_4_0_bits_store = _RANDOM[8'h21][22];
        shifterReg_4_0_bits_special = _RANDOM[8'h21][23];
        shifterReg_4_0_bits_lsWholeReg = _RANDOM[8'h21][24];
        shifterReg_4_0_bits_vs1 = _RANDOM[8'h21][29:25];
        shifterReg_4_0_bits_vs2 = {_RANDOM[8'h21][31:30], _RANDOM[8'h22][2:0]};
        shifterReg_4_0_bits_vd = _RANDOM[8'h22][7:3];
        shifterReg_4_0_bits_loadStoreEEW = _RANDOM[8'h22][9:8];
        shifterReg_4_0_bits_mask = _RANDOM[8'h22][10];
        shifterReg_4_0_bits_segment = _RANDOM[8'h22][13:11];
        shifterReg_4_0_bits_readFromScalar = {_RANDOM[8'h22][31:14], _RANDOM[8'h23][13:0]};
        shifterReg_4_0_bits_csrInterface_vl = _RANDOM[8'h23][25:14];
        shifterReg_4_0_bits_csrInterface_vStart = {_RANDOM[8'h23][31:26], _RANDOM[8'h24][5:0]};
        shifterReg_4_0_bits_csrInterface_vlmul = _RANDOM[8'h24][8:6];
        shifterReg_4_0_bits_csrInterface_vSew = _RANDOM[8'h24][10:9];
        shifterReg_4_0_bits_csrInterface_vxrm = _RANDOM[8'h24][12:11];
        shifterReg_4_0_bits_csrInterface_vta = _RANDOM[8'h24][13];
        shifterReg_4_0_bits_csrInterface_vma = _RANDOM[8'h24][14];
        releasePipe_pipe_v_5 = _RANDOM[8'h24][15];
        tokenCheck_counter_5 = _RANDOM[8'h24][18:16];
        shifterReg_5_0_valid = _RANDOM[8'h24][19];
        shifterReg_5_0_bits_instructionIndex = _RANDOM[8'h24][22:20];
        shifterReg_5_0_bits_decodeResult_specialSlot = _RANDOM[8'h24][23];
        shifterReg_5_0_bits_decodeResult_topUop = _RANDOM[8'h24][28:24];
        shifterReg_5_0_bits_decodeResult_popCount = _RANDOM[8'h24][29];
        shifterReg_5_0_bits_decodeResult_ffo = _RANDOM[8'h24][30];
        shifterReg_5_0_bits_decodeResult_average = _RANDOM[8'h24][31];
        shifterReg_5_0_bits_decodeResult_reverse = _RANDOM[8'h25][0];
        shifterReg_5_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[8'h25][1];
        shifterReg_5_0_bits_decodeResult_scheduler = _RANDOM[8'h25][2];
        shifterReg_5_0_bits_decodeResult_sReadVD = _RANDOM[8'h25][3];
        shifterReg_5_0_bits_decodeResult_vtype = _RANDOM[8'h25][4];
        shifterReg_5_0_bits_decodeResult_sWrite = _RANDOM[8'h25][5];
        shifterReg_5_0_bits_decodeResult_crossRead = _RANDOM[8'h25][6];
        shifterReg_5_0_bits_decodeResult_crossWrite = _RANDOM[8'h25][7];
        shifterReg_5_0_bits_decodeResult_maskUnit = _RANDOM[8'h25][8];
        shifterReg_5_0_bits_decodeResult_special = _RANDOM[8'h25][9];
        shifterReg_5_0_bits_decodeResult_saturate = _RANDOM[8'h25][10];
        shifterReg_5_0_bits_decodeResult_vwmacc = _RANDOM[8'h25][11];
        shifterReg_5_0_bits_decodeResult_readOnly = _RANDOM[8'h25][12];
        shifterReg_5_0_bits_decodeResult_maskSource = _RANDOM[8'h25][13];
        shifterReg_5_0_bits_decodeResult_maskDestination = _RANDOM[8'h25][14];
        shifterReg_5_0_bits_decodeResult_maskLogic = _RANDOM[8'h25][15];
        shifterReg_5_0_bits_decodeResult_uop = _RANDOM[8'h25][19:16];
        shifterReg_5_0_bits_decodeResult_iota = _RANDOM[8'h25][20];
        shifterReg_5_0_bits_decodeResult_mv = _RANDOM[8'h25][21];
        shifterReg_5_0_bits_decodeResult_extend = _RANDOM[8'h25][22];
        shifterReg_5_0_bits_decodeResult_unOrderWrite = _RANDOM[8'h25][23];
        shifterReg_5_0_bits_decodeResult_compress = _RANDOM[8'h25][24];
        shifterReg_5_0_bits_decodeResult_gather16 = _RANDOM[8'h25][25];
        shifterReg_5_0_bits_decodeResult_gather = _RANDOM[8'h25][26];
        shifterReg_5_0_bits_decodeResult_slid = _RANDOM[8'h25][27];
        shifterReg_5_0_bits_decodeResult_targetRd = _RANDOM[8'h25][28];
        shifterReg_5_0_bits_decodeResult_widenReduce = _RANDOM[8'h25][29];
        shifterReg_5_0_bits_decodeResult_red = _RANDOM[8'h25][30];
        shifterReg_5_0_bits_decodeResult_nr = _RANDOM[8'h25][31];
        shifterReg_5_0_bits_decodeResult_itype = _RANDOM[8'h26][0];
        shifterReg_5_0_bits_decodeResult_unsigned1 = _RANDOM[8'h26][1];
        shifterReg_5_0_bits_decodeResult_unsigned0 = _RANDOM[8'h26][2];
        shifterReg_5_0_bits_decodeResult_other = _RANDOM[8'h26][3];
        shifterReg_5_0_bits_decodeResult_multiCycle = _RANDOM[8'h26][4];
        shifterReg_5_0_bits_decodeResult_divider = _RANDOM[8'h26][5];
        shifterReg_5_0_bits_decodeResult_multiplier = _RANDOM[8'h26][6];
        shifterReg_5_0_bits_decodeResult_shift = _RANDOM[8'h26][7];
        shifterReg_5_0_bits_decodeResult_adder = _RANDOM[8'h26][8];
        shifterReg_5_0_bits_decodeResult_logic = _RANDOM[8'h26][9];
        shifterReg_5_0_bits_loadStore = _RANDOM[8'h26][10];
        shifterReg_5_0_bits_issueInst = _RANDOM[8'h26][11];
        shifterReg_5_0_bits_store = _RANDOM[8'h26][12];
        shifterReg_5_0_bits_special = _RANDOM[8'h26][13];
        shifterReg_5_0_bits_lsWholeReg = _RANDOM[8'h26][14];
        shifterReg_5_0_bits_vs1 = _RANDOM[8'h26][19:15];
        shifterReg_5_0_bits_vs2 = _RANDOM[8'h26][24:20];
        shifterReg_5_0_bits_vd = _RANDOM[8'h26][29:25];
        shifterReg_5_0_bits_loadStoreEEW = _RANDOM[8'h26][31:30];
        shifterReg_5_0_bits_mask = _RANDOM[8'h27][0];
        shifterReg_5_0_bits_segment = _RANDOM[8'h27][3:1];
        shifterReg_5_0_bits_readFromScalar = {_RANDOM[8'h27][31:4], _RANDOM[8'h28][3:0]};
        shifterReg_5_0_bits_csrInterface_vl = _RANDOM[8'h28][15:4];
        shifterReg_5_0_bits_csrInterface_vStart = _RANDOM[8'h28][27:16];
        shifterReg_5_0_bits_csrInterface_vlmul = _RANDOM[8'h28][30:28];
        shifterReg_5_0_bits_csrInterface_vSew = {_RANDOM[8'h28][31], _RANDOM[8'h29][0]};
        shifterReg_5_0_bits_csrInterface_vxrm = _RANDOM[8'h29][2:1];
        shifterReg_5_0_bits_csrInterface_vta = _RANDOM[8'h29][3];
        shifterReg_5_0_bits_csrInterface_vma = _RANDOM[8'h29][4];
        releasePipe_pipe_v_6 = _RANDOM[8'h29][5];
        tokenCheck_counter_6 = _RANDOM[8'h29][8:6];
        shifterReg_6_0_valid = _RANDOM[8'h29][9];
        shifterReg_6_0_bits_instructionIndex = _RANDOM[8'h29][12:10];
        shifterReg_6_0_bits_decodeResult_specialSlot = _RANDOM[8'h29][13];
        shifterReg_6_0_bits_decodeResult_topUop = _RANDOM[8'h29][18:14];
        shifterReg_6_0_bits_decodeResult_popCount = _RANDOM[8'h29][19];
        shifterReg_6_0_bits_decodeResult_ffo = _RANDOM[8'h29][20];
        shifterReg_6_0_bits_decodeResult_average = _RANDOM[8'h29][21];
        shifterReg_6_0_bits_decodeResult_reverse = _RANDOM[8'h29][22];
        shifterReg_6_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[8'h29][23];
        shifterReg_6_0_bits_decodeResult_scheduler = _RANDOM[8'h29][24];
        shifterReg_6_0_bits_decodeResult_sReadVD = _RANDOM[8'h29][25];
        shifterReg_6_0_bits_decodeResult_vtype = _RANDOM[8'h29][26];
        shifterReg_6_0_bits_decodeResult_sWrite = _RANDOM[8'h29][27];
        shifterReg_6_0_bits_decodeResult_crossRead = _RANDOM[8'h29][28];
        shifterReg_6_0_bits_decodeResult_crossWrite = _RANDOM[8'h29][29];
        shifterReg_6_0_bits_decodeResult_maskUnit = _RANDOM[8'h29][30];
        shifterReg_6_0_bits_decodeResult_special = _RANDOM[8'h29][31];
        shifterReg_6_0_bits_decodeResult_saturate = _RANDOM[8'h2A][0];
        shifterReg_6_0_bits_decodeResult_vwmacc = _RANDOM[8'h2A][1];
        shifterReg_6_0_bits_decodeResult_readOnly = _RANDOM[8'h2A][2];
        shifterReg_6_0_bits_decodeResult_maskSource = _RANDOM[8'h2A][3];
        shifterReg_6_0_bits_decodeResult_maskDestination = _RANDOM[8'h2A][4];
        shifterReg_6_0_bits_decodeResult_maskLogic = _RANDOM[8'h2A][5];
        shifterReg_6_0_bits_decodeResult_uop = _RANDOM[8'h2A][9:6];
        shifterReg_6_0_bits_decodeResult_iota = _RANDOM[8'h2A][10];
        shifterReg_6_0_bits_decodeResult_mv = _RANDOM[8'h2A][11];
        shifterReg_6_0_bits_decodeResult_extend = _RANDOM[8'h2A][12];
        shifterReg_6_0_bits_decodeResult_unOrderWrite = _RANDOM[8'h2A][13];
        shifterReg_6_0_bits_decodeResult_compress = _RANDOM[8'h2A][14];
        shifterReg_6_0_bits_decodeResult_gather16 = _RANDOM[8'h2A][15];
        shifterReg_6_0_bits_decodeResult_gather = _RANDOM[8'h2A][16];
        shifterReg_6_0_bits_decodeResult_slid = _RANDOM[8'h2A][17];
        shifterReg_6_0_bits_decodeResult_targetRd = _RANDOM[8'h2A][18];
        shifterReg_6_0_bits_decodeResult_widenReduce = _RANDOM[8'h2A][19];
        shifterReg_6_0_bits_decodeResult_red = _RANDOM[8'h2A][20];
        shifterReg_6_0_bits_decodeResult_nr = _RANDOM[8'h2A][21];
        shifterReg_6_0_bits_decodeResult_itype = _RANDOM[8'h2A][22];
        shifterReg_6_0_bits_decodeResult_unsigned1 = _RANDOM[8'h2A][23];
        shifterReg_6_0_bits_decodeResult_unsigned0 = _RANDOM[8'h2A][24];
        shifterReg_6_0_bits_decodeResult_other = _RANDOM[8'h2A][25];
        shifterReg_6_0_bits_decodeResult_multiCycle = _RANDOM[8'h2A][26];
        shifterReg_6_0_bits_decodeResult_divider = _RANDOM[8'h2A][27];
        shifterReg_6_0_bits_decodeResult_multiplier = _RANDOM[8'h2A][28];
        shifterReg_6_0_bits_decodeResult_shift = _RANDOM[8'h2A][29];
        shifterReg_6_0_bits_decodeResult_adder = _RANDOM[8'h2A][30];
        shifterReg_6_0_bits_decodeResult_logic = _RANDOM[8'h2A][31];
        shifterReg_6_0_bits_loadStore = _RANDOM[8'h2B][0];
        shifterReg_6_0_bits_issueInst = _RANDOM[8'h2B][1];
        shifterReg_6_0_bits_store = _RANDOM[8'h2B][2];
        shifterReg_6_0_bits_special = _RANDOM[8'h2B][3];
        shifterReg_6_0_bits_lsWholeReg = _RANDOM[8'h2B][4];
        shifterReg_6_0_bits_vs1 = _RANDOM[8'h2B][9:5];
        shifterReg_6_0_bits_vs2 = _RANDOM[8'h2B][14:10];
        shifterReg_6_0_bits_vd = _RANDOM[8'h2B][19:15];
        shifterReg_6_0_bits_loadStoreEEW = _RANDOM[8'h2B][21:20];
        shifterReg_6_0_bits_mask = _RANDOM[8'h2B][22];
        shifterReg_6_0_bits_segment = _RANDOM[8'h2B][25:23];
        shifterReg_6_0_bits_readFromScalar = {_RANDOM[8'h2B][31:26], _RANDOM[8'h2C][25:0]};
        shifterReg_6_0_bits_csrInterface_vl = {_RANDOM[8'h2C][31:26], _RANDOM[8'h2D][5:0]};
        shifterReg_6_0_bits_csrInterface_vStart = _RANDOM[8'h2D][17:6];
        shifterReg_6_0_bits_csrInterface_vlmul = _RANDOM[8'h2D][20:18];
        shifterReg_6_0_bits_csrInterface_vSew = _RANDOM[8'h2D][22:21];
        shifterReg_6_0_bits_csrInterface_vxrm = _RANDOM[8'h2D][24:23];
        shifterReg_6_0_bits_csrInterface_vta = _RANDOM[8'h2D][25];
        shifterReg_6_0_bits_csrInterface_vma = _RANDOM[8'h2D][26];
        releasePipe_pipe_v_7 = _RANDOM[8'h2D][27];
        tokenCheck_counter_7 = _RANDOM[8'h2D][30:28];
        shifterReg_7_0_valid = _RANDOM[8'h2D][31];
        shifterReg_7_0_bits_instructionIndex = _RANDOM[8'h2E][2:0];
        shifterReg_7_0_bits_decodeResult_specialSlot = _RANDOM[8'h2E][3];
        shifterReg_7_0_bits_decodeResult_topUop = _RANDOM[8'h2E][8:4];
        shifterReg_7_0_bits_decodeResult_popCount = _RANDOM[8'h2E][9];
        shifterReg_7_0_bits_decodeResult_ffo = _RANDOM[8'h2E][10];
        shifterReg_7_0_bits_decodeResult_average = _RANDOM[8'h2E][11];
        shifterReg_7_0_bits_decodeResult_reverse = _RANDOM[8'h2E][12];
        shifterReg_7_0_bits_decodeResult_dontNeedExecuteInLane = _RANDOM[8'h2E][13];
        shifterReg_7_0_bits_decodeResult_scheduler = _RANDOM[8'h2E][14];
        shifterReg_7_0_bits_decodeResult_sReadVD = _RANDOM[8'h2E][15];
        shifterReg_7_0_bits_decodeResult_vtype = _RANDOM[8'h2E][16];
        shifterReg_7_0_bits_decodeResult_sWrite = _RANDOM[8'h2E][17];
        shifterReg_7_0_bits_decodeResult_crossRead = _RANDOM[8'h2E][18];
        shifterReg_7_0_bits_decodeResult_crossWrite = _RANDOM[8'h2E][19];
        shifterReg_7_0_bits_decodeResult_maskUnit = _RANDOM[8'h2E][20];
        shifterReg_7_0_bits_decodeResult_special = _RANDOM[8'h2E][21];
        shifterReg_7_0_bits_decodeResult_saturate = _RANDOM[8'h2E][22];
        shifterReg_7_0_bits_decodeResult_vwmacc = _RANDOM[8'h2E][23];
        shifterReg_7_0_bits_decodeResult_readOnly = _RANDOM[8'h2E][24];
        shifterReg_7_0_bits_decodeResult_maskSource = _RANDOM[8'h2E][25];
        shifterReg_7_0_bits_decodeResult_maskDestination = _RANDOM[8'h2E][26];
        shifterReg_7_0_bits_decodeResult_maskLogic = _RANDOM[8'h2E][27];
        shifterReg_7_0_bits_decodeResult_uop = _RANDOM[8'h2E][31:28];
        shifterReg_7_0_bits_decodeResult_iota = _RANDOM[8'h2F][0];
        shifterReg_7_0_bits_decodeResult_mv = _RANDOM[8'h2F][1];
        shifterReg_7_0_bits_decodeResult_extend = _RANDOM[8'h2F][2];
        shifterReg_7_0_bits_decodeResult_unOrderWrite = _RANDOM[8'h2F][3];
        shifterReg_7_0_bits_decodeResult_compress = _RANDOM[8'h2F][4];
        shifterReg_7_0_bits_decodeResult_gather16 = _RANDOM[8'h2F][5];
        shifterReg_7_0_bits_decodeResult_gather = _RANDOM[8'h2F][6];
        shifterReg_7_0_bits_decodeResult_slid = _RANDOM[8'h2F][7];
        shifterReg_7_0_bits_decodeResult_targetRd = _RANDOM[8'h2F][8];
        shifterReg_7_0_bits_decodeResult_widenReduce = _RANDOM[8'h2F][9];
        shifterReg_7_0_bits_decodeResult_red = _RANDOM[8'h2F][10];
        shifterReg_7_0_bits_decodeResult_nr = _RANDOM[8'h2F][11];
        shifterReg_7_0_bits_decodeResult_itype = _RANDOM[8'h2F][12];
        shifterReg_7_0_bits_decodeResult_unsigned1 = _RANDOM[8'h2F][13];
        shifterReg_7_0_bits_decodeResult_unsigned0 = _RANDOM[8'h2F][14];
        shifterReg_7_0_bits_decodeResult_other = _RANDOM[8'h2F][15];
        shifterReg_7_0_bits_decodeResult_multiCycle = _RANDOM[8'h2F][16];
        shifterReg_7_0_bits_decodeResult_divider = _RANDOM[8'h2F][17];
        shifterReg_7_0_bits_decodeResult_multiplier = _RANDOM[8'h2F][18];
        shifterReg_7_0_bits_decodeResult_shift = _RANDOM[8'h2F][19];
        shifterReg_7_0_bits_decodeResult_adder = _RANDOM[8'h2F][20];
        shifterReg_7_0_bits_decodeResult_logic = _RANDOM[8'h2F][21];
        shifterReg_7_0_bits_loadStore = _RANDOM[8'h2F][22];
        shifterReg_7_0_bits_issueInst = _RANDOM[8'h2F][23];
        shifterReg_7_0_bits_store = _RANDOM[8'h2F][24];
        shifterReg_7_0_bits_special = _RANDOM[8'h2F][25];
        shifterReg_7_0_bits_lsWholeReg = _RANDOM[8'h2F][26];
        shifterReg_7_0_bits_vs1 = _RANDOM[8'h2F][31:27];
        shifterReg_7_0_bits_vs2 = _RANDOM[8'h30][4:0];
        shifterReg_7_0_bits_vd = _RANDOM[8'h30][9:5];
        shifterReg_7_0_bits_loadStoreEEW = _RANDOM[8'h30][11:10];
        shifterReg_7_0_bits_mask = _RANDOM[8'h30][12];
        shifterReg_7_0_bits_segment = _RANDOM[8'h30][15:13];
        shifterReg_7_0_bits_readFromScalar = {_RANDOM[8'h30][31:16], _RANDOM[8'h31][15:0]};
        shifterReg_7_0_bits_csrInterface_vl = _RANDOM[8'h31][27:16];
        shifterReg_7_0_bits_csrInterface_vStart = {_RANDOM[8'h31][31:28], _RANDOM[8'h32][7:0]};
        shifterReg_7_0_bits_csrInterface_vlmul = _RANDOM[8'h32][10:8];
        shifterReg_7_0_bits_csrInterface_vSew = _RANDOM[8'h32][12:11];
        shifterReg_7_0_bits_csrInterface_vxrm = _RANDOM[8'h32][14:13];
        shifterReg_7_0_bits_csrInterface_vta = _RANDOM[8'h32][15];
        shifterReg_7_0_bits_csrInterface_vma = _RANDOM[8'h32][16];
        sinkVec_releasePipe_pipe_v = _RANDOM[8'h32][17];
        sinkVec_tokenCheck_counter = _RANDOM[8'h32][20:18];
        sinkVec_shifterReg_0_valid = _RANDOM[8'h32][21];
        sinkVec_shifterReg_0_bits_vs = _RANDOM[8'h32][26:22];
        sinkVec_shifterReg_0_bits_readSource = _RANDOM[8'h32][28:27];
        sinkVec_shifterReg_0_bits_offset = _RANDOM[8'h32][31:29];
        sinkVec_shifterReg_0_bits_instructionIndex = _RANDOM[8'h33][2:0];
        sinkVec_releasePipe_pipe_v_1 = _RANDOM[8'h33][3];
        sinkVec_tokenCheck_counter_1 = _RANDOM[8'h33][6:4];
        sinkVec_shifterReg_1_0_valid = _RANDOM[8'h33][7];
        sinkVec_shifterReg_1_0_bits_vs = _RANDOM[8'h33][12:8];
        sinkVec_shifterReg_1_0_bits_readSource = _RANDOM[8'h33][14:13];
        sinkVec_shifterReg_1_0_bits_offset = _RANDOM[8'h33][17:15];
        sinkVec_shifterReg_1_0_bits_instructionIndex = _RANDOM[8'h33][20:18];
        maskUnitFirst = _RANDOM[8'h33][21];
        accessDataValid_pipe_v = _RANDOM[8'h33][22];
        accessDataValid_pipe_pipe_v = _RANDOM[8'h33][23];
        shifterReg_8_0_valid = _RANDOM[8'h33][24];
        shifterReg_8_0_bits = {_RANDOM[8'h33][31:25], _RANDOM[8'h34][24:0]};
        accessDataValid_pipe_v_1 = _RANDOM[8'h34][25];
        accessDataValid_pipe_pipe_v_1 = _RANDOM[8'h34][26];
        shifterReg_9_0_valid = _RANDOM[8'h34][27];
        shifterReg_9_0_bits = {_RANDOM[8'h34][31:28], _RANDOM[8'h35][27:0]};
        sinkVec_releasePipe_pipe_v_2 = _RANDOM[8'h35][28];
        sinkVec_tokenCheck_counter_2 = _RANDOM[8'h35][31:29];
        sinkVec_shifterReg_2_0_valid = _RANDOM[8'h36][0];
        sinkVec_shifterReg_2_0_bits_vd = _RANDOM[8'h36][5:1];
        sinkVec_shifterReg_2_0_bits_offset = _RANDOM[8'h36][8:6];
        sinkVec_shifterReg_2_0_bits_mask = _RANDOM[8'h36][12:9];
        sinkVec_shifterReg_2_0_bits_data = {_RANDOM[8'h36][31:13], _RANDOM[8'h37][12:0]};
        sinkVec_shifterReg_2_0_bits_instructionIndex = _RANDOM[8'h37][16:14];
        sinkVec_releasePipe_pipe_v_3 = _RANDOM[8'h37][17];
        sinkVec_tokenCheck_counter_3 = _RANDOM[8'h37][20:18];
        sinkVec_shifterReg_3_0_valid = _RANDOM[8'h37][21];
        sinkVec_shifterReg_3_0_bits_vd = _RANDOM[8'h37][26:22];
        sinkVec_shifterReg_3_0_bits_offset = _RANDOM[8'h37][29:27];
        sinkVec_shifterReg_3_0_bits_mask = {_RANDOM[8'h37][31:30], _RANDOM[8'h38][1:0]};
        sinkVec_shifterReg_3_0_bits_data = {_RANDOM[8'h38][31:2], _RANDOM[8'h39][1:0]};
        sinkVec_shifterReg_3_0_bits_last = _RANDOM[8'h39][2];
        sinkVec_shifterReg_3_0_bits_instructionIndex = _RANDOM[8'h39][5:3];
        maskUnitFirst_1 = _RANDOM[8'h39][6];
        view__writeRelease_0_pipe_v = _RANDOM[8'h39][7];
        pipe_v = _RANDOM[8'h39][8];
        instructionFinishedPipe_pipe_v = _RANDOM[8'h39][9];
        instructionFinishedPipe_pipe_b = _RANDOM[8'h39][17:10];
        pipe_v_1 = _RANDOM[8'h39][18];
        pipe_b_1 = {_RANDOM[8'h39][31:19], _RANDOM[8'h3A][18:0]};
        pipe_pipe_v = _RANDOM[8'h3A][19];
        pipe_pipe_b = {_RANDOM[8'h3A][31:20], _RANDOM[8'h3B][19:0]};
        view__laneMaskSelect_0_pipe_v = _RANDOM[8'h3B][20];
        view__laneMaskSelect_0_pipe_b = _RANDOM[8'h3B][26:21];
        view__laneMaskSelect_0_pipe_pipe_v = _RANDOM[8'h3B][27];
        view__laneMaskSelect_0_pipe_pipe_b = {_RANDOM[8'h3B][31:28], _RANDOM[8'h3C][1:0]};
        view__laneMaskSewSelect_0_pipe_v = _RANDOM[8'h3C][2];
        view__laneMaskSewSelect_0_pipe_b = _RANDOM[8'h3C][4:3];
        view__laneMaskSewSelect_0_pipe_pipe_v = _RANDOM[8'h3C][5];
        view__laneMaskSewSelect_0_pipe_pipe_b = _RANDOM[8'h3C][7:6];
        lsuLastPipe_pipe_v = _RANDOM[8'h3C][8];
        lsuLastPipe_pipe_b = _RANDOM[8'h3C][16:9];
        maskLastPipe_pipe_v = _RANDOM[8'h3C][17];
        maskLastPipe_pipe_b = _RANDOM[8'h3C][25:18];
        pipe_v_2 = _RANDOM[8'h3C][26];
        pipe_b_2 = {_RANDOM[8'h3C][31:27], _RANDOM[8'h3D][1:0]};
        sinkVec_releasePipe_pipe_v_4 = _RANDOM[8'h3D][2];
        sinkVec_tokenCheck_counter_4 = _RANDOM[8'h3D][5:3];
        sinkVec_shifterReg_4_0_valid = _RANDOM[8'h3D][6];
        sinkVec_shifterReg_4_0_bits_vs = _RANDOM[8'h3D][11:7];
        sinkVec_shifterReg_4_0_bits_readSource = _RANDOM[8'h3D][13:12];
        sinkVec_shifterReg_4_0_bits_offset = _RANDOM[8'h3D][16:14];
        sinkVec_shifterReg_4_0_bits_instructionIndex = _RANDOM[8'h3D][19:17];
        sinkVec_releasePipe_pipe_v_5 = _RANDOM[8'h3D][20];
        sinkVec_tokenCheck_counter_5 = _RANDOM[8'h3D][23:21];
        sinkVec_shifterReg_5_0_valid = _RANDOM[8'h3D][24];
        sinkVec_shifterReg_5_0_bits_vs = _RANDOM[8'h3D][29:25];
        sinkVec_shifterReg_5_0_bits_readSource = _RANDOM[8'h3D][31:30];
        sinkVec_shifterReg_5_0_bits_offset = _RANDOM[8'h3E][2:0];
        sinkVec_shifterReg_5_0_bits_instructionIndex = _RANDOM[8'h3E][5:3];
        maskUnitFirst_2 = _RANDOM[8'h3E][6];
        accessDataValid_pipe_v_2 = _RANDOM[8'h3E][7];
        accessDataValid_pipe_pipe_v_2 = _RANDOM[8'h3E][8];
        shifterReg_10_0_valid = _RANDOM[8'h3E][9];
        shifterReg_10_0_bits = {_RANDOM[8'h3E][31:10], _RANDOM[8'h3F][9:0]};
        accessDataValid_pipe_v_3 = _RANDOM[8'h3F][10];
        accessDataValid_pipe_pipe_v_3 = _RANDOM[8'h3F][11];
        shifterReg_11_0_valid = _RANDOM[8'h3F][12];
        shifterReg_11_0_bits = {_RANDOM[8'h3F][31:13], _RANDOM[8'h40][12:0]};
        sinkVec_releasePipe_pipe_v_6 = _RANDOM[8'h40][13];
        sinkVec_tokenCheck_counter_6 = _RANDOM[8'h40][16:14];
        sinkVec_shifterReg_6_0_valid = _RANDOM[8'h40][17];
        sinkVec_shifterReg_6_0_bits_vd = _RANDOM[8'h40][22:18];
        sinkVec_shifterReg_6_0_bits_offset = _RANDOM[8'h40][25:23];
        sinkVec_shifterReg_6_0_bits_mask = _RANDOM[8'h40][29:26];
        sinkVec_shifterReg_6_0_bits_data = {_RANDOM[8'h40][31:30], _RANDOM[8'h41][29:0]};
        sinkVec_shifterReg_6_0_bits_instructionIndex = {_RANDOM[8'h41][31], _RANDOM[8'h42][1:0]};
        sinkVec_releasePipe_pipe_v_7 = _RANDOM[8'h42][2];
        sinkVec_tokenCheck_counter_7 = _RANDOM[8'h42][5:3];
        sinkVec_shifterReg_7_0_valid = _RANDOM[8'h42][6];
        sinkVec_shifterReg_7_0_bits_vd = _RANDOM[8'h42][11:7];
        sinkVec_shifterReg_7_0_bits_offset = _RANDOM[8'h42][14:12];
        sinkVec_shifterReg_7_0_bits_mask = _RANDOM[8'h42][18:15];
        sinkVec_shifterReg_7_0_bits_data = {_RANDOM[8'h42][31:19], _RANDOM[8'h43][18:0]};
        sinkVec_shifterReg_7_0_bits_last = _RANDOM[8'h43][19];
        sinkVec_shifterReg_7_0_bits_instructionIndex = _RANDOM[8'h43][22:20];
        maskUnitFirst_3 = _RANDOM[8'h43][23];
        view__writeRelease_1_pipe_v = _RANDOM[8'h43][24];
        pipe_v_3 = _RANDOM[8'h43][25];
        instructionFinishedPipe_pipe_v_1 = _RANDOM[8'h43][26];
        instructionFinishedPipe_pipe_b_1 = {_RANDOM[8'h43][31:27], _RANDOM[8'h44][2:0]};
        pipe_v_4 = _RANDOM[8'h44][3];
        pipe_b_4 = {_RANDOM[8'h44][31:4], _RANDOM[8'h45][3:0]};
        pipe_pipe_v_1 = _RANDOM[8'h45][4];
        pipe_pipe_b_1 = {_RANDOM[8'h45][31:5], _RANDOM[8'h46][4:0]};
        view__laneMaskSelect_1_pipe_v = _RANDOM[8'h46][5];
        view__laneMaskSelect_1_pipe_b = _RANDOM[8'h46][11:6];
        view__laneMaskSelect_1_pipe_pipe_v = _RANDOM[8'h46][12];
        view__laneMaskSelect_1_pipe_pipe_b = _RANDOM[8'h46][18:13];
        view__laneMaskSewSelect_1_pipe_v = _RANDOM[8'h46][19];
        view__laneMaskSewSelect_1_pipe_b = _RANDOM[8'h46][21:20];
        view__laneMaskSewSelect_1_pipe_pipe_v = _RANDOM[8'h46][22];
        view__laneMaskSewSelect_1_pipe_pipe_b = _RANDOM[8'h46][24:23];
        lsuLastPipe_pipe_v_1 = _RANDOM[8'h46][25];
        lsuLastPipe_pipe_b_1 = {_RANDOM[8'h46][31:26], _RANDOM[8'h47][1:0]};
        maskLastPipe_pipe_v_1 = _RANDOM[8'h47][2];
        maskLastPipe_pipe_b_1 = _RANDOM[8'h47][10:3];
        pipe_v_5 = _RANDOM[8'h47][11];
        pipe_b_5 = _RANDOM[8'h47][18:12];
        sinkVec_releasePipe_pipe_v_8 = _RANDOM[8'h47][19];
        sinkVec_tokenCheck_counter_8 = _RANDOM[8'h47][22:20];
        sinkVec_shifterReg_8_0_valid = _RANDOM[8'h47][23];
        sinkVec_shifterReg_8_0_bits_vs = _RANDOM[8'h47][28:24];
        sinkVec_shifterReg_8_0_bits_readSource = _RANDOM[8'h47][30:29];
        sinkVec_shifterReg_8_0_bits_offset = {_RANDOM[8'h47][31], _RANDOM[8'h48][1:0]};
        sinkVec_shifterReg_8_0_bits_instructionIndex = _RANDOM[8'h48][4:2];
        sinkVec_releasePipe_pipe_v_9 = _RANDOM[8'h48][5];
        sinkVec_tokenCheck_counter_9 = _RANDOM[8'h48][8:6];
        sinkVec_shifterReg_9_0_valid = _RANDOM[8'h48][9];
        sinkVec_shifterReg_9_0_bits_vs = _RANDOM[8'h48][14:10];
        sinkVec_shifterReg_9_0_bits_readSource = _RANDOM[8'h48][16:15];
        sinkVec_shifterReg_9_0_bits_offset = _RANDOM[8'h48][19:17];
        sinkVec_shifterReg_9_0_bits_instructionIndex = _RANDOM[8'h48][22:20];
        maskUnitFirst_4 = _RANDOM[8'h48][23];
        accessDataValid_pipe_v_4 = _RANDOM[8'h48][24];
        accessDataValid_pipe_pipe_v_4 = _RANDOM[8'h48][25];
        shifterReg_12_0_valid = _RANDOM[8'h48][26];
        shifterReg_12_0_bits = {_RANDOM[8'h48][31:27], _RANDOM[8'h49][26:0]};
        accessDataValid_pipe_v_5 = _RANDOM[8'h49][27];
        accessDataValid_pipe_pipe_v_5 = _RANDOM[8'h49][28];
        shifterReg_13_0_valid = _RANDOM[8'h49][29];
        shifterReg_13_0_bits = {_RANDOM[8'h49][31:30], _RANDOM[8'h4A][29:0]};
        sinkVec_releasePipe_pipe_v_10 = _RANDOM[8'h4A][30];
        sinkVec_tokenCheck_counter_10 = {_RANDOM[8'h4A][31], _RANDOM[8'h4B][1:0]};
        sinkVec_shifterReg_10_0_valid = _RANDOM[8'h4B][2];
        sinkVec_shifterReg_10_0_bits_vd = _RANDOM[8'h4B][7:3];
        sinkVec_shifterReg_10_0_bits_offset = _RANDOM[8'h4B][10:8];
        sinkVec_shifterReg_10_0_bits_mask = _RANDOM[8'h4B][14:11];
        sinkVec_shifterReg_10_0_bits_data = {_RANDOM[8'h4B][31:15], _RANDOM[8'h4C][14:0]};
        sinkVec_shifterReg_10_0_bits_instructionIndex = _RANDOM[8'h4C][18:16];
        sinkVec_releasePipe_pipe_v_11 = _RANDOM[8'h4C][19];
        sinkVec_tokenCheck_counter_11 = _RANDOM[8'h4C][22:20];
        sinkVec_shifterReg_11_0_valid = _RANDOM[8'h4C][23];
        sinkVec_shifterReg_11_0_bits_vd = _RANDOM[8'h4C][28:24];
        sinkVec_shifterReg_11_0_bits_offset = _RANDOM[8'h4C][31:29];
        sinkVec_shifterReg_11_0_bits_mask = _RANDOM[8'h4D][3:0];
        sinkVec_shifterReg_11_0_bits_data = {_RANDOM[8'h4D][31:4], _RANDOM[8'h4E][3:0]};
        sinkVec_shifterReg_11_0_bits_last = _RANDOM[8'h4E][4];
        sinkVec_shifterReg_11_0_bits_instructionIndex = _RANDOM[8'h4E][7:5];
        maskUnitFirst_5 = _RANDOM[8'h4E][8];
        view__writeRelease_2_pipe_v = _RANDOM[8'h4E][9];
        pipe_v_6 = _RANDOM[8'h4E][10];
        instructionFinishedPipe_pipe_v_2 = _RANDOM[8'h4E][11];
        instructionFinishedPipe_pipe_b_2 = _RANDOM[8'h4E][19:12];
        pipe_v_7 = _RANDOM[8'h4E][20];
        pipe_b_7 = {_RANDOM[8'h4E][31:21], _RANDOM[8'h4F][20:0]};
        pipe_pipe_v_2 = _RANDOM[8'h4F][21];
        pipe_pipe_b_2 = {_RANDOM[8'h4F][31:22], _RANDOM[8'h50][21:0]};
        view__laneMaskSelect_2_pipe_v = _RANDOM[8'h50][22];
        view__laneMaskSelect_2_pipe_b = _RANDOM[8'h50][28:23];
        view__laneMaskSelect_2_pipe_pipe_v = _RANDOM[8'h50][29];
        view__laneMaskSelect_2_pipe_pipe_b = {_RANDOM[8'h50][31:30], _RANDOM[8'h51][3:0]};
        view__laneMaskSewSelect_2_pipe_v = _RANDOM[8'h51][4];
        view__laneMaskSewSelect_2_pipe_b = _RANDOM[8'h51][6:5];
        view__laneMaskSewSelect_2_pipe_pipe_v = _RANDOM[8'h51][7];
        view__laneMaskSewSelect_2_pipe_pipe_b = _RANDOM[8'h51][9:8];
        lsuLastPipe_pipe_v_2 = _RANDOM[8'h51][10];
        lsuLastPipe_pipe_b_2 = _RANDOM[8'h51][18:11];
        maskLastPipe_pipe_v_2 = _RANDOM[8'h51][19];
        maskLastPipe_pipe_b_2 = _RANDOM[8'h51][27:20];
        pipe_v_8 = _RANDOM[8'h51][28];
        pipe_b_8 = {_RANDOM[8'h51][31:29], _RANDOM[8'h52][3:0]};
        sinkVec_releasePipe_pipe_v_12 = _RANDOM[8'h52][4];
        sinkVec_tokenCheck_counter_12 = _RANDOM[8'h52][7:5];
        sinkVec_shifterReg_12_0_valid = _RANDOM[8'h52][8];
        sinkVec_shifterReg_12_0_bits_vs = _RANDOM[8'h52][13:9];
        sinkVec_shifterReg_12_0_bits_readSource = _RANDOM[8'h52][15:14];
        sinkVec_shifterReg_12_0_bits_offset = _RANDOM[8'h52][18:16];
        sinkVec_shifterReg_12_0_bits_instructionIndex = _RANDOM[8'h52][21:19];
        sinkVec_releasePipe_pipe_v_13 = _RANDOM[8'h52][22];
        sinkVec_tokenCheck_counter_13 = _RANDOM[8'h52][25:23];
        sinkVec_shifterReg_13_0_valid = _RANDOM[8'h52][26];
        sinkVec_shifterReg_13_0_bits_vs = _RANDOM[8'h52][31:27];
        sinkVec_shifterReg_13_0_bits_readSource = _RANDOM[8'h53][1:0];
        sinkVec_shifterReg_13_0_bits_offset = _RANDOM[8'h53][4:2];
        sinkVec_shifterReg_13_0_bits_instructionIndex = _RANDOM[8'h53][7:5];
        maskUnitFirst_6 = _RANDOM[8'h53][8];
        accessDataValid_pipe_v_6 = _RANDOM[8'h53][9];
        accessDataValid_pipe_pipe_v_6 = _RANDOM[8'h53][10];
        shifterReg_14_0_valid = _RANDOM[8'h53][11];
        shifterReg_14_0_bits = {_RANDOM[8'h53][31:12], _RANDOM[8'h54][11:0]};
        accessDataValid_pipe_v_7 = _RANDOM[8'h54][12];
        accessDataValid_pipe_pipe_v_7 = _RANDOM[8'h54][13];
        shifterReg_15_0_valid = _RANDOM[8'h54][14];
        shifterReg_15_0_bits = {_RANDOM[8'h54][31:15], _RANDOM[8'h55][14:0]};
        sinkVec_releasePipe_pipe_v_14 = _RANDOM[8'h55][15];
        sinkVec_tokenCheck_counter_14 = _RANDOM[8'h55][18:16];
        sinkVec_shifterReg_14_0_valid = _RANDOM[8'h55][19];
        sinkVec_shifterReg_14_0_bits_vd = _RANDOM[8'h55][24:20];
        sinkVec_shifterReg_14_0_bits_offset = _RANDOM[8'h55][27:25];
        sinkVec_shifterReg_14_0_bits_mask = _RANDOM[8'h55][31:28];
        sinkVec_shifterReg_14_0_bits_data = _RANDOM[8'h56];
        sinkVec_shifterReg_14_0_bits_instructionIndex = _RANDOM[8'h57][3:1];
        sinkVec_releasePipe_pipe_v_15 = _RANDOM[8'h57][4];
        sinkVec_tokenCheck_counter_15 = _RANDOM[8'h57][7:5];
        sinkVec_shifterReg_15_0_valid = _RANDOM[8'h57][8];
        sinkVec_shifterReg_15_0_bits_vd = _RANDOM[8'h57][13:9];
        sinkVec_shifterReg_15_0_bits_offset = _RANDOM[8'h57][16:14];
        sinkVec_shifterReg_15_0_bits_mask = _RANDOM[8'h57][20:17];
        sinkVec_shifterReg_15_0_bits_data = {_RANDOM[8'h57][31:21], _RANDOM[8'h58][20:0]};
        sinkVec_shifterReg_15_0_bits_last = _RANDOM[8'h58][21];
        sinkVec_shifterReg_15_0_bits_instructionIndex = _RANDOM[8'h58][24:22];
        maskUnitFirst_7 = _RANDOM[8'h58][25];
        view__writeRelease_3_pipe_v = _RANDOM[8'h58][26];
        pipe_v_9 = _RANDOM[8'h58][27];
        instructionFinishedPipe_pipe_v_3 = _RANDOM[8'h58][28];
        instructionFinishedPipe_pipe_b_3 = {_RANDOM[8'h58][31:29], _RANDOM[8'h59][4:0]};
        pipe_v_10 = _RANDOM[8'h59][5];
        pipe_b_10 = {_RANDOM[8'h59][31:6], _RANDOM[8'h5A][5:0]};
        pipe_pipe_v_3 = _RANDOM[8'h5A][6];
        pipe_pipe_b_3 = {_RANDOM[8'h5A][31:7], _RANDOM[8'h5B][6:0]};
        view__laneMaskSelect_3_pipe_v = _RANDOM[8'h5B][7];
        view__laneMaskSelect_3_pipe_b = _RANDOM[8'h5B][13:8];
        view__laneMaskSelect_3_pipe_pipe_v = _RANDOM[8'h5B][14];
        view__laneMaskSelect_3_pipe_pipe_b = _RANDOM[8'h5B][20:15];
        view__laneMaskSewSelect_3_pipe_v = _RANDOM[8'h5B][21];
        view__laneMaskSewSelect_3_pipe_b = _RANDOM[8'h5B][23:22];
        view__laneMaskSewSelect_3_pipe_pipe_v = _RANDOM[8'h5B][24];
        view__laneMaskSewSelect_3_pipe_pipe_b = _RANDOM[8'h5B][26:25];
        lsuLastPipe_pipe_v_3 = _RANDOM[8'h5B][27];
        lsuLastPipe_pipe_b_3 = {_RANDOM[8'h5B][31:28], _RANDOM[8'h5C][3:0]};
        maskLastPipe_pipe_v_3 = _RANDOM[8'h5C][4];
        maskLastPipe_pipe_b_3 = _RANDOM[8'h5C][12:5];
        pipe_v_11 = _RANDOM[8'h5C][13];
        pipe_b_11 = _RANDOM[8'h5C][20:14];
        sinkVec_releasePipe_pipe_v_16 = _RANDOM[8'h5C][21];
        sinkVec_tokenCheck_counter_16 = _RANDOM[8'h5C][24:22];
        sinkVec_shifterReg_16_0_valid = _RANDOM[8'h5C][25];
        sinkVec_shifterReg_16_0_bits_vs = _RANDOM[8'h5C][30:26];
        sinkVec_shifterReg_16_0_bits_readSource = {_RANDOM[8'h5C][31], _RANDOM[8'h5D][0]};
        sinkVec_shifterReg_16_0_bits_offset = _RANDOM[8'h5D][3:1];
        sinkVec_shifterReg_16_0_bits_instructionIndex = _RANDOM[8'h5D][6:4];
        sinkVec_releasePipe_pipe_v_17 = _RANDOM[8'h5D][7];
        sinkVec_tokenCheck_counter_17 = _RANDOM[8'h5D][10:8];
        sinkVec_shifterReg_17_0_valid = _RANDOM[8'h5D][11];
        sinkVec_shifterReg_17_0_bits_vs = _RANDOM[8'h5D][16:12];
        sinkVec_shifterReg_17_0_bits_readSource = _RANDOM[8'h5D][18:17];
        sinkVec_shifterReg_17_0_bits_offset = _RANDOM[8'h5D][21:19];
        sinkVec_shifterReg_17_0_bits_instructionIndex = _RANDOM[8'h5D][24:22];
        maskUnitFirst_8 = _RANDOM[8'h5D][25];
        accessDataValid_pipe_v_8 = _RANDOM[8'h5D][26];
        accessDataValid_pipe_pipe_v_8 = _RANDOM[8'h5D][27];
        shifterReg_16_0_valid = _RANDOM[8'h5D][28];
        shifterReg_16_0_bits = {_RANDOM[8'h5D][31:29], _RANDOM[8'h5E][28:0]};
        accessDataValid_pipe_v_9 = _RANDOM[8'h5E][29];
        accessDataValid_pipe_pipe_v_9 = _RANDOM[8'h5E][30];
        shifterReg_17_0_valid = _RANDOM[8'h5E][31];
        shifterReg_17_0_bits = _RANDOM[8'h5F];
        sinkVec_releasePipe_pipe_v_18 = _RANDOM[8'h60][0];
        sinkVec_tokenCheck_counter_18 = _RANDOM[8'h60][3:1];
        sinkVec_shifterReg_18_0_valid = _RANDOM[8'h60][4];
        sinkVec_shifterReg_18_0_bits_vd = _RANDOM[8'h60][9:5];
        sinkVec_shifterReg_18_0_bits_offset = _RANDOM[8'h60][12:10];
        sinkVec_shifterReg_18_0_bits_mask = _RANDOM[8'h60][16:13];
        sinkVec_shifterReg_18_0_bits_data = {_RANDOM[8'h60][31:17], _RANDOM[8'h61][16:0]};
        sinkVec_shifterReg_18_0_bits_instructionIndex = _RANDOM[8'h61][20:18];
        sinkVec_releasePipe_pipe_v_19 = _RANDOM[8'h61][21];
        sinkVec_tokenCheck_counter_19 = _RANDOM[8'h61][24:22];
        sinkVec_shifterReg_19_0_valid = _RANDOM[8'h61][25];
        sinkVec_shifterReg_19_0_bits_vd = _RANDOM[8'h61][30:26];
        sinkVec_shifterReg_19_0_bits_offset = {_RANDOM[8'h61][31], _RANDOM[8'h62][1:0]};
        sinkVec_shifterReg_19_0_bits_mask = _RANDOM[8'h62][5:2];
        sinkVec_shifterReg_19_0_bits_data = {_RANDOM[8'h62][31:6], _RANDOM[8'h63][5:0]};
        sinkVec_shifterReg_19_0_bits_last = _RANDOM[8'h63][6];
        sinkVec_shifterReg_19_0_bits_instructionIndex = _RANDOM[8'h63][9:7];
        maskUnitFirst_9 = _RANDOM[8'h63][10];
        view__writeRelease_4_pipe_v = _RANDOM[8'h63][11];
        pipe_v_12 = _RANDOM[8'h63][12];
        instructionFinishedPipe_pipe_v_4 = _RANDOM[8'h63][13];
        instructionFinishedPipe_pipe_b_4 = _RANDOM[8'h63][21:14];
        pipe_v_13 = _RANDOM[8'h63][22];
        pipe_b_13 = {_RANDOM[8'h63][31:23], _RANDOM[8'h64][22:0]};
        pipe_pipe_v_4 = _RANDOM[8'h64][23];
        pipe_pipe_b_4 = {_RANDOM[8'h64][31:24], _RANDOM[8'h65][23:0]};
        view__laneMaskSelect_4_pipe_v = _RANDOM[8'h65][24];
        view__laneMaskSelect_4_pipe_b = _RANDOM[8'h65][30:25];
        view__laneMaskSelect_4_pipe_pipe_v = _RANDOM[8'h65][31];
        view__laneMaskSelect_4_pipe_pipe_b = _RANDOM[8'h66][5:0];
        view__laneMaskSewSelect_4_pipe_v = _RANDOM[8'h66][6];
        view__laneMaskSewSelect_4_pipe_b = _RANDOM[8'h66][8:7];
        view__laneMaskSewSelect_4_pipe_pipe_v = _RANDOM[8'h66][9];
        view__laneMaskSewSelect_4_pipe_pipe_b = _RANDOM[8'h66][11:10];
        lsuLastPipe_pipe_v_4 = _RANDOM[8'h66][12];
        lsuLastPipe_pipe_b_4 = _RANDOM[8'h66][20:13];
        maskLastPipe_pipe_v_4 = _RANDOM[8'h66][21];
        maskLastPipe_pipe_b_4 = _RANDOM[8'h66][29:22];
        pipe_v_14 = _RANDOM[8'h66][30];
        pipe_b_14 = {_RANDOM[8'h66][31], _RANDOM[8'h67][5:0]};
        sinkVec_releasePipe_pipe_v_20 = _RANDOM[8'h67][6];
        sinkVec_tokenCheck_counter_20 = _RANDOM[8'h67][9:7];
        sinkVec_shifterReg_20_0_valid = _RANDOM[8'h67][10];
        sinkVec_shifterReg_20_0_bits_vs = _RANDOM[8'h67][15:11];
        sinkVec_shifterReg_20_0_bits_readSource = _RANDOM[8'h67][17:16];
        sinkVec_shifterReg_20_0_bits_offset = _RANDOM[8'h67][20:18];
        sinkVec_shifterReg_20_0_bits_instructionIndex = _RANDOM[8'h67][23:21];
        sinkVec_releasePipe_pipe_v_21 = _RANDOM[8'h67][24];
        sinkVec_tokenCheck_counter_21 = _RANDOM[8'h67][27:25];
        sinkVec_shifterReg_21_0_valid = _RANDOM[8'h67][28];
        sinkVec_shifterReg_21_0_bits_vs = {_RANDOM[8'h67][31:29], _RANDOM[8'h68][1:0]};
        sinkVec_shifterReg_21_0_bits_readSource = _RANDOM[8'h68][3:2];
        sinkVec_shifterReg_21_0_bits_offset = _RANDOM[8'h68][6:4];
        sinkVec_shifterReg_21_0_bits_instructionIndex = _RANDOM[8'h68][9:7];
        maskUnitFirst_10 = _RANDOM[8'h68][10];
        accessDataValid_pipe_v_10 = _RANDOM[8'h68][11];
        accessDataValid_pipe_pipe_v_10 = _RANDOM[8'h68][12];
        shifterReg_18_0_valid = _RANDOM[8'h68][13];
        shifterReg_18_0_bits = {_RANDOM[8'h68][31:14], _RANDOM[8'h69][13:0]};
        accessDataValid_pipe_v_11 = _RANDOM[8'h69][14];
        accessDataValid_pipe_pipe_v_11 = _RANDOM[8'h69][15];
        shifterReg_19_0_valid = _RANDOM[8'h69][16];
        shifterReg_19_0_bits = {_RANDOM[8'h69][31:17], _RANDOM[8'h6A][16:0]};
        sinkVec_releasePipe_pipe_v_22 = _RANDOM[8'h6A][17];
        sinkVec_tokenCheck_counter_22 = _RANDOM[8'h6A][20:18];
        sinkVec_shifterReg_22_0_valid = _RANDOM[8'h6A][21];
        sinkVec_shifterReg_22_0_bits_vd = _RANDOM[8'h6A][26:22];
        sinkVec_shifterReg_22_0_bits_offset = _RANDOM[8'h6A][29:27];
        sinkVec_shifterReg_22_0_bits_mask = {_RANDOM[8'h6A][31:30], _RANDOM[8'h6B][1:0]};
        sinkVec_shifterReg_22_0_bits_data = {_RANDOM[8'h6B][31:2], _RANDOM[8'h6C][1:0]};
        sinkVec_shifterReg_22_0_bits_instructionIndex = _RANDOM[8'h6C][5:3];
        sinkVec_releasePipe_pipe_v_23 = _RANDOM[8'h6C][6];
        sinkVec_tokenCheck_counter_23 = _RANDOM[8'h6C][9:7];
        sinkVec_shifterReg_23_0_valid = _RANDOM[8'h6C][10];
        sinkVec_shifterReg_23_0_bits_vd = _RANDOM[8'h6C][15:11];
        sinkVec_shifterReg_23_0_bits_offset = _RANDOM[8'h6C][18:16];
        sinkVec_shifterReg_23_0_bits_mask = _RANDOM[8'h6C][22:19];
        sinkVec_shifterReg_23_0_bits_data = {_RANDOM[8'h6C][31:23], _RANDOM[8'h6D][22:0]};
        sinkVec_shifterReg_23_0_bits_last = _RANDOM[8'h6D][23];
        sinkVec_shifterReg_23_0_bits_instructionIndex = _RANDOM[8'h6D][26:24];
        maskUnitFirst_11 = _RANDOM[8'h6D][27];
        view__writeRelease_5_pipe_v = _RANDOM[8'h6D][28];
        pipe_v_15 = _RANDOM[8'h6D][29];
        instructionFinishedPipe_pipe_v_5 = _RANDOM[8'h6D][30];
        instructionFinishedPipe_pipe_b_5 = {_RANDOM[8'h6D][31], _RANDOM[8'h6E][6:0]};
        pipe_v_16 = _RANDOM[8'h6E][7];
        pipe_b_16 = {_RANDOM[8'h6E][31:8], _RANDOM[8'h6F][7:0]};
        pipe_pipe_v_5 = _RANDOM[8'h6F][8];
        pipe_pipe_b_5 = {_RANDOM[8'h6F][31:9], _RANDOM[8'h70][8:0]};
        view__laneMaskSelect_5_pipe_v = _RANDOM[8'h70][9];
        view__laneMaskSelect_5_pipe_b = _RANDOM[8'h70][15:10];
        view__laneMaskSelect_5_pipe_pipe_v = _RANDOM[8'h70][16];
        view__laneMaskSelect_5_pipe_pipe_b = _RANDOM[8'h70][22:17];
        view__laneMaskSewSelect_5_pipe_v = _RANDOM[8'h70][23];
        view__laneMaskSewSelect_5_pipe_b = _RANDOM[8'h70][25:24];
        view__laneMaskSewSelect_5_pipe_pipe_v = _RANDOM[8'h70][26];
        view__laneMaskSewSelect_5_pipe_pipe_b = _RANDOM[8'h70][28:27];
        lsuLastPipe_pipe_v_5 = _RANDOM[8'h70][29];
        lsuLastPipe_pipe_b_5 = {_RANDOM[8'h70][31:30], _RANDOM[8'h71][5:0]};
        maskLastPipe_pipe_v_5 = _RANDOM[8'h71][6];
        maskLastPipe_pipe_b_5 = _RANDOM[8'h71][14:7];
        pipe_v_17 = _RANDOM[8'h71][15];
        pipe_b_17 = _RANDOM[8'h71][22:16];
        sinkVec_releasePipe_pipe_v_24 = _RANDOM[8'h71][23];
        sinkVec_tokenCheck_counter_24 = _RANDOM[8'h71][26:24];
        sinkVec_shifterReg_24_0_valid = _RANDOM[8'h71][27];
        sinkVec_shifterReg_24_0_bits_vs = {_RANDOM[8'h71][31:28], _RANDOM[8'h72][0]};
        sinkVec_shifterReg_24_0_bits_readSource = _RANDOM[8'h72][2:1];
        sinkVec_shifterReg_24_0_bits_offset = _RANDOM[8'h72][5:3];
        sinkVec_shifterReg_24_0_bits_instructionIndex = _RANDOM[8'h72][8:6];
        sinkVec_releasePipe_pipe_v_25 = _RANDOM[8'h72][9];
        sinkVec_tokenCheck_counter_25 = _RANDOM[8'h72][12:10];
        sinkVec_shifterReg_25_0_valid = _RANDOM[8'h72][13];
        sinkVec_shifterReg_25_0_bits_vs = _RANDOM[8'h72][18:14];
        sinkVec_shifterReg_25_0_bits_readSource = _RANDOM[8'h72][20:19];
        sinkVec_shifterReg_25_0_bits_offset = _RANDOM[8'h72][23:21];
        sinkVec_shifterReg_25_0_bits_instructionIndex = _RANDOM[8'h72][26:24];
        maskUnitFirst_12 = _RANDOM[8'h72][27];
        accessDataValid_pipe_v_12 = _RANDOM[8'h72][28];
        accessDataValid_pipe_pipe_v_12 = _RANDOM[8'h72][29];
        shifterReg_20_0_valid = _RANDOM[8'h72][30];
        shifterReg_20_0_bits = {_RANDOM[8'h72][31], _RANDOM[8'h73][30:0]};
        accessDataValid_pipe_v_13 = _RANDOM[8'h73][31];
        accessDataValid_pipe_pipe_v_13 = _RANDOM[8'h74][0];
        shifterReg_21_0_valid = _RANDOM[8'h74][1];
        shifterReg_21_0_bits = {_RANDOM[8'h74][31:2], _RANDOM[8'h75][1:0]};
        sinkVec_releasePipe_pipe_v_26 = _RANDOM[8'h75][2];
        sinkVec_tokenCheck_counter_26 = _RANDOM[8'h75][5:3];
        sinkVec_shifterReg_26_0_valid = _RANDOM[8'h75][6];
        sinkVec_shifterReg_26_0_bits_vd = _RANDOM[8'h75][11:7];
        sinkVec_shifterReg_26_0_bits_offset = _RANDOM[8'h75][14:12];
        sinkVec_shifterReg_26_0_bits_mask = _RANDOM[8'h75][18:15];
        sinkVec_shifterReg_26_0_bits_data = {_RANDOM[8'h75][31:19], _RANDOM[8'h76][18:0]};
        sinkVec_shifterReg_26_0_bits_instructionIndex = _RANDOM[8'h76][22:20];
        sinkVec_releasePipe_pipe_v_27 = _RANDOM[8'h76][23];
        sinkVec_tokenCheck_counter_27 = _RANDOM[8'h76][26:24];
        sinkVec_shifterReg_27_0_valid = _RANDOM[8'h76][27];
        sinkVec_shifterReg_27_0_bits_vd = {_RANDOM[8'h76][31:28], _RANDOM[8'h77][0]};
        sinkVec_shifterReg_27_0_bits_offset = _RANDOM[8'h77][3:1];
        sinkVec_shifterReg_27_0_bits_mask = _RANDOM[8'h77][7:4];
        sinkVec_shifterReg_27_0_bits_data = {_RANDOM[8'h77][31:8], _RANDOM[8'h78][7:0]};
        sinkVec_shifterReg_27_0_bits_last = _RANDOM[8'h78][8];
        sinkVec_shifterReg_27_0_bits_instructionIndex = _RANDOM[8'h78][11:9];
        maskUnitFirst_13 = _RANDOM[8'h78][12];
        view__writeRelease_6_pipe_v = _RANDOM[8'h78][13];
        pipe_v_18 = _RANDOM[8'h78][14];
        instructionFinishedPipe_pipe_v_6 = _RANDOM[8'h78][15];
        instructionFinishedPipe_pipe_b_6 = _RANDOM[8'h78][23:16];
        pipe_v_19 = _RANDOM[8'h78][24];
        pipe_b_19 = {_RANDOM[8'h78][31:25], _RANDOM[8'h79][24:0]};
        pipe_pipe_v_6 = _RANDOM[8'h79][25];
        pipe_pipe_b_6 = {_RANDOM[8'h79][31:26], _RANDOM[8'h7A][25:0]};
        view__laneMaskSelect_6_pipe_v = _RANDOM[8'h7A][26];
        view__laneMaskSelect_6_pipe_b = {_RANDOM[8'h7A][31:27], _RANDOM[8'h7B][0]};
        view__laneMaskSelect_6_pipe_pipe_v = _RANDOM[8'h7B][1];
        view__laneMaskSelect_6_pipe_pipe_b = _RANDOM[8'h7B][7:2];
        view__laneMaskSewSelect_6_pipe_v = _RANDOM[8'h7B][8];
        view__laneMaskSewSelect_6_pipe_b = _RANDOM[8'h7B][10:9];
        view__laneMaskSewSelect_6_pipe_pipe_v = _RANDOM[8'h7B][11];
        view__laneMaskSewSelect_6_pipe_pipe_b = _RANDOM[8'h7B][13:12];
        lsuLastPipe_pipe_v_6 = _RANDOM[8'h7B][14];
        lsuLastPipe_pipe_b_6 = _RANDOM[8'h7B][22:15];
        maskLastPipe_pipe_v_6 = _RANDOM[8'h7B][23];
        maskLastPipe_pipe_b_6 = _RANDOM[8'h7B][31:24];
        pipe_v_20 = _RANDOM[8'h7C][0];
        pipe_b_20 = _RANDOM[8'h7C][7:1];
        sinkVec_releasePipe_pipe_v_28 = _RANDOM[8'h7C][8];
        sinkVec_tokenCheck_counter_28 = _RANDOM[8'h7C][11:9];
        sinkVec_shifterReg_28_0_valid = _RANDOM[8'h7C][12];
        sinkVec_shifterReg_28_0_bits_vs = _RANDOM[8'h7C][17:13];
        sinkVec_shifterReg_28_0_bits_readSource = _RANDOM[8'h7C][19:18];
        sinkVec_shifterReg_28_0_bits_offset = _RANDOM[8'h7C][22:20];
        sinkVec_shifterReg_28_0_bits_instructionIndex = _RANDOM[8'h7C][25:23];
        sinkVec_releasePipe_pipe_v_29 = _RANDOM[8'h7C][26];
        sinkVec_tokenCheck_counter_29 = _RANDOM[8'h7C][29:27];
        sinkVec_shifterReg_29_0_valid = _RANDOM[8'h7C][30];
        sinkVec_shifterReg_29_0_bits_vs = {_RANDOM[8'h7C][31], _RANDOM[8'h7D][3:0]};
        sinkVec_shifterReg_29_0_bits_readSource = _RANDOM[8'h7D][5:4];
        sinkVec_shifterReg_29_0_bits_offset = _RANDOM[8'h7D][8:6];
        sinkVec_shifterReg_29_0_bits_instructionIndex = _RANDOM[8'h7D][11:9];
        maskUnitFirst_14 = _RANDOM[8'h7D][12];
        accessDataValid_pipe_v_14 = _RANDOM[8'h7D][13];
        accessDataValid_pipe_pipe_v_14 = _RANDOM[8'h7D][14];
        shifterReg_22_0_valid = _RANDOM[8'h7D][15];
        shifterReg_22_0_bits = {_RANDOM[8'h7D][31:16], _RANDOM[8'h7E][15:0]};
        accessDataValid_pipe_v_15 = _RANDOM[8'h7E][16];
        accessDataValid_pipe_pipe_v_15 = _RANDOM[8'h7E][17];
        shifterReg_23_0_valid = _RANDOM[8'h7E][18];
        shifterReg_23_0_bits = {_RANDOM[8'h7E][31:19], _RANDOM[8'h7F][18:0]};
        sinkVec_releasePipe_pipe_v_30 = _RANDOM[8'h7F][19];
        sinkVec_tokenCheck_counter_30 = _RANDOM[8'h7F][22:20];
        sinkVec_shifterReg_30_0_valid = _RANDOM[8'h7F][23];
        sinkVec_shifterReg_30_0_bits_vd = _RANDOM[8'h7F][28:24];
        sinkVec_shifterReg_30_0_bits_offset = _RANDOM[8'h7F][31:29];
        sinkVec_shifterReg_30_0_bits_mask = _RANDOM[8'h80][3:0];
        sinkVec_shifterReg_30_0_bits_data = {_RANDOM[8'h80][31:4], _RANDOM[8'h81][3:0]};
        sinkVec_shifterReg_30_0_bits_instructionIndex = _RANDOM[8'h81][7:5];
        sinkVec_releasePipe_pipe_v_31 = _RANDOM[8'h81][8];
        sinkVec_tokenCheck_counter_31 = _RANDOM[8'h81][11:9];
        sinkVec_shifterReg_31_0_valid = _RANDOM[8'h81][12];
        sinkVec_shifterReg_31_0_bits_vd = _RANDOM[8'h81][17:13];
        sinkVec_shifterReg_31_0_bits_offset = _RANDOM[8'h81][20:18];
        sinkVec_shifterReg_31_0_bits_mask = _RANDOM[8'h81][24:21];
        sinkVec_shifterReg_31_0_bits_data = {_RANDOM[8'h81][31:25], _RANDOM[8'h82][24:0]};
        sinkVec_shifterReg_31_0_bits_last = _RANDOM[8'h82][25];
        sinkVec_shifterReg_31_0_bits_instructionIndex = _RANDOM[8'h82][28:26];
        maskUnitFirst_15 = _RANDOM[8'h82][29];
        view__writeRelease_7_pipe_v = _RANDOM[8'h82][30];
        pipe_v_21 = _RANDOM[8'h82][31];
        instructionFinishedPipe_pipe_v_7 = _RANDOM[8'h83][0];
        instructionFinishedPipe_pipe_b_7 = _RANDOM[8'h83][8:1];
        pipe_v_22 = _RANDOM[8'h83][9];
        pipe_b_22 = {_RANDOM[8'h83][31:10], _RANDOM[8'h84][9:0]};
        pipe_pipe_v_7 = _RANDOM[8'h84][10];
        pipe_pipe_b_7 = {_RANDOM[8'h84][31:11], _RANDOM[8'h85][10:0]};
        view__laneMaskSelect_7_pipe_v = _RANDOM[8'h85][11];
        view__laneMaskSelect_7_pipe_b = _RANDOM[8'h85][17:12];
        view__laneMaskSelect_7_pipe_pipe_v = _RANDOM[8'h85][18];
        view__laneMaskSelect_7_pipe_pipe_b = _RANDOM[8'h85][24:19];
        view__laneMaskSewSelect_7_pipe_v = _RANDOM[8'h85][25];
        view__laneMaskSewSelect_7_pipe_b = _RANDOM[8'h85][27:26];
        view__laneMaskSewSelect_7_pipe_pipe_v = _RANDOM[8'h85][28];
        view__laneMaskSewSelect_7_pipe_pipe_b = _RANDOM[8'h85][30:29];
        lsuLastPipe_pipe_v_7 = _RANDOM[8'h85][31];
        lsuLastPipe_pipe_b_7 = _RANDOM[8'h86][7:0];
        maskLastPipe_pipe_v_7 = _RANDOM[8'h86][8];
        maskLastPipe_pipe_b_7 = _RANDOM[8'h86][16:9];
        pipe_v_23 = _RANDOM[8'h86][17];
        pipe_b_23 = _RANDOM[8'h86][24:18];
        pipe_v_24 = _RANDOM[8'h86][25];
        shifterReg_24_0_valid = _RANDOM[8'h86][26];
        shifterReg_24_0_bits_data = {_RANDOM[8'h86][31:27], _RANDOM[8'h87][26:0]};
        pipe_v_25 = _RANDOM[8'h87][27];
        shifterReg_25_0_valid = _RANDOM[8'h87][28];
        shifterReg_25_0_bits_data = {_RANDOM[8'h87][31:29], _RANDOM[8'h88][28:0]};
        shifterReg_25_0_bits_mask = _RANDOM[8'h88][30:29];
        shifterReg_25_0_bits_instructionIndex = {_RANDOM[8'h88][31], _RANDOM[8'h89][1:0]};
        shifterReg_25_0_bits_counter = _RANDOM[8'h89][8:2];
        pipe_v_26 = _RANDOM[8'h89][9];
        shifterReg_26_0_valid = _RANDOM[8'h89][10];
        shifterReg_26_0_bits_data = {_RANDOM[8'h89][31:11], _RANDOM[8'h8A][10:0]};
        pipe_v_27 = _RANDOM[8'h8A][11];
        shifterReg_27_0_valid = _RANDOM[8'h8A][12];
        shifterReg_27_0_bits_data = {_RANDOM[8'h8A][31:13], _RANDOM[8'h8B][12:0]};
        shifterReg_27_0_bits_mask = _RANDOM[8'h8B][14:13];
        shifterReg_27_0_bits_instructionIndex = _RANDOM[8'h8B][17:15];
        shifterReg_27_0_bits_counter = _RANDOM[8'h8B][24:18];
        pipe_v_28 = _RANDOM[8'h8B][25];
        shifterReg_28_0_valid = _RANDOM[8'h8B][26];
        shifterReg_28_0_bits_data = {_RANDOM[8'h8B][31:27], _RANDOM[8'h8C][26:0]};
        pipe_v_29 = _RANDOM[8'h8C][27];
        shifterReg_29_0_valid = _RANDOM[8'h8C][28];
        shifterReg_29_0_bits_data = {_RANDOM[8'h8C][31:29], _RANDOM[8'h8D][28:0]};
        shifterReg_29_0_bits_mask = _RANDOM[8'h8D][30:29];
        shifterReg_29_0_bits_instructionIndex = {_RANDOM[8'h8D][31], _RANDOM[8'h8E][1:0]};
        shifterReg_29_0_bits_counter = _RANDOM[8'h8E][8:2];
        pipe_v_30 = _RANDOM[8'h8E][9];
        shifterReg_30_0_valid = _RANDOM[8'h8E][10];
        shifterReg_30_0_bits_data = {_RANDOM[8'h8E][31:11], _RANDOM[8'h8F][10:0]};
        pipe_v_31 = _RANDOM[8'h8F][11];
        shifterReg_31_0_valid = _RANDOM[8'h8F][12];
        shifterReg_31_0_bits_data = {_RANDOM[8'h8F][31:13], _RANDOM[8'h90][12:0]};
        shifterReg_31_0_bits_mask = _RANDOM[8'h90][14:13];
        shifterReg_31_0_bits_instructionIndex = _RANDOM[8'h90][17:15];
        shifterReg_31_0_bits_counter = _RANDOM[8'h90][24:18];
        pipe_v_32 = _RANDOM[8'h90][25];
        shifterReg_32_0_valid = _RANDOM[8'h90][26];
        shifterReg_32_0_bits_data = {_RANDOM[8'h90][31:27], _RANDOM[8'h91][26:0]};
        pipe_v_33 = _RANDOM[8'h91][27];
        shifterReg_33_0_valid = _RANDOM[8'h91][28];
        shifterReg_33_0_bits_data = {_RANDOM[8'h91][31:29], _RANDOM[8'h92][28:0]};
        shifterReg_33_0_bits_mask = _RANDOM[8'h92][30:29];
        shifterReg_33_0_bits_instructionIndex = {_RANDOM[8'h92][31], _RANDOM[8'h93][1:0]};
        shifterReg_33_0_bits_counter = _RANDOM[8'h93][8:2];
        pipe_v_34 = _RANDOM[8'h93][9];
        shifterReg_34_0_valid = _RANDOM[8'h93][10];
        shifterReg_34_0_bits_data = {_RANDOM[8'h93][31:11], _RANDOM[8'h94][10:0]};
        pipe_v_35 = _RANDOM[8'h94][11];
        shifterReg_35_0_valid = _RANDOM[8'h94][12];
        shifterReg_35_0_bits_data = {_RANDOM[8'h94][31:13], _RANDOM[8'h95][12:0]};
        shifterReg_35_0_bits_mask = _RANDOM[8'h95][14:13];
        shifterReg_35_0_bits_instructionIndex = _RANDOM[8'h95][17:15];
        shifterReg_35_0_bits_counter = _RANDOM[8'h95][24:18];
        pipe_v_36 = _RANDOM[8'h95][25];
        shifterReg_36_0_valid = _RANDOM[8'h95][26];
        shifterReg_36_0_bits_data = {_RANDOM[8'h95][31:27], _RANDOM[8'h96][26:0]};
        pipe_v_37 = _RANDOM[8'h96][27];
        shifterReg_37_0_valid = _RANDOM[8'h96][28];
        shifterReg_37_0_bits_data = {_RANDOM[8'h96][31:29], _RANDOM[8'h97][28:0]};
        shifterReg_37_0_bits_mask = _RANDOM[8'h97][30:29];
        shifterReg_37_0_bits_instructionIndex = {_RANDOM[8'h97][31], _RANDOM[8'h98][1:0]};
        shifterReg_37_0_bits_counter = _RANDOM[8'h98][8:2];
        pipe_v_38 = _RANDOM[8'h98][9];
        shifterReg_38_0_valid = _RANDOM[8'h98][10];
        shifterReg_38_0_bits_data = {_RANDOM[8'h98][31:11], _RANDOM[8'h99][10:0]};
        pipe_v_39 = _RANDOM[8'h99][11];
        shifterReg_39_0_valid = _RANDOM[8'h99][12];
        shifterReg_39_0_bits_data = {_RANDOM[8'h99][31:13], _RANDOM[8'h9A][12:0]};
        shifterReg_39_0_bits_mask = _RANDOM[8'h9A][14:13];
        shifterReg_39_0_bits_instructionIndex = _RANDOM[8'h9A][17:15];
        shifterReg_39_0_bits_counter = _RANDOM[8'h9A][24:18];
        pipe_v_40 = _RANDOM[8'h9A][25];
        shifterReg_40_0_valid = _RANDOM[8'h9A][26];
        shifterReg_40_0_bits_data = {_RANDOM[8'h9A][31:27], _RANDOM[8'h9B][26:0]};
        pipe_v_41 = _RANDOM[8'h9B][27];
        shifterReg_41_0_valid = _RANDOM[8'h9B][28];
        shifterReg_41_0_bits_data = {_RANDOM[8'h9B][31:29], _RANDOM[8'h9C][28:0]};
        shifterReg_41_0_bits_mask = _RANDOM[8'h9C][30:29];
        shifterReg_41_0_bits_instructionIndex = {_RANDOM[8'h9C][31], _RANDOM[8'h9D][1:0]};
        shifterReg_41_0_bits_counter = _RANDOM[8'h9D][8:2];
        pipe_v_42 = _RANDOM[8'h9D][9];
        shifterReg_42_0_valid = _RANDOM[8'h9D][10];
        shifterReg_42_0_bits_data = {_RANDOM[8'h9D][31:11], _RANDOM[8'h9E][10:0]};
        pipe_v_43 = _RANDOM[8'h9E][11];
        shifterReg_43_0_valid = _RANDOM[8'h9E][12];
        shifterReg_43_0_bits_data = {_RANDOM[8'h9E][31:13], _RANDOM[8'h9F][12:0]};
        shifterReg_43_0_bits_mask = _RANDOM[8'h9F][14:13];
        shifterReg_43_0_bits_instructionIndex = _RANDOM[8'h9F][17:15];
        shifterReg_43_0_bits_counter = _RANDOM[8'h9F][24:18];
        pipe_v_44 = _RANDOM[8'h9F][25];
        shifterReg_44_0_valid = _RANDOM[8'h9F][26];
        shifterReg_44_0_bits_data = {_RANDOM[8'h9F][31:27], _RANDOM[8'hA0][26:0]};
        pipe_v_45 = _RANDOM[8'hA0][27];
        shifterReg_45_0_valid = _RANDOM[8'hA0][28];
        shifterReg_45_0_bits_data = {_RANDOM[8'hA0][31:29], _RANDOM[8'hA1][28:0]};
        shifterReg_45_0_bits_mask = _RANDOM[8'hA1][30:29];
        shifterReg_45_0_bits_instructionIndex = {_RANDOM[8'hA1][31], _RANDOM[8'hA2][1:0]};
        shifterReg_45_0_bits_counter = _RANDOM[8'hA2][8:2];
        pipe_v_46 = _RANDOM[8'hA2][9];
        shifterReg_46_0_valid = _RANDOM[8'hA2][10];
        shifterReg_46_0_bits_data = {_RANDOM[8'hA2][31:11], _RANDOM[8'hA3][10:0]};
        pipe_v_47 = _RANDOM[8'hA3][11];
        shifterReg_47_0_valid = _RANDOM[8'hA3][12];
        shifterReg_47_0_bits_data = {_RANDOM[8'hA3][31:13], _RANDOM[8'hA4][12:0]};
        shifterReg_47_0_bits_mask = _RANDOM[8'hA4][14:13];
        shifterReg_47_0_bits_instructionIndex = _RANDOM[8'hA4][17:15];
        shifterReg_47_0_bits_counter = _RANDOM[8'hA4][24:18];
        pipe_v_48 = _RANDOM[8'hA4][25];
        shifterReg_48_0_valid = _RANDOM[8'hA4][26];
        shifterReg_48_0_bits_data = {_RANDOM[8'hA4][31:27], _RANDOM[8'hA5][26:0]};
        pipe_v_49 = _RANDOM[8'hA5][27];
        shifterReg_49_0_valid = _RANDOM[8'hA5][28];
        shifterReg_49_0_bits_data = {_RANDOM[8'hA5][31:29], _RANDOM[8'hA6][28:0]};
        shifterReg_49_0_bits_mask = _RANDOM[8'hA6][30:29];
        shifterReg_49_0_bits_instructionIndex = {_RANDOM[8'hA6][31], _RANDOM[8'hA7][1:0]};
        shifterReg_49_0_bits_counter = _RANDOM[8'hA7][8:2];
        pipe_v_50 = _RANDOM[8'hA7][9];
        shifterReg_50_0_valid = _RANDOM[8'hA7][10];
        shifterReg_50_0_bits_data = {_RANDOM[8'hA7][31:11], _RANDOM[8'hA8][10:0]};
        pipe_v_51 = _RANDOM[8'hA8][11];
        shifterReg_51_0_valid = _RANDOM[8'hA8][12];
        shifterReg_51_0_bits_data = {_RANDOM[8'hA8][31:13], _RANDOM[8'hA9][12:0]};
        shifterReg_51_0_bits_mask = _RANDOM[8'hA9][14:13];
        shifterReg_51_0_bits_instructionIndex = _RANDOM[8'hA9][17:15];
        shifterReg_51_0_bits_counter = _RANDOM[8'hA9][24:18];
        pipe_v_52 = _RANDOM[8'hA9][25];
        shifterReg_52_0_valid = _RANDOM[8'hA9][26];
        shifterReg_52_0_bits_data = {_RANDOM[8'hA9][31:27], _RANDOM[8'hAA][26:0]};
        pipe_v_53 = _RANDOM[8'hAA][27];
        shifterReg_53_0_valid = _RANDOM[8'hAA][28];
        shifterReg_53_0_bits_data = {_RANDOM[8'hAA][31:29], _RANDOM[8'hAB][28:0]};
        shifterReg_53_0_bits_mask = _RANDOM[8'hAB][30:29];
        shifterReg_53_0_bits_instructionIndex = {_RANDOM[8'hAB][31], _RANDOM[8'hAC][1:0]};
        shifterReg_53_0_bits_counter = _RANDOM[8'hAC][8:2];
        pipe_v_54 = _RANDOM[8'hAC][9];
        shifterReg_54_0_valid = _RANDOM[8'hAC][10];
        shifterReg_54_0_bits_data = {_RANDOM[8'hAC][31:11], _RANDOM[8'hAD][10:0]};
        pipe_v_55 = _RANDOM[8'hAD][11];
        shifterReg_55_0_valid = _RANDOM[8'hAD][12];
        shifterReg_55_0_bits_data = {_RANDOM[8'hAD][31:13], _RANDOM[8'hAE][12:0]};
        shifterReg_55_0_bits_mask = _RANDOM[8'hAE][14:13];
        shifterReg_55_0_bits_instructionIndex = _RANDOM[8'hAE][17:15];
        shifterReg_55_0_bits_counter = _RANDOM[8'hAE][24:18];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  assign x22_1_valid = _lsu_vrfWritePort_0_valid;
  assign x22_1_bits_vd = _lsu_vrfWritePort_0_bits_vd;
  assign x22_1_bits_mask = _lsu_vrfWritePort_0_bits_mask;
  assign x22_1_bits_instructionIndex = _lsu_vrfWritePort_0_bits_instructionIndex;
  assign x22_1_1_valid = _lsu_vrfWritePort_1_valid;
  assign x22_1_1_bits_vd = _lsu_vrfWritePort_1_bits_vd;
  assign x22_1_1_bits_mask = _lsu_vrfWritePort_1_bits_mask;
  assign x22_1_1_bits_instructionIndex = _lsu_vrfWritePort_1_bits_instructionIndex;
  assign x22_2_1_valid = _lsu_vrfWritePort_2_valid;
  assign x22_2_1_bits_vd = _lsu_vrfWritePort_2_bits_vd;
  assign x22_2_1_bits_mask = _lsu_vrfWritePort_2_bits_mask;
  assign x22_2_1_bits_instructionIndex = _lsu_vrfWritePort_2_bits_instructionIndex;
  assign x22_3_1_valid = _lsu_vrfWritePort_3_valid;
  assign x22_3_1_bits_vd = _lsu_vrfWritePort_3_bits_vd;
  assign x22_3_1_bits_mask = _lsu_vrfWritePort_3_bits_mask;
  assign x22_3_1_bits_instructionIndex = _lsu_vrfWritePort_3_bits_instructionIndex;
  assign x22_4_1_valid = _lsu_vrfWritePort_4_valid;
  assign x22_4_1_bits_vd = _lsu_vrfWritePort_4_bits_vd;
  assign x22_4_1_bits_mask = _lsu_vrfWritePort_4_bits_mask;
  assign x22_4_1_bits_instructionIndex = _lsu_vrfWritePort_4_bits_instructionIndex;
  assign x22_5_1_valid = _lsu_vrfWritePort_5_valid;
  assign x22_5_1_bits_vd = _lsu_vrfWritePort_5_bits_vd;
  assign x22_5_1_bits_mask = _lsu_vrfWritePort_5_bits_mask;
  assign x22_5_1_bits_instructionIndex = _lsu_vrfWritePort_5_bits_instructionIndex;
  assign x22_6_1_valid = _lsu_vrfWritePort_6_valid;
  assign x22_6_1_bits_vd = _lsu_vrfWritePort_6_bits_vd;
  assign x22_6_1_bits_mask = _lsu_vrfWritePort_6_bits_mask;
  assign x22_6_1_bits_instructionIndex = _lsu_vrfWritePort_6_bits_instructionIndex;
  assign x22_7_1_valid = _lsu_vrfWritePort_7_valid;
  assign x22_7_1_bits_vd = _lsu_vrfWritePort_7_bits_vd;
  assign x22_7_1_bits_mask = _lsu_vrfWritePort_7_bits_mask;
  assign x22_7_1_bits_instructionIndex = _lsu_vrfWritePort_7_bits_instructionIndex;
  assign x22_0_valid = _maskUnit_exeResp_0_valid;
  assign x22_0_bits_mask = _maskUnit_exeResp_0_bits_mask;
  assign x22_0_bits_instructionIndex = _maskUnit_exeResp_0_bits_instructionIndex;
  assign x22_1_0_valid = _maskUnit_exeResp_1_valid;
  assign x22_1_0_bits_mask = _maskUnit_exeResp_1_bits_mask;
  assign x22_1_0_bits_instructionIndex = _maskUnit_exeResp_1_bits_instructionIndex;
  assign x22_2_0_valid = _maskUnit_exeResp_2_valid;
  assign x22_2_0_bits_mask = _maskUnit_exeResp_2_bits_mask;
  assign x22_2_0_bits_instructionIndex = _maskUnit_exeResp_2_bits_instructionIndex;
  assign x22_3_0_valid = _maskUnit_exeResp_3_valid;
  assign x22_3_0_bits_mask = _maskUnit_exeResp_3_bits_mask;
  assign x22_3_0_bits_instructionIndex = _maskUnit_exeResp_3_bits_instructionIndex;
  assign x22_4_0_valid = _maskUnit_exeResp_4_valid;
  assign x22_4_0_bits_mask = _maskUnit_exeResp_4_bits_mask;
  assign x22_4_0_bits_instructionIndex = _maskUnit_exeResp_4_bits_instructionIndex;
  assign x22_5_0_valid = _maskUnit_exeResp_5_valid;
  assign x22_5_0_bits_mask = _maskUnit_exeResp_5_bits_mask;
  assign x22_5_0_bits_instructionIndex = _maskUnit_exeResp_5_bits_instructionIndex;
  assign x22_6_0_valid = _maskUnit_exeResp_6_valid;
  assign x22_6_0_bits_mask = _maskUnit_exeResp_6_bits_mask;
  assign x22_6_0_bits_instructionIndex = _maskUnit_exeResp_6_bits_instructionIndex;
  assign x22_7_0_valid = _maskUnit_exeResp_7_valid;
  assign x22_7_0_bits_mask = _maskUnit_exeResp_7_bits_mask;
  assign x22_7_0_bits_instructionIndex = _maskUnit_exeResp_7_bits_instructionIndex;
  wire         queue_empty;
  assign queue_empty = _queue_fifo_empty;
  wire         queue_full;
  assign queue_full = _queue_fifo_full;
  wire         queue_1_empty;
  assign queue_1_empty = _queue_fifo_1_empty;
  wire         queue_1_full;
  assign queue_1_full = _queue_fifo_1_full;
  wire         queue_2_empty;
  assign queue_2_empty = _queue_fifo_2_empty;
  wire         queue_2_full;
  assign queue_2_full = _queue_fifo_2_full;
  wire         queue_3_empty;
  assign queue_3_empty = _queue_fifo_3_empty;
  wire         queue_3_full;
  assign queue_3_full = _queue_fifo_3_full;
  wire         queue_4_empty;
  assign queue_4_empty = _queue_fifo_4_empty;
  wire         queue_4_full;
  assign queue_4_full = _queue_fifo_4_full;
  wire         queue_5_empty;
  assign queue_5_empty = _queue_fifo_5_empty;
  wire         queue_5_full;
  assign queue_5_full = _queue_fifo_5_full;
  wire         queue_6_empty;
  assign queue_6_empty = _queue_fifo_6_empty;
  wire         queue_6_full;
  assign queue_6_full = _queue_fifo_6_full;
  wire         queue_7_empty;
  assign queue_7_empty = _queue_fifo_7_empty;
  wire         queue_7_full;
  assign queue_7_full = _queue_fifo_7_full;
  assign accessDataSource_bits = _laneVec_0_vrfReadDataChannel;
  assign accessDataSource_1_bits = _laneVec_0_vrfReadDataChannel;
  wire         sinkVec_queue_empty;
  assign sinkVec_queue_empty = _sinkVec_queue_fifo_empty;
  wire         sinkVec_queue_full;
  assign sinkVec_queue_full = _sinkVec_queue_fifo_full;
  wire         sinkVec_queue_1_empty;
  assign sinkVec_queue_1_empty = _sinkVec_queue_fifo_1_empty;
  wire         sinkVec_queue_1_full;
  assign sinkVec_queue_1_full = _sinkVec_queue_fifo_1_full;
  wire         sinkVec_queue_2_empty;
  assign sinkVec_queue_2_empty = _sinkVec_queue_fifo_2_empty;
  wire         sinkVec_queue_2_full;
  assign sinkVec_queue_2_full = _sinkVec_queue_fifo_2_full;
  wire         sinkVec_queue_3_empty;
  assign sinkVec_queue_3_empty = _sinkVec_queue_fifo_3_empty;
  wire         sinkVec_queue_3_full;
  assign sinkVec_queue_3_full = _sinkVec_queue_fifo_3_full;
  assign accessDataSource_2_bits = _laneVec_1_vrfReadDataChannel;
  assign accessDataSource_3_bits = _laneVec_1_vrfReadDataChannel;
  wire         sinkVec_queue_4_empty;
  assign sinkVec_queue_4_empty = _sinkVec_queue_fifo_4_empty;
  wire         sinkVec_queue_4_full;
  assign sinkVec_queue_4_full = _sinkVec_queue_fifo_4_full;
  wire         sinkVec_queue_5_empty;
  assign sinkVec_queue_5_empty = _sinkVec_queue_fifo_5_empty;
  wire         sinkVec_queue_5_full;
  assign sinkVec_queue_5_full = _sinkVec_queue_fifo_5_full;
  wire         sinkVec_queue_6_empty;
  assign sinkVec_queue_6_empty = _sinkVec_queue_fifo_6_empty;
  wire         sinkVec_queue_6_full;
  assign sinkVec_queue_6_full = _sinkVec_queue_fifo_6_full;
  wire         sinkVec_queue_7_empty;
  assign sinkVec_queue_7_empty = _sinkVec_queue_fifo_7_empty;
  wire         sinkVec_queue_7_full;
  assign sinkVec_queue_7_full = _sinkVec_queue_fifo_7_full;
  assign accessDataSource_4_bits = _laneVec_2_vrfReadDataChannel;
  assign accessDataSource_5_bits = _laneVec_2_vrfReadDataChannel;
  wire         sinkVec_queue_8_empty;
  assign sinkVec_queue_8_empty = _sinkVec_queue_fifo_8_empty;
  wire         sinkVec_queue_8_full;
  assign sinkVec_queue_8_full = _sinkVec_queue_fifo_8_full;
  wire         sinkVec_queue_9_empty;
  assign sinkVec_queue_9_empty = _sinkVec_queue_fifo_9_empty;
  wire         sinkVec_queue_9_full;
  assign sinkVec_queue_9_full = _sinkVec_queue_fifo_9_full;
  wire         sinkVec_queue_10_empty;
  assign sinkVec_queue_10_empty = _sinkVec_queue_fifo_10_empty;
  wire         sinkVec_queue_10_full;
  assign sinkVec_queue_10_full = _sinkVec_queue_fifo_10_full;
  wire         sinkVec_queue_11_empty;
  assign sinkVec_queue_11_empty = _sinkVec_queue_fifo_11_empty;
  wire         sinkVec_queue_11_full;
  assign sinkVec_queue_11_full = _sinkVec_queue_fifo_11_full;
  assign accessDataSource_6_bits = _laneVec_3_vrfReadDataChannel;
  assign accessDataSource_7_bits = _laneVec_3_vrfReadDataChannel;
  wire         sinkVec_queue_12_empty;
  assign sinkVec_queue_12_empty = _sinkVec_queue_fifo_12_empty;
  wire         sinkVec_queue_12_full;
  assign sinkVec_queue_12_full = _sinkVec_queue_fifo_12_full;
  wire         sinkVec_queue_13_empty;
  assign sinkVec_queue_13_empty = _sinkVec_queue_fifo_13_empty;
  wire         sinkVec_queue_13_full;
  assign sinkVec_queue_13_full = _sinkVec_queue_fifo_13_full;
  wire         sinkVec_queue_14_empty;
  assign sinkVec_queue_14_empty = _sinkVec_queue_fifo_14_empty;
  wire         sinkVec_queue_14_full;
  assign sinkVec_queue_14_full = _sinkVec_queue_fifo_14_full;
  wire         sinkVec_queue_15_empty;
  assign sinkVec_queue_15_empty = _sinkVec_queue_fifo_15_empty;
  wire         sinkVec_queue_15_full;
  assign sinkVec_queue_15_full = _sinkVec_queue_fifo_15_full;
  assign accessDataSource_8_bits = _laneVec_4_vrfReadDataChannel;
  assign accessDataSource_9_bits = _laneVec_4_vrfReadDataChannel;
  wire         sinkVec_queue_16_empty;
  assign sinkVec_queue_16_empty = _sinkVec_queue_fifo_16_empty;
  wire         sinkVec_queue_16_full;
  assign sinkVec_queue_16_full = _sinkVec_queue_fifo_16_full;
  wire         sinkVec_queue_17_empty;
  assign sinkVec_queue_17_empty = _sinkVec_queue_fifo_17_empty;
  wire         sinkVec_queue_17_full;
  assign sinkVec_queue_17_full = _sinkVec_queue_fifo_17_full;
  wire         sinkVec_queue_18_empty;
  assign sinkVec_queue_18_empty = _sinkVec_queue_fifo_18_empty;
  wire         sinkVec_queue_18_full;
  assign sinkVec_queue_18_full = _sinkVec_queue_fifo_18_full;
  wire         sinkVec_queue_19_empty;
  assign sinkVec_queue_19_empty = _sinkVec_queue_fifo_19_empty;
  wire         sinkVec_queue_19_full;
  assign sinkVec_queue_19_full = _sinkVec_queue_fifo_19_full;
  assign accessDataSource_10_bits = _laneVec_5_vrfReadDataChannel;
  assign accessDataSource_11_bits = _laneVec_5_vrfReadDataChannel;
  wire         sinkVec_queue_20_empty;
  assign sinkVec_queue_20_empty = _sinkVec_queue_fifo_20_empty;
  wire         sinkVec_queue_20_full;
  assign sinkVec_queue_20_full = _sinkVec_queue_fifo_20_full;
  wire         sinkVec_queue_21_empty;
  assign sinkVec_queue_21_empty = _sinkVec_queue_fifo_21_empty;
  wire         sinkVec_queue_21_full;
  assign sinkVec_queue_21_full = _sinkVec_queue_fifo_21_full;
  wire         sinkVec_queue_22_empty;
  assign sinkVec_queue_22_empty = _sinkVec_queue_fifo_22_empty;
  wire         sinkVec_queue_22_full;
  assign sinkVec_queue_22_full = _sinkVec_queue_fifo_22_full;
  wire         sinkVec_queue_23_empty;
  assign sinkVec_queue_23_empty = _sinkVec_queue_fifo_23_empty;
  wire         sinkVec_queue_23_full;
  assign sinkVec_queue_23_full = _sinkVec_queue_fifo_23_full;
  assign accessDataSource_12_bits = _laneVec_6_vrfReadDataChannel;
  assign accessDataSource_13_bits = _laneVec_6_vrfReadDataChannel;
  wire         sinkVec_queue_24_empty;
  assign sinkVec_queue_24_empty = _sinkVec_queue_fifo_24_empty;
  wire         sinkVec_queue_24_full;
  assign sinkVec_queue_24_full = _sinkVec_queue_fifo_24_full;
  wire         sinkVec_queue_25_empty;
  assign sinkVec_queue_25_empty = _sinkVec_queue_fifo_25_empty;
  wire         sinkVec_queue_25_full;
  assign sinkVec_queue_25_full = _sinkVec_queue_fifo_25_full;
  wire         sinkVec_queue_26_empty;
  assign sinkVec_queue_26_empty = _sinkVec_queue_fifo_26_empty;
  wire         sinkVec_queue_26_full;
  assign sinkVec_queue_26_full = _sinkVec_queue_fifo_26_full;
  wire         sinkVec_queue_27_empty;
  assign sinkVec_queue_27_empty = _sinkVec_queue_fifo_27_empty;
  wire         sinkVec_queue_27_full;
  assign sinkVec_queue_27_full = _sinkVec_queue_fifo_27_full;
  assign accessDataSource_14_bits = _laneVec_7_vrfReadDataChannel;
  assign accessDataSource_15_bits = _laneVec_7_vrfReadDataChannel;
  wire         sinkVec_queue_28_empty;
  assign sinkVec_queue_28_empty = _sinkVec_queue_fifo_28_empty;
  wire         sinkVec_queue_28_full;
  assign sinkVec_queue_28_full = _sinkVec_queue_fifo_28_full;
  wire         sinkVec_queue_29_empty;
  assign sinkVec_queue_29_empty = _sinkVec_queue_fifo_29_empty;
  wire         sinkVec_queue_29_full;
  assign sinkVec_queue_29_full = _sinkVec_queue_fifo_29_full;
  wire         sinkVec_queue_30_empty;
  assign sinkVec_queue_30_empty = _sinkVec_queue_fifo_30_empty;
  wire         sinkVec_queue_30_full;
  assign sinkVec_queue_30_full = _sinkVec_queue_fifo_30_full;
  wire         sinkVec_queue_31_empty;
  assign sinkVec_queue_31_empty = _sinkVec_queue_fifo_31_empty;
  wire         sinkVec_queue_31_full;
  assign sinkVec_queue_31_full = _sinkVec_queue_fifo_31_full;
  LSU lsu (
    .clock                                               (clock),
    .reset                                               (reset),
    .request_ready                                       (_lsu_request_ready),
    .request_valid                                       (maskUnit_gatherData_ready & isLoadStoreType),
    .request_bits_instructionInformation_nf              (requestRegDequeue_bits_instruction[31:29]),
    .request_bits_instructionInformation_mew             (requestRegDequeue_bits_instruction[28]),
    .request_bits_instructionInformation_mop             (requestRegDequeue_bits_instruction[27:26]),
    .request_bits_instructionInformation_lumop           (requestRegDequeue_bits_instruction[24:20]),
    .request_bits_instructionInformation_eew             (vSewForLsu),
    .request_bits_instructionInformation_vs3             (requestRegDequeue_bits_instruction[11:7]),
    .request_bits_instructionInformation_isStore         (isStoreType),
    .request_bits_instructionInformation_maskedLoadStore (maskType),
    .request_bits_rs1Data                                (requestRegDequeue_bits_rs1Data),
    .request_bits_rs2Data                                (requestRegDequeue_bits_rs2Data),
    .request_bits_instructionIndex                       (requestReg_bits_instructionIndex),
    .v0UpdateVec_0_valid                                 (_laneVec_0_v0Update_valid),
    .v0UpdateVec_0_bits_data                             (_laneVec_0_v0Update_bits_data),
    .v0UpdateVec_0_bits_offset                           (_laneVec_0_v0Update_bits_offset),
    .v0UpdateVec_0_bits_mask                             (_laneVec_0_v0Update_bits_mask),
    .v0UpdateVec_1_valid                                 (_laneVec_1_v0Update_valid),
    .v0UpdateVec_1_bits_data                             (_laneVec_1_v0Update_bits_data),
    .v0UpdateVec_1_bits_offset                           (_laneVec_1_v0Update_bits_offset),
    .v0UpdateVec_1_bits_mask                             (_laneVec_1_v0Update_bits_mask),
    .v0UpdateVec_2_valid                                 (_laneVec_2_v0Update_valid),
    .v0UpdateVec_2_bits_data                             (_laneVec_2_v0Update_bits_data),
    .v0UpdateVec_2_bits_offset                           (_laneVec_2_v0Update_bits_offset),
    .v0UpdateVec_2_bits_mask                             (_laneVec_2_v0Update_bits_mask),
    .v0UpdateVec_3_valid                                 (_laneVec_3_v0Update_valid),
    .v0UpdateVec_3_bits_data                             (_laneVec_3_v0Update_bits_data),
    .v0UpdateVec_3_bits_offset                           (_laneVec_3_v0Update_bits_offset),
    .v0UpdateVec_3_bits_mask                             (_laneVec_3_v0Update_bits_mask),
    .v0UpdateVec_4_valid                                 (_laneVec_4_v0Update_valid),
    .v0UpdateVec_4_bits_data                             (_laneVec_4_v0Update_bits_data),
    .v0UpdateVec_4_bits_offset                           (_laneVec_4_v0Update_bits_offset),
    .v0UpdateVec_4_bits_mask                             (_laneVec_4_v0Update_bits_mask),
    .v0UpdateVec_5_valid                                 (_laneVec_5_v0Update_valid),
    .v0UpdateVec_5_bits_data                             (_laneVec_5_v0Update_bits_data),
    .v0UpdateVec_5_bits_offset                           (_laneVec_5_v0Update_bits_offset),
    .v0UpdateVec_5_bits_mask                             (_laneVec_5_v0Update_bits_mask),
    .v0UpdateVec_6_valid                                 (_laneVec_6_v0Update_valid),
    .v0UpdateVec_6_bits_data                             (_laneVec_6_v0Update_bits_data),
    .v0UpdateVec_6_bits_offset                           (_laneVec_6_v0Update_bits_offset),
    .v0UpdateVec_6_bits_mask                             (_laneVec_6_v0Update_bits_mask),
    .v0UpdateVec_7_valid                                 (_laneVec_7_v0Update_valid),
    .v0UpdateVec_7_bits_data                             (_laneVec_7_v0Update_bits_data),
    .v0UpdateVec_7_bits_offset                           (_laneVec_7_v0Update_bits_offset),
    .v0UpdateVec_7_bits_mask                             (_laneVec_7_v0Update_bits_mask),
    .axi4Port_aw_ready                                   (highBandwidthLoadStorePort_aw_ready_0),
    .axi4Port_aw_valid                                   (highBandwidthLoadStorePort_aw_valid_0),
    .axi4Port_aw_bits_id                                 (highBandwidthLoadStorePort_aw_bits_id_0),
    .axi4Port_aw_bits_addr                               (highBandwidthLoadStorePort_aw_bits_addr_0),
    .axi4Port_w_ready                                    (highBandwidthLoadStorePort_w_ready_0),
    .axi4Port_w_valid                                    (highBandwidthLoadStorePort_w_valid_0),
    .axi4Port_w_bits_data                                (highBandwidthLoadStorePort_w_bits_data_0),
    .axi4Port_w_bits_strb                                (highBandwidthLoadStorePort_w_bits_strb_0),
    .axi4Port_b_valid                                    (highBandwidthLoadStorePort_b_valid_0),
    .axi4Port_b_bits_id                                  (highBandwidthLoadStorePort_b_bits_id_0),
    .axi4Port_b_bits_resp                                (highBandwidthLoadStorePort_b_bits_resp_0),
    .axi4Port_ar_ready                                   (highBandwidthLoadStorePort_ar_ready_0),
    .axi4Port_ar_valid                                   (highBandwidthLoadStorePort_ar_valid_0),
    .axi4Port_ar_bits_addr                               (highBandwidthLoadStorePort_ar_bits_addr_0),
    .axi4Port_r_ready                                    (highBandwidthLoadStorePort_r_ready_0),
    .axi4Port_r_valid                                    (highBandwidthLoadStorePort_r_valid_0),
    .axi4Port_r_bits_id                                  (highBandwidthLoadStorePort_r_bits_id_0),
    .axi4Port_r_bits_data                                (highBandwidthLoadStorePort_r_bits_data_0),
    .axi4Port_r_bits_resp                                (highBandwidthLoadStorePort_r_bits_resp_0),
    .axi4Port_r_bits_last                                (highBandwidthLoadStorePort_r_bits_last_0),
    .simpleAccessPorts_aw_ready                          (indexedLoadStorePort_aw_ready_0),
    .simpleAccessPorts_aw_valid                          (indexedLoadStorePort_aw_valid_0),
    .simpleAccessPorts_aw_bits_id                        (indexedLoadStorePort_aw_bits_id_0),
    .simpleAccessPorts_aw_bits_addr                      (indexedLoadStorePort_aw_bits_addr_0),
    .simpleAccessPorts_aw_bits_size                      (indexedLoadStorePort_aw_bits_size_0),
    .simpleAccessPorts_w_ready                           (indexedLoadStorePort_w_ready_0),
    .simpleAccessPorts_w_valid                           (indexedLoadStorePort_w_valid_0),
    .simpleAccessPorts_w_bits_data                       (indexedLoadStorePort_w_bits_data_0),
    .simpleAccessPorts_w_bits_strb                       (indexedLoadStorePort_w_bits_strb_0),
    .simpleAccessPorts_b_valid                           (indexedLoadStorePort_b_valid_0),
    .simpleAccessPorts_b_bits_id                         (indexedLoadStorePort_b_bits_id_0),
    .simpleAccessPorts_b_bits_resp                       (indexedLoadStorePort_b_bits_resp_0),
    .simpleAccessPorts_ar_ready                          (indexedLoadStorePort_ar_ready_0),
    .simpleAccessPorts_ar_valid                          (indexedLoadStorePort_ar_valid_0),
    .simpleAccessPorts_ar_bits_addr                      (indexedLoadStorePort_ar_bits_addr_0),
    .simpleAccessPorts_r_ready                           (indexedLoadStorePort_r_ready_0),
    .simpleAccessPorts_r_valid                           (indexedLoadStorePort_r_valid_0),
    .simpleAccessPorts_r_bits_id                         (indexedLoadStorePort_r_bits_id_0),
    .simpleAccessPorts_r_bits_data                       (indexedLoadStorePort_r_bits_data_0),
    .simpleAccessPorts_r_bits_resp                       (indexedLoadStorePort_r_bits_resp_0),
    .simpleAccessPorts_r_bits_last                       (indexedLoadStorePort_r_bits_last_0),
    .vrfReadDataPorts_0_ready                            (x13_1_ready),
    .vrfReadDataPorts_0_valid                            (x13_1_valid),
    .vrfReadDataPorts_0_bits_vs                          (x13_1_bits_vs),
    .vrfReadDataPorts_0_bits_offset                      (x13_1_bits_offset),
    .vrfReadDataPorts_0_bits_instructionIndex            (x13_1_bits_instructionIndex),
    .vrfReadDataPorts_1_ready                            (x13_1_1_ready),
    .vrfReadDataPorts_1_valid                            (x13_1_1_valid),
    .vrfReadDataPorts_1_bits_vs                          (x13_1_1_bits_vs),
    .vrfReadDataPorts_1_bits_offset                      (x13_1_1_bits_offset),
    .vrfReadDataPorts_1_bits_instructionIndex            (x13_1_1_bits_instructionIndex),
    .vrfReadDataPorts_2_ready                            (x13_2_1_ready),
    .vrfReadDataPorts_2_valid                            (x13_2_1_valid),
    .vrfReadDataPorts_2_bits_vs                          (x13_2_1_bits_vs),
    .vrfReadDataPorts_2_bits_offset                      (x13_2_1_bits_offset),
    .vrfReadDataPorts_2_bits_instructionIndex            (x13_2_1_bits_instructionIndex),
    .vrfReadDataPorts_3_ready                            (x13_3_1_ready),
    .vrfReadDataPorts_3_valid                            (x13_3_1_valid),
    .vrfReadDataPorts_3_bits_vs                          (x13_3_1_bits_vs),
    .vrfReadDataPorts_3_bits_offset                      (x13_3_1_bits_offset),
    .vrfReadDataPorts_3_bits_instructionIndex            (x13_3_1_bits_instructionIndex),
    .vrfReadDataPorts_4_ready                            (x13_4_1_ready),
    .vrfReadDataPorts_4_valid                            (x13_4_1_valid),
    .vrfReadDataPorts_4_bits_vs                          (x13_4_1_bits_vs),
    .vrfReadDataPorts_4_bits_offset                      (x13_4_1_bits_offset),
    .vrfReadDataPorts_4_bits_instructionIndex            (x13_4_1_bits_instructionIndex),
    .vrfReadDataPorts_5_ready                            (x13_5_1_ready),
    .vrfReadDataPorts_5_valid                            (x13_5_1_valid),
    .vrfReadDataPorts_5_bits_vs                          (x13_5_1_bits_vs),
    .vrfReadDataPorts_5_bits_offset                      (x13_5_1_bits_offset),
    .vrfReadDataPorts_5_bits_instructionIndex            (x13_5_1_bits_instructionIndex),
    .vrfReadDataPorts_6_ready                            (x13_6_1_ready),
    .vrfReadDataPorts_6_valid                            (x13_6_1_valid),
    .vrfReadDataPorts_6_bits_vs                          (x13_6_1_bits_vs),
    .vrfReadDataPorts_6_bits_offset                      (x13_6_1_bits_offset),
    .vrfReadDataPorts_6_bits_instructionIndex            (x13_6_1_bits_instructionIndex),
    .vrfReadDataPorts_7_ready                            (x13_7_1_ready),
    .vrfReadDataPorts_7_valid                            (x13_7_1_valid),
    .vrfReadDataPorts_7_bits_vs                          (x13_7_1_bits_vs),
    .vrfReadDataPorts_7_bits_offset                      (x13_7_1_bits_offset),
    .vrfReadDataPorts_7_bits_instructionIndex            (x13_7_1_bits_instructionIndex),
    .vrfReadResults_0_valid                              (shifterReg_9_0_valid),
    .vrfReadResults_0_bits                               (shifterReg_9_0_bits),
    .vrfReadResults_1_valid                              (shifterReg_11_0_valid),
    .vrfReadResults_1_bits                               (shifterReg_11_0_bits),
    .vrfReadResults_2_valid                              (shifterReg_13_0_valid),
    .vrfReadResults_2_bits                               (shifterReg_13_0_bits),
    .vrfReadResults_3_valid                              (shifterReg_15_0_valid),
    .vrfReadResults_3_bits                               (shifterReg_15_0_bits),
    .vrfReadResults_4_valid                              (shifterReg_17_0_valid),
    .vrfReadResults_4_bits                               (shifterReg_17_0_bits),
    .vrfReadResults_5_valid                              (shifterReg_19_0_valid),
    .vrfReadResults_5_bits                               (shifterReg_19_0_bits),
    .vrfReadResults_6_valid                              (shifterReg_21_0_valid),
    .vrfReadResults_6_bits                               (shifterReg_21_0_bits),
    .vrfReadResults_7_valid                              (shifterReg_23_0_valid),
    .vrfReadResults_7_bits                               (shifterReg_23_0_bits),
    .vrfWritePort_0_ready                                (x22_1_ready),
    .vrfWritePort_0_valid                                (_lsu_vrfWritePort_0_valid),
    .vrfWritePort_0_bits_vd                              (_lsu_vrfWritePort_0_bits_vd),
    .vrfWritePort_0_bits_offset                          (x22_1_bits_offset),
    .vrfWritePort_0_bits_mask                            (_lsu_vrfWritePort_0_bits_mask),
    .vrfWritePort_0_bits_data                            (x22_1_bits_data),
    .vrfWritePort_0_bits_last                            (x22_1_bits_last),
    .vrfWritePort_0_bits_instructionIndex                (_lsu_vrfWritePort_0_bits_instructionIndex),
    .vrfWritePort_1_ready                                (x22_1_1_ready),
    .vrfWritePort_1_valid                                (_lsu_vrfWritePort_1_valid),
    .vrfWritePort_1_bits_vd                              (_lsu_vrfWritePort_1_bits_vd),
    .vrfWritePort_1_bits_offset                          (x22_1_1_bits_offset),
    .vrfWritePort_1_bits_mask                            (_lsu_vrfWritePort_1_bits_mask),
    .vrfWritePort_1_bits_data                            (x22_1_1_bits_data),
    .vrfWritePort_1_bits_last                            (x22_1_1_bits_last),
    .vrfWritePort_1_bits_instructionIndex                (_lsu_vrfWritePort_1_bits_instructionIndex),
    .vrfWritePort_2_ready                                (x22_2_1_ready),
    .vrfWritePort_2_valid                                (_lsu_vrfWritePort_2_valid),
    .vrfWritePort_2_bits_vd                              (_lsu_vrfWritePort_2_bits_vd),
    .vrfWritePort_2_bits_offset                          (x22_2_1_bits_offset),
    .vrfWritePort_2_bits_mask                            (_lsu_vrfWritePort_2_bits_mask),
    .vrfWritePort_2_bits_data                            (x22_2_1_bits_data),
    .vrfWritePort_2_bits_last                            (x22_2_1_bits_last),
    .vrfWritePort_2_bits_instructionIndex                (_lsu_vrfWritePort_2_bits_instructionIndex),
    .vrfWritePort_3_ready                                (x22_3_1_ready),
    .vrfWritePort_3_valid                                (_lsu_vrfWritePort_3_valid),
    .vrfWritePort_3_bits_vd                              (_lsu_vrfWritePort_3_bits_vd),
    .vrfWritePort_3_bits_offset                          (x22_3_1_bits_offset),
    .vrfWritePort_3_bits_mask                            (_lsu_vrfWritePort_3_bits_mask),
    .vrfWritePort_3_bits_data                            (x22_3_1_bits_data),
    .vrfWritePort_3_bits_last                            (x22_3_1_bits_last),
    .vrfWritePort_3_bits_instructionIndex                (_lsu_vrfWritePort_3_bits_instructionIndex),
    .vrfWritePort_4_ready                                (x22_4_1_ready),
    .vrfWritePort_4_valid                                (_lsu_vrfWritePort_4_valid),
    .vrfWritePort_4_bits_vd                              (_lsu_vrfWritePort_4_bits_vd),
    .vrfWritePort_4_bits_offset                          (x22_4_1_bits_offset),
    .vrfWritePort_4_bits_mask                            (_lsu_vrfWritePort_4_bits_mask),
    .vrfWritePort_4_bits_data                            (x22_4_1_bits_data),
    .vrfWritePort_4_bits_last                            (x22_4_1_bits_last),
    .vrfWritePort_4_bits_instructionIndex                (_lsu_vrfWritePort_4_bits_instructionIndex),
    .vrfWritePort_5_ready                                (x22_5_1_ready),
    .vrfWritePort_5_valid                                (_lsu_vrfWritePort_5_valid),
    .vrfWritePort_5_bits_vd                              (_lsu_vrfWritePort_5_bits_vd),
    .vrfWritePort_5_bits_offset                          (x22_5_1_bits_offset),
    .vrfWritePort_5_bits_mask                            (_lsu_vrfWritePort_5_bits_mask),
    .vrfWritePort_5_bits_data                            (x22_5_1_bits_data),
    .vrfWritePort_5_bits_last                            (x22_5_1_bits_last),
    .vrfWritePort_5_bits_instructionIndex                (_lsu_vrfWritePort_5_bits_instructionIndex),
    .vrfWritePort_6_ready                                (x22_6_1_ready),
    .vrfWritePort_6_valid                                (_lsu_vrfWritePort_6_valid),
    .vrfWritePort_6_bits_vd                              (_lsu_vrfWritePort_6_bits_vd),
    .vrfWritePort_6_bits_offset                          (x22_6_1_bits_offset),
    .vrfWritePort_6_bits_mask                            (_lsu_vrfWritePort_6_bits_mask),
    .vrfWritePort_6_bits_data                            (x22_6_1_bits_data),
    .vrfWritePort_6_bits_last                            (x22_6_1_bits_last),
    .vrfWritePort_6_bits_instructionIndex                (_lsu_vrfWritePort_6_bits_instructionIndex),
    .vrfWritePort_7_ready                                (x22_7_1_ready),
    .vrfWritePort_7_valid                                (_lsu_vrfWritePort_7_valid),
    .vrfWritePort_7_bits_vd                              (_lsu_vrfWritePort_7_bits_vd),
    .vrfWritePort_7_bits_offset                          (x22_7_1_bits_offset),
    .vrfWritePort_7_bits_mask                            (_lsu_vrfWritePort_7_bits_mask),
    .vrfWritePort_7_bits_data                            (x22_7_1_bits_data),
    .vrfWritePort_7_bits_last                            (x22_7_1_bits_last),
    .vrfWritePort_7_bits_instructionIndex                (_lsu_vrfWritePort_7_bits_instructionIndex),
    .writeRelease_0                                      (pipe_out_valid),
    .writeRelease_1                                      (pipe_out_2_valid),
    .writeRelease_2                                      (pipe_out_4_valid),
    .writeRelease_3                                      (pipe_out_6_valid),
    .writeRelease_4                                      (pipe_out_8_valid),
    .writeRelease_5                                      (pipe_out_10_valid),
    .writeRelease_6                                      (pipe_out_12_valid),
    .writeRelease_7                                      (pipe_out_14_valid),
    .dataInWriteQueue_0                                  (_lsu_dataInWriteQueue_0),
    .dataInWriteQueue_1                                  (_lsu_dataInWriteQueue_1),
    .dataInWriteQueue_2                                  (_lsu_dataInWriteQueue_2),
    .dataInWriteQueue_3                                  (_lsu_dataInWriteQueue_3),
    .dataInWriteQueue_4                                  (_lsu_dataInWriteQueue_4),
    .dataInWriteQueue_5                                  (_lsu_dataInWriteQueue_5),
    .dataInWriteQueue_6                                  (_lsu_dataInWriteQueue_6),
    .dataInWriteQueue_7                                  (_lsu_dataInWriteQueue_7),
    .csrInterface_vl                                     (evlForLsu[11:0]),
    .csrInterface_vStart                                 (requestRegCSR_vStart),
    .csrInterface_vlmul                                  (requestRegCSR_vlmul),
    .csrInterface_vSew                                   (requestRegCSR_vSew),
    .csrInterface_vxrm                                   (requestRegCSR_vxrm),
    .csrInterface_vta                                    (requestRegCSR_vta),
    .csrInterface_vma                                    (requestRegCSR_vma),
    .offsetReadResult_0_valid                            (_laneVec_0_maskUnitRequest_valid & _laneVec_0_maskRequestToLSU),
    .offsetReadResult_0_bits                             (_laneVec_0_maskUnitRequest_bits_source2),
    .offsetReadResult_1_valid                            (_laneVec_1_maskUnitRequest_valid & _laneVec_1_maskRequestToLSU),
    .offsetReadResult_1_bits                             (_laneVec_1_maskUnitRequest_bits_source2),
    .offsetReadResult_2_valid                            (_laneVec_2_maskUnitRequest_valid & _laneVec_2_maskRequestToLSU),
    .offsetReadResult_2_bits                             (_laneVec_2_maskUnitRequest_bits_source2),
    .offsetReadResult_3_valid                            (_laneVec_3_maskUnitRequest_valid & _laneVec_3_maskRequestToLSU),
    .offsetReadResult_3_bits                             (_laneVec_3_maskUnitRequest_bits_source2),
    .offsetReadResult_4_valid                            (_laneVec_4_maskUnitRequest_valid & _laneVec_4_maskRequestToLSU),
    .offsetReadResult_4_bits                             (_laneVec_4_maskUnitRequest_bits_source2),
    .offsetReadResult_5_valid                            (_laneVec_5_maskUnitRequest_valid & _laneVec_5_maskRequestToLSU),
    .offsetReadResult_5_bits                             (_laneVec_5_maskUnitRequest_bits_source2),
    .offsetReadResult_6_valid                            (_laneVec_6_maskUnitRequest_valid & _laneVec_6_maskRequestToLSU),
    .offsetReadResult_6_bits                             (_laneVec_6_maskUnitRequest_bits_source2),
    .offsetReadResult_7_valid                            (_laneVec_7_maskUnitRequest_valid & _laneVec_7_maskRequestToLSU),
    .offsetReadResult_7_bits                             (_laneVec_7_maskUnitRequest_bits_source2),
    .lastReport                                          (_lsu_lastReport),
    .tokenIO_offsetGroupRelease                          (_lsu_tokenIO_offsetGroupRelease)
  );
  VectorDecoder decode (
    .decodeInput                        (issue_bits_instruction_0),
    .decodeResult_specialSlot           (_decode_decodeResult_specialSlot),
    .decodeResult_topUop                (_decode_decodeResult_topUop),
    .decodeResult_popCount              (_decode_decodeResult_popCount),
    .decodeResult_ffo                   (_decode_decodeResult_ffo),
    .decodeResult_average               (_decode_decodeResult_average),
    .decodeResult_reverse               (_decode_decodeResult_reverse),
    .decodeResult_dontNeedExecuteInLane (_decode_decodeResult_dontNeedExecuteInLane),
    .decodeResult_scheduler             (_decode_decodeResult_scheduler),
    .decodeResult_sReadVD               (_decode_decodeResult_sReadVD),
    .decodeResult_vtype                 (_decode_decodeResult_vtype),
    .decodeResult_sWrite                (_decode_decodeResult_sWrite),
    .decodeResult_crossRead             (_decode_decodeResult_crossRead),
    .decodeResult_crossWrite            (_decode_decodeResult_crossWrite),
    .decodeResult_maskUnit              (_decode_decodeResult_maskUnit),
    .decodeResult_special               (_decode_decodeResult_special),
    .decodeResult_saturate              (_decode_decodeResult_saturate),
    .decodeResult_vwmacc                (_decode_decodeResult_vwmacc),
    .decodeResult_readOnly              (_decode_decodeResult_readOnly),
    .decodeResult_maskSource            (_decode_decodeResult_maskSource),
    .decodeResult_maskDestination       (_decode_decodeResult_maskDestination),
    .decodeResult_maskLogic             (_decode_decodeResult_maskLogic),
    .decodeResult_uop                   (_decode_decodeResult_uop),
    .decodeResult_iota                  (_decode_decodeResult_iota),
    .decodeResult_mv                    (_decode_decodeResult_mv),
    .decodeResult_extend                (_decode_decodeResult_extend),
    .decodeResult_unOrderWrite          (_decode_decodeResult_unOrderWrite),
    .decodeResult_compress              (_decode_decodeResult_compress),
    .decodeResult_gather16              (_decode_decodeResult_gather16),
    .decodeResult_gather                (_decode_decodeResult_gather),
    .decodeResult_slid                  (_decode_decodeResult_slid),
    .decodeResult_targetRd              (_decode_decodeResult_targetRd),
    .decodeResult_widenReduce           (_decode_decodeResult_widenReduce),
    .decodeResult_red                   (_decode_decodeResult_red),
    .decodeResult_nr                    (_decode_decodeResult_nr),
    .decodeResult_itype                 (_decode_decodeResult_itype),
    .decodeResult_unsigned1             (_decode_decodeResult_unsigned1),
    .decodeResult_unsigned0             (_decode_decodeResult_unsigned0),
    .decodeResult_other                 (_decode_decodeResult_other),
    .decodeResult_multiCycle            (_decode_decodeResult_multiCycle),
    .decodeResult_divider               (_decode_decodeResult_divider),
    .decodeResult_multiplier            (_decode_decodeResult_multiplier),
    .decodeResult_shift                 (_decode_decodeResult_shift),
    .decodeResult_adder                 (_decode_decodeResult_adder),
    .decodeResult_logic                 (_decode_decodeResult_logic)
  );
  MaskUnit maskUnit (
    .clock                                           (clock),
    .reset                                           (reset),
    .instReq_valid                                   (maskUnit_gatherData_ready & requestReg_bits_decodeResult_maskUnit),
    .instReq_bits_instructionIndex                   (requestReg_bits_instructionIndex),
    .instReq_bits_decodeResult_specialSlot           (requestReg_bits_decodeResult_specialSlot),
    .instReq_bits_decodeResult_topUop                (requestReg_bits_decodeResult_topUop),
    .instReq_bits_decodeResult_popCount              (requestReg_bits_decodeResult_popCount),
    .instReq_bits_decodeResult_ffo                   (requestReg_bits_decodeResult_ffo),
    .instReq_bits_decodeResult_average               (requestReg_bits_decodeResult_average),
    .instReq_bits_decodeResult_reverse               (requestReg_bits_decodeResult_reverse),
    .instReq_bits_decodeResult_dontNeedExecuteInLane (requestReg_bits_decodeResult_dontNeedExecuteInLane),
    .instReq_bits_decodeResult_scheduler             (requestReg_bits_decodeResult_scheduler),
    .instReq_bits_decodeResult_sReadVD               (requestReg_bits_decodeResult_sReadVD),
    .instReq_bits_decodeResult_vtype                 (requestReg_bits_decodeResult_vtype),
    .instReq_bits_decodeResult_sWrite                (requestReg_bits_decodeResult_sWrite),
    .instReq_bits_decodeResult_crossRead             (requestReg_bits_decodeResult_crossRead),
    .instReq_bits_decodeResult_crossWrite            (requestReg_bits_decodeResult_crossWrite),
    .instReq_bits_decodeResult_maskUnit              (requestReg_bits_decodeResult_maskUnit),
    .instReq_bits_decodeResult_special               (requestReg_bits_decodeResult_special),
    .instReq_bits_decodeResult_saturate              (requestReg_bits_decodeResult_saturate),
    .instReq_bits_decodeResult_vwmacc                (requestReg_bits_decodeResult_vwmacc),
    .instReq_bits_decodeResult_readOnly              (requestReg_bits_decodeResult_readOnly),
    .instReq_bits_decodeResult_maskSource            (requestReg_bits_decodeResult_maskSource),
    .instReq_bits_decodeResult_maskDestination       (requestReg_bits_decodeResult_maskDestination),
    .instReq_bits_decodeResult_maskLogic             (requestReg_bits_decodeResult_maskLogic),
    .instReq_bits_decodeResult_uop                   (requestReg_bits_decodeResult_uop),
    .instReq_bits_decodeResult_iota                  (requestReg_bits_decodeResult_iota),
    .instReq_bits_decodeResult_mv                    (requestReg_bits_decodeResult_mv),
    .instReq_bits_decodeResult_extend                (requestReg_bits_decodeResult_extend),
    .instReq_bits_decodeResult_unOrderWrite          (requestReg_bits_decodeResult_unOrderWrite),
    .instReq_bits_decodeResult_compress              (requestReg_bits_decodeResult_compress),
    .instReq_bits_decodeResult_gather16              (requestReg_bits_decodeResult_gather16),
    .instReq_bits_decodeResult_gather                (requestReg_bits_decodeResult_gather),
    .instReq_bits_decodeResult_slid                  (requestReg_bits_decodeResult_slid),
    .instReq_bits_decodeResult_targetRd              (requestReg_bits_decodeResult_targetRd),
    .instReq_bits_decodeResult_widenReduce           (requestReg_bits_decodeResult_widenReduce),
    .instReq_bits_decodeResult_red                   (requestReg_bits_decodeResult_red),
    .instReq_bits_decodeResult_nr                    (requestReg_bits_decodeResult_nr),
    .instReq_bits_decodeResult_itype                 (requestReg_bits_decodeResult_itype),
    .instReq_bits_decodeResult_unsigned1             (requestReg_bits_decodeResult_unsigned1),
    .instReq_bits_decodeResult_unsigned0             (requestReg_bits_decodeResult_unsigned0),
    .instReq_bits_decodeResult_other                 (requestReg_bits_decodeResult_other),
    .instReq_bits_decodeResult_multiCycle            (requestReg_bits_decodeResult_multiCycle),
    .instReq_bits_decodeResult_divider               (requestReg_bits_decodeResult_divider),
    .instReq_bits_decodeResult_multiplier            (requestReg_bits_decodeResult_multiplier),
    .instReq_bits_decodeResult_shift                 (requestReg_bits_decodeResult_shift),
    .instReq_bits_decodeResult_adder                 (requestReg_bits_decodeResult_adder),
    .instReq_bits_decodeResult_logic                 (requestReg_bits_decodeResult_logic),
    .instReq_bits_readFromScala                      (requestReg_bits_decodeResult_itype ? {27'h0, imm} : requestRegDequeue_bits_rs1Data),
    .instReq_bits_sew                                (requestRegCSR_vSew),
    .instReq_bits_vlmul                              (requestRegCSR_vlmul),
    .instReq_bits_maskType                           (maskType),
    .instReq_bits_vxrm                               ({1'h0, requestRegCSR_vxrm}),
    .instReq_bits_vs2                                (requestRegDequeue_bits_instruction[24:20]),
    .instReq_bits_vs1                                (requestRegDequeue_bits_instruction[19:15]),
    .instReq_bits_vd                                 (requestRegDequeue_bits_instruction[11:7]),
    .instReq_bits_vl                                 (requestRegCSR_vl),
    .exeReq_0_valid                                  (_laneVec_0_maskUnitRequest_valid & ~_laneVec_0_maskRequestToLSU),
    .exeReq_0_bits_source1                           (_laneVec_0_maskUnitRequest_bits_source1),
    .exeReq_0_bits_source2                           (_laneVec_0_maskUnitRequest_bits_source2),
    .exeReq_0_bits_index                             (_laneVec_0_maskUnitRequest_bits_index),
    .exeReq_0_bits_ffo                               (_laneVec_0_maskUnitRequest_bits_ffo),
    .exeReq_1_valid                                  (_laneVec_1_maskUnitRequest_valid & ~_laneVec_1_maskRequestToLSU),
    .exeReq_1_bits_source1                           (_laneVec_1_maskUnitRequest_bits_source1),
    .exeReq_1_bits_source2                           (_laneVec_1_maskUnitRequest_bits_source2),
    .exeReq_1_bits_index                             (_laneVec_1_maskUnitRequest_bits_index),
    .exeReq_1_bits_ffo                               (_laneVec_1_maskUnitRequest_bits_ffo),
    .exeReq_2_valid                                  (_laneVec_2_maskUnitRequest_valid & ~_laneVec_2_maskRequestToLSU),
    .exeReq_2_bits_source1                           (_laneVec_2_maskUnitRequest_bits_source1),
    .exeReq_2_bits_source2                           (_laneVec_2_maskUnitRequest_bits_source2),
    .exeReq_2_bits_index                             (_laneVec_2_maskUnitRequest_bits_index),
    .exeReq_2_bits_ffo                               (_laneVec_2_maskUnitRequest_bits_ffo),
    .exeReq_3_valid                                  (_laneVec_3_maskUnitRequest_valid & ~_laneVec_3_maskRequestToLSU),
    .exeReq_3_bits_source1                           (_laneVec_3_maskUnitRequest_bits_source1),
    .exeReq_3_bits_source2                           (_laneVec_3_maskUnitRequest_bits_source2),
    .exeReq_3_bits_index                             (_laneVec_3_maskUnitRequest_bits_index),
    .exeReq_3_bits_ffo                               (_laneVec_3_maskUnitRequest_bits_ffo),
    .exeReq_4_valid                                  (_laneVec_4_maskUnitRequest_valid & ~_laneVec_4_maskRequestToLSU),
    .exeReq_4_bits_source1                           (_laneVec_4_maskUnitRequest_bits_source1),
    .exeReq_4_bits_source2                           (_laneVec_4_maskUnitRequest_bits_source2),
    .exeReq_4_bits_index                             (_laneVec_4_maskUnitRequest_bits_index),
    .exeReq_4_bits_ffo                               (_laneVec_4_maskUnitRequest_bits_ffo),
    .exeReq_5_valid                                  (_laneVec_5_maskUnitRequest_valid & ~_laneVec_5_maskRequestToLSU),
    .exeReq_5_bits_source1                           (_laneVec_5_maskUnitRequest_bits_source1),
    .exeReq_5_bits_source2                           (_laneVec_5_maskUnitRequest_bits_source2),
    .exeReq_5_bits_index                             (_laneVec_5_maskUnitRequest_bits_index),
    .exeReq_5_bits_ffo                               (_laneVec_5_maskUnitRequest_bits_ffo),
    .exeReq_6_valid                                  (_laneVec_6_maskUnitRequest_valid & ~_laneVec_6_maskRequestToLSU),
    .exeReq_6_bits_source1                           (_laneVec_6_maskUnitRequest_bits_source1),
    .exeReq_6_bits_source2                           (_laneVec_6_maskUnitRequest_bits_source2),
    .exeReq_6_bits_index                             (_laneVec_6_maskUnitRequest_bits_index),
    .exeReq_6_bits_ffo                               (_laneVec_6_maskUnitRequest_bits_ffo),
    .exeReq_7_valid                                  (_laneVec_7_maskUnitRequest_valid & ~_laneVec_7_maskRequestToLSU),
    .exeReq_7_bits_source1                           (_laneVec_7_maskUnitRequest_bits_source1),
    .exeReq_7_bits_source2                           (_laneVec_7_maskUnitRequest_bits_source2),
    .exeReq_7_bits_index                             (_laneVec_7_maskUnitRequest_bits_index),
    .exeReq_7_bits_ffo                               (_laneVec_7_maskUnitRequest_bits_ffo),
    .exeResp_0_ready                                 (x22_0_ready),
    .exeResp_0_valid                                 (_maskUnit_exeResp_0_valid),
    .exeResp_0_bits_vd                               (x22_0_bits_vd),
    .exeResp_0_bits_offset                           (x22_0_bits_offset),
    .exeResp_0_bits_mask                             (_maskUnit_exeResp_0_bits_mask),
    .exeResp_0_bits_data                             (x22_0_bits_data),
    .exeResp_0_bits_instructionIndex                 (_maskUnit_exeResp_0_bits_instructionIndex),
    .exeResp_1_ready                                 (x22_1_0_ready),
    .exeResp_1_valid                                 (_maskUnit_exeResp_1_valid),
    .exeResp_1_bits_vd                               (x22_1_0_bits_vd),
    .exeResp_1_bits_offset                           (x22_1_0_bits_offset),
    .exeResp_1_bits_mask                             (_maskUnit_exeResp_1_bits_mask),
    .exeResp_1_bits_data                             (x22_1_0_bits_data),
    .exeResp_1_bits_instructionIndex                 (_maskUnit_exeResp_1_bits_instructionIndex),
    .exeResp_2_ready                                 (x22_2_0_ready),
    .exeResp_2_valid                                 (_maskUnit_exeResp_2_valid),
    .exeResp_2_bits_vd                               (x22_2_0_bits_vd),
    .exeResp_2_bits_offset                           (x22_2_0_bits_offset),
    .exeResp_2_bits_mask                             (_maskUnit_exeResp_2_bits_mask),
    .exeResp_2_bits_data                             (x22_2_0_bits_data),
    .exeResp_2_bits_instructionIndex                 (_maskUnit_exeResp_2_bits_instructionIndex),
    .exeResp_3_ready                                 (x22_3_0_ready),
    .exeResp_3_valid                                 (_maskUnit_exeResp_3_valid),
    .exeResp_3_bits_vd                               (x22_3_0_bits_vd),
    .exeResp_3_bits_offset                           (x22_3_0_bits_offset),
    .exeResp_3_bits_mask                             (_maskUnit_exeResp_3_bits_mask),
    .exeResp_3_bits_data                             (x22_3_0_bits_data),
    .exeResp_3_bits_instructionIndex                 (_maskUnit_exeResp_3_bits_instructionIndex),
    .exeResp_4_ready                                 (x22_4_0_ready),
    .exeResp_4_valid                                 (_maskUnit_exeResp_4_valid),
    .exeResp_4_bits_vd                               (x22_4_0_bits_vd),
    .exeResp_4_bits_offset                           (x22_4_0_bits_offset),
    .exeResp_4_bits_mask                             (_maskUnit_exeResp_4_bits_mask),
    .exeResp_4_bits_data                             (x22_4_0_bits_data),
    .exeResp_4_bits_instructionIndex                 (_maskUnit_exeResp_4_bits_instructionIndex),
    .exeResp_5_ready                                 (x22_5_0_ready),
    .exeResp_5_valid                                 (_maskUnit_exeResp_5_valid),
    .exeResp_5_bits_vd                               (x22_5_0_bits_vd),
    .exeResp_5_bits_offset                           (x22_5_0_bits_offset),
    .exeResp_5_bits_mask                             (_maskUnit_exeResp_5_bits_mask),
    .exeResp_5_bits_data                             (x22_5_0_bits_data),
    .exeResp_5_bits_instructionIndex                 (_maskUnit_exeResp_5_bits_instructionIndex),
    .exeResp_6_ready                                 (x22_6_0_ready),
    .exeResp_6_valid                                 (_maskUnit_exeResp_6_valid),
    .exeResp_6_bits_vd                               (x22_6_0_bits_vd),
    .exeResp_6_bits_offset                           (x22_6_0_bits_offset),
    .exeResp_6_bits_mask                             (_maskUnit_exeResp_6_bits_mask),
    .exeResp_6_bits_data                             (x22_6_0_bits_data),
    .exeResp_6_bits_instructionIndex                 (_maskUnit_exeResp_6_bits_instructionIndex),
    .exeResp_7_ready                                 (x22_7_0_ready),
    .exeResp_7_valid                                 (_maskUnit_exeResp_7_valid),
    .exeResp_7_bits_vd                               (x22_7_0_bits_vd),
    .exeResp_7_bits_offset                           (x22_7_0_bits_offset),
    .exeResp_7_bits_mask                             (_maskUnit_exeResp_7_bits_mask),
    .exeResp_7_bits_data                             (x22_7_0_bits_data),
    .exeResp_7_bits_instructionIndex                 (_maskUnit_exeResp_7_bits_instructionIndex),
    .writeRelease_0                                  (view__writeRelease_0_pipe_out_valid),
    .writeRelease_1                                  (view__writeRelease_1_pipe_out_valid),
    .writeRelease_2                                  (view__writeRelease_2_pipe_out_valid),
    .writeRelease_3                                  (view__writeRelease_3_pipe_out_valid),
    .writeRelease_4                                  (view__writeRelease_4_pipe_out_valid),
    .writeRelease_5                                  (view__writeRelease_5_pipe_out_valid),
    .writeRelease_6                                  (view__writeRelease_6_pipe_out_valid),
    .writeRelease_7                                  (view__writeRelease_7_pipe_out_valid),
    .tokenIO_0_maskRequestRelease                    (_maskUnit_tokenIO_0_maskRequestRelease),
    .tokenIO_1_maskRequestRelease                    (_maskUnit_tokenIO_1_maskRequestRelease),
    .tokenIO_2_maskRequestRelease                    (_maskUnit_tokenIO_2_maskRequestRelease),
    .tokenIO_3_maskRequestRelease                    (_maskUnit_tokenIO_3_maskRequestRelease),
    .tokenIO_4_maskRequestRelease                    (_maskUnit_tokenIO_4_maskRequestRelease),
    .tokenIO_5_maskRequestRelease                    (_maskUnit_tokenIO_5_maskRequestRelease),
    .tokenIO_6_maskRequestRelease                    (_maskUnit_tokenIO_6_maskRequestRelease),
    .tokenIO_7_maskRequestRelease                    (_maskUnit_tokenIO_7_maskRequestRelease),
    .readChannel_0_ready                             (x13_0_ready),
    .readChannel_0_valid                             (x13_0_valid),
    .readChannel_0_bits_vs                           (x13_0_bits_vs),
    .readChannel_0_bits_offset                       (x13_0_bits_offset),
    .readChannel_0_bits_instructionIndex             (x13_0_bits_instructionIndex),
    .readChannel_1_ready                             (x13_1_0_ready),
    .readChannel_1_valid                             (x13_1_0_valid),
    .readChannel_1_bits_vs                           (x13_1_0_bits_vs),
    .readChannel_1_bits_offset                       (x13_1_0_bits_offset),
    .readChannel_1_bits_instructionIndex             (x13_1_0_bits_instructionIndex),
    .readChannel_2_ready                             (x13_2_0_ready),
    .readChannel_2_valid                             (x13_2_0_valid),
    .readChannel_2_bits_vs                           (x13_2_0_bits_vs),
    .readChannel_2_bits_offset                       (x13_2_0_bits_offset),
    .readChannel_2_bits_instructionIndex             (x13_2_0_bits_instructionIndex),
    .readChannel_3_ready                             (x13_3_0_ready),
    .readChannel_3_valid                             (x13_3_0_valid),
    .readChannel_3_bits_vs                           (x13_3_0_bits_vs),
    .readChannel_3_bits_offset                       (x13_3_0_bits_offset),
    .readChannel_3_bits_instructionIndex             (x13_3_0_bits_instructionIndex),
    .readChannel_4_ready                             (x13_4_0_ready),
    .readChannel_4_valid                             (x13_4_0_valid),
    .readChannel_4_bits_vs                           (x13_4_0_bits_vs),
    .readChannel_4_bits_offset                       (x13_4_0_bits_offset),
    .readChannel_4_bits_instructionIndex             (x13_4_0_bits_instructionIndex),
    .readChannel_5_ready                             (x13_5_0_ready),
    .readChannel_5_valid                             (x13_5_0_valid),
    .readChannel_5_bits_vs                           (x13_5_0_bits_vs),
    .readChannel_5_bits_offset                       (x13_5_0_bits_offset),
    .readChannel_5_bits_instructionIndex             (x13_5_0_bits_instructionIndex),
    .readChannel_6_ready                             (x13_6_0_ready),
    .readChannel_6_valid                             (x13_6_0_valid),
    .readChannel_6_bits_vs                           (x13_6_0_bits_vs),
    .readChannel_6_bits_offset                       (x13_6_0_bits_offset),
    .readChannel_6_bits_instructionIndex             (x13_6_0_bits_instructionIndex),
    .readChannel_7_ready                             (x13_7_0_ready),
    .readChannel_7_valid                             (x13_7_0_valid),
    .readChannel_7_bits_vs                           (x13_7_0_bits_vs),
    .readChannel_7_bits_offset                       (x13_7_0_bits_offset),
    .readChannel_7_bits_instructionIndex             (x13_7_0_bits_instructionIndex),
    .readResult_0_valid                              (shifterReg_8_0_valid),
    .readResult_0_bits                               (shifterReg_8_0_bits),
    .readResult_1_valid                              (shifterReg_10_0_valid),
    .readResult_1_bits                               (shifterReg_10_0_bits),
    .readResult_2_valid                              (shifterReg_12_0_valid),
    .readResult_2_bits                               (shifterReg_12_0_bits),
    .readResult_3_valid                              (shifterReg_14_0_valid),
    .readResult_3_bits                               (shifterReg_14_0_bits),
    .readResult_4_valid                              (shifterReg_16_0_valid),
    .readResult_4_bits                               (shifterReg_16_0_bits),
    .readResult_5_valid                              (shifterReg_18_0_valid),
    .readResult_5_bits                               (shifterReg_18_0_bits),
    .readResult_6_valid                              (shifterReg_20_0_valid),
    .readResult_6_bits                               (shifterReg_20_0_bits),
    .readResult_7_valid                              (shifterReg_22_0_valid),
    .readResult_7_bits                               (shifterReg_22_0_bits),
    .lastReport                                      (_maskUnit_lastReport),
    .laneMaskInput_0                                 (_maskUnit_laneMaskInput_0),
    .laneMaskInput_1                                 (_maskUnit_laneMaskInput_1),
    .laneMaskInput_2                                 (_maskUnit_laneMaskInput_2),
    .laneMaskInput_3                                 (_maskUnit_laneMaskInput_3),
    .laneMaskInput_4                                 (_maskUnit_laneMaskInput_4),
    .laneMaskInput_5                                 (_maskUnit_laneMaskInput_5),
    .laneMaskInput_6                                 (_maskUnit_laneMaskInput_6),
    .laneMaskInput_7                                 (_maskUnit_laneMaskInput_7),
    .laneMaskSelect_0                                (view__laneMaskSelect_0_pipe_pipe_out_bits),
    .laneMaskSelect_1                                (view__laneMaskSelect_1_pipe_pipe_out_bits),
    .laneMaskSelect_2                                (view__laneMaskSelect_2_pipe_pipe_out_bits),
    .laneMaskSelect_3                                (view__laneMaskSelect_3_pipe_pipe_out_bits),
    .laneMaskSelect_4                                (view__laneMaskSelect_4_pipe_pipe_out_bits),
    .laneMaskSelect_5                                (view__laneMaskSelect_5_pipe_pipe_out_bits),
    .laneMaskSelect_6                                (view__laneMaskSelect_6_pipe_pipe_out_bits),
    .laneMaskSelect_7                                (view__laneMaskSelect_7_pipe_pipe_out_bits),
    .laneMaskSewSelect_0                             (view__laneMaskSewSelect_0_pipe_pipe_out_bits),
    .laneMaskSewSelect_1                             (view__laneMaskSewSelect_1_pipe_pipe_out_bits),
    .laneMaskSewSelect_2                             (view__laneMaskSewSelect_2_pipe_pipe_out_bits),
    .laneMaskSewSelect_3                             (view__laneMaskSewSelect_3_pipe_pipe_out_bits),
    .laneMaskSewSelect_4                             (view__laneMaskSewSelect_4_pipe_pipe_out_bits),
    .laneMaskSewSelect_5                             (view__laneMaskSewSelect_5_pipe_pipe_out_bits),
    .laneMaskSewSelect_6                             (view__laneMaskSewSelect_6_pipe_pipe_out_bits),
    .laneMaskSewSelect_7                             (view__laneMaskSewSelect_7_pipe_pipe_out_bits),
    .v0UpdateVec_0_valid                             (_laneVec_0_v0Update_valid),
    .v0UpdateVec_0_bits_data                         (_laneVec_0_v0Update_bits_data),
    .v0UpdateVec_0_bits_offset                       (_laneVec_0_v0Update_bits_offset),
    .v0UpdateVec_0_bits_mask                         (_laneVec_0_v0Update_bits_mask),
    .v0UpdateVec_1_valid                             (_laneVec_1_v0Update_valid),
    .v0UpdateVec_1_bits_data                         (_laneVec_1_v0Update_bits_data),
    .v0UpdateVec_1_bits_offset                       (_laneVec_1_v0Update_bits_offset),
    .v0UpdateVec_1_bits_mask                         (_laneVec_1_v0Update_bits_mask),
    .v0UpdateVec_2_valid                             (_laneVec_2_v0Update_valid),
    .v0UpdateVec_2_bits_data                         (_laneVec_2_v0Update_bits_data),
    .v0UpdateVec_2_bits_offset                       (_laneVec_2_v0Update_bits_offset),
    .v0UpdateVec_2_bits_mask                         (_laneVec_2_v0Update_bits_mask),
    .v0UpdateVec_3_valid                             (_laneVec_3_v0Update_valid),
    .v0UpdateVec_3_bits_data                         (_laneVec_3_v0Update_bits_data),
    .v0UpdateVec_3_bits_offset                       (_laneVec_3_v0Update_bits_offset),
    .v0UpdateVec_3_bits_mask                         (_laneVec_3_v0Update_bits_mask),
    .v0UpdateVec_4_valid                             (_laneVec_4_v0Update_valid),
    .v0UpdateVec_4_bits_data                         (_laneVec_4_v0Update_bits_data),
    .v0UpdateVec_4_bits_offset                       (_laneVec_4_v0Update_bits_offset),
    .v0UpdateVec_4_bits_mask                         (_laneVec_4_v0Update_bits_mask),
    .v0UpdateVec_5_valid                             (_laneVec_5_v0Update_valid),
    .v0UpdateVec_5_bits_data                         (_laneVec_5_v0Update_bits_data),
    .v0UpdateVec_5_bits_offset                       (_laneVec_5_v0Update_bits_offset),
    .v0UpdateVec_5_bits_mask                         (_laneVec_5_v0Update_bits_mask),
    .v0UpdateVec_6_valid                             (_laneVec_6_v0Update_valid),
    .v0UpdateVec_6_bits_data                         (_laneVec_6_v0Update_bits_data),
    .v0UpdateVec_6_bits_offset                       (_laneVec_6_v0Update_bits_offset),
    .v0UpdateVec_6_bits_mask                         (_laneVec_6_v0Update_bits_mask),
    .v0UpdateVec_7_valid                             (_laneVec_7_v0Update_valid),
    .v0UpdateVec_7_bits_data                         (_laneVec_7_v0Update_bits_data),
    .v0UpdateVec_7_bits_offset                       (_laneVec_7_v0Update_bits_offset),
    .v0UpdateVec_7_bits_mask                         (_laneVec_7_v0Update_bits_mask),
    .writeRDData                                     (retire_rd_bits_rdData_0),
    .gatherData_ready                                (maskUnit_gatherData_ready),
    .gatherData_valid                                (_maskUnit_gatherData_valid),
    .gatherData_bits                                 (_maskUnit_gatherData_bits),
    .gatherRead                                      (gatherNeedRead)
  );
  T1TokenManager tokenManager (
    .clock                                  (clock),
    .reset                                  (reset),
    .instructionIssue_valid                 (maskUnit_gatherData_ready),
    .instructionIssue_bits_instructionIndex (requestReg_bits_instructionIndex),
    .instructionIssue_bits_writeV0          (~requestReg_bits_decodeResult_targetRd & ~isStoreType & requestReg_bits_vdIsV0),
    .instructionIssue_bits_useV0AsMask      (maskType),
    .instructionIssue_bits_toLane           (~noOffsetReadLoadStore & ~maskUnitInstruction),
    .instructionIssue_bits_toMask           (requestReg_bits_decodeResult_maskUnit),
    .lsuWriteV0_0_valid                     (x22_1_ready & _lsu_vrfWritePort_0_valid & _lsu_vrfWritePort_0_bits_vd == 5'h0 & (|_lsu_vrfWritePort_0_bits_mask)),
    .lsuWriteV0_0_bits                      (_lsu_vrfWritePort_0_bits_instructionIndex),
    .lsuWriteV0_1_valid                     (x22_1_1_ready & _lsu_vrfWritePort_1_valid & _lsu_vrfWritePort_1_bits_vd == 5'h0 & (|_lsu_vrfWritePort_1_bits_mask)),
    .lsuWriteV0_1_bits                      (_lsu_vrfWritePort_1_bits_instructionIndex),
    .lsuWriteV0_2_valid                     (x22_2_1_ready & _lsu_vrfWritePort_2_valid & _lsu_vrfWritePort_2_bits_vd == 5'h0 & (|_lsu_vrfWritePort_2_bits_mask)),
    .lsuWriteV0_2_bits                      (_lsu_vrfWritePort_2_bits_instructionIndex),
    .lsuWriteV0_3_valid                     (x22_3_1_ready & _lsu_vrfWritePort_3_valid & _lsu_vrfWritePort_3_bits_vd == 5'h0 & (|_lsu_vrfWritePort_3_bits_mask)),
    .lsuWriteV0_3_bits                      (_lsu_vrfWritePort_3_bits_instructionIndex),
    .lsuWriteV0_4_valid                     (x22_4_1_ready & _lsu_vrfWritePort_4_valid & _lsu_vrfWritePort_4_bits_vd == 5'h0 & (|_lsu_vrfWritePort_4_bits_mask)),
    .lsuWriteV0_4_bits                      (_lsu_vrfWritePort_4_bits_instructionIndex),
    .lsuWriteV0_5_valid                     (x22_5_1_ready & _lsu_vrfWritePort_5_valid & _lsu_vrfWritePort_5_bits_vd == 5'h0 & (|_lsu_vrfWritePort_5_bits_mask)),
    .lsuWriteV0_5_bits                      (_lsu_vrfWritePort_5_bits_instructionIndex),
    .lsuWriteV0_6_valid                     (x22_6_1_ready & _lsu_vrfWritePort_6_valid & _lsu_vrfWritePort_6_bits_vd == 5'h0 & (|_lsu_vrfWritePort_6_bits_mask)),
    .lsuWriteV0_6_bits                      (_lsu_vrfWritePort_6_bits_instructionIndex),
    .lsuWriteV0_7_valid                     (x22_7_1_ready & _lsu_vrfWritePort_7_valid & _lsu_vrfWritePort_7_bits_vd == 5'h0 & (|_lsu_vrfWritePort_7_bits_mask)),
    .lsuWriteV0_7_bits                      (_lsu_vrfWritePort_7_bits_instructionIndex),
    .issueAllow                             (_tokenManager_issueAllow),
    .instructionFinish_0                    (instructionFinishedPipe_pipe_out_bits),
    .instructionFinish_1                    (instructionFinishedPipe_pipe_out_1_bits),
    .instructionFinish_2                    (instructionFinishedPipe_pipe_out_2_bits),
    .instructionFinish_3                    (instructionFinishedPipe_pipe_out_3_bits),
    .instructionFinish_4                    (instructionFinishedPipe_pipe_out_4_bits),
    .instructionFinish_5                    (instructionFinishedPipe_pipe_out_5_bits),
    .instructionFinish_6                    (instructionFinishedPipe_pipe_out_6_bits),
    .instructionFinish_7                    (instructionFinishedPipe_pipe_out_7_bits),
    .v0WriteValid                           (_tokenManager_v0WriteValid),
    .maskUnitFree                           (slots_3_state_idle)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(145)
  ) queue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_enq_ready & queue_enq_valid & ~(_queue_fifo_empty & queue_deq_ready))),
    .pop_req_n    (~(queue_deq_ready & ~_queue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn),
    .empty        (_queue_fifo_empty),
    .almost_empty (queue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_almostFull),
    .full         (_queue_fifo_full),
    .error        (_queue_fifo_error),
    .data_out     (_queue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(145)
  ) queue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_1_enq_ready & queue_1_enq_valid & ~(_queue_fifo_1_empty & queue_1_deq_ready))),
    .pop_req_n    (~(queue_1_deq_ready & ~_queue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn_1),
    .empty        (_queue_fifo_1_empty),
    .almost_empty (queue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_1_almostFull),
    .full         (_queue_fifo_1_full),
    .error        (_queue_fifo_1_error),
    .data_out     (_queue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(145)
  ) queue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_2_enq_ready & queue_2_enq_valid & ~(_queue_fifo_2_empty & queue_2_deq_ready))),
    .pop_req_n    (~(queue_2_deq_ready & ~_queue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn_2),
    .empty        (_queue_fifo_2_empty),
    .almost_empty (queue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_2_almostFull),
    .full         (_queue_fifo_2_full),
    .error        (_queue_fifo_2_error),
    .data_out     (_queue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(145)
  ) queue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_3_enq_ready & queue_3_enq_valid & ~(_queue_fifo_3_empty & queue_3_deq_ready))),
    .pop_req_n    (~(queue_3_deq_ready & ~_queue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn_3),
    .empty        (_queue_fifo_3_empty),
    .almost_empty (queue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_3_almostFull),
    .full         (_queue_fifo_3_full),
    .error        (_queue_fifo_3_error),
    .data_out     (_queue_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(145)
  ) queue_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_4_enq_ready & queue_4_enq_valid & ~(_queue_fifo_4_empty & queue_4_deq_ready))),
    .pop_req_n    (~(queue_4_deq_ready & ~_queue_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn_4),
    .empty        (_queue_fifo_4_empty),
    .almost_empty (queue_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_4_almostFull),
    .full         (_queue_fifo_4_full),
    .error        (_queue_fifo_4_error),
    .data_out     (_queue_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(145)
  ) queue_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_5_enq_ready & queue_5_enq_valid & ~(_queue_fifo_5_empty & queue_5_deq_ready))),
    .pop_req_n    (~(queue_5_deq_ready & ~_queue_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn_5),
    .empty        (_queue_fifo_5_empty),
    .almost_empty (queue_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_5_almostFull),
    .full         (_queue_fifo_5_full),
    .error        (_queue_fifo_5_error),
    .data_out     (_queue_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(145)
  ) queue_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_6_enq_ready & queue_6_enq_valid & ~(_queue_fifo_6_empty & queue_6_deq_ready))),
    .pop_req_n    (~(queue_6_deq_ready & ~_queue_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn_6),
    .empty        (_queue_fifo_6_empty),
    .almost_empty (queue_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_6_almostFull),
    .full         (_queue_fifo_6_full),
    .error        (_queue_fifo_6_error),
    .data_out     (_queue_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(145)
  ) queue_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_7_enq_ready & queue_7_enq_valid & ~(_queue_fifo_7_empty & queue_7_deq_ready))),
    .pop_req_n    (~(queue_7_deq_ready & ~_queue_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_dataIn_7),
    .empty        (_queue_fifo_7_empty),
    .almost_empty (queue_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_7_almostFull),
    .full         (_queue_fifo_7_full),
    .error        (_queue_fifo_7_error),
    .data_out     (_queue_fifo_7_data_out)
  );
  Lane laneVec_0 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (3'h0),
    .readBusPort_0_enq_valid                             (shifterReg_24_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_24_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_0_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_0_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_0_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_16_valid),
    .readBusPort_1_enq_valid                             (shifterReg_26_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_26_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_0_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_0_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_0_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_32_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_25_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_25_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_25_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_25_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_25_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_0_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_0_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_0_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_0_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_0_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_0_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_17_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_41_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_41_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_41_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_41_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_41_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_0_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_0_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_0_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_0_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_0_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_0_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_19_valid),
    .laneRequest_ready                                   (_laneVec_0_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_0_valid & laneRequestSinkWire_0_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_0_bits_instructionIndex),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_0_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_0_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_0_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_0_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_0_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_0_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_0_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_0_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_0_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_0_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_0_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_0_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_0_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_0_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_0_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_0_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_0_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_0_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_0_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_0_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_0_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_0_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_0_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_0_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_0_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_0_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_0_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_0_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_0_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_0_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_0_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_0_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_0_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_0_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_0_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_0_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_0_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_0_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_0_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_0_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_0_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_0_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_0_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_0_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_0_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_0_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_0_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_0_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_0_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_0_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_0_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_0_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_0_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_0_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_0_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_0_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_0_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_0_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_0_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_0_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_0_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_0_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_0_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_0_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_0_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_0_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_0_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_0_maskUnitRequest_bits_ffo),
    .maskRequestToLSU                                    (_laneVec_0_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_0_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[0]),
    .vrfReadAddressChannel_ready                         (sinkWire_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_0_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_1_ready),
    .vrfWriteChannel_valid                               (sinkWire_1_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_1_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_1_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_1_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_1_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_1_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_1_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_0_valid_T),
    .instructionFinished                                 (_laneVec_0_instructionFinished),
    .vxsatReport                                         (_laneVec_0_vxsatReport),
    .v0Update_valid                                      (_laneVec_0_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_0_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_0_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_0_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_bits),
    .maskSelect                                          (_laneVec_0_maskSelect),
    .maskSelectSew                                       (_laneVec_0_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_bits | maskLastPipe_pipe_out_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_0),
    .writeCount                                          (pipe_out_1_bits),
    .writeQueueValid                                     (dataInWritePipeVec_0)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(13)
  ) sinkVec_queue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_enq_ready & sinkVec_queue_enq_valid & ~(_sinkVec_queue_fifo_empty & sinkVec_queue_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_deq_ready & ~_sinkVec_queue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn),
    .empty        (_sinkVec_queue_fifo_empty),
    .almost_empty (sinkVec_queue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_almostFull),
    .full         (_sinkVec_queue_fifo_full),
    .error        (_sinkVec_queue_fifo_error),
    .data_out     (_sinkVec_queue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(13)
  ) sinkVec_queue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_1_enq_ready & sinkVec_queue_1_enq_valid & ~(_sinkVec_queue_fifo_1_empty & sinkVec_queue_1_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_1_deq_ready & ~_sinkVec_queue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_1),
    .empty        (_sinkVec_queue_fifo_1_empty),
    .almost_empty (sinkVec_queue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_1_almostFull),
    .full         (_sinkVec_queue_fifo_1_full),
    .error        (_sinkVec_queue_fifo_1_error),
    .data_out     (_sinkVec_queue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) sinkVec_queue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_2_enq_ready & sinkVec_queue_2_enq_valid & ~(_sinkVec_queue_fifo_2_empty & sinkVec_queue_2_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_2_deq_ready & ~_sinkVec_queue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_2),
    .empty        (_sinkVec_queue_fifo_2_empty),
    .almost_empty (sinkVec_queue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_2_almostFull),
    .full         (_sinkVec_queue_fifo_2_full),
    .error        (_sinkVec_queue_fifo_2_error),
    .data_out     (_sinkVec_queue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) sinkVec_queue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_3_enq_ready & sinkVec_queue_3_enq_valid & ~(_sinkVec_queue_fifo_3_empty & sinkVec_queue_3_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_3_deq_ready & ~_sinkVec_queue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_3),
    .empty        (_sinkVec_queue_fifo_3_empty),
    .almost_empty (sinkVec_queue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_3_almostFull),
    .full         (_sinkVec_queue_fifo_3_full),
    .error        (_sinkVec_queue_fifo_3_error),
    .data_out     (_sinkVec_queue_fifo_3_data_out)
  );
  Lane laneVec_1 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (3'h1),
    .readBusPort_0_enq_valid                             (shifterReg_28_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_28_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_1_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_1_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_1_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_18_valid),
    .readBusPort_1_enq_valid                             (shifterReg_30_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_30_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_1_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_1_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_1_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_34_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_27_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_27_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_27_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_27_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_27_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_1_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_1_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_1_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_1_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_1_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_1_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_21_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_43_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_43_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_43_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_43_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_43_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_1_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_1_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_1_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_1_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_1_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_1_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_23_valid),
    .laneRequest_ready                                   (_laneVec_1_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_1_valid & laneRequestSinkWire_1_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_1_bits_instructionIndex),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_1_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_1_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_1_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_1_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_1_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_1_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_1_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_1_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_1_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_1_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_1_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_1_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_1_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_1_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_1_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_1_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_1_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_1_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_1_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_1_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_1_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_1_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_1_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_1_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_1_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_1_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_1_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_1_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_1_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_1_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_1_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_1_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_1_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_1_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_1_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_1_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_1_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_1_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_1_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_1_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_1_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_1_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_1_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_1_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_1_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_1_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_1_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_1_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_1_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_1_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_1_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_1_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_1_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_1_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_1_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_1_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_1_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_1_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_1_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_1_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_1_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_1_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_1_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_1_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_1_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_1_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_1_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_1_maskUnitRequest_bits_ffo),
    .maskRequestToLSU                                    (_laneVec_1_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_1_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[1]),
    .vrfReadAddressChannel_ready                         (sinkWire_2_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_2_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_2_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_2_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_2_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_2_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_1_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_3_ready),
    .vrfWriteChannel_valid                               (sinkWire_3_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_3_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_3_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_3_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_3_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_3_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_3_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_1_valid_T),
    .instructionFinished                                 (_laneVec_1_instructionFinished),
    .vxsatReport                                         (_laneVec_1_vxsatReport),
    .v0Update_valid                                      (_laneVec_1_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_1_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_1_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_1_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_1_bits),
    .maskSelect                                          (_laneVec_1_maskSelect),
    .maskSelectSew                                       (_laneVec_1_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_1_bits | maskLastPipe_pipe_out_1_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_1),
    .writeCount                                          (pipe_out_3_bits),
    .writeQueueValid                                     (dataInWritePipeVec_1)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(13)
  ) sinkVec_queue_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_4_enq_ready & sinkVec_queue_4_enq_valid & ~(_sinkVec_queue_fifo_4_empty & sinkVec_queue_4_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_4_deq_ready & ~_sinkVec_queue_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_4),
    .empty        (_sinkVec_queue_fifo_4_empty),
    .almost_empty (sinkVec_queue_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_4_almostFull),
    .full         (_sinkVec_queue_fifo_4_full),
    .error        (_sinkVec_queue_fifo_4_error),
    .data_out     (_sinkVec_queue_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(13)
  ) sinkVec_queue_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_5_enq_ready & sinkVec_queue_5_enq_valid & ~(_sinkVec_queue_fifo_5_empty & sinkVec_queue_5_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_5_deq_ready & ~_sinkVec_queue_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_5),
    .empty        (_sinkVec_queue_fifo_5_empty),
    .almost_empty (sinkVec_queue_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_5_almostFull),
    .full         (_sinkVec_queue_fifo_5_full),
    .error        (_sinkVec_queue_fifo_5_error),
    .data_out     (_sinkVec_queue_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) sinkVec_queue_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_6_enq_ready & sinkVec_queue_6_enq_valid & ~(_sinkVec_queue_fifo_6_empty & sinkVec_queue_6_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_6_deq_ready & ~_sinkVec_queue_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_6),
    .empty        (_sinkVec_queue_fifo_6_empty),
    .almost_empty (sinkVec_queue_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_6_almostFull),
    .full         (_sinkVec_queue_fifo_6_full),
    .error        (_sinkVec_queue_fifo_6_error),
    .data_out     (_sinkVec_queue_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) sinkVec_queue_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_7_enq_ready & sinkVec_queue_7_enq_valid & ~(_sinkVec_queue_fifo_7_empty & sinkVec_queue_7_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_7_deq_ready & ~_sinkVec_queue_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_7),
    .empty        (_sinkVec_queue_fifo_7_empty),
    .almost_empty (sinkVec_queue_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_7_almostFull),
    .full         (_sinkVec_queue_fifo_7_full),
    .error        (_sinkVec_queue_fifo_7_error),
    .data_out     (_sinkVec_queue_fifo_7_data_out)
  );
  Lane laneVec_2 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (3'h2),
    .readBusPort_0_enq_valid                             (shifterReg_32_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_32_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_2_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_2_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_2_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_20_valid),
    .readBusPort_1_enq_valid                             (shifterReg_34_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_34_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_2_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_2_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_2_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_36_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_29_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_29_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_29_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_29_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_29_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_2_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_2_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_2_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_2_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_2_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_2_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_25_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_45_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_45_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_45_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_45_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_45_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_2_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_2_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_2_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_2_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_2_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_2_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_27_valid),
    .laneRequest_ready                                   (_laneVec_2_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_2_valid & laneRequestSinkWire_2_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_2_bits_instructionIndex),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_2_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_2_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_2_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_2_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_2_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_2_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_2_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_2_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_2_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_2_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_2_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_2_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_2_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_2_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_2_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_2_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_2_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_2_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_2_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_2_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_2_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_2_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_2_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_2_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_2_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_2_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_2_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_2_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_2_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_2_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_2_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_2_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_2_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_2_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_2_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_2_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_2_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_2_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_2_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_2_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_2_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_2_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_2_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_2_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_2_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_2_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_2_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_2_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_2_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_2_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_2_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_2_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_2_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_2_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_2_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_2_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_2_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_2_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_2_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_2_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_2_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_2_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_2_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_2_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_2_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_2_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_2_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_2_maskUnitRequest_bits_ffo),
    .maskRequestToLSU                                    (_laneVec_2_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_2_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[2]),
    .vrfReadAddressChannel_ready                         (sinkWire_4_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_4_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_4_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_4_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_4_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_4_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_2_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_5_ready),
    .vrfWriteChannel_valid                               (sinkWire_5_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_5_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_5_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_5_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_5_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_5_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_5_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_2_valid_T),
    .instructionFinished                                 (_laneVec_2_instructionFinished),
    .vxsatReport                                         (_laneVec_2_vxsatReport),
    .v0Update_valid                                      (_laneVec_2_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_2_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_2_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_2_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_2_bits),
    .maskSelect                                          (_laneVec_2_maskSelect),
    .maskSelectSew                                       (_laneVec_2_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_2_bits | maskLastPipe_pipe_out_2_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_2),
    .writeCount                                          (pipe_out_5_bits),
    .writeQueueValid                                     (dataInWritePipeVec_2)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(13)
  ) sinkVec_queue_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_8_enq_ready & sinkVec_queue_8_enq_valid & ~(_sinkVec_queue_fifo_8_empty & sinkVec_queue_8_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_8_deq_ready & ~_sinkVec_queue_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_8),
    .empty        (_sinkVec_queue_fifo_8_empty),
    .almost_empty (sinkVec_queue_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_8_almostFull),
    .full         (_sinkVec_queue_fifo_8_full),
    .error        (_sinkVec_queue_fifo_8_error),
    .data_out     (_sinkVec_queue_fifo_8_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(13)
  ) sinkVec_queue_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_9_enq_ready & sinkVec_queue_9_enq_valid & ~(_sinkVec_queue_fifo_9_empty & sinkVec_queue_9_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_9_deq_ready & ~_sinkVec_queue_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_9),
    .empty        (_sinkVec_queue_fifo_9_empty),
    .almost_empty (sinkVec_queue_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_9_almostFull),
    .full         (_sinkVec_queue_fifo_9_full),
    .error        (_sinkVec_queue_fifo_9_error),
    .data_out     (_sinkVec_queue_fifo_9_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) sinkVec_queue_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_10_enq_ready & sinkVec_queue_10_enq_valid & ~(_sinkVec_queue_fifo_10_empty & sinkVec_queue_10_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_10_deq_ready & ~_sinkVec_queue_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_10),
    .empty        (_sinkVec_queue_fifo_10_empty),
    .almost_empty (sinkVec_queue_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_10_almostFull),
    .full         (_sinkVec_queue_fifo_10_full),
    .error        (_sinkVec_queue_fifo_10_error),
    .data_out     (_sinkVec_queue_fifo_10_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) sinkVec_queue_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_11_enq_ready & sinkVec_queue_11_enq_valid & ~(_sinkVec_queue_fifo_11_empty & sinkVec_queue_11_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_11_deq_ready & ~_sinkVec_queue_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_11),
    .empty        (_sinkVec_queue_fifo_11_empty),
    .almost_empty (sinkVec_queue_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_11_almostFull),
    .full         (_sinkVec_queue_fifo_11_full),
    .error        (_sinkVec_queue_fifo_11_error),
    .data_out     (_sinkVec_queue_fifo_11_data_out)
  );
  Lane laneVec_3 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (3'h3),
    .readBusPort_0_enq_valid                             (shifterReg_36_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_36_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_3_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_3_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_3_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_22_valid),
    .readBusPort_1_enq_valid                             (shifterReg_38_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_38_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_3_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_3_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_3_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_38_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_31_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_31_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_31_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_31_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_31_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_3_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_3_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_3_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_3_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_3_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_3_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_29_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_47_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_47_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_47_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_47_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_47_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_3_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_3_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_3_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_3_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_3_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_3_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_31_valid),
    .laneRequest_ready                                   (_laneVec_3_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_3_valid & laneRequestSinkWire_3_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_3_bits_instructionIndex),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_3_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_3_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_3_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_3_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_3_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_3_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_3_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_3_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_3_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_3_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_3_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_3_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_3_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_3_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_3_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_3_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_3_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_3_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_3_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_3_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_3_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_3_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_3_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_3_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_3_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_3_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_3_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_3_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_3_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_3_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_3_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_3_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_3_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_3_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_3_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_3_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_3_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_3_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_3_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_3_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_3_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_3_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_3_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_3_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_3_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_3_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_3_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_3_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_3_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_3_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_3_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_3_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_3_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_3_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_3_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_3_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_3_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_3_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_3_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_3_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_3_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_3_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_3_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_3_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_3_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_3_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_3_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_3_maskUnitRequest_bits_ffo),
    .maskRequestToLSU                                    (_laneVec_3_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_3_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[3]),
    .vrfReadAddressChannel_ready                         (sinkWire_6_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_6_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_6_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_6_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_6_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_6_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_3_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_7_ready),
    .vrfWriteChannel_valid                               (sinkWire_7_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_7_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_7_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_7_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_7_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_7_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_7_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_3_valid_T),
    .instructionFinished                                 (_laneVec_3_instructionFinished),
    .vxsatReport                                         (_laneVec_3_vxsatReport),
    .v0Update_valid                                      (_laneVec_3_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_3_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_3_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_3_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_3_bits),
    .maskSelect                                          (_laneVec_3_maskSelect),
    .maskSelectSew                                       (_laneVec_3_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_3_bits | maskLastPipe_pipe_out_3_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_3),
    .writeCount                                          (pipe_out_7_bits),
    .writeQueueValid                                     (dataInWritePipeVec_3)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(13)
  ) sinkVec_queue_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_12_enq_ready & sinkVec_queue_12_enq_valid & ~(_sinkVec_queue_fifo_12_empty & sinkVec_queue_12_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_12_deq_ready & ~_sinkVec_queue_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_12),
    .empty        (_sinkVec_queue_fifo_12_empty),
    .almost_empty (sinkVec_queue_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_12_almostFull),
    .full         (_sinkVec_queue_fifo_12_full),
    .error        (_sinkVec_queue_fifo_12_error),
    .data_out     (_sinkVec_queue_fifo_12_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(13)
  ) sinkVec_queue_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_13_enq_ready & sinkVec_queue_13_enq_valid & ~(_sinkVec_queue_fifo_13_empty & sinkVec_queue_13_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_13_deq_ready & ~_sinkVec_queue_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_13),
    .empty        (_sinkVec_queue_fifo_13_empty),
    .almost_empty (sinkVec_queue_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_13_almostFull),
    .full         (_sinkVec_queue_fifo_13_full),
    .error        (_sinkVec_queue_fifo_13_error),
    .data_out     (_sinkVec_queue_fifo_13_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) sinkVec_queue_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_14_enq_ready & sinkVec_queue_14_enq_valid & ~(_sinkVec_queue_fifo_14_empty & sinkVec_queue_14_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_14_deq_ready & ~_sinkVec_queue_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_14),
    .empty        (_sinkVec_queue_fifo_14_empty),
    .almost_empty (sinkVec_queue_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_14_almostFull),
    .full         (_sinkVec_queue_fifo_14_full),
    .error        (_sinkVec_queue_fifo_14_error),
    .data_out     (_sinkVec_queue_fifo_14_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) sinkVec_queue_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_15_enq_ready & sinkVec_queue_15_enq_valid & ~(_sinkVec_queue_fifo_15_empty & sinkVec_queue_15_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_15_deq_ready & ~_sinkVec_queue_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_15),
    .empty        (_sinkVec_queue_fifo_15_empty),
    .almost_empty (sinkVec_queue_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_15_almostFull),
    .full         (_sinkVec_queue_fifo_15_full),
    .error        (_sinkVec_queue_fifo_15_error),
    .data_out     (_sinkVec_queue_fifo_15_data_out)
  );
  Lane laneVec_4 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (3'h4),
    .readBusPort_0_enq_valid                             (shifterReg_40_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_40_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_4_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_4_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_4_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_24_valid),
    .readBusPort_1_enq_valid                             (shifterReg_42_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_42_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_4_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_4_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_4_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_40_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_33_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_33_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_33_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_33_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_33_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_4_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_4_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_4_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_4_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_4_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_4_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_33_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_49_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_49_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_49_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_49_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_49_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_4_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_4_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_4_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_4_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_4_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_4_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_35_valid),
    .laneRequest_ready                                   (_laneVec_4_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_4_valid & laneRequestSinkWire_4_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_4_bits_instructionIndex),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_4_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_4_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_4_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_4_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_4_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_4_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_4_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_4_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_4_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_4_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_4_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_4_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_4_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_4_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_4_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_4_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_4_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_4_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_4_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_4_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_4_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_4_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_4_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_4_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_4_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_4_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_4_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_4_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_4_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_4_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_4_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_4_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_4_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_4_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_4_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_4_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_4_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_4_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_4_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_4_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_4_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_4_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_4_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_4_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_4_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_4_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_4_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_4_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_4_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_4_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_4_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_4_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_4_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_4_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_4_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_4_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_4_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_4_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_4_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_4_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_4_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_4_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_4_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_4_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_4_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_4_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_4_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_4_maskUnitRequest_bits_ffo),
    .maskRequestToLSU                                    (_laneVec_4_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_4_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[4]),
    .vrfReadAddressChannel_ready                         (sinkWire_8_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_8_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_8_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_8_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_8_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_8_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_4_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_9_ready),
    .vrfWriteChannel_valid                               (sinkWire_9_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_9_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_9_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_9_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_9_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_9_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_9_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_4_valid_T),
    .instructionFinished                                 (_laneVec_4_instructionFinished),
    .vxsatReport                                         (_laneVec_4_vxsatReport),
    .v0Update_valid                                      (_laneVec_4_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_4_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_4_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_4_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_4_bits),
    .maskSelect                                          (_laneVec_4_maskSelect),
    .maskSelectSew                                       (_laneVec_4_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_4_bits | maskLastPipe_pipe_out_4_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_4),
    .writeCount                                          (pipe_out_9_bits),
    .writeQueueValid                                     (dataInWritePipeVec_4)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(13)
  ) sinkVec_queue_fifo_16 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_16_enq_ready & sinkVec_queue_16_enq_valid & ~(_sinkVec_queue_fifo_16_empty & sinkVec_queue_16_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_16_deq_ready & ~_sinkVec_queue_fifo_16_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_16),
    .empty        (_sinkVec_queue_fifo_16_empty),
    .almost_empty (sinkVec_queue_16_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_16_almostFull),
    .full         (_sinkVec_queue_fifo_16_full),
    .error        (_sinkVec_queue_fifo_16_error),
    .data_out     (_sinkVec_queue_fifo_16_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(13)
  ) sinkVec_queue_fifo_17 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_17_enq_ready & sinkVec_queue_17_enq_valid & ~(_sinkVec_queue_fifo_17_empty & sinkVec_queue_17_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_17_deq_ready & ~_sinkVec_queue_fifo_17_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_17),
    .empty        (_sinkVec_queue_fifo_17_empty),
    .almost_empty (sinkVec_queue_17_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_17_almostFull),
    .full         (_sinkVec_queue_fifo_17_full),
    .error        (_sinkVec_queue_fifo_17_error),
    .data_out     (_sinkVec_queue_fifo_17_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) sinkVec_queue_fifo_18 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_18_enq_ready & sinkVec_queue_18_enq_valid & ~(_sinkVec_queue_fifo_18_empty & sinkVec_queue_18_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_18_deq_ready & ~_sinkVec_queue_fifo_18_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_18),
    .empty        (_sinkVec_queue_fifo_18_empty),
    .almost_empty (sinkVec_queue_18_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_18_almostFull),
    .full         (_sinkVec_queue_fifo_18_full),
    .error        (_sinkVec_queue_fifo_18_error),
    .data_out     (_sinkVec_queue_fifo_18_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) sinkVec_queue_fifo_19 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_19_enq_ready & sinkVec_queue_19_enq_valid & ~(_sinkVec_queue_fifo_19_empty & sinkVec_queue_19_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_19_deq_ready & ~_sinkVec_queue_fifo_19_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_19),
    .empty        (_sinkVec_queue_fifo_19_empty),
    .almost_empty (sinkVec_queue_19_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_19_almostFull),
    .full         (_sinkVec_queue_fifo_19_full),
    .error        (_sinkVec_queue_fifo_19_error),
    .data_out     (_sinkVec_queue_fifo_19_data_out)
  );
  Lane laneVec_5 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (3'h5),
    .readBusPort_0_enq_valid                             (shifterReg_44_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_44_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_5_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_5_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_5_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_26_valid),
    .readBusPort_1_enq_valid                             (shifterReg_46_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_46_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_5_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_5_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_5_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_42_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_35_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_35_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_35_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_35_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_35_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_5_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_5_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_5_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_5_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_5_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_5_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_37_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_51_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_51_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_51_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_51_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_51_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_5_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_5_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_5_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_5_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_5_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_5_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_39_valid),
    .laneRequest_ready                                   (_laneVec_5_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_5_valid & laneRequestSinkWire_5_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_5_bits_instructionIndex),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_5_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_5_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_5_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_5_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_5_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_5_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_5_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_5_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_5_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_5_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_5_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_5_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_5_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_5_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_5_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_5_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_5_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_5_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_5_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_5_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_5_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_5_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_5_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_5_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_5_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_5_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_5_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_5_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_5_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_5_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_5_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_5_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_5_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_5_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_5_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_5_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_5_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_5_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_5_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_5_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_5_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_5_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_5_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_5_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_5_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_5_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_5_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_5_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_5_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_5_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_5_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_5_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_5_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_5_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_5_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_5_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_5_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_5_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_5_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_5_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_5_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_5_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_5_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_5_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_5_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_5_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_5_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_5_maskUnitRequest_bits_ffo),
    .maskRequestToLSU                                    (_laneVec_5_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_5_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[5]),
    .vrfReadAddressChannel_ready                         (sinkWire_10_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_10_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_10_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_10_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_10_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_10_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_5_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_11_ready),
    .vrfWriteChannel_valid                               (sinkWire_11_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_11_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_11_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_11_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_11_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_11_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_11_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_5_valid_T),
    .instructionFinished                                 (_laneVec_5_instructionFinished),
    .vxsatReport                                         (_laneVec_5_vxsatReport),
    .v0Update_valid                                      (_laneVec_5_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_5_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_5_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_5_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_5_bits),
    .maskSelect                                          (_laneVec_5_maskSelect),
    .maskSelectSew                                       (_laneVec_5_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_5_bits | maskLastPipe_pipe_out_5_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_5),
    .writeCount                                          (pipe_out_11_bits),
    .writeQueueValid                                     (dataInWritePipeVec_5)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(13)
  ) sinkVec_queue_fifo_20 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_20_enq_ready & sinkVec_queue_20_enq_valid & ~(_sinkVec_queue_fifo_20_empty & sinkVec_queue_20_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_20_deq_ready & ~_sinkVec_queue_fifo_20_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_20),
    .empty        (_sinkVec_queue_fifo_20_empty),
    .almost_empty (sinkVec_queue_20_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_20_almostFull),
    .full         (_sinkVec_queue_fifo_20_full),
    .error        (_sinkVec_queue_fifo_20_error),
    .data_out     (_sinkVec_queue_fifo_20_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(13)
  ) sinkVec_queue_fifo_21 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_21_enq_ready & sinkVec_queue_21_enq_valid & ~(_sinkVec_queue_fifo_21_empty & sinkVec_queue_21_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_21_deq_ready & ~_sinkVec_queue_fifo_21_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_21),
    .empty        (_sinkVec_queue_fifo_21_empty),
    .almost_empty (sinkVec_queue_21_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_21_almostFull),
    .full         (_sinkVec_queue_fifo_21_full),
    .error        (_sinkVec_queue_fifo_21_error),
    .data_out     (_sinkVec_queue_fifo_21_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) sinkVec_queue_fifo_22 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_22_enq_ready & sinkVec_queue_22_enq_valid & ~(_sinkVec_queue_fifo_22_empty & sinkVec_queue_22_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_22_deq_ready & ~_sinkVec_queue_fifo_22_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_22),
    .empty        (_sinkVec_queue_fifo_22_empty),
    .almost_empty (sinkVec_queue_22_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_22_almostFull),
    .full         (_sinkVec_queue_fifo_22_full),
    .error        (_sinkVec_queue_fifo_22_error),
    .data_out     (_sinkVec_queue_fifo_22_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) sinkVec_queue_fifo_23 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_23_enq_ready & sinkVec_queue_23_enq_valid & ~(_sinkVec_queue_fifo_23_empty & sinkVec_queue_23_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_23_deq_ready & ~_sinkVec_queue_fifo_23_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_23),
    .empty        (_sinkVec_queue_fifo_23_empty),
    .almost_empty (sinkVec_queue_23_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_23_almostFull),
    .full         (_sinkVec_queue_fifo_23_full),
    .error        (_sinkVec_queue_fifo_23_error),
    .data_out     (_sinkVec_queue_fifo_23_data_out)
  );
  Lane laneVec_6 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (3'h6),
    .readBusPort_0_enq_valid                             (shifterReg_48_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_48_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_6_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_6_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_6_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_28_valid),
    .readBusPort_1_enq_valid                             (shifterReg_50_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_50_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_6_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_6_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_6_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_44_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_37_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_37_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_37_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_37_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_37_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_6_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_6_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_6_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_6_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_6_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_6_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_41_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_53_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_53_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_53_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_53_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_53_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_6_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_6_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_6_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_6_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_6_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_6_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_43_valid),
    .laneRequest_ready                                   (_laneVec_6_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_6_valid & laneRequestSinkWire_6_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_6_bits_instructionIndex),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_6_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_6_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_6_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_6_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_6_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_6_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_6_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_6_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_6_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_6_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_6_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_6_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_6_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_6_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_6_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_6_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_6_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_6_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_6_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_6_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_6_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_6_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_6_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_6_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_6_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_6_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_6_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_6_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_6_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_6_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_6_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_6_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_6_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_6_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_6_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_6_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_6_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_6_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_6_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_6_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_6_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_6_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_6_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_6_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_6_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_6_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_6_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_6_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_6_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_6_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_6_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_6_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_6_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_6_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_6_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_6_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_6_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_6_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_6_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_6_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_6_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_6_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_6_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_6_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_6_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_6_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_6_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_6_maskUnitRequest_bits_ffo),
    .maskRequestToLSU                                    (_laneVec_6_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_6_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[6]),
    .vrfReadAddressChannel_ready                         (sinkWire_12_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_12_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_12_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_12_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_12_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_12_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_6_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_13_ready),
    .vrfWriteChannel_valid                               (sinkWire_13_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_13_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_13_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_13_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_13_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_13_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_13_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_6_valid_T),
    .instructionFinished                                 (_laneVec_6_instructionFinished),
    .vxsatReport                                         (_laneVec_6_vxsatReport),
    .v0Update_valid                                      (_laneVec_6_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_6_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_6_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_6_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_6_bits),
    .maskSelect                                          (_laneVec_6_maskSelect),
    .maskSelectSew                                       (_laneVec_6_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_6_bits | maskLastPipe_pipe_out_6_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_6),
    .writeCount                                          (pipe_out_13_bits),
    .writeQueueValid                                     (dataInWritePipeVec_6)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(13)
  ) sinkVec_queue_fifo_24 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_24_enq_ready & sinkVec_queue_24_enq_valid & ~(_sinkVec_queue_fifo_24_empty & sinkVec_queue_24_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_24_deq_ready & ~_sinkVec_queue_fifo_24_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_24),
    .empty        (_sinkVec_queue_fifo_24_empty),
    .almost_empty (sinkVec_queue_24_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_24_almostFull),
    .full         (_sinkVec_queue_fifo_24_full),
    .error        (_sinkVec_queue_fifo_24_error),
    .data_out     (_sinkVec_queue_fifo_24_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(13)
  ) sinkVec_queue_fifo_25 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_25_enq_ready & sinkVec_queue_25_enq_valid & ~(_sinkVec_queue_fifo_25_empty & sinkVec_queue_25_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_25_deq_ready & ~_sinkVec_queue_fifo_25_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_25),
    .empty        (_sinkVec_queue_fifo_25_empty),
    .almost_empty (sinkVec_queue_25_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_25_almostFull),
    .full         (_sinkVec_queue_fifo_25_full),
    .error        (_sinkVec_queue_fifo_25_error),
    .data_out     (_sinkVec_queue_fifo_25_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) sinkVec_queue_fifo_26 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_26_enq_ready & sinkVec_queue_26_enq_valid & ~(_sinkVec_queue_fifo_26_empty & sinkVec_queue_26_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_26_deq_ready & ~_sinkVec_queue_fifo_26_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_26),
    .empty        (_sinkVec_queue_fifo_26_empty),
    .almost_empty (sinkVec_queue_26_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_26_almostFull),
    .full         (_sinkVec_queue_fifo_26_full),
    .error        (_sinkVec_queue_fifo_26_error),
    .data_out     (_sinkVec_queue_fifo_26_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) sinkVec_queue_fifo_27 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_27_enq_ready & sinkVec_queue_27_enq_valid & ~(_sinkVec_queue_fifo_27_empty & sinkVec_queue_27_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_27_deq_ready & ~_sinkVec_queue_fifo_27_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_27),
    .empty        (_sinkVec_queue_fifo_27_empty),
    .almost_empty (sinkVec_queue_27_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_27_almostFull),
    .full         (_sinkVec_queue_fifo_27_full),
    .error        (_sinkVec_queue_fifo_27_error),
    .data_out     (_sinkVec_queue_fifo_27_data_out)
  );
  Lane laneVec_7 (
    .clock                                               (clock),
    .reset                                               (reset),
    .laneIndex                                           (3'h7),
    .readBusPort_0_enq_valid                             (shifterReg_52_0_valid),
    .readBusPort_0_enq_bits_data                         (shifterReg_52_0_bits_data),
    .readBusPort_0_enqRelease                            (_laneVec_7_readBusPort_0_enqRelease),
    .readBusPort_0_deq_valid                             (_laneVec_7_readBusPort_0_deq_valid),
    .readBusPort_0_deq_bits_data                         (_laneVec_7_readBusPort_0_deq_bits_data),
    .readBusPort_0_deqRelease                            (pipe_out_30_valid),
    .readBusPort_1_enq_valid                             (shifterReg_54_0_valid),
    .readBusPort_1_enq_bits_data                         (shifterReg_54_0_bits_data),
    .readBusPort_1_enqRelease                            (_laneVec_7_readBusPort_1_enqRelease),
    .readBusPort_1_deq_valid                             (_laneVec_7_readBusPort_1_deq_valid),
    .readBusPort_1_deq_bits_data                         (_laneVec_7_readBusPort_1_deq_bits_data),
    .readBusPort_1_deqRelease                            (pipe_out_46_valid),
    .writeBusPort_0_enq_valid                            (shifterReg_39_0_valid),
    .writeBusPort_0_enq_bits_data                        (shifterReg_39_0_bits_data),
    .writeBusPort_0_enq_bits_mask                        (shifterReg_39_0_bits_mask),
    .writeBusPort_0_enq_bits_instructionIndex            (shifterReg_39_0_bits_instructionIndex),
    .writeBusPort_0_enq_bits_counter                     (shifterReg_39_0_bits_counter),
    .writeBusPort_0_enqRelease                           (_laneVec_7_writeBusPort_0_enqRelease),
    .writeBusPort_0_deq_valid                            (_laneVec_7_writeBusPort_0_deq_valid),
    .writeBusPort_0_deq_bits_data                        (_laneVec_7_writeBusPort_0_deq_bits_data),
    .writeBusPort_0_deq_bits_mask                        (_laneVec_7_writeBusPort_0_deq_bits_mask),
    .writeBusPort_0_deq_bits_instructionIndex            (_laneVec_7_writeBusPort_0_deq_bits_instructionIndex),
    .writeBusPort_0_deq_bits_counter                     (_laneVec_7_writeBusPort_0_deq_bits_counter),
    .writeBusPort_0_deqRelease                           (pipe_out_45_valid),
    .writeBusPort_1_enq_valid                            (shifterReg_55_0_valid),
    .writeBusPort_1_enq_bits_data                        (shifterReg_55_0_bits_data),
    .writeBusPort_1_enq_bits_mask                        (shifterReg_55_0_bits_mask),
    .writeBusPort_1_enq_bits_instructionIndex            (shifterReg_55_0_bits_instructionIndex),
    .writeBusPort_1_enq_bits_counter                     (shifterReg_55_0_bits_counter),
    .writeBusPort_1_enqRelease                           (_laneVec_7_writeBusPort_1_enqRelease),
    .writeBusPort_1_deq_valid                            (_laneVec_7_writeBusPort_1_deq_valid),
    .writeBusPort_1_deq_bits_data                        (_laneVec_7_writeBusPort_1_deq_bits_data),
    .writeBusPort_1_deq_bits_mask                        (_laneVec_7_writeBusPort_1_deq_bits_mask),
    .writeBusPort_1_deq_bits_instructionIndex            (_laneVec_7_writeBusPort_1_deq_bits_instructionIndex),
    .writeBusPort_1_deq_bits_counter                     (_laneVec_7_writeBusPort_1_deq_bits_counter),
    .writeBusPort_1_deqRelease                           (pipe_out_47_valid),
    .laneRequest_ready                                   (_laneVec_7_laneRequest_ready),
    .laneRequest_valid                                   (laneRequestSinkWire_7_valid & laneRequestSinkWire_7_bits_issueInst),
    .laneRequest_bits_instructionIndex                   (laneRequestSinkWire_7_bits_instructionIndex),
    .laneRequest_bits_decodeResult_specialSlot           (laneRequestSinkWire_7_bits_decodeResult_specialSlot),
    .laneRequest_bits_decodeResult_topUop                (laneRequestSinkWire_7_bits_decodeResult_topUop),
    .laneRequest_bits_decodeResult_popCount              (laneRequestSinkWire_7_bits_decodeResult_popCount),
    .laneRequest_bits_decodeResult_ffo                   (laneRequestSinkWire_7_bits_decodeResult_ffo),
    .laneRequest_bits_decodeResult_average               (laneRequestSinkWire_7_bits_decodeResult_average),
    .laneRequest_bits_decodeResult_reverse               (laneRequestSinkWire_7_bits_decodeResult_reverse),
    .laneRequest_bits_decodeResult_dontNeedExecuteInLane (laneRequestSinkWire_7_bits_decodeResult_dontNeedExecuteInLane),
    .laneRequest_bits_decodeResult_scheduler             (laneRequestSinkWire_7_bits_decodeResult_scheduler),
    .laneRequest_bits_decodeResult_sReadVD               (laneRequestSinkWire_7_bits_decodeResult_sReadVD),
    .laneRequest_bits_decodeResult_vtype                 (laneRequestSinkWire_7_bits_decodeResult_vtype),
    .laneRequest_bits_decodeResult_sWrite                (laneRequestSinkWire_7_bits_decodeResult_sWrite),
    .laneRequest_bits_decodeResult_crossRead             (laneRequestSinkWire_7_bits_decodeResult_crossRead),
    .laneRequest_bits_decodeResult_crossWrite            (laneRequestSinkWire_7_bits_decodeResult_crossWrite),
    .laneRequest_bits_decodeResult_maskUnit              (laneRequestSinkWire_7_bits_decodeResult_maskUnit),
    .laneRequest_bits_decodeResult_special               (laneRequestSinkWire_7_bits_decodeResult_special),
    .laneRequest_bits_decodeResult_saturate              (laneRequestSinkWire_7_bits_decodeResult_saturate),
    .laneRequest_bits_decodeResult_vwmacc                (laneRequestSinkWire_7_bits_decodeResult_vwmacc),
    .laneRequest_bits_decodeResult_readOnly              (laneRequestSinkWire_7_bits_decodeResult_readOnly),
    .laneRequest_bits_decodeResult_maskSource            (laneRequestSinkWire_7_bits_decodeResult_maskSource),
    .laneRequest_bits_decodeResult_maskDestination       (laneRequestSinkWire_7_bits_decodeResult_maskDestination),
    .laneRequest_bits_decodeResult_maskLogic             (laneRequestSinkWire_7_bits_decodeResult_maskLogic),
    .laneRequest_bits_decodeResult_uop                   (laneRequestSinkWire_7_bits_decodeResult_uop),
    .laneRequest_bits_decodeResult_iota                  (laneRequestSinkWire_7_bits_decodeResult_iota),
    .laneRequest_bits_decodeResult_mv                    (laneRequestSinkWire_7_bits_decodeResult_mv),
    .laneRequest_bits_decodeResult_extend                (laneRequestSinkWire_7_bits_decodeResult_extend),
    .laneRequest_bits_decodeResult_unOrderWrite          (laneRequestSinkWire_7_bits_decodeResult_unOrderWrite),
    .laneRequest_bits_decodeResult_compress              (laneRequestSinkWire_7_bits_decodeResult_compress),
    .laneRequest_bits_decodeResult_gather16              (laneRequestSinkWire_7_bits_decodeResult_gather16),
    .laneRequest_bits_decodeResult_gather                (laneRequestSinkWire_7_bits_decodeResult_gather),
    .laneRequest_bits_decodeResult_slid                  (laneRequestSinkWire_7_bits_decodeResult_slid),
    .laneRequest_bits_decodeResult_targetRd              (laneRequestSinkWire_7_bits_decodeResult_targetRd),
    .laneRequest_bits_decodeResult_widenReduce           (laneRequestSinkWire_7_bits_decodeResult_widenReduce),
    .laneRequest_bits_decodeResult_red                   (laneRequestSinkWire_7_bits_decodeResult_red),
    .laneRequest_bits_decodeResult_nr                    (laneRequestSinkWire_7_bits_decodeResult_nr),
    .laneRequest_bits_decodeResult_itype                 (laneRequestSinkWire_7_bits_decodeResult_itype),
    .laneRequest_bits_decodeResult_unsigned1             (laneRequestSinkWire_7_bits_decodeResult_unsigned1),
    .laneRequest_bits_decodeResult_unsigned0             (laneRequestSinkWire_7_bits_decodeResult_unsigned0),
    .laneRequest_bits_decodeResult_other                 (laneRequestSinkWire_7_bits_decodeResult_other),
    .laneRequest_bits_decodeResult_multiCycle            (laneRequestSinkWire_7_bits_decodeResult_multiCycle),
    .laneRequest_bits_decodeResult_divider               (laneRequestSinkWire_7_bits_decodeResult_divider),
    .laneRequest_bits_decodeResult_multiplier            (laneRequestSinkWire_7_bits_decodeResult_multiplier),
    .laneRequest_bits_decodeResult_shift                 (laneRequestSinkWire_7_bits_decodeResult_shift),
    .laneRequest_bits_decodeResult_adder                 (laneRequestSinkWire_7_bits_decodeResult_adder),
    .laneRequest_bits_decodeResult_logic                 (laneRequestSinkWire_7_bits_decodeResult_logic),
    .laneRequest_bits_loadStore                          (laneRequestSinkWire_7_bits_loadStore),
    .laneRequest_bits_issueInst                          (laneVec_7_laneRequest_bits_issueInst),
    .laneRequest_bits_store                              (laneRequestSinkWire_7_bits_store),
    .laneRequest_bits_special                            (laneRequestSinkWire_7_bits_special),
    .laneRequest_bits_lsWholeReg                         (laneRequestSinkWire_7_bits_lsWholeReg),
    .laneRequest_bits_vs1                                (laneRequestSinkWire_7_bits_vs1),
    .laneRequest_bits_vs2                                (laneRequestSinkWire_7_bits_vs2),
    .laneRequest_bits_vd                                 (laneRequestSinkWire_7_bits_vd),
    .laneRequest_bits_loadStoreEEW                       (laneRequestSinkWire_7_bits_loadStoreEEW),
    .laneRequest_bits_mask                               (laneRequestSinkWire_7_bits_mask),
    .laneRequest_bits_segment                            (laneRequestSinkWire_7_bits_segment),
    .laneRequest_bits_readFromScalar                     (laneRequestSinkWire_7_bits_readFromScalar),
    .laneRequest_bits_csrInterface_vl                    (laneRequestSinkWire_7_bits_csrInterface_vl),
    .laneRequest_bits_csrInterface_vStart                (laneRequestSinkWire_7_bits_csrInterface_vStart),
    .laneRequest_bits_csrInterface_vlmul                 (laneRequestSinkWire_7_bits_csrInterface_vlmul),
    .laneRequest_bits_csrInterface_vSew                  (laneRequestSinkWire_7_bits_csrInterface_vSew),
    .laneRequest_bits_csrInterface_vxrm                  (laneRequestSinkWire_7_bits_csrInterface_vxrm),
    .laneRequest_bits_csrInterface_vta                   (laneRequestSinkWire_7_bits_csrInterface_vta),
    .laneRequest_bits_csrInterface_vma                   (laneRequestSinkWire_7_bits_csrInterface_vma),
    .maskUnitRequest_valid                               (_laneVec_7_maskUnitRequest_valid),
    .maskUnitRequest_bits_source1                        (_laneVec_7_maskUnitRequest_bits_source1),
    .maskUnitRequest_bits_source2                        (_laneVec_7_maskUnitRequest_bits_source2),
    .maskUnitRequest_bits_index                          (_laneVec_7_maskUnitRequest_bits_index),
    .maskUnitRequest_bits_ffo                            (_laneVec_7_maskUnitRequest_bits_ffo),
    .maskRequestToLSU                                    (_laneVec_7_maskRequestToLSU),
    .tokenIO_maskRequestRelease                          (_maskUnit_tokenIO_7_maskRequestRelease | _lsu_tokenIO_offsetGroupRelease[7]),
    .vrfReadAddressChannel_ready                         (sinkWire_14_ready),
    .vrfReadAddressChannel_valid                         (sinkWire_14_valid),
    .vrfReadAddressChannel_bits_vs                       (sinkWire_14_bits_vs),
    .vrfReadAddressChannel_bits_readSource               (sinkWire_14_bits_readSource),
    .vrfReadAddressChannel_bits_offset                   (sinkWire_14_bits_offset),
    .vrfReadAddressChannel_bits_instructionIndex         (sinkWire_14_bits_instructionIndex),
    .vrfReadDataChannel                                  (_laneVec_7_vrfReadDataChannel),
    .vrfWriteChannel_ready                               (sinkWire_15_ready),
    .vrfWriteChannel_valid                               (sinkWire_15_valid),
    .vrfWriteChannel_bits_vd                             (sinkWire_15_bits_vd),
    .vrfWriteChannel_bits_offset                         (sinkWire_15_bits_offset),
    .vrfWriteChannel_bits_mask                           (sinkWire_15_bits_mask),
    .vrfWriteChannel_bits_data                           (sinkWire_15_bits_data),
    .vrfWriteChannel_bits_last                           (sinkWire_15_bits_last),
    .vrfWriteChannel_bits_instructionIndex               (sinkWire_15_bits_instructionIndex),
    .writeFromMask                                       (_probeWire_writeQueueEnqVec_7_valid_T),
    .instructionFinished                                 (_laneVec_7_instructionFinished),
    .vxsatReport                                         (_laneVec_7_vxsatReport),
    .v0Update_valid                                      (_laneVec_7_v0Update_valid),
    .v0Update_bits_data                                  (_laneVec_7_v0Update_bits_data),
    .v0Update_bits_offset                                (_laneVec_7_v0Update_bits_offset),
    .v0Update_bits_mask                                  (_laneVec_7_v0Update_bits_mask),
    .maskInput                                           (pipe_pipe_out_7_bits),
    .maskSelect                                          (_laneVec_7_maskSelect),
    .maskSelectSew                                       (_laneVec_7_maskSelectSew),
    .lsuLastReport                                       (lsuLastPipe_pipe_out_7_bits | maskLastPipe_pipe_out_7_bits),
    .loadDataInLSUWriteQueue                             (_lsu_dataInWriteQueue_7),
    .writeCount                                          (pipe_out_15_bits),
    .writeQueueValid                                     (dataInWritePipeVec_7)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(13)
  ) sinkVec_queue_fifo_28 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_28_enq_ready & sinkVec_queue_28_enq_valid & ~(_sinkVec_queue_fifo_28_empty & sinkVec_queue_28_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_28_deq_ready & ~_sinkVec_queue_fifo_28_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_28),
    .empty        (_sinkVec_queue_fifo_28_empty),
    .almost_empty (sinkVec_queue_28_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_28_almostFull),
    .full         (_sinkVec_queue_fifo_28_full),
    .error        (_sinkVec_queue_fifo_28_error),
    .data_out     (_sinkVec_queue_fifo_28_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(13)
  ) sinkVec_queue_fifo_29 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_29_enq_ready & sinkVec_queue_29_enq_valid & ~(_sinkVec_queue_fifo_29_empty & sinkVec_queue_29_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_29_deq_ready & ~_sinkVec_queue_fifo_29_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_29),
    .empty        (_sinkVec_queue_fifo_29_empty),
    .almost_empty (sinkVec_queue_29_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_29_almostFull),
    .full         (_sinkVec_queue_fifo_29_full),
    .error        (_sinkVec_queue_fifo_29_error),
    .data_out     (_sinkVec_queue_fifo_29_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) sinkVec_queue_fifo_30 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_30_enq_ready & sinkVec_queue_30_enq_valid & ~(_sinkVec_queue_fifo_30_empty & sinkVec_queue_30_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_30_deq_ready & ~_sinkVec_queue_fifo_30_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_30),
    .empty        (_sinkVec_queue_fifo_30_empty),
    .almost_empty (sinkVec_queue_30_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_30_almostFull),
    .full         (_sinkVec_queue_fifo_30_full),
    .error        (_sinkVec_queue_fifo_30_error),
    .data_out     (_sinkVec_queue_fifo_30_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) sinkVec_queue_fifo_31 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sinkVec_queue_31_enq_ready & sinkVec_queue_31_enq_valid & ~(_sinkVec_queue_fifo_31_empty & sinkVec_queue_31_deq_ready))),
    .pop_req_n    (~(sinkVec_queue_31_deq_ready & ~_sinkVec_queue_fifo_31_empty)),
    .diag_n       (1'h1),
    .data_in      (sinkVec_queue_dataIn_31),
    .empty        (_sinkVec_queue_fifo_31_empty),
    .almost_empty (sinkVec_queue_31_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sinkVec_queue_31_almostFull),
    .full         (_sinkVec_queue_fifo_31_full),
    .error        (_sinkVec_queue_fifo_31_error),
    .data_out     (_sinkVec_queue_fifo_31_data_out)
  );
  assign indexedLoadStorePort_aw_valid = indexedLoadStorePort_aw_valid_0;
  assign indexedLoadStorePort_aw_bits_id = indexedLoadStorePort_aw_bits_id_0;
  assign indexedLoadStorePort_aw_bits_addr = indexedLoadStorePort_aw_bits_addr_0;
  assign indexedLoadStorePort_aw_bits_len = 8'h0;
  assign indexedLoadStorePort_aw_bits_size = indexedLoadStorePort_aw_bits_size_0;
  assign indexedLoadStorePort_aw_bits_burst = 2'h1;
  assign indexedLoadStorePort_aw_bits_lock = 1'h0;
  assign indexedLoadStorePort_aw_bits_cache = 4'h0;
  assign indexedLoadStorePort_aw_bits_prot = 3'h0;
  assign indexedLoadStorePort_aw_bits_qos = 4'h0;
  assign indexedLoadStorePort_aw_bits_region = 4'h0;
  assign indexedLoadStorePort_w_valid = indexedLoadStorePort_w_valid_0;
  assign indexedLoadStorePort_w_bits_data = indexedLoadStorePort_w_bits_data_0;
  assign indexedLoadStorePort_w_bits_strb = indexedLoadStorePort_w_bits_strb_0;
  assign indexedLoadStorePort_w_bits_last = 1'h1;
  assign indexedLoadStorePort_b_ready = 1'h1;
  assign indexedLoadStorePort_ar_valid = indexedLoadStorePort_ar_valid_0;
  assign indexedLoadStorePort_ar_bits_id = 2'h0;
  assign indexedLoadStorePort_ar_bits_addr = indexedLoadStorePort_ar_bits_addr_0;
  assign indexedLoadStorePort_ar_bits_len = 8'h0;
  assign indexedLoadStorePort_ar_bits_size = 3'h2;
  assign indexedLoadStorePort_ar_bits_burst = 2'h1;
  assign indexedLoadStorePort_ar_bits_lock = 1'h0;
  assign indexedLoadStorePort_ar_bits_cache = 4'h0;
  assign indexedLoadStorePort_ar_bits_prot = 3'h0;
  assign indexedLoadStorePort_ar_bits_qos = 4'h0;
  assign indexedLoadStorePort_ar_bits_region = 4'h0;
  assign indexedLoadStorePort_r_ready = indexedLoadStorePort_r_ready_0;
  assign highBandwidthLoadStorePort_aw_valid = highBandwidthLoadStorePort_aw_valid_0;
  assign highBandwidthLoadStorePort_aw_bits_id = highBandwidthLoadStorePort_aw_bits_id_0;
  assign highBandwidthLoadStorePort_aw_bits_addr = highBandwidthLoadStorePort_aw_bits_addr_0;
  assign highBandwidthLoadStorePort_aw_bits_len = 8'h0;
  assign highBandwidthLoadStorePort_aw_bits_size = 3'h5;
  assign highBandwidthLoadStorePort_aw_bits_burst = 2'h1;
  assign highBandwidthLoadStorePort_aw_bits_lock = 1'h0;
  assign highBandwidthLoadStorePort_aw_bits_cache = 4'h0;
  assign highBandwidthLoadStorePort_aw_bits_prot = 3'h0;
  assign highBandwidthLoadStorePort_aw_bits_qos = 4'h0;
  assign highBandwidthLoadStorePort_aw_bits_region = 4'h0;
  assign highBandwidthLoadStorePort_w_valid = highBandwidthLoadStorePort_w_valid_0;
  assign highBandwidthLoadStorePort_w_bits_data = highBandwidthLoadStorePort_w_bits_data_0;
  assign highBandwidthLoadStorePort_w_bits_strb = highBandwidthLoadStorePort_w_bits_strb_0;
  assign highBandwidthLoadStorePort_w_bits_last = 1'h1;
  assign highBandwidthLoadStorePort_b_ready = 1'h1;
  assign highBandwidthLoadStorePort_ar_valid = highBandwidthLoadStorePort_ar_valid_0;
  assign highBandwidthLoadStorePort_ar_bits_id = 2'h0;
  assign highBandwidthLoadStorePort_ar_bits_addr = highBandwidthLoadStorePort_ar_bits_addr_0;
  assign highBandwidthLoadStorePort_ar_bits_len = 8'h0;
  assign highBandwidthLoadStorePort_ar_bits_size = 3'h5;
  assign highBandwidthLoadStorePort_ar_bits_burst = 2'h1;
  assign highBandwidthLoadStorePort_ar_bits_lock = 1'h0;
  assign highBandwidthLoadStorePort_ar_bits_cache = 4'h0;
  assign highBandwidthLoadStorePort_ar_bits_prot = 3'h0;
  assign highBandwidthLoadStorePort_ar_bits_qos = 4'h0;
  assign highBandwidthLoadStorePort_ar_bits_region = 4'h0;
  assign highBandwidthLoadStorePort_r_ready = highBandwidthLoadStorePort_r_ready_0;
  assign retire_rd_valid = retire_rd_valid_0;
  assign retire_rd_bits_rdAddress = retire_rd_bits_rdAddress_0;
  assign retire_rd_bits_rdData = retire_rd_bits_rdData_0;
  assign retire_rd_bits_isFp = 1'h0;
  assign retire_csr_valid = 1'h0;
  assign retire_csr_bits_vxsat = retire_csr_bits_vxsat_0;
  assign retire_csr_bits_fflag = 32'h0;
  assign retire_mem_valid = retire_mem_valid_0;
  assign issue_ready = issue_ready_0;
endmodule

