
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module LSU(
  input           clock,
                  reset,
  output          request_ready,
  input           request_valid,
  input  [2:0]    request_bits_instructionInformation_nf,
  input           request_bits_instructionInformation_mew,
  input  [1:0]    request_bits_instructionInformation_mop,
  input  [4:0]    request_bits_instructionInformation_lumop,
  input  [1:0]    request_bits_instructionInformation_eew,
  input  [4:0]    request_bits_instructionInformation_vs3,
  input           request_bits_instructionInformation_isStore,
                  request_bits_instructionInformation_maskedLoadStore,
  input  [31:0]   request_bits_rs1Data,
                  request_bits_rs2Data,
  input  [2:0]    request_bits_instructionIndex,
  input           v0UpdateVec_0_valid,
  input  [31:0]   v0UpdateVec_0_bits_data,
  input  [3:0]    v0UpdateVec_0_bits_mask,
  input           v0UpdateVec_1_valid,
  input  [31:0]   v0UpdateVec_1_bits_data,
  input  [3:0]    v0UpdateVec_1_bits_mask,
  input           v0UpdateVec_2_valid,
  input  [31:0]   v0UpdateVec_2_bits_data,
  input  [3:0]    v0UpdateVec_2_bits_mask,
  input           v0UpdateVec_3_valid,
  input  [31:0]   v0UpdateVec_3_bits_data,
  input  [3:0]    v0UpdateVec_3_bits_mask,
  input           v0UpdateVec_4_valid,
  input  [31:0]   v0UpdateVec_4_bits_data,
  input  [3:0]    v0UpdateVec_4_bits_mask,
  input           v0UpdateVec_5_valid,
  input  [31:0]   v0UpdateVec_5_bits_data,
  input  [3:0]    v0UpdateVec_5_bits_mask,
  input           v0UpdateVec_6_valid,
  input  [31:0]   v0UpdateVec_6_bits_data,
  input  [3:0]    v0UpdateVec_6_bits_mask,
  input           v0UpdateVec_7_valid,
  input  [31:0]   v0UpdateVec_7_bits_data,
  input  [3:0]    v0UpdateVec_7_bits_mask,
  input           v0UpdateVec_8_valid,
  input  [31:0]   v0UpdateVec_8_bits_data,
  input  [3:0]    v0UpdateVec_8_bits_mask,
  input           v0UpdateVec_9_valid,
  input  [31:0]   v0UpdateVec_9_bits_data,
  input  [3:0]    v0UpdateVec_9_bits_mask,
  input           v0UpdateVec_10_valid,
  input  [31:0]   v0UpdateVec_10_bits_data,
  input  [3:0]    v0UpdateVec_10_bits_mask,
  input           v0UpdateVec_11_valid,
  input  [31:0]   v0UpdateVec_11_bits_data,
  input  [3:0]    v0UpdateVec_11_bits_mask,
  input           v0UpdateVec_12_valid,
  input  [31:0]   v0UpdateVec_12_bits_data,
  input  [3:0]    v0UpdateVec_12_bits_mask,
  input           v0UpdateVec_13_valid,
  input  [31:0]   v0UpdateVec_13_bits_data,
  input  [3:0]    v0UpdateVec_13_bits_mask,
  input           v0UpdateVec_14_valid,
  input  [31:0]   v0UpdateVec_14_bits_data,
  input  [3:0]    v0UpdateVec_14_bits_mask,
  input           v0UpdateVec_15_valid,
  input  [31:0]   v0UpdateVec_15_bits_data,
  input  [3:0]    v0UpdateVec_15_bits_mask,
  input           v0UpdateVec_16_valid,
  input  [31:0]   v0UpdateVec_16_bits_data,
  input  [3:0]    v0UpdateVec_16_bits_mask,
  input           v0UpdateVec_17_valid,
  input  [31:0]   v0UpdateVec_17_bits_data,
  input  [3:0]    v0UpdateVec_17_bits_mask,
  input           v0UpdateVec_18_valid,
  input  [31:0]   v0UpdateVec_18_bits_data,
  input  [3:0]    v0UpdateVec_18_bits_mask,
  input           v0UpdateVec_19_valid,
  input  [31:0]   v0UpdateVec_19_bits_data,
  input  [3:0]    v0UpdateVec_19_bits_mask,
  input           v0UpdateVec_20_valid,
  input  [31:0]   v0UpdateVec_20_bits_data,
  input  [3:0]    v0UpdateVec_20_bits_mask,
  input           v0UpdateVec_21_valid,
  input  [31:0]   v0UpdateVec_21_bits_data,
  input  [3:0]    v0UpdateVec_21_bits_mask,
  input           v0UpdateVec_22_valid,
  input  [31:0]   v0UpdateVec_22_bits_data,
  input  [3:0]    v0UpdateVec_22_bits_mask,
  input           v0UpdateVec_23_valid,
  input  [31:0]   v0UpdateVec_23_bits_data,
  input  [3:0]    v0UpdateVec_23_bits_mask,
  input           v0UpdateVec_24_valid,
  input  [31:0]   v0UpdateVec_24_bits_data,
  input  [3:0]    v0UpdateVec_24_bits_mask,
  input           v0UpdateVec_25_valid,
  input  [31:0]   v0UpdateVec_25_bits_data,
  input  [3:0]    v0UpdateVec_25_bits_mask,
  input           v0UpdateVec_26_valid,
  input  [31:0]   v0UpdateVec_26_bits_data,
  input  [3:0]    v0UpdateVec_26_bits_mask,
  input           v0UpdateVec_27_valid,
  input  [31:0]   v0UpdateVec_27_bits_data,
  input  [3:0]    v0UpdateVec_27_bits_mask,
  input           v0UpdateVec_28_valid,
  input  [31:0]   v0UpdateVec_28_bits_data,
  input  [3:0]    v0UpdateVec_28_bits_mask,
  input           v0UpdateVec_29_valid,
  input  [31:0]   v0UpdateVec_29_bits_data,
  input  [3:0]    v0UpdateVec_29_bits_mask,
  input           v0UpdateVec_30_valid,
  input  [31:0]   v0UpdateVec_30_bits_data,
  input  [3:0]    v0UpdateVec_30_bits_mask,
  input           v0UpdateVec_31_valid,
  input  [31:0]   v0UpdateVec_31_bits_data,
  input  [3:0]    v0UpdateVec_31_bits_mask,
  input           axi4Port_aw_ready,
  output          axi4Port_aw_valid,
  output [1:0]    axi4Port_aw_bits_id,
  output [31:0]   axi4Port_aw_bits_addr,
  input           axi4Port_w_ready,
  output          axi4Port_w_valid,
  output [1023:0] axi4Port_w_bits_data,
  output [127:0]  axi4Port_w_bits_strb,
  input           axi4Port_b_valid,
  input  [1:0]    axi4Port_b_bits_id,
                  axi4Port_b_bits_resp,
  input           axi4Port_ar_ready,
  output          axi4Port_ar_valid,
  output [31:0]   axi4Port_ar_bits_addr,
  output          axi4Port_r_ready,
  input           axi4Port_r_valid,
  input  [1:0]    axi4Port_r_bits_id,
  input  [1023:0] axi4Port_r_bits_data,
  input  [1:0]    axi4Port_r_bits_resp,
  input           axi4Port_r_bits_last,
                  simpleAccessPorts_aw_ready,
  output          simpleAccessPorts_aw_valid,
  output [1:0]    simpleAccessPorts_aw_bits_id,
  output [31:0]   simpleAccessPorts_aw_bits_addr,
  output [2:0]    simpleAccessPorts_aw_bits_size,
  input           simpleAccessPorts_w_ready,
  output          simpleAccessPorts_w_valid,
  output [31:0]   simpleAccessPorts_w_bits_data,
  output [3:0]    simpleAccessPorts_w_bits_strb,
  input           simpleAccessPorts_b_valid,
  input  [1:0]    simpleAccessPorts_b_bits_id,
                  simpleAccessPorts_b_bits_resp,
  input           simpleAccessPorts_ar_ready,
  output          simpleAccessPorts_ar_valid,
  output [31:0]   simpleAccessPorts_ar_bits_addr,
  output          simpleAccessPorts_r_ready,
  input           simpleAccessPorts_r_valid,
  input  [1:0]    simpleAccessPorts_r_bits_id,
  input  [31:0]   simpleAccessPorts_r_bits_data,
  input  [1:0]    simpleAccessPorts_r_bits_resp,
  input           simpleAccessPorts_r_bits_last,
                  vrfReadDataPorts_0_ready,
  output          vrfReadDataPorts_0_valid,
  output [4:0]    vrfReadDataPorts_0_bits_vs,
  output [2:0]    vrfReadDataPorts_0_bits_instructionIndex,
  input           vrfReadDataPorts_1_ready,
  output          vrfReadDataPorts_1_valid,
  output [4:0]    vrfReadDataPorts_1_bits_vs,
  output [2:0]    vrfReadDataPorts_1_bits_instructionIndex,
  input           vrfReadDataPorts_2_ready,
  output          vrfReadDataPorts_2_valid,
  output [4:0]    vrfReadDataPorts_2_bits_vs,
  output [2:0]    vrfReadDataPorts_2_bits_instructionIndex,
  input           vrfReadDataPorts_3_ready,
  output          vrfReadDataPorts_3_valid,
  output [4:0]    vrfReadDataPorts_3_bits_vs,
  output [2:0]    vrfReadDataPorts_3_bits_instructionIndex,
  input           vrfReadDataPorts_4_ready,
  output          vrfReadDataPorts_4_valid,
  output [4:0]    vrfReadDataPorts_4_bits_vs,
  output [2:0]    vrfReadDataPorts_4_bits_instructionIndex,
  input           vrfReadDataPorts_5_ready,
  output          vrfReadDataPorts_5_valid,
  output [4:0]    vrfReadDataPorts_5_bits_vs,
  output [2:0]    vrfReadDataPorts_5_bits_instructionIndex,
  input           vrfReadDataPorts_6_ready,
  output          vrfReadDataPorts_6_valid,
  output [4:0]    vrfReadDataPorts_6_bits_vs,
  output [2:0]    vrfReadDataPorts_6_bits_instructionIndex,
  input           vrfReadDataPorts_7_ready,
  output          vrfReadDataPorts_7_valid,
  output [4:0]    vrfReadDataPorts_7_bits_vs,
  output [2:0]    vrfReadDataPorts_7_bits_instructionIndex,
  input           vrfReadDataPorts_8_ready,
  output          vrfReadDataPorts_8_valid,
  output [4:0]    vrfReadDataPorts_8_bits_vs,
  output [2:0]    vrfReadDataPorts_8_bits_instructionIndex,
  input           vrfReadDataPorts_9_ready,
  output          vrfReadDataPorts_9_valid,
  output [4:0]    vrfReadDataPorts_9_bits_vs,
  output [2:0]    vrfReadDataPorts_9_bits_instructionIndex,
  input           vrfReadDataPorts_10_ready,
  output          vrfReadDataPorts_10_valid,
  output [4:0]    vrfReadDataPorts_10_bits_vs,
  output [2:0]    vrfReadDataPorts_10_bits_instructionIndex,
  input           vrfReadDataPorts_11_ready,
  output          vrfReadDataPorts_11_valid,
  output [4:0]    vrfReadDataPorts_11_bits_vs,
  output [2:0]    vrfReadDataPorts_11_bits_instructionIndex,
  input           vrfReadDataPorts_12_ready,
  output          vrfReadDataPorts_12_valid,
  output [4:0]    vrfReadDataPorts_12_bits_vs,
  output [2:0]    vrfReadDataPorts_12_bits_instructionIndex,
  input           vrfReadDataPorts_13_ready,
  output          vrfReadDataPorts_13_valid,
  output [4:0]    vrfReadDataPorts_13_bits_vs,
  output [2:0]    vrfReadDataPorts_13_bits_instructionIndex,
  input           vrfReadDataPorts_14_ready,
  output          vrfReadDataPorts_14_valid,
  output [4:0]    vrfReadDataPorts_14_bits_vs,
  output [2:0]    vrfReadDataPorts_14_bits_instructionIndex,
  input           vrfReadDataPorts_15_ready,
  output          vrfReadDataPorts_15_valid,
  output [4:0]    vrfReadDataPorts_15_bits_vs,
  output [2:0]    vrfReadDataPorts_15_bits_instructionIndex,
  input           vrfReadDataPorts_16_ready,
  output          vrfReadDataPorts_16_valid,
  output [4:0]    vrfReadDataPorts_16_bits_vs,
  output [2:0]    vrfReadDataPorts_16_bits_instructionIndex,
  input           vrfReadDataPorts_17_ready,
  output          vrfReadDataPorts_17_valid,
  output [4:0]    vrfReadDataPorts_17_bits_vs,
  output [2:0]    vrfReadDataPorts_17_bits_instructionIndex,
  input           vrfReadDataPorts_18_ready,
  output          vrfReadDataPorts_18_valid,
  output [4:0]    vrfReadDataPorts_18_bits_vs,
  output [2:0]    vrfReadDataPorts_18_bits_instructionIndex,
  input           vrfReadDataPorts_19_ready,
  output          vrfReadDataPorts_19_valid,
  output [4:0]    vrfReadDataPorts_19_bits_vs,
  output [2:0]    vrfReadDataPorts_19_bits_instructionIndex,
  input           vrfReadDataPorts_20_ready,
  output          vrfReadDataPorts_20_valid,
  output [4:0]    vrfReadDataPorts_20_bits_vs,
  output [2:0]    vrfReadDataPorts_20_bits_instructionIndex,
  input           vrfReadDataPorts_21_ready,
  output          vrfReadDataPorts_21_valid,
  output [4:0]    vrfReadDataPorts_21_bits_vs,
  output [2:0]    vrfReadDataPorts_21_bits_instructionIndex,
  input           vrfReadDataPorts_22_ready,
  output          vrfReadDataPorts_22_valid,
  output [4:0]    vrfReadDataPorts_22_bits_vs,
  output [2:0]    vrfReadDataPorts_22_bits_instructionIndex,
  input           vrfReadDataPorts_23_ready,
  output          vrfReadDataPorts_23_valid,
  output [4:0]    vrfReadDataPorts_23_bits_vs,
  output [2:0]    vrfReadDataPorts_23_bits_instructionIndex,
  input           vrfReadDataPorts_24_ready,
  output          vrfReadDataPorts_24_valid,
  output [4:0]    vrfReadDataPorts_24_bits_vs,
  output [2:0]    vrfReadDataPorts_24_bits_instructionIndex,
  input           vrfReadDataPorts_25_ready,
  output          vrfReadDataPorts_25_valid,
  output [4:0]    vrfReadDataPorts_25_bits_vs,
  output [2:0]    vrfReadDataPorts_25_bits_instructionIndex,
  input           vrfReadDataPorts_26_ready,
  output          vrfReadDataPorts_26_valid,
  output [4:0]    vrfReadDataPorts_26_bits_vs,
  output [2:0]    vrfReadDataPorts_26_bits_instructionIndex,
  input           vrfReadDataPorts_27_ready,
  output          vrfReadDataPorts_27_valid,
  output [4:0]    vrfReadDataPorts_27_bits_vs,
  output [2:0]    vrfReadDataPorts_27_bits_instructionIndex,
  input           vrfReadDataPorts_28_ready,
  output          vrfReadDataPorts_28_valid,
  output [4:0]    vrfReadDataPorts_28_bits_vs,
  output [2:0]    vrfReadDataPorts_28_bits_instructionIndex,
  input           vrfReadDataPorts_29_ready,
  output          vrfReadDataPorts_29_valid,
  output [4:0]    vrfReadDataPorts_29_bits_vs,
  output [2:0]    vrfReadDataPorts_29_bits_instructionIndex,
  input           vrfReadDataPorts_30_ready,
  output          vrfReadDataPorts_30_valid,
  output [4:0]    vrfReadDataPorts_30_bits_vs,
  output [2:0]    vrfReadDataPorts_30_bits_instructionIndex,
  input           vrfReadDataPorts_31_ready,
  output          vrfReadDataPorts_31_valid,
  output [4:0]    vrfReadDataPorts_31_bits_vs,
  output [2:0]    vrfReadDataPorts_31_bits_instructionIndex,
  input           vrfReadResults_0_valid,
  input  [31:0]   vrfReadResults_0_bits,
  input           vrfReadResults_1_valid,
  input  [31:0]   vrfReadResults_1_bits,
  input           vrfReadResults_2_valid,
  input  [31:0]   vrfReadResults_2_bits,
  input           vrfReadResults_3_valid,
  input  [31:0]   vrfReadResults_3_bits,
  input           vrfReadResults_4_valid,
  input  [31:0]   vrfReadResults_4_bits,
  input           vrfReadResults_5_valid,
  input  [31:0]   vrfReadResults_5_bits,
  input           vrfReadResults_6_valid,
  input  [31:0]   vrfReadResults_6_bits,
  input           vrfReadResults_7_valid,
  input  [31:0]   vrfReadResults_7_bits,
  input           vrfReadResults_8_valid,
  input  [31:0]   vrfReadResults_8_bits,
  input           vrfReadResults_9_valid,
  input  [31:0]   vrfReadResults_9_bits,
  input           vrfReadResults_10_valid,
  input  [31:0]   vrfReadResults_10_bits,
  input           vrfReadResults_11_valid,
  input  [31:0]   vrfReadResults_11_bits,
  input           vrfReadResults_12_valid,
  input  [31:0]   vrfReadResults_12_bits,
  input           vrfReadResults_13_valid,
  input  [31:0]   vrfReadResults_13_bits,
  input           vrfReadResults_14_valid,
  input  [31:0]   vrfReadResults_14_bits,
  input           vrfReadResults_15_valid,
  input  [31:0]   vrfReadResults_15_bits,
  input           vrfReadResults_16_valid,
  input  [31:0]   vrfReadResults_16_bits,
  input           vrfReadResults_17_valid,
  input  [31:0]   vrfReadResults_17_bits,
  input           vrfReadResults_18_valid,
  input  [31:0]   vrfReadResults_18_bits,
  input           vrfReadResults_19_valid,
  input  [31:0]   vrfReadResults_19_bits,
  input           vrfReadResults_20_valid,
  input  [31:0]   vrfReadResults_20_bits,
  input           vrfReadResults_21_valid,
  input  [31:0]   vrfReadResults_21_bits,
  input           vrfReadResults_22_valid,
  input  [31:0]   vrfReadResults_22_bits,
  input           vrfReadResults_23_valid,
  input  [31:0]   vrfReadResults_23_bits,
  input           vrfReadResults_24_valid,
  input  [31:0]   vrfReadResults_24_bits,
  input           vrfReadResults_25_valid,
  input  [31:0]   vrfReadResults_25_bits,
  input           vrfReadResults_26_valid,
  input  [31:0]   vrfReadResults_26_bits,
  input           vrfReadResults_27_valid,
  input  [31:0]   vrfReadResults_27_bits,
  input           vrfReadResults_28_valid,
  input  [31:0]   vrfReadResults_28_bits,
  input           vrfReadResults_29_valid,
  input  [31:0]   vrfReadResults_29_bits,
  input           vrfReadResults_30_valid,
  input  [31:0]   vrfReadResults_30_bits,
  input           vrfReadResults_31_valid,
  input  [31:0]   vrfReadResults_31_bits,
  input           vrfWritePort_0_ready,
  output          vrfWritePort_0_valid,
  output [4:0]    vrfWritePort_0_bits_vd,
  output [3:0]    vrfWritePort_0_bits_mask,
  output [31:0]   vrfWritePort_0_bits_data,
  output          vrfWritePort_0_bits_last,
  output [2:0]    vrfWritePort_0_bits_instructionIndex,
  input           vrfWritePort_1_ready,
  output          vrfWritePort_1_valid,
  output [4:0]    vrfWritePort_1_bits_vd,
  output [3:0]    vrfWritePort_1_bits_mask,
  output [31:0]   vrfWritePort_1_bits_data,
  output          vrfWritePort_1_bits_last,
  output [2:0]    vrfWritePort_1_bits_instructionIndex,
  input           vrfWritePort_2_ready,
  output          vrfWritePort_2_valid,
  output [4:0]    vrfWritePort_2_bits_vd,
  output [3:0]    vrfWritePort_2_bits_mask,
  output [31:0]   vrfWritePort_2_bits_data,
  output          vrfWritePort_2_bits_last,
  output [2:0]    vrfWritePort_2_bits_instructionIndex,
  input           vrfWritePort_3_ready,
  output          vrfWritePort_3_valid,
  output [4:0]    vrfWritePort_3_bits_vd,
  output [3:0]    vrfWritePort_3_bits_mask,
  output [31:0]   vrfWritePort_3_bits_data,
  output          vrfWritePort_3_bits_last,
  output [2:0]    vrfWritePort_3_bits_instructionIndex,
  input           vrfWritePort_4_ready,
  output          vrfWritePort_4_valid,
  output [4:0]    vrfWritePort_4_bits_vd,
  output [3:0]    vrfWritePort_4_bits_mask,
  output [31:0]   vrfWritePort_4_bits_data,
  output          vrfWritePort_4_bits_last,
  output [2:0]    vrfWritePort_4_bits_instructionIndex,
  input           vrfWritePort_5_ready,
  output          vrfWritePort_5_valid,
  output [4:0]    vrfWritePort_5_bits_vd,
  output [3:0]    vrfWritePort_5_bits_mask,
  output [31:0]   vrfWritePort_5_bits_data,
  output          vrfWritePort_5_bits_last,
  output [2:0]    vrfWritePort_5_bits_instructionIndex,
  input           vrfWritePort_6_ready,
  output          vrfWritePort_6_valid,
  output [4:0]    vrfWritePort_6_bits_vd,
  output [3:0]    vrfWritePort_6_bits_mask,
  output [31:0]   vrfWritePort_6_bits_data,
  output          vrfWritePort_6_bits_last,
  output [2:0]    vrfWritePort_6_bits_instructionIndex,
  input           vrfWritePort_7_ready,
  output          vrfWritePort_7_valid,
  output [4:0]    vrfWritePort_7_bits_vd,
  output [3:0]    vrfWritePort_7_bits_mask,
  output [31:0]   vrfWritePort_7_bits_data,
  output          vrfWritePort_7_bits_last,
  output [2:0]    vrfWritePort_7_bits_instructionIndex,
  input           vrfWritePort_8_ready,
  output          vrfWritePort_8_valid,
  output [4:0]    vrfWritePort_8_bits_vd,
  output [3:0]    vrfWritePort_8_bits_mask,
  output [31:0]   vrfWritePort_8_bits_data,
  output          vrfWritePort_8_bits_last,
  output [2:0]    vrfWritePort_8_bits_instructionIndex,
  input           vrfWritePort_9_ready,
  output          vrfWritePort_9_valid,
  output [4:0]    vrfWritePort_9_bits_vd,
  output [3:0]    vrfWritePort_9_bits_mask,
  output [31:0]   vrfWritePort_9_bits_data,
  output          vrfWritePort_9_bits_last,
  output [2:0]    vrfWritePort_9_bits_instructionIndex,
  input           vrfWritePort_10_ready,
  output          vrfWritePort_10_valid,
  output [4:0]    vrfWritePort_10_bits_vd,
  output [3:0]    vrfWritePort_10_bits_mask,
  output [31:0]   vrfWritePort_10_bits_data,
  output          vrfWritePort_10_bits_last,
  output [2:0]    vrfWritePort_10_bits_instructionIndex,
  input           vrfWritePort_11_ready,
  output          vrfWritePort_11_valid,
  output [4:0]    vrfWritePort_11_bits_vd,
  output [3:0]    vrfWritePort_11_bits_mask,
  output [31:0]   vrfWritePort_11_bits_data,
  output          vrfWritePort_11_bits_last,
  output [2:0]    vrfWritePort_11_bits_instructionIndex,
  input           vrfWritePort_12_ready,
  output          vrfWritePort_12_valid,
  output [4:0]    vrfWritePort_12_bits_vd,
  output [3:0]    vrfWritePort_12_bits_mask,
  output [31:0]   vrfWritePort_12_bits_data,
  output          vrfWritePort_12_bits_last,
  output [2:0]    vrfWritePort_12_bits_instructionIndex,
  input           vrfWritePort_13_ready,
  output          vrfWritePort_13_valid,
  output [4:0]    vrfWritePort_13_bits_vd,
  output [3:0]    vrfWritePort_13_bits_mask,
  output [31:0]   vrfWritePort_13_bits_data,
  output          vrfWritePort_13_bits_last,
  output [2:0]    vrfWritePort_13_bits_instructionIndex,
  input           vrfWritePort_14_ready,
  output          vrfWritePort_14_valid,
  output [4:0]    vrfWritePort_14_bits_vd,
  output [3:0]    vrfWritePort_14_bits_mask,
  output [31:0]   vrfWritePort_14_bits_data,
  output          vrfWritePort_14_bits_last,
  output [2:0]    vrfWritePort_14_bits_instructionIndex,
  input           vrfWritePort_15_ready,
  output          vrfWritePort_15_valid,
  output [4:0]    vrfWritePort_15_bits_vd,
  output [3:0]    vrfWritePort_15_bits_mask,
  output [31:0]   vrfWritePort_15_bits_data,
  output          vrfWritePort_15_bits_last,
  output [2:0]    vrfWritePort_15_bits_instructionIndex,
  input           vrfWritePort_16_ready,
  output          vrfWritePort_16_valid,
  output [4:0]    vrfWritePort_16_bits_vd,
  output [3:0]    vrfWritePort_16_bits_mask,
  output [31:0]   vrfWritePort_16_bits_data,
  output          vrfWritePort_16_bits_last,
  output [2:0]    vrfWritePort_16_bits_instructionIndex,
  input           vrfWritePort_17_ready,
  output          vrfWritePort_17_valid,
  output [4:0]    vrfWritePort_17_bits_vd,
  output [3:0]    vrfWritePort_17_bits_mask,
  output [31:0]   vrfWritePort_17_bits_data,
  output          vrfWritePort_17_bits_last,
  output [2:0]    vrfWritePort_17_bits_instructionIndex,
  input           vrfWritePort_18_ready,
  output          vrfWritePort_18_valid,
  output [4:0]    vrfWritePort_18_bits_vd,
  output [3:0]    vrfWritePort_18_bits_mask,
  output [31:0]   vrfWritePort_18_bits_data,
  output          vrfWritePort_18_bits_last,
  output [2:0]    vrfWritePort_18_bits_instructionIndex,
  input           vrfWritePort_19_ready,
  output          vrfWritePort_19_valid,
  output [4:0]    vrfWritePort_19_bits_vd,
  output [3:0]    vrfWritePort_19_bits_mask,
  output [31:0]   vrfWritePort_19_bits_data,
  output          vrfWritePort_19_bits_last,
  output [2:0]    vrfWritePort_19_bits_instructionIndex,
  input           vrfWritePort_20_ready,
  output          vrfWritePort_20_valid,
  output [4:0]    vrfWritePort_20_bits_vd,
  output [3:0]    vrfWritePort_20_bits_mask,
  output [31:0]   vrfWritePort_20_bits_data,
  output          vrfWritePort_20_bits_last,
  output [2:0]    vrfWritePort_20_bits_instructionIndex,
  input           vrfWritePort_21_ready,
  output          vrfWritePort_21_valid,
  output [4:0]    vrfWritePort_21_bits_vd,
  output [3:0]    vrfWritePort_21_bits_mask,
  output [31:0]   vrfWritePort_21_bits_data,
  output          vrfWritePort_21_bits_last,
  output [2:0]    vrfWritePort_21_bits_instructionIndex,
  input           vrfWritePort_22_ready,
  output          vrfWritePort_22_valid,
  output [4:0]    vrfWritePort_22_bits_vd,
  output [3:0]    vrfWritePort_22_bits_mask,
  output [31:0]   vrfWritePort_22_bits_data,
  output          vrfWritePort_22_bits_last,
  output [2:0]    vrfWritePort_22_bits_instructionIndex,
  input           vrfWritePort_23_ready,
  output          vrfWritePort_23_valid,
  output [4:0]    vrfWritePort_23_bits_vd,
  output [3:0]    vrfWritePort_23_bits_mask,
  output [31:0]   vrfWritePort_23_bits_data,
  output          vrfWritePort_23_bits_last,
  output [2:0]    vrfWritePort_23_bits_instructionIndex,
  input           vrfWritePort_24_ready,
  output          vrfWritePort_24_valid,
  output [4:0]    vrfWritePort_24_bits_vd,
  output [3:0]    vrfWritePort_24_bits_mask,
  output [31:0]   vrfWritePort_24_bits_data,
  output          vrfWritePort_24_bits_last,
  output [2:0]    vrfWritePort_24_bits_instructionIndex,
  input           vrfWritePort_25_ready,
  output          vrfWritePort_25_valid,
  output [4:0]    vrfWritePort_25_bits_vd,
  output [3:0]    vrfWritePort_25_bits_mask,
  output [31:0]   vrfWritePort_25_bits_data,
  output          vrfWritePort_25_bits_last,
  output [2:0]    vrfWritePort_25_bits_instructionIndex,
  input           vrfWritePort_26_ready,
  output          vrfWritePort_26_valid,
  output [4:0]    vrfWritePort_26_bits_vd,
  output [3:0]    vrfWritePort_26_bits_mask,
  output [31:0]   vrfWritePort_26_bits_data,
  output          vrfWritePort_26_bits_last,
  output [2:0]    vrfWritePort_26_bits_instructionIndex,
  input           vrfWritePort_27_ready,
  output          vrfWritePort_27_valid,
  output [4:0]    vrfWritePort_27_bits_vd,
  output [3:0]    vrfWritePort_27_bits_mask,
  output [31:0]   vrfWritePort_27_bits_data,
  output          vrfWritePort_27_bits_last,
  output [2:0]    vrfWritePort_27_bits_instructionIndex,
  input           vrfWritePort_28_ready,
  output          vrfWritePort_28_valid,
  output [4:0]    vrfWritePort_28_bits_vd,
  output [3:0]    vrfWritePort_28_bits_mask,
  output [31:0]   vrfWritePort_28_bits_data,
  output          vrfWritePort_28_bits_last,
  output [2:0]    vrfWritePort_28_bits_instructionIndex,
  input           vrfWritePort_29_ready,
  output          vrfWritePort_29_valid,
  output [4:0]    vrfWritePort_29_bits_vd,
  output [3:0]    vrfWritePort_29_bits_mask,
  output [31:0]   vrfWritePort_29_bits_data,
  output          vrfWritePort_29_bits_last,
  output [2:0]    vrfWritePort_29_bits_instructionIndex,
  input           vrfWritePort_30_ready,
  output          vrfWritePort_30_valid,
  output [4:0]    vrfWritePort_30_bits_vd,
  output [3:0]    vrfWritePort_30_bits_mask,
  output [31:0]   vrfWritePort_30_bits_data,
  output          vrfWritePort_30_bits_last,
  output [2:0]    vrfWritePort_30_bits_instructionIndex,
  input           vrfWritePort_31_ready,
  output          vrfWritePort_31_valid,
  output [4:0]    vrfWritePort_31_bits_vd,
  output [3:0]    vrfWritePort_31_bits_mask,
  output [31:0]   vrfWritePort_31_bits_data,
  output          vrfWritePort_31_bits_last,
  output [2:0]    vrfWritePort_31_bits_instructionIndex,
  input           writeRelease_0,
                  writeRelease_1,
                  writeRelease_2,
                  writeRelease_3,
                  writeRelease_4,
                  writeRelease_5,
                  writeRelease_6,
                  writeRelease_7,
                  writeRelease_8,
                  writeRelease_9,
                  writeRelease_10,
                  writeRelease_11,
                  writeRelease_12,
                  writeRelease_13,
                  writeRelease_14,
                  writeRelease_15,
                  writeRelease_16,
                  writeRelease_17,
                  writeRelease_18,
                  writeRelease_19,
                  writeRelease_20,
                  writeRelease_21,
                  writeRelease_22,
                  writeRelease_23,
                  writeRelease_24,
                  writeRelease_25,
                  writeRelease_26,
                  writeRelease_27,
                  writeRelease_28,
                  writeRelease_29,
                  writeRelease_30,
                  writeRelease_31,
  output [7:0]    dataInWriteQueue_0,
                  dataInWriteQueue_1,
                  dataInWriteQueue_2,
                  dataInWriteQueue_3,
                  dataInWriteQueue_4,
                  dataInWriteQueue_5,
                  dataInWriteQueue_6,
                  dataInWriteQueue_7,
                  dataInWriteQueue_8,
                  dataInWriteQueue_9,
                  dataInWriteQueue_10,
                  dataInWriteQueue_11,
                  dataInWriteQueue_12,
                  dataInWriteQueue_13,
                  dataInWriteQueue_14,
                  dataInWriteQueue_15,
                  dataInWriteQueue_16,
                  dataInWriteQueue_17,
                  dataInWriteQueue_18,
                  dataInWriteQueue_19,
                  dataInWriteQueue_20,
                  dataInWriteQueue_21,
                  dataInWriteQueue_22,
                  dataInWriteQueue_23,
                  dataInWriteQueue_24,
                  dataInWriteQueue_25,
                  dataInWriteQueue_26,
                  dataInWriteQueue_27,
                  dataInWriteQueue_28,
                  dataInWriteQueue_29,
                  dataInWriteQueue_30,
                  dataInWriteQueue_31,
  input  [10:0]   csrInterface_vl,
                  csrInterface_vStart,
  input  [2:0]    csrInterface_vlmul,
  input  [1:0]    csrInterface_vSew,
                  csrInterface_vxrm,
  input           csrInterface_vta,
                  csrInterface_vma,
                  offsetReadResult_0_valid,
  input  [31:0]   offsetReadResult_0_bits,
  input           offsetReadResult_1_valid,
  input  [31:0]   offsetReadResult_1_bits,
  input           offsetReadResult_2_valid,
  input  [31:0]   offsetReadResult_2_bits,
  input           offsetReadResult_3_valid,
  input  [31:0]   offsetReadResult_3_bits,
  input           offsetReadResult_4_valid,
  input  [31:0]   offsetReadResult_4_bits,
  input           offsetReadResult_5_valid,
  input  [31:0]   offsetReadResult_5_bits,
  input           offsetReadResult_6_valid,
  input  [31:0]   offsetReadResult_6_bits,
  input           offsetReadResult_7_valid,
  input  [31:0]   offsetReadResult_7_bits,
  input           offsetReadResult_8_valid,
  input  [31:0]   offsetReadResult_8_bits,
  input           offsetReadResult_9_valid,
  input  [31:0]   offsetReadResult_9_bits,
  input           offsetReadResult_10_valid,
  input  [31:0]   offsetReadResult_10_bits,
  input           offsetReadResult_11_valid,
  input  [31:0]   offsetReadResult_11_bits,
  input           offsetReadResult_12_valid,
  input  [31:0]   offsetReadResult_12_bits,
  input           offsetReadResult_13_valid,
  input  [31:0]   offsetReadResult_13_bits,
  input           offsetReadResult_14_valid,
  input  [31:0]   offsetReadResult_14_bits,
  input           offsetReadResult_15_valid,
  input  [31:0]   offsetReadResult_15_bits,
  input           offsetReadResult_16_valid,
  input  [31:0]   offsetReadResult_16_bits,
  input           offsetReadResult_17_valid,
  input  [31:0]   offsetReadResult_17_bits,
  input           offsetReadResult_18_valid,
  input  [31:0]   offsetReadResult_18_bits,
  input           offsetReadResult_19_valid,
  input  [31:0]   offsetReadResult_19_bits,
  input           offsetReadResult_20_valid,
  input  [31:0]   offsetReadResult_20_bits,
  input           offsetReadResult_21_valid,
  input  [31:0]   offsetReadResult_21_bits,
  input           offsetReadResult_22_valid,
  input  [31:0]   offsetReadResult_22_bits,
  input           offsetReadResult_23_valid,
  input  [31:0]   offsetReadResult_23_bits,
  input           offsetReadResult_24_valid,
  input  [31:0]   offsetReadResult_24_bits,
  input           offsetReadResult_25_valid,
  input  [31:0]   offsetReadResult_25_bits,
  input           offsetReadResult_26_valid,
  input  [31:0]   offsetReadResult_26_bits,
  input           offsetReadResult_27_valid,
  input  [31:0]   offsetReadResult_27_bits,
  input           offsetReadResult_28_valid,
  input  [31:0]   offsetReadResult_28_bits,
  input           offsetReadResult_29_valid,
  input  [31:0]   offsetReadResult_29_bits,
  input           offsetReadResult_30_valid,
  input  [31:0]   offsetReadResult_30_bits,
  input           offsetReadResult_31_valid,
  input  [31:0]   offsetReadResult_31_bits,
  output [7:0]    lastReport,
  output [31:0]   tokenIO_offsetGroupRelease
);

  wire              _simpleDataQueue_fifo_empty;
  wire              _simpleDataQueue_fifo_full;
  wire              _simpleDataQueue_fifo_error;
  wire [77:0]       _simpleDataQueue_fifo_data_out;
  wire              _simpleSourceQueue_fifo_empty;
  wire              _simpleSourceQueue_fifo_full;
  wire              _simpleSourceQueue_fifo_error;
  wire              _dataQueue_fifo_empty;
  wire              _dataQueue_fifo_full;
  wire              _dataQueue_fifo_error;
  wire [1187:0]     _dataQueue_fifo_data_out;
  wire              _sourceQueue_fifo_empty;
  wire              _sourceQueue_fifo_full;
  wire              _sourceQueue_fifo_error;
  wire              _writeIndexQueue_fifo_31_empty;
  wire              _writeIndexQueue_fifo_31_full;
  wire              _writeIndexQueue_fifo_31_error;
  wire              _writeIndexQueue_fifo_30_empty;
  wire              _writeIndexQueue_fifo_30_full;
  wire              _writeIndexQueue_fifo_30_error;
  wire              _writeIndexQueue_fifo_29_empty;
  wire              _writeIndexQueue_fifo_29_full;
  wire              _writeIndexQueue_fifo_29_error;
  wire              _writeIndexQueue_fifo_28_empty;
  wire              _writeIndexQueue_fifo_28_full;
  wire              _writeIndexQueue_fifo_28_error;
  wire              _writeIndexQueue_fifo_27_empty;
  wire              _writeIndexQueue_fifo_27_full;
  wire              _writeIndexQueue_fifo_27_error;
  wire              _writeIndexQueue_fifo_26_empty;
  wire              _writeIndexQueue_fifo_26_full;
  wire              _writeIndexQueue_fifo_26_error;
  wire              _writeIndexQueue_fifo_25_empty;
  wire              _writeIndexQueue_fifo_25_full;
  wire              _writeIndexQueue_fifo_25_error;
  wire              _writeIndexQueue_fifo_24_empty;
  wire              _writeIndexQueue_fifo_24_full;
  wire              _writeIndexQueue_fifo_24_error;
  wire              _writeIndexQueue_fifo_23_empty;
  wire              _writeIndexQueue_fifo_23_full;
  wire              _writeIndexQueue_fifo_23_error;
  wire              _writeIndexQueue_fifo_22_empty;
  wire              _writeIndexQueue_fifo_22_full;
  wire              _writeIndexQueue_fifo_22_error;
  wire              _writeIndexQueue_fifo_21_empty;
  wire              _writeIndexQueue_fifo_21_full;
  wire              _writeIndexQueue_fifo_21_error;
  wire              _writeIndexQueue_fifo_20_empty;
  wire              _writeIndexQueue_fifo_20_full;
  wire              _writeIndexQueue_fifo_20_error;
  wire              _writeIndexQueue_fifo_19_empty;
  wire              _writeIndexQueue_fifo_19_full;
  wire              _writeIndexQueue_fifo_19_error;
  wire              _writeIndexQueue_fifo_18_empty;
  wire              _writeIndexQueue_fifo_18_full;
  wire              _writeIndexQueue_fifo_18_error;
  wire              _writeIndexQueue_fifo_17_empty;
  wire              _writeIndexQueue_fifo_17_full;
  wire              _writeIndexQueue_fifo_17_error;
  wire              _writeIndexQueue_fifo_16_empty;
  wire              _writeIndexQueue_fifo_16_full;
  wire              _writeIndexQueue_fifo_16_error;
  wire              _writeIndexQueue_fifo_15_empty;
  wire              _writeIndexQueue_fifo_15_full;
  wire              _writeIndexQueue_fifo_15_error;
  wire              _writeIndexQueue_fifo_14_empty;
  wire              _writeIndexQueue_fifo_14_full;
  wire              _writeIndexQueue_fifo_14_error;
  wire              _writeIndexQueue_fifo_13_empty;
  wire              _writeIndexQueue_fifo_13_full;
  wire              _writeIndexQueue_fifo_13_error;
  wire              _writeIndexQueue_fifo_12_empty;
  wire              _writeIndexQueue_fifo_12_full;
  wire              _writeIndexQueue_fifo_12_error;
  wire              _writeIndexQueue_fifo_11_empty;
  wire              _writeIndexQueue_fifo_11_full;
  wire              _writeIndexQueue_fifo_11_error;
  wire              _writeIndexQueue_fifo_10_empty;
  wire              _writeIndexQueue_fifo_10_full;
  wire              _writeIndexQueue_fifo_10_error;
  wire              _writeIndexQueue_fifo_9_empty;
  wire              _writeIndexQueue_fifo_9_full;
  wire              _writeIndexQueue_fifo_9_error;
  wire              _writeIndexQueue_fifo_8_empty;
  wire              _writeIndexQueue_fifo_8_full;
  wire              _writeIndexQueue_fifo_8_error;
  wire              _writeIndexQueue_fifo_7_empty;
  wire              _writeIndexQueue_fifo_7_full;
  wire              _writeIndexQueue_fifo_7_error;
  wire              _writeIndexQueue_fifo_6_empty;
  wire              _writeIndexQueue_fifo_6_full;
  wire              _writeIndexQueue_fifo_6_error;
  wire              _writeIndexQueue_fifo_5_empty;
  wire              _writeIndexQueue_fifo_5_full;
  wire              _writeIndexQueue_fifo_5_error;
  wire              _writeIndexQueue_fifo_4_empty;
  wire              _writeIndexQueue_fifo_4_full;
  wire              _writeIndexQueue_fifo_4_error;
  wire              _writeIndexQueue_fifo_3_empty;
  wire              _writeIndexQueue_fifo_3_full;
  wire              _writeIndexQueue_fifo_3_error;
  wire              _writeIndexQueue_fifo_2_empty;
  wire              _writeIndexQueue_fifo_2_full;
  wire              _writeIndexQueue_fifo_2_error;
  wire              _writeIndexQueue_fifo_1_empty;
  wire              _writeIndexQueue_fifo_1_full;
  wire              _writeIndexQueue_fifo_1_error;
  wire              _writeIndexQueue_fifo_empty;
  wire              _writeIndexQueue_fifo_full;
  wire              _writeIndexQueue_fifo_error;
  wire              _otherUnitDataQueueVec_fifo_31_empty;
  wire              _otherUnitDataQueueVec_fifo_31_full;
  wire              _otherUnitDataQueueVec_fifo_31_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_31_data_out;
  wire              _otherUnitDataQueueVec_fifo_30_empty;
  wire              _otherUnitDataQueueVec_fifo_30_full;
  wire              _otherUnitDataQueueVec_fifo_30_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_30_data_out;
  wire              _otherUnitDataQueueVec_fifo_29_empty;
  wire              _otherUnitDataQueueVec_fifo_29_full;
  wire              _otherUnitDataQueueVec_fifo_29_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_29_data_out;
  wire              _otherUnitDataQueueVec_fifo_28_empty;
  wire              _otherUnitDataQueueVec_fifo_28_full;
  wire              _otherUnitDataQueueVec_fifo_28_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_28_data_out;
  wire              _otherUnitDataQueueVec_fifo_27_empty;
  wire              _otherUnitDataQueueVec_fifo_27_full;
  wire              _otherUnitDataQueueVec_fifo_27_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_27_data_out;
  wire              _otherUnitDataQueueVec_fifo_26_empty;
  wire              _otherUnitDataQueueVec_fifo_26_full;
  wire              _otherUnitDataQueueVec_fifo_26_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_26_data_out;
  wire              _otherUnitDataQueueVec_fifo_25_empty;
  wire              _otherUnitDataQueueVec_fifo_25_full;
  wire              _otherUnitDataQueueVec_fifo_25_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_25_data_out;
  wire              _otherUnitDataQueueVec_fifo_24_empty;
  wire              _otherUnitDataQueueVec_fifo_24_full;
  wire              _otherUnitDataQueueVec_fifo_24_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_24_data_out;
  wire              _otherUnitDataQueueVec_fifo_23_empty;
  wire              _otherUnitDataQueueVec_fifo_23_full;
  wire              _otherUnitDataQueueVec_fifo_23_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_23_data_out;
  wire              _otherUnitDataQueueVec_fifo_22_empty;
  wire              _otherUnitDataQueueVec_fifo_22_full;
  wire              _otherUnitDataQueueVec_fifo_22_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_22_data_out;
  wire              _otherUnitDataQueueVec_fifo_21_empty;
  wire              _otherUnitDataQueueVec_fifo_21_full;
  wire              _otherUnitDataQueueVec_fifo_21_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_21_data_out;
  wire              _otherUnitDataQueueVec_fifo_20_empty;
  wire              _otherUnitDataQueueVec_fifo_20_full;
  wire              _otherUnitDataQueueVec_fifo_20_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_20_data_out;
  wire              _otherUnitDataQueueVec_fifo_19_empty;
  wire              _otherUnitDataQueueVec_fifo_19_full;
  wire              _otherUnitDataQueueVec_fifo_19_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_19_data_out;
  wire              _otherUnitDataQueueVec_fifo_18_empty;
  wire              _otherUnitDataQueueVec_fifo_18_full;
  wire              _otherUnitDataQueueVec_fifo_18_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_18_data_out;
  wire              _otherUnitDataQueueVec_fifo_17_empty;
  wire              _otherUnitDataQueueVec_fifo_17_full;
  wire              _otherUnitDataQueueVec_fifo_17_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_17_data_out;
  wire              _otherUnitDataQueueVec_fifo_16_empty;
  wire              _otherUnitDataQueueVec_fifo_16_full;
  wire              _otherUnitDataQueueVec_fifo_16_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_16_data_out;
  wire              _otherUnitDataQueueVec_fifo_15_empty;
  wire              _otherUnitDataQueueVec_fifo_15_full;
  wire              _otherUnitDataQueueVec_fifo_15_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_15_data_out;
  wire              _otherUnitDataQueueVec_fifo_14_empty;
  wire              _otherUnitDataQueueVec_fifo_14_full;
  wire              _otherUnitDataQueueVec_fifo_14_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_14_data_out;
  wire              _otherUnitDataQueueVec_fifo_13_empty;
  wire              _otherUnitDataQueueVec_fifo_13_full;
  wire              _otherUnitDataQueueVec_fifo_13_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_13_data_out;
  wire              _otherUnitDataQueueVec_fifo_12_empty;
  wire              _otherUnitDataQueueVec_fifo_12_full;
  wire              _otherUnitDataQueueVec_fifo_12_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_12_data_out;
  wire              _otherUnitDataQueueVec_fifo_11_empty;
  wire              _otherUnitDataQueueVec_fifo_11_full;
  wire              _otherUnitDataQueueVec_fifo_11_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_11_data_out;
  wire              _otherUnitDataQueueVec_fifo_10_empty;
  wire              _otherUnitDataQueueVec_fifo_10_full;
  wire              _otherUnitDataQueueVec_fifo_10_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_10_data_out;
  wire              _otherUnitDataQueueVec_fifo_9_empty;
  wire              _otherUnitDataQueueVec_fifo_9_full;
  wire              _otherUnitDataQueueVec_fifo_9_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_9_data_out;
  wire              _otherUnitDataQueueVec_fifo_8_empty;
  wire              _otherUnitDataQueueVec_fifo_8_full;
  wire              _otherUnitDataQueueVec_fifo_8_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_8_data_out;
  wire              _otherUnitDataQueueVec_fifo_7_empty;
  wire              _otherUnitDataQueueVec_fifo_7_full;
  wire              _otherUnitDataQueueVec_fifo_7_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_7_data_out;
  wire              _otherUnitDataQueueVec_fifo_6_empty;
  wire              _otherUnitDataQueueVec_fifo_6_full;
  wire              _otherUnitDataQueueVec_fifo_6_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_6_data_out;
  wire              _otherUnitDataQueueVec_fifo_5_empty;
  wire              _otherUnitDataQueueVec_fifo_5_full;
  wire              _otherUnitDataQueueVec_fifo_5_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_5_data_out;
  wire              _otherUnitDataQueueVec_fifo_4_empty;
  wire              _otherUnitDataQueueVec_fifo_4_full;
  wire              _otherUnitDataQueueVec_fifo_4_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_4_data_out;
  wire              _otherUnitDataQueueVec_fifo_3_empty;
  wire              _otherUnitDataQueueVec_fifo_3_full;
  wire              _otherUnitDataQueueVec_fifo_3_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_3_data_out;
  wire              _otherUnitDataQueueVec_fifo_2_empty;
  wire              _otherUnitDataQueueVec_fifo_2_full;
  wire              _otherUnitDataQueueVec_fifo_2_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_2_data_out;
  wire              _otherUnitDataQueueVec_fifo_1_empty;
  wire              _otherUnitDataQueueVec_fifo_1_full;
  wire              _otherUnitDataQueueVec_fifo_1_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_1_data_out;
  wire              _otherUnitDataQueueVec_fifo_empty;
  wire              _otherUnitDataQueueVec_fifo_full;
  wire              _otherUnitDataQueueVec_fifo_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_data_out;
  wire              _otherUnitTargetQueue_fifo_empty;
  wire              _otherUnitTargetQueue_fifo_full;
  wire              _otherUnitTargetQueue_fifo_error;
  wire              _writeQueueVec_fifo_31_empty;
  wire              _writeQueueVec_fifo_31_full;
  wire              _writeQueueVec_fifo_31_error;
  wire [76:0]       _writeQueueVec_fifo_31_data_out;
  wire              _writeQueueVec_fifo_30_empty;
  wire              _writeQueueVec_fifo_30_full;
  wire              _writeQueueVec_fifo_30_error;
  wire [76:0]       _writeQueueVec_fifo_30_data_out;
  wire              _writeQueueVec_fifo_29_empty;
  wire              _writeQueueVec_fifo_29_full;
  wire              _writeQueueVec_fifo_29_error;
  wire [76:0]       _writeQueueVec_fifo_29_data_out;
  wire              _writeQueueVec_fifo_28_empty;
  wire              _writeQueueVec_fifo_28_full;
  wire              _writeQueueVec_fifo_28_error;
  wire [76:0]       _writeQueueVec_fifo_28_data_out;
  wire              _writeQueueVec_fifo_27_empty;
  wire              _writeQueueVec_fifo_27_full;
  wire              _writeQueueVec_fifo_27_error;
  wire [76:0]       _writeQueueVec_fifo_27_data_out;
  wire              _writeQueueVec_fifo_26_empty;
  wire              _writeQueueVec_fifo_26_full;
  wire              _writeQueueVec_fifo_26_error;
  wire [76:0]       _writeQueueVec_fifo_26_data_out;
  wire              _writeQueueVec_fifo_25_empty;
  wire              _writeQueueVec_fifo_25_full;
  wire              _writeQueueVec_fifo_25_error;
  wire [76:0]       _writeQueueVec_fifo_25_data_out;
  wire              _writeQueueVec_fifo_24_empty;
  wire              _writeQueueVec_fifo_24_full;
  wire              _writeQueueVec_fifo_24_error;
  wire [76:0]       _writeQueueVec_fifo_24_data_out;
  wire              _writeQueueVec_fifo_23_empty;
  wire              _writeQueueVec_fifo_23_full;
  wire              _writeQueueVec_fifo_23_error;
  wire [76:0]       _writeQueueVec_fifo_23_data_out;
  wire              _writeQueueVec_fifo_22_empty;
  wire              _writeQueueVec_fifo_22_full;
  wire              _writeQueueVec_fifo_22_error;
  wire [76:0]       _writeQueueVec_fifo_22_data_out;
  wire              _writeQueueVec_fifo_21_empty;
  wire              _writeQueueVec_fifo_21_full;
  wire              _writeQueueVec_fifo_21_error;
  wire [76:0]       _writeQueueVec_fifo_21_data_out;
  wire              _writeQueueVec_fifo_20_empty;
  wire              _writeQueueVec_fifo_20_full;
  wire              _writeQueueVec_fifo_20_error;
  wire [76:0]       _writeQueueVec_fifo_20_data_out;
  wire              _writeQueueVec_fifo_19_empty;
  wire              _writeQueueVec_fifo_19_full;
  wire              _writeQueueVec_fifo_19_error;
  wire [76:0]       _writeQueueVec_fifo_19_data_out;
  wire              _writeQueueVec_fifo_18_empty;
  wire              _writeQueueVec_fifo_18_full;
  wire              _writeQueueVec_fifo_18_error;
  wire [76:0]       _writeQueueVec_fifo_18_data_out;
  wire              _writeQueueVec_fifo_17_empty;
  wire              _writeQueueVec_fifo_17_full;
  wire              _writeQueueVec_fifo_17_error;
  wire [76:0]       _writeQueueVec_fifo_17_data_out;
  wire              _writeQueueVec_fifo_16_empty;
  wire              _writeQueueVec_fifo_16_full;
  wire              _writeQueueVec_fifo_16_error;
  wire [76:0]       _writeQueueVec_fifo_16_data_out;
  wire              _writeQueueVec_fifo_15_empty;
  wire              _writeQueueVec_fifo_15_full;
  wire              _writeQueueVec_fifo_15_error;
  wire [76:0]       _writeQueueVec_fifo_15_data_out;
  wire              _writeQueueVec_fifo_14_empty;
  wire              _writeQueueVec_fifo_14_full;
  wire              _writeQueueVec_fifo_14_error;
  wire [76:0]       _writeQueueVec_fifo_14_data_out;
  wire              _writeQueueVec_fifo_13_empty;
  wire              _writeQueueVec_fifo_13_full;
  wire              _writeQueueVec_fifo_13_error;
  wire [76:0]       _writeQueueVec_fifo_13_data_out;
  wire              _writeQueueVec_fifo_12_empty;
  wire              _writeQueueVec_fifo_12_full;
  wire              _writeQueueVec_fifo_12_error;
  wire [76:0]       _writeQueueVec_fifo_12_data_out;
  wire              _writeQueueVec_fifo_11_empty;
  wire              _writeQueueVec_fifo_11_full;
  wire              _writeQueueVec_fifo_11_error;
  wire [76:0]       _writeQueueVec_fifo_11_data_out;
  wire              _writeQueueVec_fifo_10_empty;
  wire              _writeQueueVec_fifo_10_full;
  wire              _writeQueueVec_fifo_10_error;
  wire [76:0]       _writeQueueVec_fifo_10_data_out;
  wire              _writeQueueVec_fifo_9_empty;
  wire              _writeQueueVec_fifo_9_full;
  wire              _writeQueueVec_fifo_9_error;
  wire [76:0]       _writeQueueVec_fifo_9_data_out;
  wire              _writeQueueVec_fifo_8_empty;
  wire              _writeQueueVec_fifo_8_full;
  wire              _writeQueueVec_fifo_8_error;
  wire [76:0]       _writeQueueVec_fifo_8_data_out;
  wire              _writeQueueVec_fifo_7_empty;
  wire              _writeQueueVec_fifo_7_full;
  wire              _writeQueueVec_fifo_7_error;
  wire [76:0]       _writeQueueVec_fifo_7_data_out;
  wire              _writeQueueVec_fifo_6_empty;
  wire              _writeQueueVec_fifo_6_full;
  wire              _writeQueueVec_fifo_6_error;
  wire [76:0]       _writeQueueVec_fifo_6_data_out;
  wire              _writeQueueVec_fifo_5_empty;
  wire              _writeQueueVec_fifo_5_full;
  wire              _writeQueueVec_fifo_5_error;
  wire [76:0]       _writeQueueVec_fifo_5_data_out;
  wire              _writeQueueVec_fifo_4_empty;
  wire              _writeQueueVec_fifo_4_full;
  wire              _writeQueueVec_fifo_4_error;
  wire [76:0]       _writeQueueVec_fifo_4_data_out;
  wire              _writeQueueVec_fifo_3_empty;
  wire              _writeQueueVec_fifo_3_full;
  wire              _writeQueueVec_fifo_3_error;
  wire [76:0]       _writeQueueVec_fifo_3_data_out;
  wire              _writeQueueVec_fifo_2_empty;
  wire              _writeQueueVec_fifo_2_full;
  wire              _writeQueueVec_fifo_2_error;
  wire [76:0]       _writeQueueVec_fifo_2_data_out;
  wire              _writeQueueVec_fifo_1_empty;
  wire              _writeQueueVec_fifo_1_full;
  wire              _writeQueueVec_fifo_1_error;
  wire [76:0]       _writeQueueVec_fifo_1_data_out;
  wire              _writeQueueVec_fifo_empty;
  wire              _writeQueueVec_fifo_full;
  wire              _writeQueueVec_fifo_error;
  wire [76:0]       _writeQueueVec_fifo_data_out;
  wire              _otherUnit_vrfReadDataPorts_valid;
  wire [4:0]        _otherUnit_vrfReadDataPorts_bits_vs;
  wire [2:0]        _otherUnit_vrfReadDataPorts_bits_instructionIndex;
  wire              _otherUnit_maskSelect_valid;
  wire [2:0]        _otherUnit_maskSelect_bits;
  wire              _otherUnit_memReadRequest_valid;
  wire              _otherUnit_memWriteRequest_valid;
  wire [7:0]        _otherUnit_memWriteRequest_bits_source;
  wire [31:0]       _otherUnit_memWriteRequest_bits_address;
  wire [1:0]        _otherUnit_memWriteRequest_bits_size;
  wire              _otherUnit_vrfWritePort_valid;
  wire [4:0]        _otherUnit_vrfWritePort_bits_vd;
  wire [3:0]        _otherUnit_vrfWritePort_bits_mask;
  wire [31:0]       _otherUnit_vrfWritePort_bits_data;
  wire              _otherUnit_vrfWritePort_bits_last;
  wire [2:0]        _otherUnit_vrfWritePort_bits_instructionIndex;
  wire              _otherUnit_status_idle;
  wire              _otherUnit_status_last;
  wire [2:0]        _otherUnit_status_instructionIndex;
  wire [31:0]       _otherUnit_status_targetLane;
  wire              _otherUnit_status_isStore;
  wire              _otherUnit_offsetRelease_0;
  wire              _otherUnit_offsetRelease_1;
  wire              _otherUnit_offsetRelease_2;
  wire              _otherUnit_offsetRelease_3;
  wire              _otherUnit_offsetRelease_4;
  wire              _otherUnit_offsetRelease_5;
  wire              _otherUnit_offsetRelease_6;
  wire              _otherUnit_offsetRelease_7;
  wire              _otherUnit_offsetRelease_8;
  wire              _otherUnit_offsetRelease_9;
  wire              _otherUnit_offsetRelease_10;
  wire              _otherUnit_offsetRelease_11;
  wire              _otherUnit_offsetRelease_12;
  wire              _otherUnit_offsetRelease_13;
  wire              _otherUnit_offsetRelease_14;
  wire              _otherUnit_offsetRelease_15;
  wire              _otherUnit_offsetRelease_16;
  wire              _otherUnit_offsetRelease_17;
  wire              _otherUnit_offsetRelease_18;
  wire              _otherUnit_offsetRelease_19;
  wire              _otherUnit_offsetRelease_20;
  wire              _otherUnit_offsetRelease_21;
  wire              _otherUnit_offsetRelease_22;
  wire              _otherUnit_offsetRelease_23;
  wire              _otherUnit_offsetRelease_24;
  wire              _otherUnit_offsetRelease_25;
  wire              _otherUnit_offsetRelease_26;
  wire              _otherUnit_offsetRelease_27;
  wire              _otherUnit_offsetRelease_28;
  wire              _otherUnit_offsetRelease_29;
  wire              _otherUnit_offsetRelease_30;
  wire              _otherUnit_offsetRelease_31;
  wire              _storeUnit_maskSelect_valid;
  wire [2:0]        _storeUnit_maskSelect_bits;
  wire              _storeUnit_memRequest_valid;
  wire [3:0]        _storeUnit_memRequest_bits_index;
  wire [31:0]       _storeUnit_memRequest_bits_address;
  wire              _storeUnit_status_idle;
  wire              _storeUnit_status_last;
  wire [2:0]        _storeUnit_status_instructionIndex;
  wire [31:0]       _storeUnit_status_startAddress;
  wire [31:0]       _storeUnit_status_endAddress;
  wire              _storeUnit_vrfReadDataPorts_0_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_0_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_0_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_1_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_1_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_1_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_2_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_2_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_2_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_3_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_3_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_3_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_4_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_4_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_4_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_5_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_5_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_5_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_6_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_6_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_6_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_7_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_7_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_7_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_8_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_8_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_8_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_9_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_9_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_9_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_10_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_10_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_10_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_11_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_11_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_11_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_12_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_12_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_12_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_13_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_13_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_13_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_14_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_14_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_14_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_15_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_15_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_15_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_16_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_16_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_16_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_17_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_17_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_17_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_18_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_18_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_18_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_19_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_19_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_19_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_20_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_20_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_20_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_21_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_21_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_21_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_22_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_22_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_22_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_23_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_23_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_23_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_24_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_24_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_24_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_25_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_25_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_25_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_26_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_26_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_26_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_27_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_27_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_27_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_28_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_28_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_28_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_29_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_29_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_29_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_30_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_30_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_30_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_31_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_31_bits_vs;
  wire [2:0]        _storeUnit_vrfReadDataPorts_31_bits_instructionIndex;
  wire              _loadUnit_maskSelect_valid;
  wire [2:0]        _loadUnit_maskSelect_bits;
  wire              _loadUnit_memRequest_valid;
  wire              _loadUnit_status_idle;
  wire              _loadUnit_status_last;
  wire [2:0]        _loadUnit_status_instructionIndex;
  wire [31:0]       _loadUnit_status_startAddress;
  wire [31:0]       _loadUnit_status_endAddress;
  wire              _loadUnit_vrfWritePort_0_valid;
  wire [4:0]        _loadUnit_vrfWritePort_0_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_0_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_0_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_0_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_1_valid;
  wire [4:0]        _loadUnit_vrfWritePort_1_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_1_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_1_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_1_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_2_valid;
  wire [4:0]        _loadUnit_vrfWritePort_2_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_2_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_2_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_2_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_3_valid;
  wire [4:0]        _loadUnit_vrfWritePort_3_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_3_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_3_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_3_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_4_valid;
  wire [4:0]        _loadUnit_vrfWritePort_4_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_4_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_4_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_4_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_5_valid;
  wire [4:0]        _loadUnit_vrfWritePort_5_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_5_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_5_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_5_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_6_valid;
  wire [4:0]        _loadUnit_vrfWritePort_6_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_6_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_6_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_6_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_7_valid;
  wire [4:0]        _loadUnit_vrfWritePort_7_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_7_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_7_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_7_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_8_valid;
  wire [4:0]        _loadUnit_vrfWritePort_8_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_8_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_8_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_8_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_9_valid;
  wire [4:0]        _loadUnit_vrfWritePort_9_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_9_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_9_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_9_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_10_valid;
  wire [4:0]        _loadUnit_vrfWritePort_10_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_10_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_10_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_10_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_11_valid;
  wire [4:0]        _loadUnit_vrfWritePort_11_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_11_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_11_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_11_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_12_valid;
  wire [4:0]        _loadUnit_vrfWritePort_12_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_12_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_12_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_12_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_13_valid;
  wire [4:0]        _loadUnit_vrfWritePort_13_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_13_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_13_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_13_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_14_valid;
  wire [4:0]        _loadUnit_vrfWritePort_14_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_14_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_14_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_14_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_15_valid;
  wire [4:0]        _loadUnit_vrfWritePort_15_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_15_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_15_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_15_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_16_valid;
  wire [4:0]        _loadUnit_vrfWritePort_16_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_16_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_16_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_16_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_17_valid;
  wire [4:0]        _loadUnit_vrfWritePort_17_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_17_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_17_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_17_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_18_valid;
  wire [4:0]        _loadUnit_vrfWritePort_18_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_18_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_18_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_18_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_19_valid;
  wire [4:0]        _loadUnit_vrfWritePort_19_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_19_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_19_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_19_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_20_valid;
  wire [4:0]        _loadUnit_vrfWritePort_20_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_20_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_20_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_20_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_21_valid;
  wire [4:0]        _loadUnit_vrfWritePort_21_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_21_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_21_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_21_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_22_valid;
  wire [4:0]        _loadUnit_vrfWritePort_22_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_22_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_22_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_22_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_23_valid;
  wire [4:0]        _loadUnit_vrfWritePort_23_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_23_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_23_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_23_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_24_valid;
  wire [4:0]        _loadUnit_vrfWritePort_24_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_24_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_24_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_24_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_25_valid;
  wire [4:0]        _loadUnit_vrfWritePort_25_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_25_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_25_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_25_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_26_valid;
  wire [4:0]        _loadUnit_vrfWritePort_26_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_26_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_26_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_26_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_27_valid;
  wire [4:0]        _loadUnit_vrfWritePort_27_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_27_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_27_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_27_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_28_valid;
  wire [4:0]        _loadUnit_vrfWritePort_28_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_28_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_28_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_28_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_29_valid;
  wire [4:0]        _loadUnit_vrfWritePort_29_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_29_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_29_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_29_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_30_valid;
  wire [4:0]        _loadUnit_vrfWritePort_30_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_30_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_30_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_30_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_31_valid;
  wire [4:0]        _loadUnit_vrfWritePort_31_bits_vd;
  wire [3:0]        _loadUnit_vrfWritePort_31_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_31_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_31_bits_instructionIndex;
  wire              simpleDataQueue_almostFull;
  wire              simpleDataQueue_almostEmpty;
  wire              simpleSourceQueue_almostFull;
  wire              simpleSourceQueue_almostEmpty;
  wire              dataQueue_almostFull;
  wire              dataQueue_almostEmpty;
  wire              sourceQueue_almostFull;
  wire              sourceQueue_almostEmpty;
  wire              writeIndexQueue_31_almostFull;
  wire              writeIndexQueue_31_almostEmpty;
  wire              writeIndexQueue_30_almostFull;
  wire              writeIndexQueue_30_almostEmpty;
  wire              writeIndexQueue_29_almostFull;
  wire              writeIndexQueue_29_almostEmpty;
  wire              writeIndexQueue_28_almostFull;
  wire              writeIndexQueue_28_almostEmpty;
  wire              writeIndexQueue_27_almostFull;
  wire              writeIndexQueue_27_almostEmpty;
  wire              writeIndexQueue_26_almostFull;
  wire              writeIndexQueue_26_almostEmpty;
  wire              writeIndexQueue_25_almostFull;
  wire              writeIndexQueue_25_almostEmpty;
  wire              writeIndexQueue_24_almostFull;
  wire              writeIndexQueue_24_almostEmpty;
  wire              writeIndexQueue_23_almostFull;
  wire              writeIndexQueue_23_almostEmpty;
  wire              writeIndexQueue_22_almostFull;
  wire              writeIndexQueue_22_almostEmpty;
  wire              writeIndexQueue_21_almostFull;
  wire              writeIndexQueue_21_almostEmpty;
  wire              writeIndexQueue_20_almostFull;
  wire              writeIndexQueue_20_almostEmpty;
  wire              writeIndexQueue_19_almostFull;
  wire              writeIndexQueue_19_almostEmpty;
  wire              writeIndexQueue_18_almostFull;
  wire              writeIndexQueue_18_almostEmpty;
  wire              writeIndexQueue_17_almostFull;
  wire              writeIndexQueue_17_almostEmpty;
  wire              writeIndexQueue_16_almostFull;
  wire              writeIndexQueue_16_almostEmpty;
  wire              writeIndexQueue_15_almostFull;
  wire              writeIndexQueue_15_almostEmpty;
  wire              writeIndexQueue_14_almostFull;
  wire              writeIndexQueue_14_almostEmpty;
  wire              writeIndexQueue_13_almostFull;
  wire              writeIndexQueue_13_almostEmpty;
  wire              writeIndexQueue_12_almostFull;
  wire              writeIndexQueue_12_almostEmpty;
  wire              writeIndexQueue_11_almostFull;
  wire              writeIndexQueue_11_almostEmpty;
  wire              writeIndexQueue_10_almostFull;
  wire              writeIndexQueue_10_almostEmpty;
  wire              writeIndexQueue_9_almostFull;
  wire              writeIndexQueue_9_almostEmpty;
  wire              writeIndexQueue_8_almostFull;
  wire              writeIndexQueue_8_almostEmpty;
  wire              writeIndexQueue_7_almostFull;
  wire              writeIndexQueue_7_almostEmpty;
  wire              writeIndexQueue_6_almostFull;
  wire              writeIndexQueue_6_almostEmpty;
  wire              writeIndexQueue_5_almostFull;
  wire              writeIndexQueue_5_almostEmpty;
  wire              writeIndexQueue_4_almostFull;
  wire              writeIndexQueue_4_almostEmpty;
  wire              writeIndexQueue_3_almostFull;
  wire              writeIndexQueue_3_almostEmpty;
  wire              writeIndexQueue_2_almostFull;
  wire              writeIndexQueue_2_almostEmpty;
  wire              writeIndexQueue_1_almostFull;
  wire              writeIndexQueue_1_almostEmpty;
  wire              writeIndexQueue_almostFull;
  wire              writeIndexQueue_almostEmpty;
  wire              otherUnitDataQueueVec_31_almostFull;
  wire              otherUnitDataQueueVec_31_almostEmpty;
  wire              otherUnitDataQueueVec_30_almostFull;
  wire              otherUnitDataQueueVec_30_almostEmpty;
  wire              otherUnitDataQueueVec_29_almostFull;
  wire              otherUnitDataQueueVec_29_almostEmpty;
  wire              otherUnitDataQueueVec_28_almostFull;
  wire              otherUnitDataQueueVec_28_almostEmpty;
  wire              otherUnitDataQueueVec_27_almostFull;
  wire              otherUnitDataQueueVec_27_almostEmpty;
  wire              otherUnitDataQueueVec_26_almostFull;
  wire              otherUnitDataQueueVec_26_almostEmpty;
  wire              otherUnitDataQueueVec_25_almostFull;
  wire              otherUnitDataQueueVec_25_almostEmpty;
  wire              otherUnitDataQueueVec_24_almostFull;
  wire              otherUnitDataQueueVec_24_almostEmpty;
  wire              otherUnitDataQueueVec_23_almostFull;
  wire              otherUnitDataQueueVec_23_almostEmpty;
  wire              otherUnitDataQueueVec_22_almostFull;
  wire              otherUnitDataQueueVec_22_almostEmpty;
  wire              otherUnitDataQueueVec_21_almostFull;
  wire              otherUnitDataQueueVec_21_almostEmpty;
  wire              otherUnitDataQueueVec_20_almostFull;
  wire              otherUnitDataQueueVec_20_almostEmpty;
  wire              otherUnitDataQueueVec_19_almostFull;
  wire              otherUnitDataQueueVec_19_almostEmpty;
  wire              otherUnitDataQueueVec_18_almostFull;
  wire              otherUnitDataQueueVec_18_almostEmpty;
  wire              otherUnitDataQueueVec_17_almostFull;
  wire              otherUnitDataQueueVec_17_almostEmpty;
  wire              otherUnitDataQueueVec_16_almostFull;
  wire              otherUnitDataQueueVec_16_almostEmpty;
  wire              otherUnitDataQueueVec_15_almostFull;
  wire              otherUnitDataQueueVec_15_almostEmpty;
  wire              otherUnitDataQueueVec_14_almostFull;
  wire              otherUnitDataQueueVec_14_almostEmpty;
  wire              otherUnitDataQueueVec_13_almostFull;
  wire              otherUnitDataQueueVec_13_almostEmpty;
  wire              otherUnitDataQueueVec_12_almostFull;
  wire              otherUnitDataQueueVec_12_almostEmpty;
  wire              otherUnitDataQueueVec_11_almostFull;
  wire              otherUnitDataQueueVec_11_almostEmpty;
  wire              otherUnitDataQueueVec_10_almostFull;
  wire              otherUnitDataQueueVec_10_almostEmpty;
  wire              otherUnitDataQueueVec_9_almostFull;
  wire              otherUnitDataQueueVec_9_almostEmpty;
  wire              otherUnitDataQueueVec_8_almostFull;
  wire              otherUnitDataQueueVec_8_almostEmpty;
  wire              otherUnitDataQueueVec_7_almostFull;
  wire              otherUnitDataQueueVec_7_almostEmpty;
  wire              otherUnitDataQueueVec_6_almostFull;
  wire              otherUnitDataQueueVec_6_almostEmpty;
  wire              otherUnitDataQueueVec_5_almostFull;
  wire              otherUnitDataQueueVec_5_almostEmpty;
  wire              otherUnitDataQueueVec_4_almostFull;
  wire              otherUnitDataQueueVec_4_almostEmpty;
  wire              otherUnitDataQueueVec_3_almostFull;
  wire              otherUnitDataQueueVec_3_almostEmpty;
  wire              otherUnitDataQueueVec_2_almostFull;
  wire              otherUnitDataQueueVec_2_almostEmpty;
  wire              otherUnitDataQueueVec_1_almostFull;
  wire              otherUnitDataQueueVec_1_almostEmpty;
  wire              otherUnitDataQueueVec_0_almostFull;
  wire              otherUnitDataQueueVec_0_almostEmpty;
  wire              otherUnitTargetQueue_almostFull;
  wire              otherUnitTargetQueue_almostEmpty;
  wire              writeQueueVec_31_almostFull;
  wire              writeQueueVec_31_almostEmpty;
  wire              writeQueueVec_30_almostFull;
  wire              writeQueueVec_30_almostEmpty;
  wire              writeQueueVec_29_almostFull;
  wire              writeQueueVec_29_almostEmpty;
  wire              writeQueueVec_28_almostFull;
  wire              writeQueueVec_28_almostEmpty;
  wire              writeQueueVec_27_almostFull;
  wire              writeQueueVec_27_almostEmpty;
  wire              writeQueueVec_26_almostFull;
  wire              writeQueueVec_26_almostEmpty;
  wire              writeQueueVec_25_almostFull;
  wire              writeQueueVec_25_almostEmpty;
  wire              writeQueueVec_24_almostFull;
  wire              writeQueueVec_24_almostEmpty;
  wire              writeQueueVec_23_almostFull;
  wire              writeQueueVec_23_almostEmpty;
  wire              writeQueueVec_22_almostFull;
  wire              writeQueueVec_22_almostEmpty;
  wire              writeQueueVec_21_almostFull;
  wire              writeQueueVec_21_almostEmpty;
  wire              writeQueueVec_20_almostFull;
  wire              writeQueueVec_20_almostEmpty;
  wire              writeQueueVec_19_almostFull;
  wire              writeQueueVec_19_almostEmpty;
  wire              writeQueueVec_18_almostFull;
  wire              writeQueueVec_18_almostEmpty;
  wire              writeQueueVec_17_almostFull;
  wire              writeQueueVec_17_almostEmpty;
  wire              writeQueueVec_16_almostFull;
  wire              writeQueueVec_16_almostEmpty;
  wire              writeQueueVec_15_almostFull;
  wire              writeQueueVec_15_almostEmpty;
  wire              writeQueueVec_14_almostFull;
  wire              writeQueueVec_14_almostEmpty;
  wire              writeQueueVec_13_almostFull;
  wire              writeQueueVec_13_almostEmpty;
  wire              writeQueueVec_12_almostFull;
  wire              writeQueueVec_12_almostEmpty;
  wire              writeQueueVec_11_almostFull;
  wire              writeQueueVec_11_almostEmpty;
  wire              writeQueueVec_10_almostFull;
  wire              writeQueueVec_10_almostEmpty;
  wire              writeQueueVec_9_almostFull;
  wire              writeQueueVec_9_almostEmpty;
  wire              writeQueueVec_8_almostFull;
  wire              writeQueueVec_8_almostEmpty;
  wire              writeQueueVec_7_almostFull;
  wire              writeQueueVec_7_almostEmpty;
  wire              writeQueueVec_6_almostFull;
  wire              writeQueueVec_6_almostEmpty;
  wire              writeQueueVec_5_almostFull;
  wire              writeQueueVec_5_almostEmpty;
  wire              writeQueueVec_4_almostFull;
  wire              writeQueueVec_4_almostEmpty;
  wire              writeQueueVec_3_almostFull;
  wire              writeQueueVec_3_almostEmpty;
  wire              writeQueueVec_2_almostFull;
  wire              writeQueueVec_2_almostEmpty;
  wire              writeQueueVec_1_almostFull;
  wire              writeQueueVec_1_almostEmpty;
  wire              writeQueueVec_0_almostFull;
  wire              writeQueueVec_0_almostEmpty;
  wire [9:0]        simpleSourceQueue_enq_bits;
  wire [31:0]       simpleAccessPorts_ar_bits_addr_0;
  wire [3:0]        sourceQueue_enq_bits;
  wire [31:0]       axi4Port_ar_bits_addr_0;
  wire [4:0]        writeQueueVec_31_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_30_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_29_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_28_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_27_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_26_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_25_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_24_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_23_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_22_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_21_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_20_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_19_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_18_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_17_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_16_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_15_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_14_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_13_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_12_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_11_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_10_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_9_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_8_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_7_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_6_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_5_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_4_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_3_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_2_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_1_enq_bits_data_vd;
  wire [4:0]        writeQueueVec_0_enq_bits_data_vd;
  wire              request_valid_0 = request_valid;
  wire [2:0]        request_bits_instructionInformation_nf_0 = request_bits_instructionInformation_nf;
  wire              request_bits_instructionInformation_mew_0 = request_bits_instructionInformation_mew;
  wire [1:0]        request_bits_instructionInformation_mop_0 = request_bits_instructionInformation_mop;
  wire [4:0]        request_bits_instructionInformation_lumop_0 = request_bits_instructionInformation_lumop;
  wire [1:0]        request_bits_instructionInformation_eew_0 = request_bits_instructionInformation_eew;
  wire [4:0]        request_bits_instructionInformation_vs3_0 = request_bits_instructionInformation_vs3;
  wire              request_bits_instructionInformation_isStore_0 = request_bits_instructionInformation_isStore;
  wire              request_bits_instructionInformation_maskedLoadStore_0 = request_bits_instructionInformation_maskedLoadStore;
  wire [31:0]       request_bits_rs1Data_0 = request_bits_rs1Data;
  wire [31:0]       request_bits_rs2Data_0 = request_bits_rs2Data;
  wire [2:0]        request_bits_instructionIndex_0 = request_bits_instructionIndex;
  wire              axi4Port_aw_ready_0 = axi4Port_aw_ready;
  wire              axi4Port_w_ready_0 = axi4Port_w_ready;
  wire              axi4Port_b_valid_0 = axi4Port_b_valid;
  wire [1:0]        axi4Port_b_bits_id_0 = axi4Port_b_bits_id;
  wire [1:0]        axi4Port_b_bits_resp_0 = axi4Port_b_bits_resp;
  wire              axi4Port_ar_ready_0 = axi4Port_ar_ready;
  wire              axi4Port_r_valid_0 = axi4Port_r_valid;
  wire [1:0]        axi4Port_r_bits_id_0 = axi4Port_r_bits_id;
  wire [1023:0]     axi4Port_r_bits_data_0 = axi4Port_r_bits_data;
  wire [1:0]        axi4Port_r_bits_resp_0 = axi4Port_r_bits_resp;
  wire              axi4Port_r_bits_last_0 = axi4Port_r_bits_last;
  wire              simpleAccessPorts_aw_ready_0 = simpleAccessPorts_aw_ready;
  wire              simpleAccessPorts_w_ready_0 = simpleAccessPorts_w_ready;
  wire              simpleAccessPorts_b_valid_0 = simpleAccessPorts_b_valid;
  wire [1:0]        simpleAccessPorts_b_bits_id_0 = simpleAccessPorts_b_bits_id;
  wire [1:0]        simpleAccessPorts_b_bits_resp_0 = simpleAccessPorts_b_bits_resp;
  wire              simpleAccessPorts_ar_ready_0 = simpleAccessPorts_ar_ready;
  wire              simpleAccessPorts_r_valid_0 = simpleAccessPorts_r_valid;
  wire [1:0]        simpleAccessPorts_r_bits_id_0 = simpleAccessPorts_r_bits_id;
  wire [31:0]       simpleAccessPorts_r_bits_data_0 = simpleAccessPorts_r_bits_data;
  wire [1:0]        simpleAccessPorts_r_bits_resp_0 = simpleAccessPorts_r_bits_resp;
  wire              simpleAccessPorts_r_bits_last_0 = simpleAccessPorts_r_bits_last;
  wire              vrfReadDataPorts_0_ready_0 = vrfReadDataPorts_0_ready;
  wire              vrfReadDataPorts_1_ready_0 = vrfReadDataPorts_1_ready;
  wire              vrfReadDataPorts_2_ready_0 = vrfReadDataPorts_2_ready;
  wire              vrfReadDataPorts_3_ready_0 = vrfReadDataPorts_3_ready;
  wire              vrfReadDataPorts_4_ready_0 = vrfReadDataPorts_4_ready;
  wire              vrfReadDataPorts_5_ready_0 = vrfReadDataPorts_5_ready;
  wire              vrfReadDataPorts_6_ready_0 = vrfReadDataPorts_6_ready;
  wire              vrfReadDataPorts_7_ready_0 = vrfReadDataPorts_7_ready;
  wire              vrfReadDataPorts_8_ready_0 = vrfReadDataPorts_8_ready;
  wire              vrfReadDataPorts_9_ready_0 = vrfReadDataPorts_9_ready;
  wire              vrfReadDataPorts_10_ready_0 = vrfReadDataPorts_10_ready;
  wire              vrfReadDataPorts_11_ready_0 = vrfReadDataPorts_11_ready;
  wire              vrfReadDataPorts_12_ready_0 = vrfReadDataPorts_12_ready;
  wire              vrfReadDataPorts_13_ready_0 = vrfReadDataPorts_13_ready;
  wire              vrfReadDataPorts_14_ready_0 = vrfReadDataPorts_14_ready;
  wire              vrfReadDataPorts_15_ready_0 = vrfReadDataPorts_15_ready;
  wire              vrfReadDataPorts_16_ready_0 = vrfReadDataPorts_16_ready;
  wire              vrfReadDataPorts_17_ready_0 = vrfReadDataPorts_17_ready;
  wire              vrfReadDataPorts_18_ready_0 = vrfReadDataPorts_18_ready;
  wire              vrfReadDataPorts_19_ready_0 = vrfReadDataPorts_19_ready;
  wire              vrfReadDataPorts_20_ready_0 = vrfReadDataPorts_20_ready;
  wire              vrfReadDataPorts_21_ready_0 = vrfReadDataPorts_21_ready;
  wire              vrfReadDataPorts_22_ready_0 = vrfReadDataPorts_22_ready;
  wire              vrfReadDataPorts_23_ready_0 = vrfReadDataPorts_23_ready;
  wire              vrfReadDataPorts_24_ready_0 = vrfReadDataPorts_24_ready;
  wire              vrfReadDataPorts_25_ready_0 = vrfReadDataPorts_25_ready;
  wire              vrfReadDataPorts_26_ready_0 = vrfReadDataPorts_26_ready;
  wire              vrfReadDataPorts_27_ready_0 = vrfReadDataPorts_27_ready;
  wire              vrfReadDataPorts_28_ready_0 = vrfReadDataPorts_28_ready;
  wire              vrfReadDataPorts_29_ready_0 = vrfReadDataPorts_29_ready;
  wire              vrfReadDataPorts_30_ready_0 = vrfReadDataPorts_30_ready;
  wire              vrfReadDataPorts_31_ready_0 = vrfReadDataPorts_31_ready;
  wire              vrfWritePort_0_ready_0 = vrfWritePort_0_ready;
  wire              vrfWritePort_1_ready_0 = vrfWritePort_1_ready;
  wire              vrfWritePort_2_ready_0 = vrfWritePort_2_ready;
  wire              vrfWritePort_3_ready_0 = vrfWritePort_3_ready;
  wire              vrfWritePort_4_ready_0 = vrfWritePort_4_ready;
  wire              vrfWritePort_5_ready_0 = vrfWritePort_5_ready;
  wire              vrfWritePort_6_ready_0 = vrfWritePort_6_ready;
  wire              vrfWritePort_7_ready_0 = vrfWritePort_7_ready;
  wire              vrfWritePort_8_ready_0 = vrfWritePort_8_ready;
  wire              vrfWritePort_9_ready_0 = vrfWritePort_9_ready;
  wire              vrfWritePort_10_ready_0 = vrfWritePort_10_ready;
  wire              vrfWritePort_11_ready_0 = vrfWritePort_11_ready;
  wire              vrfWritePort_12_ready_0 = vrfWritePort_12_ready;
  wire              vrfWritePort_13_ready_0 = vrfWritePort_13_ready;
  wire              vrfWritePort_14_ready_0 = vrfWritePort_14_ready;
  wire              vrfWritePort_15_ready_0 = vrfWritePort_15_ready;
  wire              vrfWritePort_16_ready_0 = vrfWritePort_16_ready;
  wire              vrfWritePort_17_ready_0 = vrfWritePort_17_ready;
  wire              vrfWritePort_18_ready_0 = vrfWritePort_18_ready;
  wire              vrfWritePort_19_ready_0 = vrfWritePort_19_ready;
  wire              vrfWritePort_20_ready_0 = vrfWritePort_20_ready;
  wire              vrfWritePort_21_ready_0 = vrfWritePort_21_ready;
  wire              vrfWritePort_22_ready_0 = vrfWritePort_22_ready;
  wire              vrfWritePort_23_ready_0 = vrfWritePort_23_ready;
  wire              vrfWritePort_24_ready_0 = vrfWritePort_24_ready;
  wire              vrfWritePort_25_ready_0 = vrfWritePort_25_ready;
  wire              vrfWritePort_26_ready_0 = vrfWritePort_26_ready;
  wire              vrfWritePort_27_ready_0 = vrfWritePort_27_ready;
  wire              vrfWritePort_28_ready_0 = vrfWritePort_28_ready;
  wire              vrfWritePort_29_ready_0 = vrfWritePort_29_ready;
  wire              vrfWritePort_30_ready_0 = vrfWritePort_30_ready;
  wire              vrfWritePort_31_ready_0 = vrfWritePort_31_ready;
  wire [31:0]       otherUnitDataQueueVec_0_enq_bits = vrfReadResults_0_bits;
  wire [31:0]       otherUnitDataQueueVec_1_enq_bits = vrfReadResults_1_bits;
  wire [31:0]       otherUnitDataQueueVec_2_enq_bits = vrfReadResults_2_bits;
  wire [31:0]       otherUnitDataQueueVec_3_enq_bits = vrfReadResults_3_bits;
  wire [31:0]       otherUnitDataQueueVec_4_enq_bits = vrfReadResults_4_bits;
  wire [31:0]       otherUnitDataQueueVec_5_enq_bits = vrfReadResults_5_bits;
  wire [31:0]       otherUnitDataQueueVec_6_enq_bits = vrfReadResults_6_bits;
  wire [31:0]       otherUnitDataQueueVec_7_enq_bits = vrfReadResults_7_bits;
  wire [31:0]       otherUnitDataQueueVec_8_enq_bits = vrfReadResults_8_bits;
  wire [31:0]       otherUnitDataQueueVec_9_enq_bits = vrfReadResults_9_bits;
  wire [31:0]       otherUnitDataQueueVec_10_enq_bits = vrfReadResults_10_bits;
  wire [31:0]       otherUnitDataQueueVec_11_enq_bits = vrfReadResults_11_bits;
  wire [31:0]       otherUnitDataQueueVec_12_enq_bits = vrfReadResults_12_bits;
  wire [31:0]       otherUnitDataQueueVec_13_enq_bits = vrfReadResults_13_bits;
  wire [31:0]       otherUnitDataQueueVec_14_enq_bits = vrfReadResults_14_bits;
  wire [31:0]       otherUnitDataQueueVec_15_enq_bits = vrfReadResults_15_bits;
  wire [31:0]       otherUnitDataQueueVec_16_enq_bits = vrfReadResults_16_bits;
  wire [31:0]       otherUnitDataQueueVec_17_enq_bits = vrfReadResults_17_bits;
  wire [31:0]       otherUnitDataQueueVec_18_enq_bits = vrfReadResults_18_bits;
  wire [31:0]       otherUnitDataQueueVec_19_enq_bits = vrfReadResults_19_bits;
  wire [31:0]       otherUnitDataQueueVec_20_enq_bits = vrfReadResults_20_bits;
  wire [31:0]       otherUnitDataQueueVec_21_enq_bits = vrfReadResults_21_bits;
  wire [31:0]       otherUnitDataQueueVec_22_enq_bits = vrfReadResults_22_bits;
  wire [31:0]       otherUnitDataQueueVec_23_enq_bits = vrfReadResults_23_bits;
  wire [31:0]       otherUnitDataQueueVec_24_enq_bits = vrfReadResults_24_bits;
  wire [31:0]       otherUnitDataQueueVec_25_enq_bits = vrfReadResults_25_bits;
  wire [31:0]       otherUnitDataQueueVec_26_enq_bits = vrfReadResults_26_bits;
  wire [31:0]       otherUnitDataQueueVec_27_enq_bits = vrfReadResults_27_bits;
  wire [31:0]       otherUnitDataQueueVec_28_enq_bits = vrfReadResults_28_bits;
  wire [31:0]       otherUnitDataQueueVec_29_enq_bits = vrfReadResults_29_bits;
  wire [31:0]       otherUnitDataQueueVec_30_enq_bits = vrfReadResults_30_bits;
  wire [31:0]       otherUnitDataQueueVec_31_enq_bits = vrfReadResults_31_bits;
  wire              writeIndexQueue_deq_ready = writeRelease_0;
  wire              writeIndexQueue_1_deq_ready = writeRelease_1;
  wire              writeIndexQueue_2_deq_ready = writeRelease_2;
  wire              writeIndexQueue_3_deq_ready = writeRelease_3;
  wire              writeIndexQueue_4_deq_ready = writeRelease_4;
  wire              writeIndexQueue_5_deq_ready = writeRelease_5;
  wire              writeIndexQueue_6_deq_ready = writeRelease_6;
  wire              writeIndexQueue_7_deq_ready = writeRelease_7;
  wire              writeIndexQueue_8_deq_ready = writeRelease_8;
  wire              writeIndexQueue_9_deq_ready = writeRelease_9;
  wire              writeIndexQueue_10_deq_ready = writeRelease_10;
  wire              writeIndexQueue_11_deq_ready = writeRelease_11;
  wire              writeIndexQueue_12_deq_ready = writeRelease_12;
  wire              writeIndexQueue_13_deq_ready = writeRelease_13;
  wire              writeIndexQueue_14_deq_ready = writeRelease_14;
  wire              writeIndexQueue_15_deq_ready = writeRelease_15;
  wire              writeIndexQueue_16_deq_ready = writeRelease_16;
  wire              writeIndexQueue_17_deq_ready = writeRelease_17;
  wire              writeIndexQueue_18_deq_ready = writeRelease_18;
  wire              writeIndexQueue_19_deq_ready = writeRelease_19;
  wire              writeIndexQueue_20_deq_ready = writeRelease_20;
  wire              writeIndexQueue_21_deq_ready = writeRelease_21;
  wire              writeIndexQueue_22_deq_ready = writeRelease_22;
  wire              writeIndexQueue_23_deq_ready = writeRelease_23;
  wire              writeIndexQueue_24_deq_ready = writeRelease_24;
  wire              writeIndexQueue_25_deq_ready = writeRelease_25;
  wire              writeIndexQueue_26_deq_ready = writeRelease_26;
  wire              writeIndexQueue_27_deq_ready = writeRelease_27;
  wire              writeIndexQueue_28_deq_ready = writeRelease_28;
  wire              writeIndexQueue_29_deq_ready = writeRelease_29;
  wire              writeIndexQueue_30_deq_ready = writeRelease_30;
  wire              writeIndexQueue_31_deq_ready = writeRelease_31;
  wire [31:0]       writeQueueVec_0_enq_bits_targetLane = 32'h1;
  wire [31:0]       writeQueueVec_1_enq_bits_targetLane = 32'h2;
  wire [31:0]       writeQueueVec_2_enq_bits_targetLane = 32'h4;
  wire [31:0]       writeQueueVec_3_enq_bits_targetLane = 32'h8;
  wire [31:0]       writeQueueVec_4_enq_bits_targetLane = 32'h10;
  wire [31:0]       writeQueueVec_5_enq_bits_targetLane = 32'h20;
  wire [31:0]       writeQueueVec_6_enq_bits_targetLane = 32'h40;
  wire [31:0]       writeQueueVec_7_enq_bits_targetLane = 32'h80;
  wire [31:0]       writeQueueVec_8_enq_bits_targetLane = 32'h100;
  wire [31:0]       writeQueueVec_9_enq_bits_targetLane = 32'h200;
  wire [31:0]       writeQueueVec_10_enq_bits_targetLane = 32'h400;
  wire [31:0]       writeQueueVec_11_enq_bits_targetLane = 32'h800;
  wire [31:0]       writeQueueVec_12_enq_bits_targetLane = 32'h1000;
  wire [31:0]       writeQueueVec_13_enq_bits_targetLane = 32'h2000;
  wire [31:0]       writeQueueVec_14_enq_bits_targetLane = 32'h4000;
  wire [31:0]       writeQueueVec_15_enq_bits_targetLane = 32'h8000;
  wire [31:0]       writeQueueVec_16_enq_bits_targetLane = 32'h10000;
  wire [31:0]       writeQueueVec_17_enq_bits_targetLane = 32'h20000;
  wire [31:0]       writeQueueVec_18_enq_bits_targetLane = 32'h40000;
  wire [31:0]       writeQueueVec_19_enq_bits_targetLane = 32'h80000;
  wire [31:0]       writeQueueVec_20_enq_bits_targetLane = 32'h100000;
  wire [31:0]       writeQueueVec_21_enq_bits_targetLane = 32'h200000;
  wire [31:0]       writeQueueVec_22_enq_bits_targetLane = 32'h400000;
  wire [31:0]       writeQueueVec_23_enq_bits_targetLane = 32'h800000;
  wire [31:0]       writeQueueVec_24_enq_bits_targetLane = 32'h1000000;
  wire [31:0]       writeQueueVec_25_enq_bits_targetLane = 32'h2000000;
  wire [31:0]       writeQueueVec_26_enq_bits_targetLane = 32'h4000000;
  wire [31:0]       writeQueueVec_27_enq_bits_targetLane = 32'h8000000;
  wire [31:0]       writeQueueVec_28_enq_bits_targetLane = 32'h10000000;
  wire [31:0]       writeQueueVec_29_enq_bits_targetLane = 32'h20000000;
  wire [31:0]       writeQueueVec_30_enq_bits_targetLane = 32'h40000000;
  wire [31:0]       writeQueueVec_31_enq_bits_targetLane = 32'h80000000;
  wire [7:0]        axi4Port_aw_bits_len = 8'h0;
  wire [7:0]        axi4Port_ar_bits_len = 8'h0;
  wire [7:0]        simpleAccessPorts_aw_bits_len = 8'h0;
  wire [7:0]        simpleAccessPorts_ar_bits_len = 8'h0;
  wire [2:0]        axi4Port_aw_bits_size = 3'h7;
  wire [2:0]        axi4Port_ar_bits_size = 3'h7;
  wire [1:0]        axi4Port_aw_bits_burst = 2'h1;
  wire [1:0]        axi4Port_ar_bits_burst = 2'h1;
  wire [1:0]        simpleAccessPorts_aw_bits_burst = 2'h1;
  wire [1:0]        simpleAccessPorts_ar_bits_burst = 2'h1;
  wire              axi4Port_aw_bits_lock = 1'h0;
  wire              axi4Port_ar_bits_lock = 1'h0;
  wire              simpleAccessPorts_aw_bits_lock = 1'h0;
  wire              simpleAccessPorts_ar_bits_lock = 1'h0;
  wire [3:0]        axi4Port_aw_bits_cache = 4'h0;
  wire [3:0]        axi4Port_aw_bits_qos = 4'h0;
  wire [3:0]        axi4Port_aw_bits_region = 4'h0;
  wire [3:0]        axi4Port_ar_bits_cache = 4'h0;
  wire [3:0]        axi4Port_ar_bits_qos = 4'h0;
  wire [3:0]        axi4Port_ar_bits_region = 4'h0;
  wire [3:0]        simpleAccessPorts_aw_bits_cache = 4'h0;
  wire [3:0]        simpleAccessPorts_aw_bits_qos = 4'h0;
  wire [3:0]        simpleAccessPorts_aw_bits_region = 4'h0;
  wire [3:0]        simpleAccessPorts_ar_bits_cache = 4'h0;
  wire [3:0]        simpleAccessPorts_ar_bits_qos = 4'h0;
  wire [3:0]        simpleAccessPorts_ar_bits_region = 4'h0;
  wire [2:0]        axi4Port_aw_bits_prot = 3'h0;
  wire [2:0]        axi4Port_ar_bits_prot = 3'h0;
  wire [2:0]        simpleAccessPorts_aw_bits_prot = 3'h0;
  wire [2:0]        simpleAccessPorts_ar_bits_prot = 3'h0;
  wire              axi4Port_w_bits_last = 1'h1;
  wire              axi4Port_b_ready = 1'h1;
  wire              simpleAccessPorts_w_bits_last = 1'h1;
  wire              simpleAccessPorts_b_ready = 1'h1;
  wire [1:0]        axi4Port_ar_bits_id = 2'h0;
  wire [1:0]        simpleAccessPorts_ar_bits_id = 2'h0;
  wire [2:0]        simpleAccessPorts_ar_bits_size = 3'h2;
  wire [1:0]        vrfReadDataPorts_0_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_1_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_2_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_3_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_4_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_5_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_6_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_7_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_8_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_9_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_10_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_11_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_12_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_13_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_14_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_15_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_16_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_17_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_18_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_19_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_20_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_21_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_22_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_23_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_24_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_25_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_26_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_27_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_28_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_29_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_30_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_31_bits_readSource = 2'h2;
  wire              dataQueue_deq_ready = axi4Port_w_ready_0;
  wire              dataQueue_deq_valid;
  wire [1023:0]     dataQueue_deq_bits_data;
  wire [127:0]      dataQueue_deq_bits_mask;
  wire              simpleDataQueue_deq_ready = simpleAccessPorts_w_ready_0;
  wire              simpleDataQueue_deq_valid;
  wire [31:0]       simpleDataQueue_deq_bits_data;
  wire [3:0]        simpleDataQueue_deq_bits_mask;
  wire              writeQueueVec_0_deq_ready = vrfWritePort_0_ready_0;
  wire              writeQueueVec_0_deq_valid;
  wire [4:0]        writeQueueVec_0_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_0_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_0_deq_bits_data_data;
  wire              writeQueueVec_0_deq_bits_data_last;
  wire [2:0]        writeQueueVec_0_deq_bits_data_instructionIndex;
  wire              writeQueueVec_1_deq_ready = vrfWritePort_1_ready_0;
  wire              writeQueueVec_1_deq_valid;
  wire [4:0]        writeQueueVec_1_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_1_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_1_deq_bits_data_data;
  wire              writeQueueVec_1_deq_bits_data_last;
  wire [2:0]        writeQueueVec_1_deq_bits_data_instructionIndex;
  wire              writeQueueVec_2_deq_ready = vrfWritePort_2_ready_0;
  wire              writeQueueVec_2_deq_valid;
  wire [4:0]        writeQueueVec_2_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_2_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_2_deq_bits_data_data;
  wire              writeQueueVec_2_deq_bits_data_last;
  wire [2:0]        writeQueueVec_2_deq_bits_data_instructionIndex;
  wire              writeQueueVec_3_deq_ready = vrfWritePort_3_ready_0;
  wire              writeQueueVec_3_deq_valid;
  wire [4:0]        writeQueueVec_3_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_3_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_3_deq_bits_data_data;
  wire              writeQueueVec_3_deq_bits_data_last;
  wire [2:0]        writeQueueVec_3_deq_bits_data_instructionIndex;
  wire              writeQueueVec_4_deq_ready = vrfWritePort_4_ready_0;
  wire              writeQueueVec_4_deq_valid;
  wire [4:0]        writeQueueVec_4_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_4_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_4_deq_bits_data_data;
  wire              writeQueueVec_4_deq_bits_data_last;
  wire [2:0]        writeQueueVec_4_deq_bits_data_instructionIndex;
  wire              writeQueueVec_5_deq_ready = vrfWritePort_5_ready_0;
  wire              writeQueueVec_5_deq_valid;
  wire [4:0]        writeQueueVec_5_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_5_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_5_deq_bits_data_data;
  wire              writeQueueVec_5_deq_bits_data_last;
  wire [2:0]        writeQueueVec_5_deq_bits_data_instructionIndex;
  wire              writeQueueVec_6_deq_ready = vrfWritePort_6_ready_0;
  wire              writeQueueVec_6_deq_valid;
  wire [4:0]        writeQueueVec_6_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_6_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_6_deq_bits_data_data;
  wire              writeQueueVec_6_deq_bits_data_last;
  wire [2:0]        writeQueueVec_6_deq_bits_data_instructionIndex;
  wire              writeQueueVec_7_deq_ready = vrfWritePort_7_ready_0;
  wire              writeQueueVec_7_deq_valid;
  wire [4:0]        writeQueueVec_7_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_7_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_7_deq_bits_data_data;
  wire              writeQueueVec_7_deq_bits_data_last;
  wire [2:0]        writeQueueVec_7_deq_bits_data_instructionIndex;
  wire              writeQueueVec_8_deq_ready = vrfWritePort_8_ready_0;
  wire              writeQueueVec_8_deq_valid;
  wire [4:0]        writeQueueVec_8_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_8_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_8_deq_bits_data_data;
  wire              writeQueueVec_8_deq_bits_data_last;
  wire [2:0]        writeQueueVec_8_deq_bits_data_instructionIndex;
  wire              writeQueueVec_9_deq_ready = vrfWritePort_9_ready_0;
  wire              writeQueueVec_9_deq_valid;
  wire [4:0]        writeQueueVec_9_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_9_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_9_deq_bits_data_data;
  wire              writeQueueVec_9_deq_bits_data_last;
  wire [2:0]        writeQueueVec_9_deq_bits_data_instructionIndex;
  wire              writeQueueVec_10_deq_ready = vrfWritePort_10_ready_0;
  wire              writeQueueVec_10_deq_valid;
  wire [4:0]        writeQueueVec_10_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_10_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_10_deq_bits_data_data;
  wire              writeQueueVec_10_deq_bits_data_last;
  wire [2:0]        writeQueueVec_10_deq_bits_data_instructionIndex;
  wire              writeQueueVec_11_deq_ready = vrfWritePort_11_ready_0;
  wire              writeQueueVec_11_deq_valid;
  wire [4:0]        writeQueueVec_11_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_11_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_11_deq_bits_data_data;
  wire              writeQueueVec_11_deq_bits_data_last;
  wire [2:0]        writeQueueVec_11_deq_bits_data_instructionIndex;
  wire              writeQueueVec_12_deq_ready = vrfWritePort_12_ready_0;
  wire              writeQueueVec_12_deq_valid;
  wire [4:0]        writeQueueVec_12_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_12_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_12_deq_bits_data_data;
  wire              writeQueueVec_12_deq_bits_data_last;
  wire [2:0]        writeQueueVec_12_deq_bits_data_instructionIndex;
  wire              writeQueueVec_13_deq_ready = vrfWritePort_13_ready_0;
  wire              writeQueueVec_13_deq_valid;
  wire [4:0]        writeQueueVec_13_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_13_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_13_deq_bits_data_data;
  wire              writeQueueVec_13_deq_bits_data_last;
  wire [2:0]        writeQueueVec_13_deq_bits_data_instructionIndex;
  wire              writeQueueVec_14_deq_ready = vrfWritePort_14_ready_0;
  wire              writeQueueVec_14_deq_valid;
  wire [4:0]        writeQueueVec_14_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_14_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_14_deq_bits_data_data;
  wire              writeQueueVec_14_deq_bits_data_last;
  wire [2:0]        writeQueueVec_14_deq_bits_data_instructionIndex;
  wire              writeQueueVec_15_deq_ready = vrfWritePort_15_ready_0;
  wire              writeQueueVec_15_deq_valid;
  wire [4:0]        writeQueueVec_15_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_15_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_15_deq_bits_data_data;
  wire              writeQueueVec_15_deq_bits_data_last;
  wire [2:0]        writeQueueVec_15_deq_bits_data_instructionIndex;
  wire              writeQueueVec_16_deq_ready = vrfWritePort_16_ready_0;
  wire              writeQueueVec_16_deq_valid;
  wire [4:0]        writeQueueVec_16_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_16_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_16_deq_bits_data_data;
  wire              writeQueueVec_16_deq_bits_data_last;
  wire [2:0]        writeQueueVec_16_deq_bits_data_instructionIndex;
  wire              writeQueueVec_17_deq_ready = vrfWritePort_17_ready_0;
  wire              writeQueueVec_17_deq_valid;
  wire [4:0]        writeQueueVec_17_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_17_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_17_deq_bits_data_data;
  wire              writeQueueVec_17_deq_bits_data_last;
  wire [2:0]        writeQueueVec_17_deq_bits_data_instructionIndex;
  wire              writeQueueVec_18_deq_ready = vrfWritePort_18_ready_0;
  wire              writeQueueVec_18_deq_valid;
  wire [4:0]        writeQueueVec_18_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_18_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_18_deq_bits_data_data;
  wire              writeQueueVec_18_deq_bits_data_last;
  wire [2:0]        writeQueueVec_18_deq_bits_data_instructionIndex;
  wire              writeQueueVec_19_deq_ready = vrfWritePort_19_ready_0;
  wire              writeQueueVec_19_deq_valid;
  wire [4:0]        writeQueueVec_19_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_19_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_19_deq_bits_data_data;
  wire              writeQueueVec_19_deq_bits_data_last;
  wire [2:0]        writeQueueVec_19_deq_bits_data_instructionIndex;
  wire              writeQueueVec_20_deq_ready = vrfWritePort_20_ready_0;
  wire              writeQueueVec_20_deq_valid;
  wire [4:0]        writeQueueVec_20_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_20_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_20_deq_bits_data_data;
  wire              writeQueueVec_20_deq_bits_data_last;
  wire [2:0]        writeQueueVec_20_deq_bits_data_instructionIndex;
  wire              writeQueueVec_21_deq_ready = vrfWritePort_21_ready_0;
  wire              writeQueueVec_21_deq_valid;
  wire [4:0]        writeQueueVec_21_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_21_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_21_deq_bits_data_data;
  wire              writeQueueVec_21_deq_bits_data_last;
  wire [2:0]        writeQueueVec_21_deq_bits_data_instructionIndex;
  wire              writeQueueVec_22_deq_ready = vrfWritePort_22_ready_0;
  wire              writeQueueVec_22_deq_valid;
  wire [4:0]        writeQueueVec_22_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_22_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_22_deq_bits_data_data;
  wire              writeQueueVec_22_deq_bits_data_last;
  wire [2:0]        writeQueueVec_22_deq_bits_data_instructionIndex;
  wire              writeQueueVec_23_deq_ready = vrfWritePort_23_ready_0;
  wire              writeQueueVec_23_deq_valid;
  wire [4:0]        writeQueueVec_23_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_23_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_23_deq_bits_data_data;
  wire              writeQueueVec_23_deq_bits_data_last;
  wire [2:0]        writeQueueVec_23_deq_bits_data_instructionIndex;
  wire              writeQueueVec_24_deq_ready = vrfWritePort_24_ready_0;
  wire              writeQueueVec_24_deq_valid;
  wire [4:0]        writeQueueVec_24_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_24_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_24_deq_bits_data_data;
  wire              writeQueueVec_24_deq_bits_data_last;
  wire [2:0]        writeQueueVec_24_deq_bits_data_instructionIndex;
  wire              writeQueueVec_25_deq_ready = vrfWritePort_25_ready_0;
  wire              writeQueueVec_25_deq_valid;
  wire [4:0]        writeQueueVec_25_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_25_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_25_deq_bits_data_data;
  wire              writeQueueVec_25_deq_bits_data_last;
  wire [2:0]        writeQueueVec_25_deq_bits_data_instructionIndex;
  wire              writeQueueVec_26_deq_ready = vrfWritePort_26_ready_0;
  wire              writeQueueVec_26_deq_valid;
  wire [4:0]        writeQueueVec_26_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_26_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_26_deq_bits_data_data;
  wire              writeQueueVec_26_deq_bits_data_last;
  wire [2:0]        writeQueueVec_26_deq_bits_data_instructionIndex;
  wire              writeQueueVec_27_deq_ready = vrfWritePort_27_ready_0;
  wire              writeQueueVec_27_deq_valid;
  wire [4:0]        writeQueueVec_27_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_27_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_27_deq_bits_data_data;
  wire              writeQueueVec_27_deq_bits_data_last;
  wire [2:0]        writeQueueVec_27_deq_bits_data_instructionIndex;
  wire              writeQueueVec_28_deq_ready = vrfWritePort_28_ready_0;
  wire              writeQueueVec_28_deq_valid;
  wire [4:0]        writeQueueVec_28_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_28_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_28_deq_bits_data_data;
  wire              writeQueueVec_28_deq_bits_data_last;
  wire [2:0]        writeQueueVec_28_deq_bits_data_instructionIndex;
  wire              writeQueueVec_29_deq_ready = vrfWritePort_29_ready_0;
  wire              writeQueueVec_29_deq_valid;
  wire [4:0]        writeQueueVec_29_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_29_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_29_deq_bits_data_data;
  wire              writeQueueVec_29_deq_bits_data_last;
  wire [2:0]        writeQueueVec_29_deq_bits_data_instructionIndex;
  wire              writeQueueVec_30_deq_ready = vrfWritePort_30_ready_0;
  wire              writeQueueVec_30_deq_valid;
  wire [4:0]        writeQueueVec_30_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_30_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_30_deq_bits_data_data;
  wire              writeQueueVec_30_deq_bits_data_last;
  wire [2:0]        writeQueueVec_30_deq_bits_data_instructionIndex;
  wire              writeQueueVec_31_deq_ready = vrfWritePort_31_ready_0;
  wire              writeQueueVec_31_deq_valid;
  wire [4:0]        writeQueueVec_31_deq_bits_data_vd;
  wire [3:0]        writeQueueVec_31_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_31_deq_bits_data_data;
  wire              writeQueueVec_31_deq_bits_data_last;
  wire [2:0]        writeQueueVec_31_deq_bits_data_instructionIndex;
  reg  [31:0]       v0_0;
  reg  [31:0]       v0_1;
  reg  [31:0]       v0_2;
  reg  [31:0]       v0_3;
  reg  [31:0]       v0_4;
  reg  [31:0]       v0_5;
  reg  [31:0]       v0_6;
  reg  [31:0]       v0_7;
  reg  [31:0]       v0_8;
  reg  [31:0]       v0_9;
  reg  [31:0]       v0_10;
  reg  [31:0]       v0_11;
  reg  [31:0]       v0_12;
  reg  [31:0]       v0_13;
  reg  [31:0]       v0_14;
  reg  [31:0]       v0_15;
  reg  [31:0]       v0_16;
  reg  [31:0]       v0_17;
  reg  [31:0]       v0_18;
  reg  [31:0]       v0_19;
  reg  [31:0]       v0_20;
  reg  [31:0]       v0_21;
  reg  [31:0]       v0_22;
  reg  [31:0]       v0_23;
  reg  [31:0]       v0_24;
  reg  [31:0]       v0_25;
  reg  [31:0]       v0_26;
  reg  [31:0]       v0_27;
  reg  [31:0]       v0_28;
  reg  [31:0]       v0_29;
  reg  [31:0]       v0_30;
  reg  [31:0]       v0_31;
  wire [15:0]       maskExt_lo = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]       maskExt_hi = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]       maskExt = {maskExt_hi, maskExt_lo};
  wire [15:0]       maskExt_lo_1 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_1 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]       maskExt_1 = {maskExt_hi_1, maskExt_lo_1};
  wire [15:0]       maskExt_lo_2 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_2 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]       maskExt_2 = {maskExt_hi_2, maskExt_lo_2};
  wire [15:0]       maskExt_lo_3 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_3 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]       maskExt_3 = {maskExt_hi_3, maskExt_lo_3};
  wire [15:0]       maskExt_lo_4 = {{8{v0UpdateVec_4_bits_mask[1]}}, {8{v0UpdateVec_4_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_4 = {{8{v0UpdateVec_4_bits_mask[3]}}, {8{v0UpdateVec_4_bits_mask[2]}}};
  wire [31:0]       maskExt_4 = {maskExt_hi_4, maskExt_lo_4};
  wire [15:0]       maskExt_lo_5 = {{8{v0UpdateVec_5_bits_mask[1]}}, {8{v0UpdateVec_5_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_5 = {{8{v0UpdateVec_5_bits_mask[3]}}, {8{v0UpdateVec_5_bits_mask[2]}}};
  wire [31:0]       maskExt_5 = {maskExt_hi_5, maskExt_lo_5};
  wire [15:0]       maskExt_lo_6 = {{8{v0UpdateVec_6_bits_mask[1]}}, {8{v0UpdateVec_6_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_6 = {{8{v0UpdateVec_6_bits_mask[3]}}, {8{v0UpdateVec_6_bits_mask[2]}}};
  wire [31:0]       maskExt_6 = {maskExt_hi_6, maskExt_lo_6};
  wire [15:0]       maskExt_lo_7 = {{8{v0UpdateVec_7_bits_mask[1]}}, {8{v0UpdateVec_7_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_7 = {{8{v0UpdateVec_7_bits_mask[3]}}, {8{v0UpdateVec_7_bits_mask[2]}}};
  wire [31:0]       maskExt_7 = {maskExt_hi_7, maskExt_lo_7};
  wire [15:0]       maskExt_lo_8 = {{8{v0UpdateVec_8_bits_mask[1]}}, {8{v0UpdateVec_8_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_8 = {{8{v0UpdateVec_8_bits_mask[3]}}, {8{v0UpdateVec_8_bits_mask[2]}}};
  wire [31:0]       maskExt_8 = {maskExt_hi_8, maskExt_lo_8};
  wire [15:0]       maskExt_lo_9 = {{8{v0UpdateVec_9_bits_mask[1]}}, {8{v0UpdateVec_9_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_9 = {{8{v0UpdateVec_9_bits_mask[3]}}, {8{v0UpdateVec_9_bits_mask[2]}}};
  wire [31:0]       maskExt_9 = {maskExt_hi_9, maskExt_lo_9};
  wire [15:0]       maskExt_lo_10 = {{8{v0UpdateVec_10_bits_mask[1]}}, {8{v0UpdateVec_10_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_10 = {{8{v0UpdateVec_10_bits_mask[3]}}, {8{v0UpdateVec_10_bits_mask[2]}}};
  wire [31:0]       maskExt_10 = {maskExt_hi_10, maskExt_lo_10};
  wire [15:0]       maskExt_lo_11 = {{8{v0UpdateVec_11_bits_mask[1]}}, {8{v0UpdateVec_11_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_11 = {{8{v0UpdateVec_11_bits_mask[3]}}, {8{v0UpdateVec_11_bits_mask[2]}}};
  wire [31:0]       maskExt_11 = {maskExt_hi_11, maskExt_lo_11};
  wire [15:0]       maskExt_lo_12 = {{8{v0UpdateVec_12_bits_mask[1]}}, {8{v0UpdateVec_12_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_12 = {{8{v0UpdateVec_12_bits_mask[3]}}, {8{v0UpdateVec_12_bits_mask[2]}}};
  wire [31:0]       maskExt_12 = {maskExt_hi_12, maskExt_lo_12};
  wire [15:0]       maskExt_lo_13 = {{8{v0UpdateVec_13_bits_mask[1]}}, {8{v0UpdateVec_13_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_13 = {{8{v0UpdateVec_13_bits_mask[3]}}, {8{v0UpdateVec_13_bits_mask[2]}}};
  wire [31:0]       maskExt_13 = {maskExt_hi_13, maskExt_lo_13};
  wire [15:0]       maskExt_lo_14 = {{8{v0UpdateVec_14_bits_mask[1]}}, {8{v0UpdateVec_14_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_14 = {{8{v0UpdateVec_14_bits_mask[3]}}, {8{v0UpdateVec_14_bits_mask[2]}}};
  wire [31:0]       maskExt_14 = {maskExt_hi_14, maskExt_lo_14};
  wire [15:0]       maskExt_lo_15 = {{8{v0UpdateVec_15_bits_mask[1]}}, {8{v0UpdateVec_15_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_15 = {{8{v0UpdateVec_15_bits_mask[3]}}, {8{v0UpdateVec_15_bits_mask[2]}}};
  wire [31:0]       maskExt_15 = {maskExt_hi_15, maskExt_lo_15};
  wire [15:0]       maskExt_lo_16 = {{8{v0UpdateVec_16_bits_mask[1]}}, {8{v0UpdateVec_16_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_16 = {{8{v0UpdateVec_16_bits_mask[3]}}, {8{v0UpdateVec_16_bits_mask[2]}}};
  wire [31:0]       maskExt_16 = {maskExt_hi_16, maskExt_lo_16};
  wire [15:0]       maskExt_lo_17 = {{8{v0UpdateVec_17_bits_mask[1]}}, {8{v0UpdateVec_17_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_17 = {{8{v0UpdateVec_17_bits_mask[3]}}, {8{v0UpdateVec_17_bits_mask[2]}}};
  wire [31:0]       maskExt_17 = {maskExt_hi_17, maskExt_lo_17};
  wire [15:0]       maskExt_lo_18 = {{8{v0UpdateVec_18_bits_mask[1]}}, {8{v0UpdateVec_18_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_18 = {{8{v0UpdateVec_18_bits_mask[3]}}, {8{v0UpdateVec_18_bits_mask[2]}}};
  wire [31:0]       maskExt_18 = {maskExt_hi_18, maskExt_lo_18};
  wire [15:0]       maskExt_lo_19 = {{8{v0UpdateVec_19_bits_mask[1]}}, {8{v0UpdateVec_19_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_19 = {{8{v0UpdateVec_19_bits_mask[3]}}, {8{v0UpdateVec_19_bits_mask[2]}}};
  wire [31:0]       maskExt_19 = {maskExt_hi_19, maskExt_lo_19};
  wire [15:0]       maskExt_lo_20 = {{8{v0UpdateVec_20_bits_mask[1]}}, {8{v0UpdateVec_20_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_20 = {{8{v0UpdateVec_20_bits_mask[3]}}, {8{v0UpdateVec_20_bits_mask[2]}}};
  wire [31:0]       maskExt_20 = {maskExt_hi_20, maskExt_lo_20};
  wire [15:0]       maskExt_lo_21 = {{8{v0UpdateVec_21_bits_mask[1]}}, {8{v0UpdateVec_21_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_21 = {{8{v0UpdateVec_21_bits_mask[3]}}, {8{v0UpdateVec_21_bits_mask[2]}}};
  wire [31:0]       maskExt_21 = {maskExt_hi_21, maskExt_lo_21};
  wire [15:0]       maskExt_lo_22 = {{8{v0UpdateVec_22_bits_mask[1]}}, {8{v0UpdateVec_22_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_22 = {{8{v0UpdateVec_22_bits_mask[3]}}, {8{v0UpdateVec_22_bits_mask[2]}}};
  wire [31:0]       maskExt_22 = {maskExt_hi_22, maskExt_lo_22};
  wire [15:0]       maskExt_lo_23 = {{8{v0UpdateVec_23_bits_mask[1]}}, {8{v0UpdateVec_23_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_23 = {{8{v0UpdateVec_23_bits_mask[3]}}, {8{v0UpdateVec_23_bits_mask[2]}}};
  wire [31:0]       maskExt_23 = {maskExt_hi_23, maskExt_lo_23};
  wire [15:0]       maskExt_lo_24 = {{8{v0UpdateVec_24_bits_mask[1]}}, {8{v0UpdateVec_24_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_24 = {{8{v0UpdateVec_24_bits_mask[3]}}, {8{v0UpdateVec_24_bits_mask[2]}}};
  wire [31:0]       maskExt_24 = {maskExt_hi_24, maskExt_lo_24};
  wire [15:0]       maskExt_lo_25 = {{8{v0UpdateVec_25_bits_mask[1]}}, {8{v0UpdateVec_25_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_25 = {{8{v0UpdateVec_25_bits_mask[3]}}, {8{v0UpdateVec_25_bits_mask[2]}}};
  wire [31:0]       maskExt_25 = {maskExt_hi_25, maskExt_lo_25};
  wire [15:0]       maskExt_lo_26 = {{8{v0UpdateVec_26_bits_mask[1]}}, {8{v0UpdateVec_26_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_26 = {{8{v0UpdateVec_26_bits_mask[3]}}, {8{v0UpdateVec_26_bits_mask[2]}}};
  wire [31:0]       maskExt_26 = {maskExt_hi_26, maskExt_lo_26};
  wire [15:0]       maskExt_lo_27 = {{8{v0UpdateVec_27_bits_mask[1]}}, {8{v0UpdateVec_27_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_27 = {{8{v0UpdateVec_27_bits_mask[3]}}, {8{v0UpdateVec_27_bits_mask[2]}}};
  wire [31:0]       maskExt_27 = {maskExt_hi_27, maskExt_lo_27};
  wire [15:0]       maskExt_lo_28 = {{8{v0UpdateVec_28_bits_mask[1]}}, {8{v0UpdateVec_28_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_28 = {{8{v0UpdateVec_28_bits_mask[3]}}, {8{v0UpdateVec_28_bits_mask[2]}}};
  wire [31:0]       maskExt_28 = {maskExt_hi_28, maskExt_lo_28};
  wire [15:0]       maskExt_lo_29 = {{8{v0UpdateVec_29_bits_mask[1]}}, {8{v0UpdateVec_29_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_29 = {{8{v0UpdateVec_29_bits_mask[3]}}, {8{v0UpdateVec_29_bits_mask[2]}}};
  wire [31:0]       maskExt_29 = {maskExt_hi_29, maskExt_lo_29};
  wire [15:0]       maskExt_lo_30 = {{8{v0UpdateVec_30_bits_mask[1]}}, {8{v0UpdateVec_30_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_30 = {{8{v0UpdateVec_30_bits_mask[3]}}, {8{v0UpdateVec_30_bits_mask[2]}}};
  wire [31:0]       maskExt_30 = {maskExt_hi_30, maskExt_lo_30};
  wire [15:0]       maskExt_lo_31 = {{8{v0UpdateVec_31_bits_mask[1]}}, {8{v0UpdateVec_31_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_31 = {{8{v0UpdateVec_31_bits_mask[3]}}, {8{v0UpdateVec_31_bits_mask[2]}}};
  wire [31:0]       maskExt_31 = {maskExt_hi_31, maskExt_lo_31};
  wire              alwaysMerge = {request_bits_instructionInformation_mop_0, request_bits_instructionInformation_lumop_0[2:0], request_bits_instructionInformation_lumop_0[4]} == 6'h0;
  wire              useLoadUnit = alwaysMerge & ~request_bits_instructionInformation_isStore_0;
  wire              useStoreUnit = alwaysMerge & request_bits_instructionInformation_isStore_0;
  wire              useOtherUnit = ~alwaysMerge;
  wire              addressCheck = _otherUnit_status_idle & (~useOtherUnit | _loadUnit_status_idle & _storeUnit_status_idle);
  wire              unitReady = useLoadUnit & _loadUnit_status_idle | useStoreUnit & _storeUnit_status_idle | useOtherUnit & _otherUnit_status_idle;
  wire              request_ready_0 = unitReady & addressCheck;
  wire              requestFire = request_ready_0 & request_valid_0;
  wire              reqEnq_0 = useLoadUnit & requestFire;
  wire              reqEnq_1 = useStoreUnit & requestFire;
  wire              reqEnq_2 = useOtherUnit & requestFire;
  wire [2:0]        maskSelect = _loadUnit_maskSelect_valid ? _loadUnit_maskSelect_bits : 3'h0;
  wire [63:0]       _GEN = {v0_1, v0_0};
  wire [63:0]       loadUnit_maskInput_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo = _GEN;
  wire [63:0]       storeUnit_maskInput_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo = _GEN;
  wire [63:0]       otherUnit_maskInput_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo = _GEN;
  wire [63:0]       _GEN_0 = {v0_3, v0_2};
  wire [63:0]       loadUnit_maskInput_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi = _GEN_0;
  wire [63:0]       storeUnit_maskInput_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi = _GEN_0;
  wire [63:0]       otherUnit_maskInput_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi = _GEN_0;
  wire [127:0]      loadUnit_maskInput_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo};
  wire [63:0]       _GEN_1 = {v0_5, v0_4};
  wire [63:0]       loadUnit_maskInput_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo = _GEN_1;
  wire [63:0]       storeUnit_maskInput_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo = _GEN_1;
  wire [63:0]       otherUnit_maskInput_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo = _GEN_1;
  wire [63:0]       _GEN_2 = {v0_7, v0_6};
  wire [63:0]       loadUnit_maskInput_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi = _GEN_2;
  wire [63:0]       storeUnit_maskInput_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi = _GEN_2;
  wire [63:0]       otherUnit_maskInput_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi = _GEN_2;
  wire [127:0]      loadUnit_maskInput_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo};
  wire [255:0]      loadUnit_maskInput_lo_lo = {loadUnit_maskInput_lo_lo_hi, loadUnit_maskInput_lo_lo_lo};
  wire [63:0]       _GEN_3 = {v0_9, v0_8};
  wire [63:0]       loadUnit_maskInput_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo = _GEN_3;
  wire [63:0]       storeUnit_maskInput_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo = _GEN_3;
  wire [63:0]       otherUnit_maskInput_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo = _GEN_3;
  wire [63:0]       _GEN_4 = {v0_11, v0_10};
  wire [63:0]       loadUnit_maskInput_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi = _GEN_4;
  wire [63:0]       storeUnit_maskInput_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi = _GEN_4;
  wire [63:0]       otherUnit_maskInput_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi = _GEN_4;
  wire [127:0]      loadUnit_maskInput_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo};
  wire [63:0]       _GEN_5 = {v0_13, v0_12};
  wire [63:0]       loadUnit_maskInput_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo = _GEN_5;
  wire [63:0]       storeUnit_maskInput_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo = _GEN_5;
  wire [63:0]       otherUnit_maskInput_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo = _GEN_5;
  wire [63:0]       _GEN_6 = {v0_15, v0_14};
  wire [63:0]       loadUnit_maskInput_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi = _GEN_6;
  wire [63:0]       storeUnit_maskInput_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi = _GEN_6;
  wire [63:0]       otherUnit_maskInput_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi = _GEN_6;
  wire [127:0]      loadUnit_maskInput_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo};
  wire [255:0]      loadUnit_maskInput_lo_hi = {loadUnit_maskInput_lo_hi_hi, loadUnit_maskInput_lo_hi_lo};
  wire [511:0]      loadUnit_maskInput_lo = {loadUnit_maskInput_lo_hi, loadUnit_maskInput_lo_lo};
  wire [63:0]       _GEN_7 = {v0_17, v0_16};
  wire [63:0]       loadUnit_maskInput_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo = _GEN_7;
  wire [63:0]       storeUnit_maskInput_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo = _GEN_7;
  wire [63:0]       otherUnit_maskInput_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo = _GEN_7;
  wire [63:0]       _GEN_8 = {v0_19, v0_18};
  wire [63:0]       loadUnit_maskInput_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi = _GEN_8;
  wire [63:0]       storeUnit_maskInput_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi = _GEN_8;
  wire [63:0]       otherUnit_maskInput_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi = _GEN_8;
  wire [127:0]      loadUnit_maskInput_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo};
  wire [63:0]       _GEN_9 = {v0_21, v0_20};
  wire [63:0]       loadUnit_maskInput_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo = _GEN_9;
  wire [63:0]       storeUnit_maskInput_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo = _GEN_9;
  wire [63:0]       otherUnit_maskInput_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo = _GEN_9;
  wire [63:0]       _GEN_10 = {v0_23, v0_22};
  wire [63:0]       loadUnit_maskInput_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi = _GEN_10;
  wire [63:0]       storeUnit_maskInput_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi = _GEN_10;
  wire [63:0]       otherUnit_maskInput_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi = _GEN_10;
  wire [127:0]      loadUnit_maskInput_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo};
  wire [255:0]      loadUnit_maskInput_hi_lo = {loadUnit_maskInput_hi_lo_hi, loadUnit_maskInput_hi_lo_lo};
  wire [63:0]       _GEN_11 = {v0_25, v0_24};
  wire [63:0]       loadUnit_maskInput_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo = _GEN_11;
  wire [63:0]       storeUnit_maskInput_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo = _GEN_11;
  wire [63:0]       otherUnit_maskInput_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo = _GEN_11;
  wire [63:0]       _GEN_12 = {v0_27, v0_26};
  wire [63:0]       loadUnit_maskInput_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi = _GEN_12;
  wire [63:0]       storeUnit_maskInput_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi = _GEN_12;
  wire [63:0]       otherUnit_maskInput_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi = _GEN_12;
  wire [127:0]      loadUnit_maskInput_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo};
  wire [63:0]       _GEN_13 = {v0_29, v0_28};
  wire [63:0]       loadUnit_maskInput_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo = _GEN_13;
  wire [63:0]       storeUnit_maskInput_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo = _GEN_13;
  wire [63:0]       otherUnit_maskInput_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo = _GEN_13;
  wire [63:0]       _GEN_14 = {v0_31, v0_30};
  wire [63:0]       loadUnit_maskInput_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi = _GEN_14;
  wire [63:0]       storeUnit_maskInput_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi = _GEN_14;
  wire [63:0]       otherUnit_maskInput_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi = _GEN_14;
  wire [127:0]      loadUnit_maskInput_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo};
  wire [255:0]      loadUnit_maskInput_hi_hi = {loadUnit_maskInput_hi_hi_hi, loadUnit_maskInput_hi_hi_lo};
  wire [511:0]      loadUnit_maskInput_hi = {loadUnit_maskInput_hi_hi, loadUnit_maskInput_hi_lo};
  wire [7:0][127:0] _GEN_15 =
    {{loadUnit_maskInput_hi[511:384]},
     {loadUnit_maskInput_hi[383:256]},
     {loadUnit_maskInput_hi[255:128]},
     {loadUnit_maskInput_hi[127:0]},
     {loadUnit_maskInput_lo[511:384]},
     {loadUnit_maskInput_lo[383:256]},
     {loadUnit_maskInput_lo[255:128]},
     {loadUnit_maskInput_lo[127:0]}};
  wire [2:0]        maskSelect_1 = _storeUnit_maskSelect_valid ? _storeUnit_maskSelect_bits : 3'h0;
  wire [127:0]      storeUnit_maskInput_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo};
  wire [127:0]      storeUnit_maskInput_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo};
  wire [255:0]      storeUnit_maskInput_lo_lo = {storeUnit_maskInput_lo_lo_hi, storeUnit_maskInput_lo_lo_lo};
  wire [127:0]      storeUnit_maskInput_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo};
  wire [127:0]      storeUnit_maskInput_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo};
  wire [255:0]      storeUnit_maskInput_lo_hi = {storeUnit_maskInput_lo_hi_hi, storeUnit_maskInput_lo_hi_lo};
  wire [511:0]      storeUnit_maskInput_lo = {storeUnit_maskInput_lo_hi, storeUnit_maskInput_lo_lo};
  wire [127:0]      storeUnit_maskInput_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo};
  wire [127:0]      storeUnit_maskInput_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo};
  wire [255:0]      storeUnit_maskInput_hi_lo = {storeUnit_maskInput_hi_lo_hi, storeUnit_maskInput_hi_lo_lo};
  wire [127:0]      storeUnit_maskInput_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo};
  wire [127:0]      storeUnit_maskInput_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo};
  wire [255:0]      storeUnit_maskInput_hi_hi = {storeUnit_maskInput_hi_hi_hi, storeUnit_maskInput_hi_hi_lo};
  wire [511:0]      storeUnit_maskInput_hi = {storeUnit_maskInput_hi_hi, storeUnit_maskInput_hi_lo};
  wire [7:0][127:0] _GEN_16 =
    {{storeUnit_maskInput_hi[511:384]},
     {storeUnit_maskInput_hi[383:256]},
     {storeUnit_maskInput_hi[255:128]},
     {storeUnit_maskInput_hi[127:0]},
     {storeUnit_maskInput_lo[511:384]},
     {storeUnit_maskInput_lo[383:256]},
     {storeUnit_maskInput_lo[255:128]},
     {storeUnit_maskInput_lo[127:0]}};
  wire [2:0]        maskSelect_2 = _otherUnit_maskSelect_valid ? _otherUnit_maskSelect_bits : 3'h0;
  wire [127:0]      otherUnit_maskInput_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo};
  wire [127:0]      otherUnit_maskInput_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo};
  wire [255:0]      otherUnit_maskInput_lo_lo = {otherUnit_maskInput_lo_lo_hi, otherUnit_maskInput_lo_lo_lo};
  wire [127:0]      otherUnit_maskInput_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo};
  wire [127:0]      otherUnit_maskInput_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo};
  wire [255:0]      otherUnit_maskInput_lo_hi = {otherUnit_maskInput_lo_hi_hi, otherUnit_maskInput_lo_hi_lo};
  wire [511:0]      otherUnit_maskInput_lo = {otherUnit_maskInput_lo_hi, otherUnit_maskInput_lo_lo};
  wire [127:0]      otherUnit_maskInput_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo};
  wire [127:0]      otherUnit_maskInput_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo};
  wire [255:0]      otherUnit_maskInput_hi_lo = {otherUnit_maskInput_hi_lo_hi, otherUnit_maskInput_hi_lo_lo};
  wire [127:0]      otherUnit_maskInput_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo};
  wire [127:0]      otherUnit_maskInput_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo};
  wire [255:0]      otherUnit_maskInput_hi_hi = {otherUnit_maskInput_hi_hi_hi, otherUnit_maskInput_hi_hi_lo};
  wire [511:0]      otherUnit_maskInput_hi = {otherUnit_maskInput_hi_hi, otherUnit_maskInput_hi_lo};
  wire [7:0][127:0] _GEN_17 =
    {{otherUnit_maskInput_hi[511:384]},
     {otherUnit_maskInput_hi[383:256]},
     {otherUnit_maskInput_hi[255:128]},
     {otherUnit_maskInput_hi[127:0]},
     {otherUnit_maskInput_lo[511:384]},
     {otherUnit_maskInput_lo[383:256]},
     {otherUnit_maskInput_lo[255:128]},
     {otherUnit_maskInput_lo[127:0]}};
  wire [4:0]        writeQueueVec_dataIn_hi_hi = writeQueueVec_0_enq_bits_data_vd;
  wire              vrfWritePort_0_valid_0 = writeQueueVec_0_deq_valid;
  wire [4:0]        vrfWritePort_0_bits_vd_0 = writeQueueVec_0_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_0_bits_mask_0 = writeQueueVec_0_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_0_bits_data_0 = writeQueueVec_0_deq_bits_data_data;
  wire              vrfWritePort_0_bits_last_0 = writeQueueVec_0_deq_bits_data_last;
  wire [2:0]        vrfWritePort_0_bits_instructionIndex_0 = writeQueueVec_0_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_enq_bits = writeQueueVec_0_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_0_enq_bits_data_data;
  wire              writeQueueVec_0_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi = {writeQueueVec_0_enq_bits_data_data, writeQueueVec_0_enq_bits_data_last};
  wire [2:0]        writeQueueVec_0_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo = {writeQueueVec_dataIn_lo_hi, writeQueueVec_0_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_0_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi = {writeQueueVec_dataIn_hi_hi, writeQueueVec_0_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn = {writeQueueVec_dataIn_hi, writeQueueVec_dataIn_lo, 32'h1};
  wire [31:0]       writeQueueVec_dataOut_targetLane = _writeQueueVec_fifo_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_data_instructionIndex = _writeQueueVec_fifo_data_out[34:32];
  wire              writeQueueVec_dataOut_data_last = _writeQueueVec_fifo_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_data_data = _writeQueueVec_fifo_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_data_mask = _writeQueueVec_fifo_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_data_vd = _writeQueueVec_fifo_data_out[76:72];
  wire              writeQueueVec_0_enq_ready = ~_writeQueueVec_fifo_full;
  wire              writeQueueVec_0_enq_valid;
  wire              _probeWire_slots_0_writeValid_T = writeQueueVec_0_enq_ready & writeQueueVec_0_enq_valid;
  assign writeQueueVec_0_deq_valid = ~_writeQueueVec_fifo_empty | writeQueueVec_0_enq_valid;
  assign writeQueueVec_0_deq_bits_data_vd = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_vd : writeQueueVec_dataOut_data_vd;
  assign writeQueueVec_0_deq_bits_data_mask = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_mask : writeQueueVec_dataOut_data_mask;
  assign writeQueueVec_0_deq_bits_data_data = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_data : writeQueueVec_dataOut_data_data;
  assign writeQueueVec_0_deq_bits_data_last = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_last : writeQueueVec_dataOut_data_last;
  assign writeQueueVec_0_deq_bits_data_instructionIndex = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_instructionIndex : writeQueueVec_dataOut_data_instructionIndex;
  wire [31:0]       writeQueueVec_0_deq_bits_targetLane = _writeQueueVec_fifo_empty ? 32'h1 : writeQueueVec_dataOut_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_1 = writeQueueVec_1_enq_bits_data_vd;
  wire              vrfWritePort_1_valid_0 = writeQueueVec_1_deq_valid;
  wire [4:0]        vrfWritePort_1_bits_vd_0 = writeQueueVec_1_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_1_bits_mask_0 = writeQueueVec_1_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_1_bits_data_0 = writeQueueVec_1_deq_bits_data_data;
  wire              vrfWritePort_1_bits_last_0 = writeQueueVec_1_deq_bits_data_last;
  wire [2:0]        vrfWritePort_1_bits_instructionIndex_0 = writeQueueVec_1_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_1_enq_bits = writeQueueVec_1_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_1_enq_bits_data_data;
  wire              writeQueueVec_1_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_1 = {writeQueueVec_1_enq_bits_data_data, writeQueueVec_1_enq_bits_data_last};
  wire [2:0]        writeQueueVec_1_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_1 = {writeQueueVec_dataIn_lo_hi_1, writeQueueVec_1_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_1_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_1 = {writeQueueVec_dataIn_hi_hi_1, writeQueueVec_1_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_1 = {writeQueueVec_dataIn_hi_1, writeQueueVec_dataIn_lo_1, 32'h2};
  wire [31:0]       writeQueueVec_dataOut_1_targetLane = _writeQueueVec_fifo_1_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_1_data_instructionIndex = _writeQueueVec_fifo_1_data_out[34:32];
  wire              writeQueueVec_dataOut_1_data_last = _writeQueueVec_fifo_1_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_1_data_data = _writeQueueVec_fifo_1_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_1_data_mask = _writeQueueVec_fifo_1_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_1_data_vd = _writeQueueVec_fifo_1_data_out[76:72];
  wire              writeQueueVec_1_enq_ready = ~_writeQueueVec_fifo_1_full;
  wire              writeQueueVec_1_enq_valid;
  wire              _probeWire_slots_1_writeValid_T = writeQueueVec_1_enq_ready & writeQueueVec_1_enq_valid;
  assign writeQueueVec_1_deq_valid = ~_writeQueueVec_fifo_1_empty | writeQueueVec_1_enq_valid;
  assign writeQueueVec_1_deq_bits_data_vd = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_vd : writeQueueVec_dataOut_1_data_vd;
  assign writeQueueVec_1_deq_bits_data_mask = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_mask : writeQueueVec_dataOut_1_data_mask;
  assign writeQueueVec_1_deq_bits_data_data = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_data : writeQueueVec_dataOut_1_data_data;
  assign writeQueueVec_1_deq_bits_data_last = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_last : writeQueueVec_dataOut_1_data_last;
  assign writeQueueVec_1_deq_bits_data_instructionIndex = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_instructionIndex : writeQueueVec_dataOut_1_data_instructionIndex;
  wire [31:0]       writeQueueVec_1_deq_bits_targetLane = _writeQueueVec_fifo_1_empty ? 32'h2 : writeQueueVec_dataOut_1_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_2 = writeQueueVec_2_enq_bits_data_vd;
  wire              vrfWritePort_2_valid_0 = writeQueueVec_2_deq_valid;
  wire [4:0]        vrfWritePort_2_bits_vd_0 = writeQueueVec_2_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_2_bits_mask_0 = writeQueueVec_2_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_2_bits_data_0 = writeQueueVec_2_deq_bits_data_data;
  wire              vrfWritePort_2_bits_last_0 = writeQueueVec_2_deq_bits_data_last;
  wire [2:0]        vrfWritePort_2_bits_instructionIndex_0 = writeQueueVec_2_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_2_enq_bits = writeQueueVec_2_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_2_enq_bits_data_data;
  wire              writeQueueVec_2_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_2 = {writeQueueVec_2_enq_bits_data_data, writeQueueVec_2_enq_bits_data_last};
  wire [2:0]        writeQueueVec_2_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_2 = {writeQueueVec_dataIn_lo_hi_2, writeQueueVec_2_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_2_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_2 = {writeQueueVec_dataIn_hi_hi_2, writeQueueVec_2_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_2 = {writeQueueVec_dataIn_hi_2, writeQueueVec_dataIn_lo_2, 32'h4};
  wire [31:0]       writeQueueVec_dataOut_2_targetLane = _writeQueueVec_fifo_2_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_2_data_instructionIndex = _writeQueueVec_fifo_2_data_out[34:32];
  wire              writeQueueVec_dataOut_2_data_last = _writeQueueVec_fifo_2_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_2_data_data = _writeQueueVec_fifo_2_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_2_data_mask = _writeQueueVec_fifo_2_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_2_data_vd = _writeQueueVec_fifo_2_data_out[76:72];
  wire              writeQueueVec_2_enq_ready = ~_writeQueueVec_fifo_2_full;
  wire              writeQueueVec_2_enq_valid;
  wire              _probeWire_slots_2_writeValid_T = writeQueueVec_2_enq_ready & writeQueueVec_2_enq_valid;
  assign writeQueueVec_2_deq_valid = ~_writeQueueVec_fifo_2_empty | writeQueueVec_2_enq_valid;
  assign writeQueueVec_2_deq_bits_data_vd = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_vd : writeQueueVec_dataOut_2_data_vd;
  assign writeQueueVec_2_deq_bits_data_mask = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_mask : writeQueueVec_dataOut_2_data_mask;
  assign writeQueueVec_2_deq_bits_data_data = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_data : writeQueueVec_dataOut_2_data_data;
  assign writeQueueVec_2_deq_bits_data_last = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_last : writeQueueVec_dataOut_2_data_last;
  assign writeQueueVec_2_deq_bits_data_instructionIndex = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_instructionIndex : writeQueueVec_dataOut_2_data_instructionIndex;
  wire [31:0]       writeQueueVec_2_deq_bits_targetLane = _writeQueueVec_fifo_2_empty ? 32'h4 : writeQueueVec_dataOut_2_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_3 = writeQueueVec_3_enq_bits_data_vd;
  wire              vrfWritePort_3_valid_0 = writeQueueVec_3_deq_valid;
  wire [4:0]        vrfWritePort_3_bits_vd_0 = writeQueueVec_3_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_3_bits_mask_0 = writeQueueVec_3_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_3_bits_data_0 = writeQueueVec_3_deq_bits_data_data;
  wire              vrfWritePort_3_bits_last_0 = writeQueueVec_3_deq_bits_data_last;
  wire [2:0]        vrfWritePort_3_bits_instructionIndex_0 = writeQueueVec_3_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_3_enq_bits = writeQueueVec_3_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_3_enq_bits_data_data;
  wire              writeQueueVec_3_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_3 = {writeQueueVec_3_enq_bits_data_data, writeQueueVec_3_enq_bits_data_last};
  wire [2:0]        writeQueueVec_3_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_3 = {writeQueueVec_dataIn_lo_hi_3, writeQueueVec_3_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_3_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_3 = {writeQueueVec_dataIn_hi_hi_3, writeQueueVec_3_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_3 = {writeQueueVec_dataIn_hi_3, writeQueueVec_dataIn_lo_3, 32'h8};
  wire [31:0]       writeQueueVec_dataOut_3_targetLane = _writeQueueVec_fifo_3_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_3_data_instructionIndex = _writeQueueVec_fifo_3_data_out[34:32];
  wire              writeQueueVec_dataOut_3_data_last = _writeQueueVec_fifo_3_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_3_data_data = _writeQueueVec_fifo_3_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_3_data_mask = _writeQueueVec_fifo_3_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_3_data_vd = _writeQueueVec_fifo_3_data_out[76:72];
  wire              writeQueueVec_3_enq_ready = ~_writeQueueVec_fifo_3_full;
  wire              writeQueueVec_3_enq_valid;
  wire              _probeWire_slots_3_writeValid_T = writeQueueVec_3_enq_ready & writeQueueVec_3_enq_valid;
  assign writeQueueVec_3_deq_valid = ~_writeQueueVec_fifo_3_empty | writeQueueVec_3_enq_valid;
  assign writeQueueVec_3_deq_bits_data_vd = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_vd : writeQueueVec_dataOut_3_data_vd;
  assign writeQueueVec_3_deq_bits_data_mask = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_mask : writeQueueVec_dataOut_3_data_mask;
  assign writeQueueVec_3_deq_bits_data_data = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_data : writeQueueVec_dataOut_3_data_data;
  assign writeQueueVec_3_deq_bits_data_last = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_last : writeQueueVec_dataOut_3_data_last;
  assign writeQueueVec_3_deq_bits_data_instructionIndex = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_instructionIndex : writeQueueVec_dataOut_3_data_instructionIndex;
  wire [31:0]       writeQueueVec_3_deq_bits_targetLane = _writeQueueVec_fifo_3_empty ? 32'h8 : writeQueueVec_dataOut_3_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_4 = writeQueueVec_4_enq_bits_data_vd;
  wire              vrfWritePort_4_valid_0 = writeQueueVec_4_deq_valid;
  wire [4:0]        vrfWritePort_4_bits_vd_0 = writeQueueVec_4_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_4_bits_mask_0 = writeQueueVec_4_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_4_bits_data_0 = writeQueueVec_4_deq_bits_data_data;
  wire              vrfWritePort_4_bits_last_0 = writeQueueVec_4_deq_bits_data_last;
  wire [2:0]        vrfWritePort_4_bits_instructionIndex_0 = writeQueueVec_4_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_4_enq_bits = writeQueueVec_4_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_4_enq_bits_data_data;
  wire              writeQueueVec_4_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_4 = {writeQueueVec_4_enq_bits_data_data, writeQueueVec_4_enq_bits_data_last};
  wire [2:0]        writeQueueVec_4_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_4 = {writeQueueVec_dataIn_lo_hi_4, writeQueueVec_4_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_4_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_4 = {writeQueueVec_dataIn_hi_hi_4, writeQueueVec_4_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_4 = {writeQueueVec_dataIn_hi_4, writeQueueVec_dataIn_lo_4, 32'h10};
  wire [31:0]       writeQueueVec_dataOut_4_targetLane = _writeQueueVec_fifo_4_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_4_data_instructionIndex = _writeQueueVec_fifo_4_data_out[34:32];
  wire              writeQueueVec_dataOut_4_data_last = _writeQueueVec_fifo_4_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_4_data_data = _writeQueueVec_fifo_4_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_4_data_mask = _writeQueueVec_fifo_4_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_4_data_vd = _writeQueueVec_fifo_4_data_out[76:72];
  wire              writeQueueVec_4_enq_ready = ~_writeQueueVec_fifo_4_full;
  wire              writeQueueVec_4_enq_valid;
  wire              _probeWire_slots_4_writeValid_T = writeQueueVec_4_enq_ready & writeQueueVec_4_enq_valid;
  assign writeQueueVec_4_deq_valid = ~_writeQueueVec_fifo_4_empty | writeQueueVec_4_enq_valid;
  assign writeQueueVec_4_deq_bits_data_vd = _writeQueueVec_fifo_4_empty ? writeQueueVec_4_enq_bits_data_vd : writeQueueVec_dataOut_4_data_vd;
  assign writeQueueVec_4_deq_bits_data_mask = _writeQueueVec_fifo_4_empty ? writeQueueVec_4_enq_bits_data_mask : writeQueueVec_dataOut_4_data_mask;
  assign writeQueueVec_4_deq_bits_data_data = _writeQueueVec_fifo_4_empty ? writeQueueVec_4_enq_bits_data_data : writeQueueVec_dataOut_4_data_data;
  assign writeQueueVec_4_deq_bits_data_last = _writeQueueVec_fifo_4_empty ? writeQueueVec_4_enq_bits_data_last : writeQueueVec_dataOut_4_data_last;
  assign writeQueueVec_4_deq_bits_data_instructionIndex = _writeQueueVec_fifo_4_empty ? writeQueueVec_4_enq_bits_data_instructionIndex : writeQueueVec_dataOut_4_data_instructionIndex;
  wire [31:0]       writeQueueVec_4_deq_bits_targetLane = _writeQueueVec_fifo_4_empty ? 32'h10 : writeQueueVec_dataOut_4_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_5 = writeQueueVec_5_enq_bits_data_vd;
  wire              vrfWritePort_5_valid_0 = writeQueueVec_5_deq_valid;
  wire [4:0]        vrfWritePort_5_bits_vd_0 = writeQueueVec_5_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_5_bits_mask_0 = writeQueueVec_5_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_5_bits_data_0 = writeQueueVec_5_deq_bits_data_data;
  wire              vrfWritePort_5_bits_last_0 = writeQueueVec_5_deq_bits_data_last;
  wire [2:0]        vrfWritePort_5_bits_instructionIndex_0 = writeQueueVec_5_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_5_enq_bits = writeQueueVec_5_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_5_enq_bits_data_data;
  wire              writeQueueVec_5_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_5 = {writeQueueVec_5_enq_bits_data_data, writeQueueVec_5_enq_bits_data_last};
  wire [2:0]        writeQueueVec_5_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_5 = {writeQueueVec_dataIn_lo_hi_5, writeQueueVec_5_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_5_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_5 = {writeQueueVec_dataIn_hi_hi_5, writeQueueVec_5_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_5 = {writeQueueVec_dataIn_hi_5, writeQueueVec_dataIn_lo_5, 32'h20};
  wire [31:0]       writeQueueVec_dataOut_5_targetLane = _writeQueueVec_fifo_5_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_5_data_instructionIndex = _writeQueueVec_fifo_5_data_out[34:32];
  wire              writeQueueVec_dataOut_5_data_last = _writeQueueVec_fifo_5_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_5_data_data = _writeQueueVec_fifo_5_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_5_data_mask = _writeQueueVec_fifo_5_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_5_data_vd = _writeQueueVec_fifo_5_data_out[76:72];
  wire              writeQueueVec_5_enq_ready = ~_writeQueueVec_fifo_5_full;
  wire              writeQueueVec_5_enq_valid;
  wire              _probeWire_slots_5_writeValid_T = writeQueueVec_5_enq_ready & writeQueueVec_5_enq_valid;
  assign writeQueueVec_5_deq_valid = ~_writeQueueVec_fifo_5_empty | writeQueueVec_5_enq_valid;
  assign writeQueueVec_5_deq_bits_data_vd = _writeQueueVec_fifo_5_empty ? writeQueueVec_5_enq_bits_data_vd : writeQueueVec_dataOut_5_data_vd;
  assign writeQueueVec_5_deq_bits_data_mask = _writeQueueVec_fifo_5_empty ? writeQueueVec_5_enq_bits_data_mask : writeQueueVec_dataOut_5_data_mask;
  assign writeQueueVec_5_deq_bits_data_data = _writeQueueVec_fifo_5_empty ? writeQueueVec_5_enq_bits_data_data : writeQueueVec_dataOut_5_data_data;
  assign writeQueueVec_5_deq_bits_data_last = _writeQueueVec_fifo_5_empty ? writeQueueVec_5_enq_bits_data_last : writeQueueVec_dataOut_5_data_last;
  assign writeQueueVec_5_deq_bits_data_instructionIndex = _writeQueueVec_fifo_5_empty ? writeQueueVec_5_enq_bits_data_instructionIndex : writeQueueVec_dataOut_5_data_instructionIndex;
  wire [31:0]       writeQueueVec_5_deq_bits_targetLane = _writeQueueVec_fifo_5_empty ? 32'h20 : writeQueueVec_dataOut_5_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_6 = writeQueueVec_6_enq_bits_data_vd;
  wire              vrfWritePort_6_valid_0 = writeQueueVec_6_deq_valid;
  wire [4:0]        vrfWritePort_6_bits_vd_0 = writeQueueVec_6_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_6_bits_mask_0 = writeQueueVec_6_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_6_bits_data_0 = writeQueueVec_6_deq_bits_data_data;
  wire              vrfWritePort_6_bits_last_0 = writeQueueVec_6_deq_bits_data_last;
  wire [2:0]        vrfWritePort_6_bits_instructionIndex_0 = writeQueueVec_6_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_6_enq_bits = writeQueueVec_6_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_6_enq_bits_data_data;
  wire              writeQueueVec_6_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_6 = {writeQueueVec_6_enq_bits_data_data, writeQueueVec_6_enq_bits_data_last};
  wire [2:0]        writeQueueVec_6_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_6 = {writeQueueVec_dataIn_lo_hi_6, writeQueueVec_6_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_6_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_6 = {writeQueueVec_dataIn_hi_hi_6, writeQueueVec_6_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_6 = {writeQueueVec_dataIn_hi_6, writeQueueVec_dataIn_lo_6, 32'h40};
  wire [31:0]       writeQueueVec_dataOut_6_targetLane = _writeQueueVec_fifo_6_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_6_data_instructionIndex = _writeQueueVec_fifo_6_data_out[34:32];
  wire              writeQueueVec_dataOut_6_data_last = _writeQueueVec_fifo_6_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_6_data_data = _writeQueueVec_fifo_6_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_6_data_mask = _writeQueueVec_fifo_6_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_6_data_vd = _writeQueueVec_fifo_6_data_out[76:72];
  wire              writeQueueVec_6_enq_ready = ~_writeQueueVec_fifo_6_full;
  wire              writeQueueVec_6_enq_valid;
  wire              _probeWire_slots_6_writeValid_T = writeQueueVec_6_enq_ready & writeQueueVec_6_enq_valid;
  assign writeQueueVec_6_deq_valid = ~_writeQueueVec_fifo_6_empty | writeQueueVec_6_enq_valid;
  assign writeQueueVec_6_deq_bits_data_vd = _writeQueueVec_fifo_6_empty ? writeQueueVec_6_enq_bits_data_vd : writeQueueVec_dataOut_6_data_vd;
  assign writeQueueVec_6_deq_bits_data_mask = _writeQueueVec_fifo_6_empty ? writeQueueVec_6_enq_bits_data_mask : writeQueueVec_dataOut_6_data_mask;
  assign writeQueueVec_6_deq_bits_data_data = _writeQueueVec_fifo_6_empty ? writeQueueVec_6_enq_bits_data_data : writeQueueVec_dataOut_6_data_data;
  assign writeQueueVec_6_deq_bits_data_last = _writeQueueVec_fifo_6_empty ? writeQueueVec_6_enq_bits_data_last : writeQueueVec_dataOut_6_data_last;
  assign writeQueueVec_6_deq_bits_data_instructionIndex = _writeQueueVec_fifo_6_empty ? writeQueueVec_6_enq_bits_data_instructionIndex : writeQueueVec_dataOut_6_data_instructionIndex;
  wire [31:0]       writeQueueVec_6_deq_bits_targetLane = _writeQueueVec_fifo_6_empty ? 32'h40 : writeQueueVec_dataOut_6_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_7 = writeQueueVec_7_enq_bits_data_vd;
  wire              vrfWritePort_7_valid_0 = writeQueueVec_7_deq_valid;
  wire [4:0]        vrfWritePort_7_bits_vd_0 = writeQueueVec_7_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_7_bits_mask_0 = writeQueueVec_7_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_7_bits_data_0 = writeQueueVec_7_deq_bits_data_data;
  wire              vrfWritePort_7_bits_last_0 = writeQueueVec_7_deq_bits_data_last;
  wire [2:0]        vrfWritePort_7_bits_instructionIndex_0 = writeQueueVec_7_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_7_enq_bits = writeQueueVec_7_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_7_enq_bits_data_data;
  wire              writeQueueVec_7_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_7 = {writeQueueVec_7_enq_bits_data_data, writeQueueVec_7_enq_bits_data_last};
  wire [2:0]        writeQueueVec_7_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_7 = {writeQueueVec_dataIn_lo_hi_7, writeQueueVec_7_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_7_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_7 = {writeQueueVec_dataIn_hi_hi_7, writeQueueVec_7_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_7 = {writeQueueVec_dataIn_hi_7, writeQueueVec_dataIn_lo_7, 32'h80};
  wire [31:0]       writeQueueVec_dataOut_7_targetLane = _writeQueueVec_fifo_7_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_7_data_instructionIndex = _writeQueueVec_fifo_7_data_out[34:32];
  wire              writeQueueVec_dataOut_7_data_last = _writeQueueVec_fifo_7_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_7_data_data = _writeQueueVec_fifo_7_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_7_data_mask = _writeQueueVec_fifo_7_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_7_data_vd = _writeQueueVec_fifo_7_data_out[76:72];
  wire              writeQueueVec_7_enq_ready = ~_writeQueueVec_fifo_7_full;
  wire              writeQueueVec_7_enq_valid;
  wire              _probeWire_slots_7_writeValid_T = writeQueueVec_7_enq_ready & writeQueueVec_7_enq_valid;
  assign writeQueueVec_7_deq_valid = ~_writeQueueVec_fifo_7_empty | writeQueueVec_7_enq_valid;
  assign writeQueueVec_7_deq_bits_data_vd = _writeQueueVec_fifo_7_empty ? writeQueueVec_7_enq_bits_data_vd : writeQueueVec_dataOut_7_data_vd;
  assign writeQueueVec_7_deq_bits_data_mask = _writeQueueVec_fifo_7_empty ? writeQueueVec_7_enq_bits_data_mask : writeQueueVec_dataOut_7_data_mask;
  assign writeQueueVec_7_deq_bits_data_data = _writeQueueVec_fifo_7_empty ? writeQueueVec_7_enq_bits_data_data : writeQueueVec_dataOut_7_data_data;
  assign writeQueueVec_7_deq_bits_data_last = _writeQueueVec_fifo_7_empty ? writeQueueVec_7_enq_bits_data_last : writeQueueVec_dataOut_7_data_last;
  assign writeQueueVec_7_deq_bits_data_instructionIndex = _writeQueueVec_fifo_7_empty ? writeQueueVec_7_enq_bits_data_instructionIndex : writeQueueVec_dataOut_7_data_instructionIndex;
  wire [31:0]       writeQueueVec_7_deq_bits_targetLane = _writeQueueVec_fifo_7_empty ? 32'h80 : writeQueueVec_dataOut_7_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_8 = writeQueueVec_8_enq_bits_data_vd;
  wire              vrfWritePort_8_valid_0 = writeQueueVec_8_deq_valid;
  wire [4:0]        vrfWritePort_8_bits_vd_0 = writeQueueVec_8_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_8_bits_mask_0 = writeQueueVec_8_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_8_bits_data_0 = writeQueueVec_8_deq_bits_data_data;
  wire              vrfWritePort_8_bits_last_0 = writeQueueVec_8_deq_bits_data_last;
  wire [2:0]        vrfWritePort_8_bits_instructionIndex_0 = writeQueueVec_8_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_8_enq_bits = writeQueueVec_8_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_8_enq_bits_data_data;
  wire              writeQueueVec_8_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_8 = {writeQueueVec_8_enq_bits_data_data, writeQueueVec_8_enq_bits_data_last};
  wire [2:0]        writeQueueVec_8_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_8 = {writeQueueVec_dataIn_lo_hi_8, writeQueueVec_8_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_8_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_8 = {writeQueueVec_dataIn_hi_hi_8, writeQueueVec_8_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_8 = {writeQueueVec_dataIn_hi_8, writeQueueVec_dataIn_lo_8, 32'h100};
  wire [31:0]       writeQueueVec_dataOut_8_targetLane = _writeQueueVec_fifo_8_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_8_data_instructionIndex = _writeQueueVec_fifo_8_data_out[34:32];
  wire              writeQueueVec_dataOut_8_data_last = _writeQueueVec_fifo_8_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_8_data_data = _writeQueueVec_fifo_8_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_8_data_mask = _writeQueueVec_fifo_8_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_8_data_vd = _writeQueueVec_fifo_8_data_out[76:72];
  wire              writeQueueVec_8_enq_ready = ~_writeQueueVec_fifo_8_full;
  wire              writeQueueVec_8_enq_valid;
  wire              _probeWire_slots_8_writeValid_T = writeQueueVec_8_enq_ready & writeQueueVec_8_enq_valid;
  assign writeQueueVec_8_deq_valid = ~_writeQueueVec_fifo_8_empty | writeQueueVec_8_enq_valid;
  assign writeQueueVec_8_deq_bits_data_vd = _writeQueueVec_fifo_8_empty ? writeQueueVec_8_enq_bits_data_vd : writeQueueVec_dataOut_8_data_vd;
  assign writeQueueVec_8_deq_bits_data_mask = _writeQueueVec_fifo_8_empty ? writeQueueVec_8_enq_bits_data_mask : writeQueueVec_dataOut_8_data_mask;
  assign writeQueueVec_8_deq_bits_data_data = _writeQueueVec_fifo_8_empty ? writeQueueVec_8_enq_bits_data_data : writeQueueVec_dataOut_8_data_data;
  assign writeQueueVec_8_deq_bits_data_last = _writeQueueVec_fifo_8_empty ? writeQueueVec_8_enq_bits_data_last : writeQueueVec_dataOut_8_data_last;
  assign writeQueueVec_8_deq_bits_data_instructionIndex = _writeQueueVec_fifo_8_empty ? writeQueueVec_8_enq_bits_data_instructionIndex : writeQueueVec_dataOut_8_data_instructionIndex;
  wire [31:0]       writeQueueVec_8_deq_bits_targetLane = _writeQueueVec_fifo_8_empty ? 32'h100 : writeQueueVec_dataOut_8_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_9 = writeQueueVec_9_enq_bits_data_vd;
  wire              vrfWritePort_9_valid_0 = writeQueueVec_9_deq_valid;
  wire [4:0]        vrfWritePort_9_bits_vd_0 = writeQueueVec_9_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_9_bits_mask_0 = writeQueueVec_9_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_9_bits_data_0 = writeQueueVec_9_deq_bits_data_data;
  wire              vrfWritePort_9_bits_last_0 = writeQueueVec_9_deq_bits_data_last;
  wire [2:0]        vrfWritePort_9_bits_instructionIndex_0 = writeQueueVec_9_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_9_enq_bits = writeQueueVec_9_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_9_enq_bits_data_data;
  wire              writeQueueVec_9_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_9 = {writeQueueVec_9_enq_bits_data_data, writeQueueVec_9_enq_bits_data_last};
  wire [2:0]        writeQueueVec_9_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_9 = {writeQueueVec_dataIn_lo_hi_9, writeQueueVec_9_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_9_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_9 = {writeQueueVec_dataIn_hi_hi_9, writeQueueVec_9_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_9 = {writeQueueVec_dataIn_hi_9, writeQueueVec_dataIn_lo_9, 32'h200};
  wire [31:0]       writeQueueVec_dataOut_9_targetLane = _writeQueueVec_fifo_9_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_9_data_instructionIndex = _writeQueueVec_fifo_9_data_out[34:32];
  wire              writeQueueVec_dataOut_9_data_last = _writeQueueVec_fifo_9_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_9_data_data = _writeQueueVec_fifo_9_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_9_data_mask = _writeQueueVec_fifo_9_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_9_data_vd = _writeQueueVec_fifo_9_data_out[76:72];
  wire              writeQueueVec_9_enq_ready = ~_writeQueueVec_fifo_9_full;
  wire              writeQueueVec_9_enq_valid;
  wire              _probeWire_slots_9_writeValid_T = writeQueueVec_9_enq_ready & writeQueueVec_9_enq_valid;
  assign writeQueueVec_9_deq_valid = ~_writeQueueVec_fifo_9_empty | writeQueueVec_9_enq_valid;
  assign writeQueueVec_9_deq_bits_data_vd = _writeQueueVec_fifo_9_empty ? writeQueueVec_9_enq_bits_data_vd : writeQueueVec_dataOut_9_data_vd;
  assign writeQueueVec_9_deq_bits_data_mask = _writeQueueVec_fifo_9_empty ? writeQueueVec_9_enq_bits_data_mask : writeQueueVec_dataOut_9_data_mask;
  assign writeQueueVec_9_deq_bits_data_data = _writeQueueVec_fifo_9_empty ? writeQueueVec_9_enq_bits_data_data : writeQueueVec_dataOut_9_data_data;
  assign writeQueueVec_9_deq_bits_data_last = _writeQueueVec_fifo_9_empty ? writeQueueVec_9_enq_bits_data_last : writeQueueVec_dataOut_9_data_last;
  assign writeQueueVec_9_deq_bits_data_instructionIndex = _writeQueueVec_fifo_9_empty ? writeQueueVec_9_enq_bits_data_instructionIndex : writeQueueVec_dataOut_9_data_instructionIndex;
  wire [31:0]       writeQueueVec_9_deq_bits_targetLane = _writeQueueVec_fifo_9_empty ? 32'h200 : writeQueueVec_dataOut_9_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_10 = writeQueueVec_10_enq_bits_data_vd;
  wire              vrfWritePort_10_valid_0 = writeQueueVec_10_deq_valid;
  wire [4:0]        vrfWritePort_10_bits_vd_0 = writeQueueVec_10_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_10_bits_mask_0 = writeQueueVec_10_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_10_bits_data_0 = writeQueueVec_10_deq_bits_data_data;
  wire              vrfWritePort_10_bits_last_0 = writeQueueVec_10_deq_bits_data_last;
  wire [2:0]        vrfWritePort_10_bits_instructionIndex_0 = writeQueueVec_10_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_10_enq_bits = writeQueueVec_10_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_10_enq_bits_data_data;
  wire              writeQueueVec_10_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_10 = {writeQueueVec_10_enq_bits_data_data, writeQueueVec_10_enq_bits_data_last};
  wire [2:0]        writeQueueVec_10_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_10 = {writeQueueVec_dataIn_lo_hi_10, writeQueueVec_10_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_10_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_10 = {writeQueueVec_dataIn_hi_hi_10, writeQueueVec_10_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_10 = {writeQueueVec_dataIn_hi_10, writeQueueVec_dataIn_lo_10, 32'h400};
  wire [31:0]       writeQueueVec_dataOut_10_targetLane = _writeQueueVec_fifo_10_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_10_data_instructionIndex = _writeQueueVec_fifo_10_data_out[34:32];
  wire              writeQueueVec_dataOut_10_data_last = _writeQueueVec_fifo_10_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_10_data_data = _writeQueueVec_fifo_10_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_10_data_mask = _writeQueueVec_fifo_10_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_10_data_vd = _writeQueueVec_fifo_10_data_out[76:72];
  wire              writeQueueVec_10_enq_ready = ~_writeQueueVec_fifo_10_full;
  wire              writeQueueVec_10_enq_valid;
  wire              _probeWire_slots_10_writeValid_T = writeQueueVec_10_enq_ready & writeQueueVec_10_enq_valid;
  assign writeQueueVec_10_deq_valid = ~_writeQueueVec_fifo_10_empty | writeQueueVec_10_enq_valid;
  assign writeQueueVec_10_deq_bits_data_vd = _writeQueueVec_fifo_10_empty ? writeQueueVec_10_enq_bits_data_vd : writeQueueVec_dataOut_10_data_vd;
  assign writeQueueVec_10_deq_bits_data_mask = _writeQueueVec_fifo_10_empty ? writeQueueVec_10_enq_bits_data_mask : writeQueueVec_dataOut_10_data_mask;
  assign writeQueueVec_10_deq_bits_data_data = _writeQueueVec_fifo_10_empty ? writeQueueVec_10_enq_bits_data_data : writeQueueVec_dataOut_10_data_data;
  assign writeQueueVec_10_deq_bits_data_last = _writeQueueVec_fifo_10_empty ? writeQueueVec_10_enq_bits_data_last : writeQueueVec_dataOut_10_data_last;
  assign writeQueueVec_10_deq_bits_data_instructionIndex = _writeQueueVec_fifo_10_empty ? writeQueueVec_10_enq_bits_data_instructionIndex : writeQueueVec_dataOut_10_data_instructionIndex;
  wire [31:0]       writeQueueVec_10_deq_bits_targetLane = _writeQueueVec_fifo_10_empty ? 32'h400 : writeQueueVec_dataOut_10_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_11 = writeQueueVec_11_enq_bits_data_vd;
  wire              vrfWritePort_11_valid_0 = writeQueueVec_11_deq_valid;
  wire [4:0]        vrfWritePort_11_bits_vd_0 = writeQueueVec_11_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_11_bits_mask_0 = writeQueueVec_11_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_11_bits_data_0 = writeQueueVec_11_deq_bits_data_data;
  wire              vrfWritePort_11_bits_last_0 = writeQueueVec_11_deq_bits_data_last;
  wire [2:0]        vrfWritePort_11_bits_instructionIndex_0 = writeQueueVec_11_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_11_enq_bits = writeQueueVec_11_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_11_enq_bits_data_data;
  wire              writeQueueVec_11_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_11 = {writeQueueVec_11_enq_bits_data_data, writeQueueVec_11_enq_bits_data_last};
  wire [2:0]        writeQueueVec_11_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_11 = {writeQueueVec_dataIn_lo_hi_11, writeQueueVec_11_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_11_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_11 = {writeQueueVec_dataIn_hi_hi_11, writeQueueVec_11_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_11 = {writeQueueVec_dataIn_hi_11, writeQueueVec_dataIn_lo_11, 32'h800};
  wire [31:0]       writeQueueVec_dataOut_11_targetLane = _writeQueueVec_fifo_11_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_11_data_instructionIndex = _writeQueueVec_fifo_11_data_out[34:32];
  wire              writeQueueVec_dataOut_11_data_last = _writeQueueVec_fifo_11_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_11_data_data = _writeQueueVec_fifo_11_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_11_data_mask = _writeQueueVec_fifo_11_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_11_data_vd = _writeQueueVec_fifo_11_data_out[76:72];
  wire              writeQueueVec_11_enq_ready = ~_writeQueueVec_fifo_11_full;
  wire              writeQueueVec_11_enq_valid;
  wire              _probeWire_slots_11_writeValid_T = writeQueueVec_11_enq_ready & writeQueueVec_11_enq_valid;
  assign writeQueueVec_11_deq_valid = ~_writeQueueVec_fifo_11_empty | writeQueueVec_11_enq_valid;
  assign writeQueueVec_11_deq_bits_data_vd = _writeQueueVec_fifo_11_empty ? writeQueueVec_11_enq_bits_data_vd : writeQueueVec_dataOut_11_data_vd;
  assign writeQueueVec_11_deq_bits_data_mask = _writeQueueVec_fifo_11_empty ? writeQueueVec_11_enq_bits_data_mask : writeQueueVec_dataOut_11_data_mask;
  assign writeQueueVec_11_deq_bits_data_data = _writeQueueVec_fifo_11_empty ? writeQueueVec_11_enq_bits_data_data : writeQueueVec_dataOut_11_data_data;
  assign writeQueueVec_11_deq_bits_data_last = _writeQueueVec_fifo_11_empty ? writeQueueVec_11_enq_bits_data_last : writeQueueVec_dataOut_11_data_last;
  assign writeQueueVec_11_deq_bits_data_instructionIndex = _writeQueueVec_fifo_11_empty ? writeQueueVec_11_enq_bits_data_instructionIndex : writeQueueVec_dataOut_11_data_instructionIndex;
  wire [31:0]       writeQueueVec_11_deq_bits_targetLane = _writeQueueVec_fifo_11_empty ? 32'h800 : writeQueueVec_dataOut_11_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_12 = writeQueueVec_12_enq_bits_data_vd;
  wire              vrfWritePort_12_valid_0 = writeQueueVec_12_deq_valid;
  wire [4:0]        vrfWritePort_12_bits_vd_0 = writeQueueVec_12_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_12_bits_mask_0 = writeQueueVec_12_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_12_bits_data_0 = writeQueueVec_12_deq_bits_data_data;
  wire              vrfWritePort_12_bits_last_0 = writeQueueVec_12_deq_bits_data_last;
  wire [2:0]        vrfWritePort_12_bits_instructionIndex_0 = writeQueueVec_12_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_12_enq_bits = writeQueueVec_12_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_12_enq_bits_data_data;
  wire              writeQueueVec_12_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_12 = {writeQueueVec_12_enq_bits_data_data, writeQueueVec_12_enq_bits_data_last};
  wire [2:0]        writeQueueVec_12_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_12 = {writeQueueVec_dataIn_lo_hi_12, writeQueueVec_12_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_12_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_12 = {writeQueueVec_dataIn_hi_hi_12, writeQueueVec_12_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_12 = {writeQueueVec_dataIn_hi_12, writeQueueVec_dataIn_lo_12, 32'h1000};
  wire [31:0]       writeQueueVec_dataOut_12_targetLane = _writeQueueVec_fifo_12_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_12_data_instructionIndex = _writeQueueVec_fifo_12_data_out[34:32];
  wire              writeQueueVec_dataOut_12_data_last = _writeQueueVec_fifo_12_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_12_data_data = _writeQueueVec_fifo_12_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_12_data_mask = _writeQueueVec_fifo_12_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_12_data_vd = _writeQueueVec_fifo_12_data_out[76:72];
  wire              writeQueueVec_12_enq_ready = ~_writeQueueVec_fifo_12_full;
  wire              writeQueueVec_12_enq_valid;
  wire              _probeWire_slots_12_writeValid_T = writeQueueVec_12_enq_ready & writeQueueVec_12_enq_valid;
  assign writeQueueVec_12_deq_valid = ~_writeQueueVec_fifo_12_empty | writeQueueVec_12_enq_valid;
  assign writeQueueVec_12_deq_bits_data_vd = _writeQueueVec_fifo_12_empty ? writeQueueVec_12_enq_bits_data_vd : writeQueueVec_dataOut_12_data_vd;
  assign writeQueueVec_12_deq_bits_data_mask = _writeQueueVec_fifo_12_empty ? writeQueueVec_12_enq_bits_data_mask : writeQueueVec_dataOut_12_data_mask;
  assign writeQueueVec_12_deq_bits_data_data = _writeQueueVec_fifo_12_empty ? writeQueueVec_12_enq_bits_data_data : writeQueueVec_dataOut_12_data_data;
  assign writeQueueVec_12_deq_bits_data_last = _writeQueueVec_fifo_12_empty ? writeQueueVec_12_enq_bits_data_last : writeQueueVec_dataOut_12_data_last;
  assign writeQueueVec_12_deq_bits_data_instructionIndex = _writeQueueVec_fifo_12_empty ? writeQueueVec_12_enq_bits_data_instructionIndex : writeQueueVec_dataOut_12_data_instructionIndex;
  wire [31:0]       writeQueueVec_12_deq_bits_targetLane = _writeQueueVec_fifo_12_empty ? 32'h1000 : writeQueueVec_dataOut_12_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_13 = writeQueueVec_13_enq_bits_data_vd;
  wire              vrfWritePort_13_valid_0 = writeQueueVec_13_deq_valid;
  wire [4:0]        vrfWritePort_13_bits_vd_0 = writeQueueVec_13_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_13_bits_mask_0 = writeQueueVec_13_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_13_bits_data_0 = writeQueueVec_13_deq_bits_data_data;
  wire              vrfWritePort_13_bits_last_0 = writeQueueVec_13_deq_bits_data_last;
  wire [2:0]        vrfWritePort_13_bits_instructionIndex_0 = writeQueueVec_13_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_13_enq_bits = writeQueueVec_13_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_13_enq_bits_data_data;
  wire              writeQueueVec_13_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_13 = {writeQueueVec_13_enq_bits_data_data, writeQueueVec_13_enq_bits_data_last};
  wire [2:0]        writeQueueVec_13_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_13 = {writeQueueVec_dataIn_lo_hi_13, writeQueueVec_13_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_13_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_13 = {writeQueueVec_dataIn_hi_hi_13, writeQueueVec_13_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_13 = {writeQueueVec_dataIn_hi_13, writeQueueVec_dataIn_lo_13, 32'h2000};
  wire [31:0]       writeQueueVec_dataOut_13_targetLane = _writeQueueVec_fifo_13_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_13_data_instructionIndex = _writeQueueVec_fifo_13_data_out[34:32];
  wire              writeQueueVec_dataOut_13_data_last = _writeQueueVec_fifo_13_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_13_data_data = _writeQueueVec_fifo_13_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_13_data_mask = _writeQueueVec_fifo_13_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_13_data_vd = _writeQueueVec_fifo_13_data_out[76:72];
  wire              writeQueueVec_13_enq_ready = ~_writeQueueVec_fifo_13_full;
  wire              writeQueueVec_13_enq_valid;
  wire              _probeWire_slots_13_writeValid_T = writeQueueVec_13_enq_ready & writeQueueVec_13_enq_valid;
  assign writeQueueVec_13_deq_valid = ~_writeQueueVec_fifo_13_empty | writeQueueVec_13_enq_valid;
  assign writeQueueVec_13_deq_bits_data_vd = _writeQueueVec_fifo_13_empty ? writeQueueVec_13_enq_bits_data_vd : writeQueueVec_dataOut_13_data_vd;
  assign writeQueueVec_13_deq_bits_data_mask = _writeQueueVec_fifo_13_empty ? writeQueueVec_13_enq_bits_data_mask : writeQueueVec_dataOut_13_data_mask;
  assign writeQueueVec_13_deq_bits_data_data = _writeQueueVec_fifo_13_empty ? writeQueueVec_13_enq_bits_data_data : writeQueueVec_dataOut_13_data_data;
  assign writeQueueVec_13_deq_bits_data_last = _writeQueueVec_fifo_13_empty ? writeQueueVec_13_enq_bits_data_last : writeQueueVec_dataOut_13_data_last;
  assign writeQueueVec_13_deq_bits_data_instructionIndex = _writeQueueVec_fifo_13_empty ? writeQueueVec_13_enq_bits_data_instructionIndex : writeQueueVec_dataOut_13_data_instructionIndex;
  wire [31:0]       writeQueueVec_13_deq_bits_targetLane = _writeQueueVec_fifo_13_empty ? 32'h2000 : writeQueueVec_dataOut_13_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_14 = writeQueueVec_14_enq_bits_data_vd;
  wire              vrfWritePort_14_valid_0 = writeQueueVec_14_deq_valid;
  wire [4:0]        vrfWritePort_14_bits_vd_0 = writeQueueVec_14_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_14_bits_mask_0 = writeQueueVec_14_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_14_bits_data_0 = writeQueueVec_14_deq_bits_data_data;
  wire              vrfWritePort_14_bits_last_0 = writeQueueVec_14_deq_bits_data_last;
  wire [2:0]        vrfWritePort_14_bits_instructionIndex_0 = writeQueueVec_14_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_14_enq_bits = writeQueueVec_14_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_14_enq_bits_data_data;
  wire              writeQueueVec_14_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_14 = {writeQueueVec_14_enq_bits_data_data, writeQueueVec_14_enq_bits_data_last};
  wire [2:0]        writeQueueVec_14_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_14 = {writeQueueVec_dataIn_lo_hi_14, writeQueueVec_14_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_14_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_14 = {writeQueueVec_dataIn_hi_hi_14, writeQueueVec_14_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_14 = {writeQueueVec_dataIn_hi_14, writeQueueVec_dataIn_lo_14, 32'h4000};
  wire [31:0]       writeQueueVec_dataOut_14_targetLane = _writeQueueVec_fifo_14_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_14_data_instructionIndex = _writeQueueVec_fifo_14_data_out[34:32];
  wire              writeQueueVec_dataOut_14_data_last = _writeQueueVec_fifo_14_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_14_data_data = _writeQueueVec_fifo_14_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_14_data_mask = _writeQueueVec_fifo_14_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_14_data_vd = _writeQueueVec_fifo_14_data_out[76:72];
  wire              writeQueueVec_14_enq_ready = ~_writeQueueVec_fifo_14_full;
  wire              writeQueueVec_14_enq_valid;
  wire              _probeWire_slots_14_writeValid_T = writeQueueVec_14_enq_ready & writeQueueVec_14_enq_valid;
  assign writeQueueVec_14_deq_valid = ~_writeQueueVec_fifo_14_empty | writeQueueVec_14_enq_valid;
  assign writeQueueVec_14_deq_bits_data_vd = _writeQueueVec_fifo_14_empty ? writeQueueVec_14_enq_bits_data_vd : writeQueueVec_dataOut_14_data_vd;
  assign writeQueueVec_14_deq_bits_data_mask = _writeQueueVec_fifo_14_empty ? writeQueueVec_14_enq_bits_data_mask : writeQueueVec_dataOut_14_data_mask;
  assign writeQueueVec_14_deq_bits_data_data = _writeQueueVec_fifo_14_empty ? writeQueueVec_14_enq_bits_data_data : writeQueueVec_dataOut_14_data_data;
  assign writeQueueVec_14_deq_bits_data_last = _writeQueueVec_fifo_14_empty ? writeQueueVec_14_enq_bits_data_last : writeQueueVec_dataOut_14_data_last;
  assign writeQueueVec_14_deq_bits_data_instructionIndex = _writeQueueVec_fifo_14_empty ? writeQueueVec_14_enq_bits_data_instructionIndex : writeQueueVec_dataOut_14_data_instructionIndex;
  wire [31:0]       writeQueueVec_14_deq_bits_targetLane = _writeQueueVec_fifo_14_empty ? 32'h4000 : writeQueueVec_dataOut_14_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_15 = writeQueueVec_15_enq_bits_data_vd;
  wire              vrfWritePort_15_valid_0 = writeQueueVec_15_deq_valid;
  wire [4:0]        vrfWritePort_15_bits_vd_0 = writeQueueVec_15_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_15_bits_mask_0 = writeQueueVec_15_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_15_bits_data_0 = writeQueueVec_15_deq_bits_data_data;
  wire              vrfWritePort_15_bits_last_0 = writeQueueVec_15_deq_bits_data_last;
  wire [2:0]        vrfWritePort_15_bits_instructionIndex_0 = writeQueueVec_15_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_15_enq_bits = writeQueueVec_15_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_15_enq_bits_data_data;
  wire              writeQueueVec_15_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_15 = {writeQueueVec_15_enq_bits_data_data, writeQueueVec_15_enq_bits_data_last};
  wire [2:0]        writeQueueVec_15_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_15 = {writeQueueVec_dataIn_lo_hi_15, writeQueueVec_15_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_15_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_15 = {writeQueueVec_dataIn_hi_hi_15, writeQueueVec_15_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_15 = {writeQueueVec_dataIn_hi_15, writeQueueVec_dataIn_lo_15, 32'h8000};
  wire [31:0]       writeQueueVec_dataOut_15_targetLane = _writeQueueVec_fifo_15_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_15_data_instructionIndex = _writeQueueVec_fifo_15_data_out[34:32];
  wire              writeQueueVec_dataOut_15_data_last = _writeQueueVec_fifo_15_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_15_data_data = _writeQueueVec_fifo_15_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_15_data_mask = _writeQueueVec_fifo_15_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_15_data_vd = _writeQueueVec_fifo_15_data_out[76:72];
  wire              writeQueueVec_15_enq_ready = ~_writeQueueVec_fifo_15_full;
  wire              writeQueueVec_15_enq_valid;
  wire              _probeWire_slots_15_writeValid_T = writeQueueVec_15_enq_ready & writeQueueVec_15_enq_valid;
  assign writeQueueVec_15_deq_valid = ~_writeQueueVec_fifo_15_empty | writeQueueVec_15_enq_valid;
  assign writeQueueVec_15_deq_bits_data_vd = _writeQueueVec_fifo_15_empty ? writeQueueVec_15_enq_bits_data_vd : writeQueueVec_dataOut_15_data_vd;
  assign writeQueueVec_15_deq_bits_data_mask = _writeQueueVec_fifo_15_empty ? writeQueueVec_15_enq_bits_data_mask : writeQueueVec_dataOut_15_data_mask;
  assign writeQueueVec_15_deq_bits_data_data = _writeQueueVec_fifo_15_empty ? writeQueueVec_15_enq_bits_data_data : writeQueueVec_dataOut_15_data_data;
  assign writeQueueVec_15_deq_bits_data_last = _writeQueueVec_fifo_15_empty ? writeQueueVec_15_enq_bits_data_last : writeQueueVec_dataOut_15_data_last;
  assign writeQueueVec_15_deq_bits_data_instructionIndex = _writeQueueVec_fifo_15_empty ? writeQueueVec_15_enq_bits_data_instructionIndex : writeQueueVec_dataOut_15_data_instructionIndex;
  wire [31:0]       writeQueueVec_15_deq_bits_targetLane = _writeQueueVec_fifo_15_empty ? 32'h8000 : writeQueueVec_dataOut_15_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_16 = writeQueueVec_16_enq_bits_data_vd;
  wire              vrfWritePort_16_valid_0 = writeQueueVec_16_deq_valid;
  wire [4:0]        vrfWritePort_16_bits_vd_0 = writeQueueVec_16_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_16_bits_mask_0 = writeQueueVec_16_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_16_bits_data_0 = writeQueueVec_16_deq_bits_data_data;
  wire              vrfWritePort_16_bits_last_0 = writeQueueVec_16_deq_bits_data_last;
  wire [2:0]        vrfWritePort_16_bits_instructionIndex_0 = writeQueueVec_16_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_16_enq_bits = writeQueueVec_16_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_16_enq_bits_data_data;
  wire              writeQueueVec_16_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_16 = {writeQueueVec_16_enq_bits_data_data, writeQueueVec_16_enq_bits_data_last};
  wire [2:0]        writeQueueVec_16_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_16 = {writeQueueVec_dataIn_lo_hi_16, writeQueueVec_16_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_16_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_16 = {writeQueueVec_dataIn_hi_hi_16, writeQueueVec_16_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_16 = {writeQueueVec_dataIn_hi_16, writeQueueVec_dataIn_lo_16, 32'h10000};
  wire [31:0]       writeQueueVec_dataOut_16_targetLane = _writeQueueVec_fifo_16_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_16_data_instructionIndex = _writeQueueVec_fifo_16_data_out[34:32];
  wire              writeQueueVec_dataOut_16_data_last = _writeQueueVec_fifo_16_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_16_data_data = _writeQueueVec_fifo_16_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_16_data_mask = _writeQueueVec_fifo_16_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_16_data_vd = _writeQueueVec_fifo_16_data_out[76:72];
  wire              writeQueueVec_16_enq_ready = ~_writeQueueVec_fifo_16_full;
  wire              writeQueueVec_16_enq_valid;
  wire              _probeWire_slots_16_writeValid_T = writeQueueVec_16_enq_ready & writeQueueVec_16_enq_valid;
  assign writeQueueVec_16_deq_valid = ~_writeQueueVec_fifo_16_empty | writeQueueVec_16_enq_valid;
  assign writeQueueVec_16_deq_bits_data_vd = _writeQueueVec_fifo_16_empty ? writeQueueVec_16_enq_bits_data_vd : writeQueueVec_dataOut_16_data_vd;
  assign writeQueueVec_16_deq_bits_data_mask = _writeQueueVec_fifo_16_empty ? writeQueueVec_16_enq_bits_data_mask : writeQueueVec_dataOut_16_data_mask;
  assign writeQueueVec_16_deq_bits_data_data = _writeQueueVec_fifo_16_empty ? writeQueueVec_16_enq_bits_data_data : writeQueueVec_dataOut_16_data_data;
  assign writeQueueVec_16_deq_bits_data_last = _writeQueueVec_fifo_16_empty ? writeQueueVec_16_enq_bits_data_last : writeQueueVec_dataOut_16_data_last;
  assign writeQueueVec_16_deq_bits_data_instructionIndex = _writeQueueVec_fifo_16_empty ? writeQueueVec_16_enq_bits_data_instructionIndex : writeQueueVec_dataOut_16_data_instructionIndex;
  wire [31:0]       writeQueueVec_16_deq_bits_targetLane = _writeQueueVec_fifo_16_empty ? 32'h10000 : writeQueueVec_dataOut_16_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_17 = writeQueueVec_17_enq_bits_data_vd;
  wire              vrfWritePort_17_valid_0 = writeQueueVec_17_deq_valid;
  wire [4:0]        vrfWritePort_17_bits_vd_0 = writeQueueVec_17_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_17_bits_mask_0 = writeQueueVec_17_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_17_bits_data_0 = writeQueueVec_17_deq_bits_data_data;
  wire              vrfWritePort_17_bits_last_0 = writeQueueVec_17_deq_bits_data_last;
  wire [2:0]        vrfWritePort_17_bits_instructionIndex_0 = writeQueueVec_17_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_17_enq_bits = writeQueueVec_17_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_17_enq_bits_data_data;
  wire              writeQueueVec_17_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_17 = {writeQueueVec_17_enq_bits_data_data, writeQueueVec_17_enq_bits_data_last};
  wire [2:0]        writeQueueVec_17_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_17 = {writeQueueVec_dataIn_lo_hi_17, writeQueueVec_17_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_17_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_17 = {writeQueueVec_dataIn_hi_hi_17, writeQueueVec_17_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_17 = {writeQueueVec_dataIn_hi_17, writeQueueVec_dataIn_lo_17, 32'h20000};
  wire [31:0]       writeQueueVec_dataOut_17_targetLane = _writeQueueVec_fifo_17_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_17_data_instructionIndex = _writeQueueVec_fifo_17_data_out[34:32];
  wire              writeQueueVec_dataOut_17_data_last = _writeQueueVec_fifo_17_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_17_data_data = _writeQueueVec_fifo_17_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_17_data_mask = _writeQueueVec_fifo_17_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_17_data_vd = _writeQueueVec_fifo_17_data_out[76:72];
  wire              writeQueueVec_17_enq_ready = ~_writeQueueVec_fifo_17_full;
  wire              writeQueueVec_17_enq_valid;
  wire              _probeWire_slots_17_writeValid_T = writeQueueVec_17_enq_ready & writeQueueVec_17_enq_valid;
  assign writeQueueVec_17_deq_valid = ~_writeQueueVec_fifo_17_empty | writeQueueVec_17_enq_valid;
  assign writeQueueVec_17_deq_bits_data_vd = _writeQueueVec_fifo_17_empty ? writeQueueVec_17_enq_bits_data_vd : writeQueueVec_dataOut_17_data_vd;
  assign writeQueueVec_17_deq_bits_data_mask = _writeQueueVec_fifo_17_empty ? writeQueueVec_17_enq_bits_data_mask : writeQueueVec_dataOut_17_data_mask;
  assign writeQueueVec_17_deq_bits_data_data = _writeQueueVec_fifo_17_empty ? writeQueueVec_17_enq_bits_data_data : writeQueueVec_dataOut_17_data_data;
  assign writeQueueVec_17_deq_bits_data_last = _writeQueueVec_fifo_17_empty ? writeQueueVec_17_enq_bits_data_last : writeQueueVec_dataOut_17_data_last;
  assign writeQueueVec_17_deq_bits_data_instructionIndex = _writeQueueVec_fifo_17_empty ? writeQueueVec_17_enq_bits_data_instructionIndex : writeQueueVec_dataOut_17_data_instructionIndex;
  wire [31:0]       writeQueueVec_17_deq_bits_targetLane = _writeQueueVec_fifo_17_empty ? 32'h20000 : writeQueueVec_dataOut_17_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_18 = writeQueueVec_18_enq_bits_data_vd;
  wire              vrfWritePort_18_valid_0 = writeQueueVec_18_deq_valid;
  wire [4:0]        vrfWritePort_18_bits_vd_0 = writeQueueVec_18_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_18_bits_mask_0 = writeQueueVec_18_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_18_bits_data_0 = writeQueueVec_18_deq_bits_data_data;
  wire              vrfWritePort_18_bits_last_0 = writeQueueVec_18_deq_bits_data_last;
  wire [2:0]        vrfWritePort_18_bits_instructionIndex_0 = writeQueueVec_18_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_18_enq_bits = writeQueueVec_18_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_18_enq_bits_data_data;
  wire              writeQueueVec_18_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_18 = {writeQueueVec_18_enq_bits_data_data, writeQueueVec_18_enq_bits_data_last};
  wire [2:0]        writeQueueVec_18_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_18 = {writeQueueVec_dataIn_lo_hi_18, writeQueueVec_18_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_18_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_18 = {writeQueueVec_dataIn_hi_hi_18, writeQueueVec_18_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_18 = {writeQueueVec_dataIn_hi_18, writeQueueVec_dataIn_lo_18, 32'h40000};
  wire [31:0]       writeQueueVec_dataOut_18_targetLane = _writeQueueVec_fifo_18_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_18_data_instructionIndex = _writeQueueVec_fifo_18_data_out[34:32];
  wire              writeQueueVec_dataOut_18_data_last = _writeQueueVec_fifo_18_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_18_data_data = _writeQueueVec_fifo_18_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_18_data_mask = _writeQueueVec_fifo_18_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_18_data_vd = _writeQueueVec_fifo_18_data_out[76:72];
  wire              writeQueueVec_18_enq_ready = ~_writeQueueVec_fifo_18_full;
  wire              writeQueueVec_18_enq_valid;
  wire              _probeWire_slots_18_writeValid_T = writeQueueVec_18_enq_ready & writeQueueVec_18_enq_valid;
  assign writeQueueVec_18_deq_valid = ~_writeQueueVec_fifo_18_empty | writeQueueVec_18_enq_valid;
  assign writeQueueVec_18_deq_bits_data_vd = _writeQueueVec_fifo_18_empty ? writeQueueVec_18_enq_bits_data_vd : writeQueueVec_dataOut_18_data_vd;
  assign writeQueueVec_18_deq_bits_data_mask = _writeQueueVec_fifo_18_empty ? writeQueueVec_18_enq_bits_data_mask : writeQueueVec_dataOut_18_data_mask;
  assign writeQueueVec_18_deq_bits_data_data = _writeQueueVec_fifo_18_empty ? writeQueueVec_18_enq_bits_data_data : writeQueueVec_dataOut_18_data_data;
  assign writeQueueVec_18_deq_bits_data_last = _writeQueueVec_fifo_18_empty ? writeQueueVec_18_enq_bits_data_last : writeQueueVec_dataOut_18_data_last;
  assign writeQueueVec_18_deq_bits_data_instructionIndex = _writeQueueVec_fifo_18_empty ? writeQueueVec_18_enq_bits_data_instructionIndex : writeQueueVec_dataOut_18_data_instructionIndex;
  wire [31:0]       writeQueueVec_18_deq_bits_targetLane = _writeQueueVec_fifo_18_empty ? 32'h40000 : writeQueueVec_dataOut_18_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_19 = writeQueueVec_19_enq_bits_data_vd;
  wire              vrfWritePort_19_valid_0 = writeQueueVec_19_deq_valid;
  wire [4:0]        vrfWritePort_19_bits_vd_0 = writeQueueVec_19_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_19_bits_mask_0 = writeQueueVec_19_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_19_bits_data_0 = writeQueueVec_19_deq_bits_data_data;
  wire              vrfWritePort_19_bits_last_0 = writeQueueVec_19_deq_bits_data_last;
  wire [2:0]        vrfWritePort_19_bits_instructionIndex_0 = writeQueueVec_19_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_19_enq_bits = writeQueueVec_19_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_19_enq_bits_data_data;
  wire              writeQueueVec_19_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_19 = {writeQueueVec_19_enq_bits_data_data, writeQueueVec_19_enq_bits_data_last};
  wire [2:0]        writeQueueVec_19_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_19 = {writeQueueVec_dataIn_lo_hi_19, writeQueueVec_19_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_19_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_19 = {writeQueueVec_dataIn_hi_hi_19, writeQueueVec_19_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_19 = {writeQueueVec_dataIn_hi_19, writeQueueVec_dataIn_lo_19, 32'h80000};
  wire [31:0]       writeQueueVec_dataOut_19_targetLane = _writeQueueVec_fifo_19_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_19_data_instructionIndex = _writeQueueVec_fifo_19_data_out[34:32];
  wire              writeQueueVec_dataOut_19_data_last = _writeQueueVec_fifo_19_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_19_data_data = _writeQueueVec_fifo_19_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_19_data_mask = _writeQueueVec_fifo_19_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_19_data_vd = _writeQueueVec_fifo_19_data_out[76:72];
  wire              writeQueueVec_19_enq_ready = ~_writeQueueVec_fifo_19_full;
  wire              writeQueueVec_19_enq_valid;
  wire              _probeWire_slots_19_writeValid_T = writeQueueVec_19_enq_ready & writeQueueVec_19_enq_valid;
  assign writeQueueVec_19_deq_valid = ~_writeQueueVec_fifo_19_empty | writeQueueVec_19_enq_valid;
  assign writeQueueVec_19_deq_bits_data_vd = _writeQueueVec_fifo_19_empty ? writeQueueVec_19_enq_bits_data_vd : writeQueueVec_dataOut_19_data_vd;
  assign writeQueueVec_19_deq_bits_data_mask = _writeQueueVec_fifo_19_empty ? writeQueueVec_19_enq_bits_data_mask : writeQueueVec_dataOut_19_data_mask;
  assign writeQueueVec_19_deq_bits_data_data = _writeQueueVec_fifo_19_empty ? writeQueueVec_19_enq_bits_data_data : writeQueueVec_dataOut_19_data_data;
  assign writeQueueVec_19_deq_bits_data_last = _writeQueueVec_fifo_19_empty ? writeQueueVec_19_enq_bits_data_last : writeQueueVec_dataOut_19_data_last;
  assign writeQueueVec_19_deq_bits_data_instructionIndex = _writeQueueVec_fifo_19_empty ? writeQueueVec_19_enq_bits_data_instructionIndex : writeQueueVec_dataOut_19_data_instructionIndex;
  wire [31:0]       writeQueueVec_19_deq_bits_targetLane = _writeQueueVec_fifo_19_empty ? 32'h80000 : writeQueueVec_dataOut_19_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_20 = writeQueueVec_20_enq_bits_data_vd;
  wire              vrfWritePort_20_valid_0 = writeQueueVec_20_deq_valid;
  wire [4:0]        vrfWritePort_20_bits_vd_0 = writeQueueVec_20_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_20_bits_mask_0 = writeQueueVec_20_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_20_bits_data_0 = writeQueueVec_20_deq_bits_data_data;
  wire              vrfWritePort_20_bits_last_0 = writeQueueVec_20_deq_bits_data_last;
  wire [2:0]        vrfWritePort_20_bits_instructionIndex_0 = writeQueueVec_20_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_20_enq_bits = writeQueueVec_20_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_20_enq_bits_data_data;
  wire              writeQueueVec_20_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_20 = {writeQueueVec_20_enq_bits_data_data, writeQueueVec_20_enq_bits_data_last};
  wire [2:0]        writeQueueVec_20_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_20 = {writeQueueVec_dataIn_lo_hi_20, writeQueueVec_20_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_20_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_20 = {writeQueueVec_dataIn_hi_hi_20, writeQueueVec_20_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_20 = {writeQueueVec_dataIn_hi_20, writeQueueVec_dataIn_lo_20, 32'h100000};
  wire [31:0]       writeQueueVec_dataOut_20_targetLane = _writeQueueVec_fifo_20_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_20_data_instructionIndex = _writeQueueVec_fifo_20_data_out[34:32];
  wire              writeQueueVec_dataOut_20_data_last = _writeQueueVec_fifo_20_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_20_data_data = _writeQueueVec_fifo_20_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_20_data_mask = _writeQueueVec_fifo_20_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_20_data_vd = _writeQueueVec_fifo_20_data_out[76:72];
  wire              writeQueueVec_20_enq_ready = ~_writeQueueVec_fifo_20_full;
  wire              writeQueueVec_20_enq_valid;
  wire              _probeWire_slots_20_writeValid_T = writeQueueVec_20_enq_ready & writeQueueVec_20_enq_valid;
  assign writeQueueVec_20_deq_valid = ~_writeQueueVec_fifo_20_empty | writeQueueVec_20_enq_valid;
  assign writeQueueVec_20_deq_bits_data_vd = _writeQueueVec_fifo_20_empty ? writeQueueVec_20_enq_bits_data_vd : writeQueueVec_dataOut_20_data_vd;
  assign writeQueueVec_20_deq_bits_data_mask = _writeQueueVec_fifo_20_empty ? writeQueueVec_20_enq_bits_data_mask : writeQueueVec_dataOut_20_data_mask;
  assign writeQueueVec_20_deq_bits_data_data = _writeQueueVec_fifo_20_empty ? writeQueueVec_20_enq_bits_data_data : writeQueueVec_dataOut_20_data_data;
  assign writeQueueVec_20_deq_bits_data_last = _writeQueueVec_fifo_20_empty ? writeQueueVec_20_enq_bits_data_last : writeQueueVec_dataOut_20_data_last;
  assign writeQueueVec_20_deq_bits_data_instructionIndex = _writeQueueVec_fifo_20_empty ? writeQueueVec_20_enq_bits_data_instructionIndex : writeQueueVec_dataOut_20_data_instructionIndex;
  wire [31:0]       writeQueueVec_20_deq_bits_targetLane = _writeQueueVec_fifo_20_empty ? 32'h100000 : writeQueueVec_dataOut_20_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_21 = writeQueueVec_21_enq_bits_data_vd;
  wire              vrfWritePort_21_valid_0 = writeQueueVec_21_deq_valid;
  wire [4:0]        vrfWritePort_21_bits_vd_0 = writeQueueVec_21_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_21_bits_mask_0 = writeQueueVec_21_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_21_bits_data_0 = writeQueueVec_21_deq_bits_data_data;
  wire              vrfWritePort_21_bits_last_0 = writeQueueVec_21_deq_bits_data_last;
  wire [2:0]        vrfWritePort_21_bits_instructionIndex_0 = writeQueueVec_21_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_21_enq_bits = writeQueueVec_21_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_21_enq_bits_data_data;
  wire              writeQueueVec_21_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_21 = {writeQueueVec_21_enq_bits_data_data, writeQueueVec_21_enq_bits_data_last};
  wire [2:0]        writeQueueVec_21_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_21 = {writeQueueVec_dataIn_lo_hi_21, writeQueueVec_21_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_21_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_21 = {writeQueueVec_dataIn_hi_hi_21, writeQueueVec_21_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_21 = {writeQueueVec_dataIn_hi_21, writeQueueVec_dataIn_lo_21, 32'h200000};
  wire [31:0]       writeQueueVec_dataOut_21_targetLane = _writeQueueVec_fifo_21_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_21_data_instructionIndex = _writeQueueVec_fifo_21_data_out[34:32];
  wire              writeQueueVec_dataOut_21_data_last = _writeQueueVec_fifo_21_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_21_data_data = _writeQueueVec_fifo_21_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_21_data_mask = _writeQueueVec_fifo_21_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_21_data_vd = _writeQueueVec_fifo_21_data_out[76:72];
  wire              writeQueueVec_21_enq_ready = ~_writeQueueVec_fifo_21_full;
  wire              writeQueueVec_21_enq_valid;
  wire              _probeWire_slots_21_writeValid_T = writeQueueVec_21_enq_ready & writeQueueVec_21_enq_valid;
  assign writeQueueVec_21_deq_valid = ~_writeQueueVec_fifo_21_empty | writeQueueVec_21_enq_valid;
  assign writeQueueVec_21_deq_bits_data_vd = _writeQueueVec_fifo_21_empty ? writeQueueVec_21_enq_bits_data_vd : writeQueueVec_dataOut_21_data_vd;
  assign writeQueueVec_21_deq_bits_data_mask = _writeQueueVec_fifo_21_empty ? writeQueueVec_21_enq_bits_data_mask : writeQueueVec_dataOut_21_data_mask;
  assign writeQueueVec_21_deq_bits_data_data = _writeQueueVec_fifo_21_empty ? writeQueueVec_21_enq_bits_data_data : writeQueueVec_dataOut_21_data_data;
  assign writeQueueVec_21_deq_bits_data_last = _writeQueueVec_fifo_21_empty ? writeQueueVec_21_enq_bits_data_last : writeQueueVec_dataOut_21_data_last;
  assign writeQueueVec_21_deq_bits_data_instructionIndex = _writeQueueVec_fifo_21_empty ? writeQueueVec_21_enq_bits_data_instructionIndex : writeQueueVec_dataOut_21_data_instructionIndex;
  wire [31:0]       writeQueueVec_21_deq_bits_targetLane = _writeQueueVec_fifo_21_empty ? 32'h200000 : writeQueueVec_dataOut_21_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_22 = writeQueueVec_22_enq_bits_data_vd;
  wire              vrfWritePort_22_valid_0 = writeQueueVec_22_deq_valid;
  wire [4:0]        vrfWritePort_22_bits_vd_0 = writeQueueVec_22_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_22_bits_mask_0 = writeQueueVec_22_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_22_bits_data_0 = writeQueueVec_22_deq_bits_data_data;
  wire              vrfWritePort_22_bits_last_0 = writeQueueVec_22_deq_bits_data_last;
  wire [2:0]        vrfWritePort_22_bits_instructionIndex_0 = writeQueueVec_22_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_22_enq_bits = writeQueueVec_22_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_22_enq_bits_data_data;
  wire              writeQueueVec_22_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_22 = {writeQueueVec_22_enq_bits_data_data, writeQueueVec_22_enq_bits_data_last};
  wire [2:0]        writeQueueVec_22_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_22 = {writeQueueVec_dataIn_lo_hi_22, writeQueueVec_22_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_22_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_22 = {writeQueueVec_dataIn_hi_hi_22, writeQueueVec_22_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_22 = {writeQueueVec_dataIn_hi_22, writeQueueVec_dataIn_lo_22, 32'h400000};
  wire [31:0]       writeQueueVec_dataOut_22_targetLane = _writeQueueVec_fifo_22_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_22_data_instructionIndex = _writeQueueVec_fifo_22_data_out[34:32];
  wire              writeQueueVec_dataOut_22_data_last = _writeQueueVec_fifo_22_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_22_data_data = _writeQueueVec_fifo_22_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_22_data_mask = _writeQueueVec_fifo_22_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_22_data_vd = _writeQueueVec_fifo_22_data_out[76:72];
  wire              writeQueueVec_22_enq_ready = ~_writeQueueVec_fifo_22_full;
  wire              writeQueueVec_22_enq_valid;
  wire              _probeWire_slots_22_writeValid_T = writeQueueVec_22_enq_ready & writeQueueVec_22_enq_valid;
  assign writeQueueVec_22_deq_valid = ~_writeQueueVec_fifo_22_empty | writeQueueVec_22_enq_valid;
  assign writeQueueVec_22_deq_bits_data_vd = _writeQueueVec_fifo_22_empty ? writeQueueVec_22_enq_bits_data_vd : writeQueueVec_dataOut_22_data_vd;
  assign writeQueueVec_22_deq_bits_data_mask = _writeQueueVec_fifo_22_empty ? writeQueueVec_22_enq_bits_data_mask : writeQueueVec_dataOut_22_data_mask;
  assign writeQueueVec_22_deq_bits_data_data = _writeQueueVec_fifo_22_empty ? writeQueueVec_22_enq_bits_data_data : writeQueueVec_dataOut_22_data_data;
  assign writeQueueVec_22_deq_bits_data_last = _writeQueueVec_fifo_22_empty ? writeQueueVec_22_enq_bits_data_last : writeQueueVec_dataOut_22_data_last;
  assign writeQueueVec_22_deq_bits_data_instructionIndex = _writeQueueVec_fifo_22_empty ? writeQueueVec_22_enq_bits_data_instructionIndex : writeQueueVec_dataOut_22_data_instructionIndex;
  wire [31:0]       writeQueueVec_22_deq_bits_targetLane = _writeQueueVec_fifo_22_empty ? 32'h400000 : writeQueueVec_dataOut_22_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_23 = writeQueueVec_23_enq_bits_data_vd;
  wire              vrfWritePort_23_valid_0 = writeQueueVec_23_deq_valid;
  wire [4:0]        vrfWritePort_23_bits_vd_0 = writeQueueVec_23_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_23_bits_mask_0 = writeQueueVec_23_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_23_bits_data_0 = writeQueueVec_23_deq_bits_data_data;
  wire              vrfWritePort_23_bits_last_0 = writeQueueVec_23_deq_bits_data_last;
  wire [2:0]        vrfWritePort_23_bits_instructionIndex_0 = writeQueueVec_23_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_23_enq_bits = writeQueueVec_23_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_23_enq_bits_data_data;
  wire              writeQueueVec_23_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_23 = {writeQueueVec_23_enq_bits_data_data, writeQueueVec_23_enq_bits_data_last};
  wire [2:0]        writeQueueVec_23_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_23 = {writeQueueVec_dataIn_lo_hi_23, writeQueueVec_23_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_23_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_23 = {writeQueueVec_dataIn_hi_hi_23, writeQueueVec_23_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_23 = {writeQueueVec_dataIn_hi_23, writeQueueVec_dataIn_lo_23, 32'h800000};
  wire [31:0]       writeQueueVec_dataOut_23_targetLane = _writeQueueVec_fifo_23_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_23_data_instructionIndex = _writeQueueVec_fifo_23_data_out[34:32];
  wire              writeQueueVec_dataOut_23_data_last = _writeQueueVec_fifo_23_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_23_data_data = _writeQueueVec_fifo_23_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_23_data_mask = _writeQueueVec_fifo_23_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_23_data_vd = _writeQueueVec_fifo_23_data_out[76:72];
  wire              writeQueueVec_23_enq_ready = ~_writeQueueVec_fifo_23_full;
  wire              writeQueueVec_23_enq_valid;
  wire              _probeWire_slots_23_writeValid_T = writeQueueVec_23_enq_ready & writeQueueVec_23_enq_valid;
  assign writeQueueVec_23_deq_valid = ~_writeQueueVec_fifo_23_empty | writeQueueVec_23_enq_valid;
  assign writeQueueVec_23_deq_bits_data_vd = _writeQueueVec_fifo_23_empty ? writeQueueVec_23_enq_bits_data_vd : writeQueueVec_dataOut_23_data_vd;
  assign writeQueueVec_23_deq_bits_data_mask = _writeQueueVec_fifo_23_empty ? writeQueueVec_23_enq_bits_data_mask : writeQueueVec_dataOut_23_data_mask;
  assign writeQueueVec_23_deq_bits_data_data = _writeQueueVec_fifo_23_empty ? writeQueueVec_23_enq_bits_data_data : writeQueueVec_dataOut_23_data_data;
  assign writeQueueVec_23_deq_bits_data_last = _writeQueueVec_fifo_23_empty ? writeQueueVec_23_enq_bits_data_last : writeQueueVec_dataOut_23_data_last;
  assign writeQueueVec_23_deq_bits_data_instructionIndex = _writeQueueVec_fifo_23_empty ? writeQueueVec_23_enq_bits_data_instructionIndex : writeQueueVec_dataOut_23_data_instructionIndex;
  wire [31:0]       writeQueueVec_23_deq_bits_targetLane = _writeQueueVec_fifo_23_empty ? 32'h800000 : writeQueueVec_dataOut_23_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_24 = writeQueueVec_24_enq_bits_data_vd;
  wire              vrfWritePort_24_valid_0 = writeQueueVec_24_deq_valid;
  wire [4:0]        vrfWritePort_24_bits_vd_0 = writeQueueVec_24_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_24_bits_mask_0 = writeQueueVec_24_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_24_bits_data_0 = writeQueueVec_24_deq_bits_data_data;
  wire              vrfWritePort_24_bits_last_0 = writeQueueVec_24_deq_bits_data_last;
  wire [2:0]        vrfWritePort_24_bits_instructionIndex_0 = writeQueueVec_24_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_24_enq_bits = writeQueueVec_24_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_24_enq_bits_data_data;
  wire              writeQueueVec_24_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_24 = {writeQueueVec_24_enq_bits_data_data, writeQueueVec_24_enq_bits_data_last};
  wire [2:0]        writeQueueVec_24_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_24 = {writeQueueVec_dataIn_lo_hi_24, writeQueueVec_24_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_24_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_24 = {writeQueueVec_dataIn_hi_hi_24, writeQueueVec_24_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_24 = {writeQueueVec_dataIn_hi_24, writeQueueVec_dataIn_lo_24, 32'h1000000};
  wire [31:0]       writeQueueVec_dataOut_24_targetLane = _writeQueueVec_fifo_24_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_24_data_instructionIndex = _writeQueueVec_fifo_24_data_out[34:32];
  wire              writeQueueVec_dataOut_24_data_last = _writeQueueVec_fifo_24_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_24_data_data = _writeQueueVec_fifo_24_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_24_data_mask = _writeQueueVec_fifo_24_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_24_data_vd = _writeQueueVec_fifo_24_data_out[76:72];
  wire              writeQueueVec_24_enq_ready = ~_writeQueueVec_fifo_24_full;
  wire              writeQueueVec_24_enq_valid;
  wire              _probeWire_slots_24_writeValid_T = writeQueueVec_24_enq_ready & writeQueueVec_24_enq_valid;
  assign writeQueueVec_24_deq_valid = ~_writeQueueVec_fifo_24_empty | writeQueueVec_24_enq_valid;
  assign writeQueueVec_24_deq_bits_data_vd = _writeQueueVec_fifo_24_empty ? writeQueueVec_24_enq_bits_data_vd : writeQueueVec_dataOut_24_data_vd;
  assign writeQueueVec_24_deq_bits_data_mask = _writeQueueVec_fifo_24_empty ? writeQueueVec_24_enq_bits_data_mask : writeQueueVec_dataOut_24_data_mask;
  assign writeQueueVec_24_deq_bits_data_data = _writeQueueVec_fifo_24_empty ? writeQueueVec_24_enq_bits_data_data : writeQueueVec_dataOut_24_data_data;
  assign writeQueueVec_24_deq_bits_data_last = _writeQueueVec_fifo_24_empty ? writeQueueVec_24_enq_bits_data_last : writeQueueVec_dataOut_24_data_last;
  assign writeQueueVec_24_deq_bits_data_instructionIndex = _writeQueueVec_fifo_24_empty ? writeQueueVec_24_enq_bits_data_instructionIndex : writeQueueVec_dataOut_24_data_instructionIndex;
  wire [31:0]       writeQueueVec_24_deq_bits_targetLane = _writeQueueVec_fifo_24_empty ? 32'h1000000 : writeQueueVec_dataOut_24_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_25 = writeQueueVec_25_enq_bits_data_vd;
  wire              vrfWritePort_25_valid_0 = writeQueueVec_25_deq_valid;
  wire [4:0]        vrfWritePort_25_bits_vd_0 = writeQueueVec_25_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_25_bits_mask_0 = writeQueueVec_25_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_25_bits_data_0 = writeQueueVec_25_deq_bits_data_data;
  wire              vrfWritePort_25_bits_last_0 = writeQueueVec_25_deq_bits_data_last;
  wire [2:0]        vrfWritePort_25_bits_instructionIndex_0 = writeQueueVec_25_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_25_enq_bits = writeQueueVec_25_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_25_enq_bits_data_data;
  wire              writeQueueVec_25_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_25 = {writeQueueVec_25_enq_bits_data_data, writeQueueVec_25_enq_bits_data_last};
  wire [2:0]        writeQueueVec_25_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_25 = {writeQueueVec_dataIn_lo_hi_25, writeQueueVec_25_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_25_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_25 = {writeQueueVec_dataIn_hi_hi_25, writeQueueVec_25_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_25 = {writeQueueVec_dataIn_hi_25, writeQueueVec_dataIn_lo_25, 32'h2000000};
  wire [31:0]       writeQueueVec_dataOut_25_targetLane = _writeQueueVec_fifo_25_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_25_data_instructionIndex = _writeQueueVec_fifo_25_data_out[34:32];
  wire              writeQueueVec_dataOut_25_data_last = _writeQueueVec_fifo_25_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_25_data_data = _writeQueueVec_fifo_25_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_25_data_mask = _writeQueueVec_fifo_25_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_25_data_vd = _writeQueueVec_fifo_25_data_out[76:72];
  wire              writeQueueVec_25_enq_ready = ~_writeQueueVec_fifo_25_full;
  wire              writeQueueVec_25_enq_valid;
  wire              _probeWire_slots_25_writeValid_T = writeQueueVec_25_enq_ready & writeQueueVec_25_enq_valid;
  assign writeQueueVec_25_deq_valid = ~_writeQueueVec_fifo_25_empty | writeQueueVec_25_enq_valid;
  assign writeQueueVec_25_deq_bits_data_vd = _writeQueueVec_fifo_25_empty ? writeQueueVec_25_enq_bits_data_vd : writeQueueVec_dataOut_25_data_vd;
  assign writeQueueVec_25_deq_bits_data_mask = _writeQueueVec_fifo_25_empty ? writeQueueVec_25_enq_bits_data_mask : writeQueueVec_dataOut_25_data_mask;
  assign writeQueueVec_25_deq_bits_data_data = _writeQueueVec_fifo_25_empty ? writeQueueVec_25_enq_bits_data_data : writeQueueVec_dataOut_25_data_data;
  assign writeQueueVec_25_deq_bits_data_last = _writeQueueVec_fifo_25_empty ? writeQueueVec_25_enq_bits_data_last : writeQueueVec_dataOut_25_data_last;
  assign writeQueueVec_25_deq_bits_data_instructionIndex = _writeQueueVec_fifo_25_empty ? writeQueueVec_25_enq_bits_data_instructionIndex : writeQueueVec_dataOut_25_data_instructionIndex;
  wire [31:0]       writeQueueVec_25_deq_bits_targetLane = _writeQueueVec_fifo_25_empty ? 32'h2000000 : writeQueueVec_dataOut_25_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_26 = writeQueueVec_26_enq_bits_data_vd;
  wire              vrfWritePort_26_valid_0 = writeQueueVec_26_deq_valid;
  wire [4:0]        vrfWritePort_26_bits_vd_0 = writeQueueVec_26_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_26_bits_mask_0 = writeQueueVec_26_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_26_bits_data_0 = writeQueueVec_26_deq_bits_data_data;
  wire              vrfWritePort_26_bits_last_0 = writeQueueVec_26_deq_bits_data_last;
  wire [2:0]        vrfWritePort_26_bits_instructionIndex_0 = writeQueueVec_26_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_26_enq_bits = writeQueueVec_26_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_26_enq_bits_data_data;
  wire              writeQueueVec_26_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_26 = {writeQueueVec_26_enq_bits_data_data, writeQueueVec_26_enq_bits_data_last};
  wire [2:0]        writeQueueVec_26_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_26 = {writeQueueVec_dataIn_lo_hi_26, writeQueueVec_26_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_26_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_26 = {writeQueueVec_dataIn_hi_hi_26, writeQueueVec_26_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_26 = {writeQueueVec_dataIn_hi_26, writeQueueVec_dataIn_lo_26, 32'h4000000};
  wire [31:0]       writeQueueVec_dataOut_26_targetLane = _writeQueueVec_fifo_26_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_26_data_instructionIndex = _writeQueueVec_fifo_26_data_out[34:32];
  wire              writeQueueVec_dataOut_26_data_last = _writeQueueVec_fifo_26_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_26_data_data = _writeQueueVec_fifo_26_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_26_data_mask = _writeQueueVec_fifo_26_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_26_data_vd = _writeQueueVec_fifo_26_data_out[76:72];
  wire              writeQueueVec_26_enq_ready = ~_writeQueueVec_fifo_26_full;
  wire              writeQueueVec_26_enq_valid;
  wire              _probeWire_slots_26_writeValid_T = writeQueueVec_26_enq_ready & writeQueueVec_26_enq_valid;
  assign writeQueueVec_26_deq_valid = ~_writeQueueVec_fifo_26_empty | writeQueueVec_26_enq_valid;
  assign writeQueueVec_26_deq_bits_data_vd = _writeQueueVec_fifo_26_empty ? writeQueueVec_26_enq_bits_data_vd : writeQueueVec_dataOut_26_data_vd;
  assign writeQueueVec_26_deq_bits_data_mask = _writeQueueVec_fifo_26_empty ? writeQueueVec_26_enq_bits_data_mask : writeQueueVec_dataOut_26_data_mask;
  assign writeQueueVec_26_deq_bits_data_data = _writeQueueVec_fifo_26_empty ? writeQueueVec_26_enq_bits_data_data : writeQueueVec_dataOut_26_data_data;
  assign writeQueueVec_26_deq_bits_data_last = _writeQueueVec_fifo_26_empty ? writeQueueVec_26_enq_bits_data_last : writeQueueVec_dataOut_26_data_last;
  assign writeQueueVec_26_deq_bits_data_instructionIndex = _writeQueueVec_fifo_26_empty ? writeQueueVec_26_enq_bits_data_instructionIndex : writeQueueVec_dataOut_26_data_instructionIndex;
  wire [31:0]       writeQueueVec_26_deq_bits_targetLane = _writeQueueVec_fifo_26_empty ? 32'h4000000 : writeQueueVec_dataOut_26_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_27 = writeQueueVec_27_enq_bits_data_vd;
  wire              vrfWritePort_27_valid_0 = writeQueueVec_27_deq_valid;
  wire [4:0]        vrfWritePort_27_bits_vd_0 = writeQueueVec_27_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_27_bits_mask_0 = writeQueueVec_27_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_27_bits_data_0 = writeQueueVec_27_deq_bits_data_data;
  wire              vrfWritePort_27_bits_last_0 = writeQueueVec_27_deq_bits_data_last;
  wire [2:0]        vrfWritePort_27_bits_instructionIndex_0 = writeQueueVec_27_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_27_enq_bits = writeQueueVec_27_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_27_enq_bits_data_data;
  wire              writeQueueVec_27_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_27 = {writeQueueVec_27_enq_bits_data_data, writeQueueVec_27_enq_bits_data_last};
  wire [2:0]        writeQueueVec_27_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_27 = {writeQueueVec_dataIn_lo_hi_27, writeQueueVec_27_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_27_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_27 = {writeQueueVec_dataIn_hi_hi_27, writeQueueVec_27_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_27 = {writeQueueVec_dataIn_hi_27, writeQueueVec_dataIn_lo_27, 32'h8000000};
  wire [31:0]       writeQueueVec_dataOut_27_targetLane = _writeQueueVec_fifo_27_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_27_data_instructionIndex = _writeQueueVec_fifo_27_data_out[34:32];
  wire              writeQueueVec_dataOut_27_data_last = _writeQueueVec_fifo_27_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_27_data_data = _writeQueueVec_fifo_27_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_27_data_mask = _writeQueueVec_fifo_27_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_27_data_vd = _writeQueueVec_fifo_27_data_out[76:72];
  wire              writeQueueVec_27_enq_ready = ~_writeQueueVec_fifo_27_full;
  wire              writeQueueVec_27_enq_valid;
  wire              _probeWire_slots_27_writeValid_T = writeQueueVec_27_enq_ready & writeQueueVec_27_enq_valid;
  assign writeQueueVec_27_deq_valid = ~_writeQueueVec_fifo_27_empty | writeQueueVec_27_enq_valid;
  assign writeQueueVec_27_deq_bits_data_vd = _writeQueueVec_fifo_27_empty ? writeQueueVec_27_enq_bits_data_vd : writeQueueVec_dataOut_27_data_vd;
  assign writeQueueVec_27_deq_bits_data_mask = _writeQueueVec_fifo_27_empty ? writeQueueVec_27_enq_bits_data_mask : writeQueueVec_dataOut_27_data_mask;
  assign writeQueueVec_27_deq_bits_data_data = _writeQueueVec_fifo_27_empty ? writeQueueVec_27_enq_bits_data_data : writeQueueVec_dataOut_27_data_data;
  assign writeQueueVec_27_deq_bits_data_last = _writeQueueVec_fifo_27_empty ? writeQueueVec_27_enq_bits_data_last : writeQueueVec_dataOut_27_data_last;
  assign writeQueueVec_27_deq_bits_data_instructionIndex = _writeQueueVec_fifo_27_empty ? writeQueueVec_27_enq_bits_data_instructionIndex : writeQueueVec_dataOut_27_data_instructionIndex;
  wire [31:0]       writeQueueVec_27_deq_bits_targetLane = _writeQueueVec_fifo_27_empty ? 32'h8000000 : writeQueueVec_dataOut_27_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_28 = writeQueueVec_28_enq_bits_data_vd;
  wire              vrfWritePort_28_valid_0 = writeQueueVec_28_deq_valid;
  wire [4:0]        vrfWritePort_28_bits_vd_0 = writeQueueVec_28_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_28_bits_mask_0 = writeQueueVec_28_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_28_bits_data_0 = writeQueueVec_28_deq_bits_data_data;
  wire              vrfWritePort_28_bits_last_0 = writeQueueVec_28_deq_bits_data_last;
  wire [2:0]        vrfWritePort_28_bits_instructionIndex_0 = writeQueueVec_28_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_28_enq_bits = writeQueueVec_28_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_28_enq_bits_data_data;
  wire              writeQueueVec_28_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_28 = {writeQueueVec_28_enq_bits_data_data, writeQueueVec_28_enq_bits_data_last};
  wire [2:0]        writeQueueVec_28_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_28 = {writeQueueVec_dataIn_lo_hi_28, writeQueueVec_28_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_28_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_28 = {writeQueueVec_dataIn_hi_hi_28, writeQueueVec_28_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_28 = {writeQueueVec_dataIn_hi_28, writeQueueVec_dataIn_lo_28, 32'h10000000};
  wire [31:0]       writeQueueVec_dataOut_28_targetLane = _writeQueueVec_fifo_28_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_28_data_instructionIndex = _writeQueueVec_fifo_28_data_out[34:32];
  wire              writeQueueVec_dataOut_28_data_last = _writeQueueVec_fifo_28_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_28_data_data = _writeQueueVec_fifo_28_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_28_data_mask = _writeQueueVec_fifo_28_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_28_data_vd = _writeQueueVec_fifo_28_data_out[76:72];
  wire              writeQueueVec_28_enq_ready = ~_writeQueueVec_fifo_28_full;
  wire              writeQueueVec_28_enq_valid;
  wire              _probeWire_slots_28_writeValid_T = writeQueueVec_28_enq_ready & writeQueueVec_28_enq_valid;
  assign writeQueueVec_28_deq_valid = ~_writeQueueVec_fifo_28_empty | writeQueueVec_28_enq_valid;
  assign writeQueueVec_28_deq_bits_data_vd = _writeQueueVec_fifo_28_empty ? writeQueueVec_28_enq_bits_data_vd : writeQueueVec_dataOut_28_data_vd;
  assign writeQueueVec_28_deq_bits_data_mask = _writeQueueVec_fifo_28_empty ? writeQueueVec_28_enq_bits_data_mask : writeQueueVec_dataOut_28_data_mask;
  assign writeQueueVec_28_deq_bits_data_data = _writeQueueVec_fifo_28_empty ? writeQueueVec_28_enq_bits_data_data : writeQueueVec_dataOut_28_data_data;
  assign writeQueueVec_28_deq_bits_data_last = _writeQueueVec_fifo_28_empty ? writeQueueVec_28_enq_bits_data_last : writeQueueVec_dataOut_28_data_last;
  assign writeQueueVec_28_deq_bits_data_instructionIndex = _writeQueueVec_fifo_28_empty ? writeQueueVec_28_enq_bits_data_instructionIndex : writeQueueVec_dataOut_28_data_instructionIndex;
  wire [31:0]       writeQueueVec_28_deq_bits_targetLane = _writeQueueVec_fifo_28_empty ? 32'h10000000 : writeQueueVec_dataOut_28_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_29 = writeQueueVec_29_enq_bits_data_vd;
  wire              vrfWritePort_29_valid_0 = writeQueueVec_29_deq_valid;
  wire [4:0]        vrfWritePort_29_bits_vd_0 = writeQueueVec_29_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_29_bits_mask_0 = writeQueueVec_29_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_29_bits_data_0 = writeQueueVec_29_deq_bits_data_data;
  wire              vrfWritePort_29_bits_last_0 = writeQueueVec_29_deq_bits_data_last;
  wire [2:0]        vrfWritePort_29_bits_instructionIndex_0 = writeQueueVec_29_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_29_enq_bits = writeQueueVec_29_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_29_enq_bits_data_data;
  wire              writeQueueVec_29_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_29 = {writeQueueVec_29_enq_bits_data_data, writeQueueVec_29_enq_bits_data_last};
  wire [2:0]        writeQueueVec_29_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_29 = {writeQueueVec_dataIn_lo_hi_29, writeQueueVec_29_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_29_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_29 = {writeQueueVec_dataIn_hi_hi_29, writeQueueVec_29_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_29 = {writeQueueVec_dataIn_hi_29, writeQueueVec_dataIn_lo_29, 32'h20000000};
  wire [31:0]       writeQueueVec_dataOut_29_targetLane = _writeQueueVec_fifo_29_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_29_data_instructionIndex = _writeQueueVec_fifo_29_data_out[34:32];
  wire              writeQueueVec_dataOut_29_data_last = _writeQueueVec_fifo_29_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_29_data_data = _writeQueueVec_fifo_29_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_29_data_mask = _writeQueueVec_fifo_29_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_29_data_vd = _writeQueueVec_fifo_29_data_out[76:72];
  wire              writeQueueVec_29_enq_ready = ~_writeQueueVec_fifo_29_full;
  wire              writeQueueVec_29_enq_valid;
  wire              _probeWire_slots_29_writeValid_T = writeQueueVec_29_enq_ready & writeQueueVec_29_enq_valid;
  assign writeQueueVec_29_deq_valid = ~_writeQueueVec_fifo_29_empty | writeQueueVec_29_enq_valid;
  assign writeQueueVec_29_deq_bits_data_vd = _writeQueueVec_fifo_29_empty ? writeQueueVec_29_enq_bits_data_vd : writeQueueVec_dataOut_29_data_vd;
  assign writeQueueVec_29_deq_bits_data_mask = _writeQueueVec_fifo_29_empty ? writeQueueVec_29_enq_bits_data_mask : writeQueueVec_dataOut_29_data_mask;
  assign writeQueueVec_29_deq_bits_data_data = _writeQueueVec_fifo_29_empty ? writeQueueVec_29_enq_bits_data_data : writeQueueVec_dataOut_29_data_data;
  assign writeQueueVec_29_deq_bits_data_last = _writeQueueVec_fifo_29_empty ? writeQueueVec_29_enq_bits_data_last : writeQueueVec_dataOut_29_data_last;
  assign writeQueueVec_29_deq_bits_data_instructionIndex = _writeQueueVec_fifo_29_empty ? writeQueueVec_29_enq_bits_data_instructionIndex : writeQueueVec_dataOut_29_data_instructionIndex;
  wire [31:0]       writeQueueVec_29_deq_bits_targetLane = _writeQueueVec_fifo_29_empty ? 32'h20000000 : writeQueueVec_dataOut_29_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_30 = writeQueueVec_30_enq_bits_data_vd;
  wire              vrfWritePort_30_valid_0 = writeQueueVec_30_deq_valid;
  wire [4:0]        vrfWritePort_30_bits_vd_0 = writeQueueVec_30_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_30_bits_mask_0 = writeQueueVec_30_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_30_bits_data_0 = writeQueueVec_30_deq_bits_data_data;
  wire              vrfWritePort_30_bits_last_0 = writeQueueVec_30_deq_bits_data_last;
  wire [2:0]        vrfWritePort_30_bits_instructionIndex_0 = writeQueueVec_30_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_30_enq_bits = writeQueueVec_30_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_30_enq_bits_data_data;
  wire              writeQueueVec_30_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_30 = {writeQueueVec_30_enq_bits_data_data, writeQueueVec_30_enq_bits_data_last};
  wire [2:0]        writeQueueVec_30_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_30 = {writeQueueVec_dataIn_lo_hi_30, writeQueueVec_30_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_30_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_30 = {writeQueueVec_dataIn_hi_hi_30, writeQueueVec_30_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_30 = {writeQueueVec_dataIn_hi_30, writeQueueVec_dataIn_lo_30, 32'h40000000};
  wire [31:0]       writeQueueVec_dataOut_30_targetLane = _writeQueueVec_fifo_30_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_30_data_instructionIndex = _writeQueueVec_fifo_30_data_out[34:32];
  wire              writeQueueVec_dataOut_30_data_last = _writeQueueVec_fifo_30_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_30_data_data = _writeQueueVec_fifo_30_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_30_data_mask = _writeQueueVec_fifo_30_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_30_data_vd = _writeQueueVec_fifo_30_data_out[76:72];
  wire              writeQueueVec_30_enq_ready = ~_writeQueueVec_fifo_30_full;
  wire              writeQueueVec_30_enq_valid;
  wire              _probeWire_slots_30_writeValid_T = writeQueueVec_30_enq_ready & writeQueueVec_30_enq_valid;
  assign writeQueueVec_30_deq_valid = ~_writeQueueVec_fifo_30_empty | writeQueueVec_30_enq_valid;
  assign writeQueueVec_30_deq_bits_data_vd = _writeQueueVec_fifo_30_empty ? writeQueueVec_30_enq_bits_data_vd : writeQueueVec_dataOut_30_data_vd;
  assign writeQueueVec_30_deq_bits_data_mask = _writeQueueVec_fifo_30_empty ? writeQueueVec_30_enq_bits_data_mask : writeQueueVec_dataOut_30_data_mask;
  assign writeQueueVec_30_deq_bits_data_data = _writeQueueVec_fifo_30_empty ? writeQueueVec_30_enq_bits_data_data : writeQueueVec_dataOut_30_data_data;
  assign writeQueueVec_30_deq_bits_data_last = _writeQueueVec_fifo_30_empty ? writeQueueVec_30_enq_bits_data_last : writeQueueVec_dataOut_30_data_last;
  assign writeQueueVec_30_deq_bits_data_instructionIndex = _writeQueueVec_fifo_30_empty ? writeQueueVec_30_enq_bits_data_instructionIndex : writeQueueVec_dataOut_30_data_instructionIndex;
  wire [31:0]       writeQueueVec_30_deq_bits_targetLane = _writeQueueVec_fifo_30_empty ? 32'h40000000 : writeQueueVec_dataOut_30_targetLane;
  wire [4:0]        writeQueueVec_dataIn_hi_hi_31 = writeQueueVec_31_enq_bits_data_vd;
  wire              vrfWritePort_31_valid_0 = writeQueueVec_31_deq_valid;
  wire [4:0]        vrfWritePort_31_bits_vd_0 = writeQueueVec_31_deq_bits_data_vd;
  wire [3:0]        vrfWritePort_31_bits_mask_0 = writeQueueVec_31_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_31_bits_data_0 = writeQueueVec_31_deq_bits_data_data;
  wire              vrfWritePort_31_bits_last_0 = writeQueueVec_31_deq_bits_data_last;
  wire [2:0]        vrfWritePort_31_bits_instructionIndex_0 = writeQueueVec_31_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_31_enq_bits = writeQueueVec_31_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_31_enq_bits_data_data;
  wire              writeQueueVec_31_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_31 = {writeQueueVec_31_enq_bits_data_data, writeQueueVec_31_enq_bits_data_last};
  wire [2:0]        writeQueueVec_31_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_31 = {writeQueueVec_dataIn_lo_hi_31, writeQueueVec_31_enq_bits_data_instructionIndex};
  wire [3:0]        writeQueueVec_31_enq_bits_data_mask;
  wire [8:0]        writeQueueVec_dataIn_hi_31 = {writeQueueVec_dataIn_hi_hi_31, writeQueueVec_31_enq_bits_data_mask};
  wire [76:0]       writeQueueVec_dataIn_31 = {writeQueueVec_dataIn_hi_31, writeQueueVec_dataIn_lo_31, 32'h80000000};
  wire [31:0]       writeQueueVec_dataOut_31_targetLane = _writeQueueVec_fifo_31_data_out[31:0];
  wire [2:0]        writeQueueVec_dataOut_31_data_instructionIndex = _writeQueueVec_fifo_31_data_out[34:32];
  wire              writeQueueVec_dataOut_31_data_last = _writeQueueVec_fifo_31_data_out[35];
  wire [31:0]       writeQueueVec_dataOut_31_data_data = _writeQueueVec_fifo_31_data_out[67:36];
  wire [3:0]        writeQueueVec_dataOut_31_data_mask = _writeQueueVec_fifo_31_data_out[71:68];
  wire [4:0]        writeQueueVec_dataOut_31_data_vd = _writeQueueVec_fifo_31_data_out[76:72];
  wire              writeQueueVec_31_enq_ready = ~_writeQueueVec_fifo_31_full;
  wire              writeQueueVec_31_enq_valid;
  wire              _probeWire_slots_31_writeValid_T = writeQueueVec_31_enq_ready & writeQueueVec_31_enq_valid;
  assign writeQueueVec_31_deq_valid = ~_writeQueueVec_fifo_31_empty | writeQueueVec_31_enq_valid;
  assign writeQueueVec_31_deq_bits_data_vd = _writeQueueVec_fifo_31_empty ? writeQueueVec_31_enq_bits_data_vd : writeQueueVec_dataOut_31_data_vd;
  assign writeQueueVec_31_deq_bits_data_mask = _writeQueueVec_fifo_31_empty ? writeQueueVec_31_enq_bits_data_mask : writeQueueVec_dataOut_31_data_mask;
  assign writeQueueVec_31_deq_bits_data_data = _writeQueueVec_fifo_31_empty ? writeQueueVec_31_enq_bits_data_data : writeQueueVec_dataOut_31_data_data;
  assign writeQueueVec_31_deq_bits_data_last = _writeQueueVec_fifo_31_empty ? writeQueueVec_31_enq_bits_data_last : writeQueueVec_dataOut_31_data_last;
  assign writeQueueVec_31_deq_bits_data_instructionIndex = _writeQueueVec_fifo_31_empty ? writeQueueVec_31_enq_bits_data_instructionIndex : writeQueueVec_dataOut_31_data_instructionIndex;
  wire [31:0]       writeQueueVec_31_deq_bits_targetLane = _writeQueueVec_fifo_31_empty ? 32'h80000000 : writeQueueVec_dataOut_31_targetLane;
  wire              otherUnitTargetQueue_deq_valid;
  assign otherUnitTargetQueue_deq_valid = ~_otherUnitTargetQueue_fifo_empty;
  wire              otherUnitTargetQueue_deq_ready;
  wire              otherUnitTargetQueue_enq_ready = ~_otherUnitTargetQueue_fifo_full | otherUnitTargetQueue_deq_ready;
  wire              otherUnitTargetQueue_enq_valid;
  wire              otherUnitDataQueueVec_0_enq_ready = ~_otherUnitDataQueueVec_fifo_full;
  wire              otherUnitDataQueueVec_0_deq_ready;
  wire              otherUnitDataQueueVec_0_enq_valid;
  wire              otherUnitDataQueueVec_0_deq_valid = ~_otherUnitDataQueueVec_fifo_empty | otherUnitDataQueueVec_0_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_0_deq_bits = _otherUnitDataQueueVec_fifo_empty ? otherUnitDataQueueVec_0_enq_bits : _otherUnitDataQueueVec_fifo_data_out;
  wire              otherUnitDataQueueVec_1_enq_ready = ~_otherUnitDataQueueVec_fifo_1_full;
  wire              otherUnitDataQueueVec_1_deq_ready;
  wire              otherUnitDataQueueVec_1_enq_valid;
  wire              otherUnitDataQueueVec_1_deq_valid = ~_otherUnitDataQueueVec_fifo_1_empty | otherUnitDataQueueVec_1_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_1_deq_bits = _otherUnitDataQueueVec_fifo_1_empty ? otherUnitDataQueueVec_1_enq_bits : _otherUnitDataQueueVec_fifo_1_data_out;
  wire              otherUnitDataQueueVec_2_enq_ready = ~_otherUnitDataQueueVec_fifo_2_full;
  wire              otherUnitDataQueueVec_2_deq_ready;
  wire              otherUnitDataQueueVec_2_enq_valid;
  wire              otherUnitDataQueueVec_2_deq_valid = ~_otherUnitDataQueueVec_fifo_2_empty | otherUnitDataQueueVec_2_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_2_deq_bits = _otherUnitDataQueueVec_fifo_2_empty ? otherUnitDataQueueVec_2_enq_bits : _otherUnitDataQueueVec_fifo_2_data_out;
  wire              otherUnitDataQueueVec_3_enq_ready = ~_otherUnitDataQueueVec_fifo_3_full;
  wire              otherUnitDataQueueVec_3_deq_ready;
  wire              otherUnitDataQueueVec_3_enq_valid;
  wire              otherUnitDataQueueVec_3_deq_valid = ~_otherUnitDataQueueVec_fifo_3_empty | otherUnitDataQueueVec_3_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_3_deq_bits = _otherUnitDataQueueVec_fifo_3_empty ? otherUnitDataQueueVec_3_enq_bits : _otherUnitDataQueueVec_fifo_3_data_out;
  wire              otherUnitDataQueueVec_4_enq_ready = ~_otherUnitDataQueueVec_fifo_4_full;
  wire              otherUnitDataQueueVec_4_deq_ready;
  wire              otherUnitDataQueueVec_4_enq_valid;
  wire              otherUnitDataQueueVec_4_deq_valid = ~_otherUnitDataQueueVec_fifo_4_empty | otherUnitDataQueueVec_4_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_4_deq_bits = _otherUnitDataQueueVec_fifo_4_empty ? otherUnitDataQueueVec_4_enq_bits : _otherUnitDataQueueVec_fifo_4_data_out;
  wire              otherUnitDataQueueVec_5_enq_ready = ~_otherUnitDataQueueVec_fifo_5_full;
  wire              otherUnitDataQueueVec_5_deq_ready;
  wire              otherUnitDataQueueVec_5_enq_valid;
  wire              otherUnitDataQueueVec_5_deq_valid = ~_otherUnitDataQueueVec_fifo_5_empty | otherUnitDataQueueVec_5_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_5_deq_bits = _otherUnitDataQueueVec_fifo_5_empty ? otherUnitDataQueueVec_5_enq_bits : _otherUnitDataQueueVec_fifo_5_data_out;
  wire              otherUnitDataQueueVec_6_enq_ready = ~_otherUnitDataQueueVec_fifo_6_full;
  wire              otherUnitDataQueueVec_6_deq_ready;
  wire              otherUnitDataQueueVec_6_enq_valid;
  wire              otherUnitDataQueueVec_6_deq_valid = ~_otherUnitDataQueueVec_fifo_6_empty | otherUnitDataQueueVec_6_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_6_deq_bits = _otherUnitDataQueueVec_fifo_6_empty ? otherUnitDataQueueVec_6_enq_bits : _otherUnitDataQueueVec_fifo_6_data_out;
  wire              otherUnitDataQueueVec_7_enq_ready = ~_otherUnitDataQueueVec_fifo_7_full;
  wire              otherUnitDataQueueVec_7_deq_ready;
  wire              otherUnitDataQueueVec_7_enq_valid;
  wire              otherUnitDataQueueVec_7_deq_valid = ~_otherUnitDataQueueVec_fifo_7_empty | otherUnitDataQueueVec_7_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_7_deq_bits = _otherUnitDataQueueVec_fifo_7_empty ? otherUnitDataQueueVec_7_enq_bits : _otherUnitDataQueueVec_fifo_7_data_out;
  wire              otherUnitDataQueueVec_8_enq_ready = ~_otherUnitDataQueueVec_fifo_8_full;
  wire              otherUnitDataQueueVec_8_deq_ready;
  wire              otherUnitDataQueueVec_8_enq_valid;
  wire              otherUnitDataQueueVec_8_deq_valid = ~_otherUnitDataQueueVec_fifo_8_empty | otherUnitDataQueueVec_8_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_8_deq_bits = _otherUnitDataQueueVec_fifo_8_empty ? otherUnitDataQueueVec_8_enq_bits : _otherUnitDataQueueVec_fifo_8_data_out;
  wire              otherUnitDataQueueVec_9_enq_ready = ~_otherUnitDataQueueVec_fifo_9_full;
  wire              otherUnitDataQueueVec_9_deq_ready;
  wire              otherUnitDataQueueVec_9_enq_valid;
  wire              otherUnitDataQueueVec_9_deq_valid = ~_otherUnitDataQueueVec_fifo_9_empty | otherUnitDataQueueVec_9_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_9_deq_bits = _otherUnitDataQueueVec_fifo_9_empty ? otherUnitDataQueueVec_9_enq_bits : _otherUnitDataQueueVec_fifo_9_data_out;
  wire              otherUnitDataQueueVec_10_enq_ready = ~_otherUnitDataQueueVec_fifo_10_full;
  wire              otherUnitDataQueueVec_10_deq_ready;
  wire              otherUnitDataQueueVec_10_enq_valid;
  wire              otherUnitDataQueueVec_10_deq_valid = ~_otherUnitDataQueueVec_fifo_10_empty | otherUnitDataQueueVec_10_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_10_deq_bits = _otherUnitDataQueueVec_fifo_10_empty ? otherUnitDataQueueVec_10_enq_bits : _otherUnitDataQueueVec_fifo_10_data_out;
  wire              otherUnitDataQueueVec_11_enq_ready = ~_otherUnitDataQueueVec_fifo_11_full;
  wire              otherUnitDataQueueVec_11_deq_ready;
  wire              otherUnitDataQueueVec_11_enq_valid;
  wire              otherUnitDataQueueVec_11_deq_valid = ~_otherUnitDataQueueVec_fifo_11_empty | otherUnitDataQueueVec_11_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_11_deq_bits = _otherUnitDataQueueVec_fifo_11_empty ? otherUnitDataQueueVec_11_enq_bits : _otherUnitDataQueueVec_fifo_11_data_out;
  wire              otherUnitDataQueueVec_12_enq_ready = ~_otherUnitDataQueueVec_fifo_12_full;
  wire              otherUnitDataQueueVec_12_deq_ready;
  wire              otherUnitDataQueueVec_12_enq_valid;
  wire              otherUnitDataQueueVec_12_deq_valid = ~_otherUnitDataQueueVec_fifo_12_empty | otherUnitDataQueueVec_12_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_12_deq_bits = _otherUnitDataQueueVec_fifo_12_empty ? otherUnitDataQueueVec_12_enq_bits : _otherUnitDataQueueVec_fifo_12_data_out;
  wire              otherUnitDataQueueVec_13_enq_ready = ~_otherUnitDataQueueVec_fifo_13_full;
  wire              otherUnitDataQueueVec_13_deq_ready;
  wire              otherUnitDataQueueVec_13_enq_valid;
  wire              otherUnitDataQueueVec_13_deq_valid = ~_otherUnitDataQueueVec_fifo_13_empty | otherUnitDataQueueVec_13_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_13_deq_bits = _otherUnitDataQueueVec_fifo_13_empty ? otherUnitDataQueueVec_13_enq_bits : _otherUnitDataQueueVec_fifo_13_data_out;
  wire              otherUnitDataQueueVec_14_enq_ready = ~_otherUnitDataQueueVec_fifo_14_full;
  wire              otherUnitDataQueueVec_14_deq_ready;
  wire              otherUnitDataQueueVec_14_enq_valid;
  wire              otherUnitDataQueueVec_14_deq_valid = ~_otherUnitDataQueueVec_fifo_14_empty | otherUnitDataQueueVec_14_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_14_deq_bits = _otherUnitDataQueueVec_fifo_14_empty ? otherUnitDataQueueVec_14_enq_bits : _otherUnitDataQueueVec_fifo_14_data_out;
  wire              otherUnitDataQueueVec_15_enq_ready = ~_otherUnitDataQueueVec_fifo_15_full;
  wire              otherUnitDataQueueVec_15_deq_ready;
  wire              otherUnitDataQueueVec_15_enq_valid;
  wire              otherUnitDataQueueVec_15_deq_valid = ~_otherUnitDataQueueVec_fifo_15_empty | otherUnitDataQueueVec_15_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_15_deq_bits = _otherUnitDataQueueVec_fifo_15_empty ? otherUnitDataQueueVec_15_enq_bits : _otherUnitDataQueueVec_fifo_15_data_out;
  wire              otherUnitDataQueueVec_16_enq_ready = ~_otherUnitDataQueueVec_fifo_16_full;
  wire              otherUnitDataQueueVec_16_deq_ready;
  wire              otherUnitDataQueueVec_16_enq_valid;
  wire              otherUnitDataQueueVec_16_deq_valid = ~_otherUnitDataQueueVec_fifo_16_empty | otherUnitDataQueueVec_16_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_16_deq_bits = _otherUnitDataQueueVec_fifo_16_empty ? otherUnitDataQueueVec_16_enq_bits : _otherUnitDataQueueVec_fifo_16_data_out;
  wire              otherUnitDataQueueVec_17_enq_ready = ~_otherUnitDataQueueVec_fifo_17_full;
  wire              otherUnitDataQueueVec_17_deq_ready;
  wire              otherUnitDataQueueVec_17_enq_valid;
  wire              otherUnitDataQueueVec_17_deq_valid = ~_otherUnitDataQueueVec_fifo_17_empty | otherUnitDataQueueVec_17_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_17_deq_bits = _otherUnitDataQueueVec_fifo_17_empty ? otherUnitDataQueueVec_17_enq_bits : _otherUnitDataQueueVec_fifo_17_data_out;
  wire              otherUnitDataQueueVec_18_enq_ready = ~_otherUnitDataQueueVec_fifo_18_full;
  wire              otherUnitDataQueueVec_18_deq_ready;
  wire              otherUnitDataQueueVec_18_enq_valid;
  wire              otherUnitDataQueueVec_18_deq_valid = ~_otherUnitDataQueueVec_fifo_18_empty | otherUnitDataQueueVec_18_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_18_deq_bits = _otherUnitDataQueueVec_fifo_18_empty ? otherUnitDataQueueVec_18_enq_bits : _otherUnitDataQueueVec_fifo_18_data_out;
  wire              otherUnitDataQueueVec_19_enq_ready = ~_otherUnitDataQueueVec_fifo_19_full;
  wire              otherUnitDataQueueVec_19_deq_ready;
  wire              otherUnitDataQueueVec_19_enq_valid;
  wire              otherUnitDataQueueVec_19_deq_valid = ~_otherUnitDataQueueVec_fifo_19_empty | otherUnitDataQueueVec_19_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_19_deq_bits = _otherUnitDataQueueVec_fifo_19_empty ? otherUnitDataQueueVec_19_enq_bits : _otherUnitDataQueueVec_fifo_19_data_out;
  wire              otherUnitDataQueueVec_20_enq_ready = ~_otherUnitDataQueueVec_fifo_20_full;
  wire              otherUnitDataQueueVec_20_deq_ready;
  wire              otherUnitDataQueueVec_20_enq_valid;
  wire              otherUnitDataQueueVec_20_deq_valid = ~_otherUnitDataQueueVec_fifo_20_empty | otherUnitDataQueueVec_20_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_20_deq_bits = _otherUnitDataQueueVec_fifo_20_empty ? otherUnitDataQueueVec_20_enq_bits : _otherUnitDataQueueVec_fifo_20_data_out;
  wire              otherUnitDataQueueVec_21_enq_ready = ~_otherUnitDataQueueVec_fifo_21_full;
  wire              otherUnitDataQueueVec_21_deq_ready;
  wire              otherUnitDataQueueVec_21_enq_valid;
  wire              otherUnitDataQueueVec_21_deq_valid = ~_otherUnitDataQueueVec_fifo_21_empty | otherUnitDataQueueVec_21_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_21_deq_bits = _otherUnitDataQueueVec_fifo_21_empty ? otherUnitDataQueueVec_21_enq_bits : _otherUnitDataQueueVec_fifo_21_data_out;
  wire              otherUnitDataQueueVec_22_enq_ready = ~_otherUnitDataQueueVec_fifo_22_full;
  wire              otherUnitDataQueueVec_22_deq_ready;
  wire              otherUnitDataQueueVec_22_enq_valid;
  wire              otherUnitDataQueueVec_22_deq_valid = ~_otherUnitDataQueueVec_fifo_22_empty | otherUnitDataQueueVec_22_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_22_deq_bits = _otherUnitDataQueueVec_fifo_22_empty ? otherUnitDataQueueVec_22_enq_bits : _otherUnitDataQueueVec_fifo_22_data_out;
  wire              otherUnitDataQueueVec_23_enq_ready = ~_otherUnitDataQueueVec_fifo_23_full;
  wire              otherUnitDataQueueVec_23_deq_ready;
  wire              otherUnitDataQueueVec_23_enq_valid;
  wire              otherUnitDataQueueVec_23_deq_valid = ~_otherUnitDataQueueVec_fifo_23_empty | otherUnitDataQueueVec_23_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_23_deq_bits = _otherUnitDataQueueVec_fifo_23_empty ? otherUnitDataQueueVec_23_enq_bits : _otherUnitDataQueueVec_fifo_23_data_out;
  wire              otherUnitDataQueueVec_24_enq_ready = ~_otherUnitDataQueueVec_fifo_24_full;
  wire              otherUnitDataQueueVec_24_deq_ready;
  wire              otherUnitDataQueueVec_24_enq_valid;
  wire              otherUnitDataQueueVec_24_deq_valid = ~_otherUnitDataQueueVec_fifo_24_empty | otherUnitDataQueueVec_24_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_24_deq_bits = _otherUnitDataQueueVec_fifo_24_empty ? otherUnitDataQueueVec_24_enq_bits : _otherUnitDataQueueVec_fifo_24_data_out;
  wire              otherUnitDataQueueVec_25_enq_ready = ~_otherUnitDataQueueVec_fifo_25_full;
  wire              otherUnitDataQueueVec_25_deq_ready;
  wire              otherUnitDataQueueVec_25_enq_valid;
  wire              otherUnitDataQueueVec_25_deq_valid = ~_otherUnitDataQueueVec_fifo_25_empty | otherUnitDataQueueVec_25_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_25_deq_bits = _otherUnitDataQueueVec_fifo_25_empty ? otherUnitDataQueueVec_25_enq_bits : _otherUnitDataQueueVec_fifo_25_data_out;
  wire              otherUnitDataQueueVec_26_enq_ready = ~_otherUnitDataQueueVec_fifo_26_full;
  wire              otherUnitDataQueueVec_26_deq_ready;
  wire              otherUnitDataQueueVec_26_enq_valid;
  wire              otherUnitDataQueueVec_26_deq_valid = ~_otherUnitDataQueueVec_fifo_26_empty | otherUnitDataQueueVec_26_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_26_deq_bits = _otherUnitDataQueueVec_fifo_26_empty ? otherUnitDataQueueVec_26_enq_bits : _otherUnitDataQueueVec_fifo_26_data_out;
  wire              otherUnitDataQueueVec_27_enq_ready = ~_otherUnitDataQueueVec_fifo_27_full;
  wire              otherUnitDataQueueVec_27_deq_ready;
  wire              otherUnitDataQueueVec_27_enq_valid;
  wire              otherUnitDataQueueVec_27_deq_valid = ~_otherUnitDataQueueVec_fifo_27_empty | otherUnitDataQueueVec_27_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_27_deq_bits = _otherUnitDataQueueVec_fifo_27_empty ? otherUnitDataQueueVec_27_enq_bits : _otherUnitDataQueueVec_fifo_27_data_out;
  wire              otherUnitDataQueueVec_28_enq_ready = ~_otherUnitDataQueueVec_fifo_28_full;
  wire              otherUnitDataQueueVec_28_deq_ready;
  wire              otherUnitDataQueueVec_28_enq_valid;
  wire              otherUnitDataQueueVec_28_deq_valid = ~_otherUnitDataQueueVec_fifo_28_empty | otherUnitDataQueueVec_28_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_28_deq_bits = _otherUnitDataQueueVec_fifo_28_empty ? otherUnitDataQueueVec_28_enq_bits : _otherUnitDataQueueVec_fifo_28_data_out;
  wire              otherUnitDataQueueVec_29_enq_ready = ~_otherUnitDataQueueVec_fifo_29_full;
  wire              otherUnitDataQueueVec_29_deq_ready;
  wire              otherUnitDataQueueVec_29_enq_valid;
  wire              otherUnitDataQueueVec_29_deq_valid = ~_otherUnitDataQueueVec_fifo_29_empty | otherUnitDataQueueVec_29_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_29_deq_bits = _otherUnitDataQueueVec_fifo_29_empty ? otherUnitDataQueueVec_29_enq_bits : _otherUnitDataQueueVec_fifo_29_data_out;
  wire              otherUnitDataQueueVec_30_enq_ready = ~_otherUnitDataQueueVec_fifo_30_full;
  wire              otherUnitDataQueueVec_30_deq_ready;
  wire              otherUnitDataQueueVec_30_enq_valid;
  wire              otherUnitDataQueueVec_30_deq_valid = ~_otherUnitDataQueueVec_fifo_30_empty | otherUnitDataQueueVec_30_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_30_deq_bits = _otherUnitDataQueueVec_fifo_30_empty ? otherUnitDataQueueVec_30_enq_bits : _otherUnitDataQueueVec_fifo_30_data_out;
  wire              otherUnitDataQueueVec_31_enq_ready = ~_otherUnitDataQueueVec_fifo_31_full;
  wire              otherUnitDataQueueVec_31_deq_ready;
  wire              otherUnitDataQueueVec_31_enq_valid;
  wire              otherUnitDataQueueVec_31_deq_valid = ~_otherUnitDataQueueVec_fifo_31_empty | otherUnitDataQueueVec_31_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_31_deq_bits = _otherUnitDataQueueVec_fifo_31_empty ? otherUnitDataQueueVec_31_enq_bits : _otherUnitDataQueueVec_fifo_31_data_out;
  wire [31:0]       otherTryReadVrf = _otherUnit_vrfReadDataPorts_valid ? _otherUnit_status_targetLane : 32'h0;
  wire              vrfReadDataPorts_0_valid_0 = otherTryReadVrf[0] | _storeUnit_vrfReadDataPorts_0_valid;
  wire [4:0]        vrfReadDataPorts_0_bits_vs_0 = otherTryReadVrf[0] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_0_bits_vs;
  wire [2:0]        vrfReadDataPorts_0_bits_instructionIndex_0 = otherTryReadVrf[0] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_0_bits_instructionIndex;
  wire              otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_0_enq_valid = vrfReadResults_0_valid & ~otherUnitTargetQueue_empty;
  wire [31:0]       dataDeqFire;
  assign otherUnitDataQueueVec_0_deq_ready = dataDeqFire[0];
  wire              vrfReadDataPorts_1_valid_0 = otherTryReadVrf[1] | _storeUnit_vrfReadDataPorts_1_valid;
  wire [4:0]        vrfReadDataPorts_1_bits_vs_0 = otherTryReadVrf[1] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_1_bits_vs;
  wire [2:0]        vrfReadDataPorts_1_bits_instructionIndex_0 = otherTryReadVrf[1] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_1_bits_instructionIndex;
  assign otherUnitDataQueueVec_1_enq_valid = vrfReadResults_1_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_1_deq_ready = dataDeqFire[1];
  wire              vrfReadDataPorts_2_valid_0 = otherTryReadVrf[2] | _storeUnit_vrfReadDataPorts_2_valid;
  wire [4:0]        vrfReadDataPorts_2_bits_vs_0 = otherTryReadVrf[2] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_2_bits_vs;
  wire [2:0]        vrfReadDataPorts_2_bits_instructionIndex_0 = otherTryReadVrf[2] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_2_bits_instructionIndex;
  assign otherUnitDataQueueVec_2_enq_valid = vrfReadResults_2_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_2_deq_ready = dataDeqFire[2];
  wire              vrfReadDataPorts_3_valid_0 = otherTryReadVrf[3] | _storeUnit_vrfReadDataPorts_3_valid;
  wire [4:0]        vrfReadDataPorts_3_bits_vs_0 = otherTryReadVrf[3] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_3_bits_vs;
  wire [2:0]        vrfReadDataPorts_3_bits_instructionIndex_0 = otherTryReadVrf[3] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_3_bits_instructionIndex;
  assign otherUnitDataQueueVec_3_enq_valid = vrfReadResults_3_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_3_deq_ready = dataDeqFire[3];
  wire              vrfReadDataPorts_4_valid_0 = otherTryReadVrf[4] | _storeUnit_vrfReadDataPorts_4_valid;
  wire [4:0]        vrfReadDataPorts_4_bits_vs_0 = otherTryReadVrf[4] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_4_bits_vs;
  wire [2:0]        vrfReadDataPorts_4_bits_instructionIndex_0 = otherTryReadVrf[4] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_4_bits_instructionIndex;
  assign otherUnitDataQueueVec_4_enq_valid = vrfReadResults_4_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_4_deq_ready = dataDeqFire[4];
  wire              vrfReadDataPorts_5_valid_0 = otherTryReadVrf[5] | _storeUnit_vrfReadDataPorts_5_valid;
  wire [4:0]        vrfReadDataPorts_5_bits_vs_0 = otherTryReadVrf[5] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_5_bits_vs;
  wire [2:0]        vrfReadDataPorts_5_bits_instructionIndex_0 = otherTryReadVrf[5] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_5_bits_instructionIndex;
  assign otherUnitDataQueueVec_5_enq_valid = vrfReadResults_5_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_5_deq_ready = dataDeqFire[5];
  wire              vrfReadDataPorts_6_valid_0 = otherTryReadVrf[6] | _storeUnit_vrfReadDataPorts_6_valid;
  wire [4:0]        vrfReadDataPorts_6_bits_vs_0 = otherTryReadVrf[6] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_6_bits_vs;
  wire [2:0]        vrfReadDataPorts_6_bits_instructionIndex_0 = otherTryReadVrf[6] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_6_bits_instructionIndex;
  assign otherUnitDataQueueVec_6_enq_valid = vrfReadResults_6_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_6_deq_ready = dataDeqFire[6];
  wire              vrfReadDataPorts_7_valid_0 = otherTryReadVrf[7] | _storeUnit_vrfReadDataPorts_7_valid;
  wire [4:0]        vrfReadDataPorts_7_bits_vs_0 = otherTryReadVrf[7] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_7_bits_vs;
  wire [2:0]        vrfReadDataPorts_7_bits_instructionIndex_0 = otherTryReadVrf[7] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_7_bits_instructionIndex;
  assign otherUnitDataQueueVec_7_enq_valid = vrfReadResults_7_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_7_deq_ready = dataDeqFire[7];
  wire              vrfReadDataPorts_8_valid_0 = otherTryReadVrf[8] | _storeUnit_vrfReadDataPorts_8_valid;
  wire [4:0]        vrfReadDataPorts_8_bits_vs_0 = otherTryReadVrf[8] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_8_bits_vs;
  wire [2:0]        vrfReadDataPorts_8_bits_instructionIndex_0 = otherTryReadVrf[8] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_8_bits_instructionIndex;
  assign otherUnitDataQueueVec_8_enq_valid = vrfReadResults_8_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_8_deq_ready = dataDeqFire[8];
  wire              vrfReadDataPorts_9_valid_0 = otherTryReadVrf[9] | _storeUnit_vrfReadDataPorts_9_valid;
  wire [4:0]        vrfReadDataPorts_9_bits_vs_0 = otherTryReadVrf[9] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_9_bits_vs;
  wire [2:0]        vrfReadDataPorts_9_bits_instructionIndex_0 = otherTryReadVrf[9] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_9_bits_instructionIndex;
  assign otherUnitDataQueueVec_9_enq_valid = vrfReadResults_9_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_9_deq_ready = dataDeqFire[9];
  wire              vrfReadDataPorts_10_valid_0 = otherTryReadVrf[10] | _storeUnit_vrfReadDataPorts_10_valid;
  wire [4:0]        vrfReadDataPorts_10_bits_vs_0 = otherTryReadVrf[10] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_10_bits_vs;
  wire [2:0]        vrfReadDataPorts_10_bits_instructionIndex_0 = otherTryReadVrf[10] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_10_bits_instructionIndex;
  assign otherUnitDataQueueVec_10_enq_valid = vrfReadResults_10_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_10_deq_ready = dataDeqFire[10];
  wire              vrfReadDataPorts_11_valid_0 = otherTryReadVrf[11] | _storeUnit_vrfReadDataPorts_11_valid;
  wire [4:0]        vrfReadDataPorts_11_bits_vs_0 = otherTryReadVrf[11] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_11_bits_vs;
  wire [2:0]        vrfReadDataPorts_11_bits_instructionIndex_0 = otherTryReadVrf[11] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_11_bits_instructionIndex;
  assign otherUnitDataQueueVec_11_enq_valid = vrfReadResults_11_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_11_deq_ready = dataDeqFire[11];
  wire              vrfReadDataPorts_12_valid_0 = otherTryReadVrf[12] | _storeUnit_vrfReadDataPorts_12_valid;
  wire [4:0]        vrfReadDataPorts_12_bits_vs_0 = otherTryReadVrf[12] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_12_bits_vs;
  wire [2:0]        vrfReadDataPorts_12_bits_instructionIndex_0 = otherTryReadVrf[12] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_12_bits_instructionIndex;
  assign otherUnitDataQueueVec_12_enq_valid = vrfReadResults_12_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_12_deq_ready = dataDeqFire[12];
  wire              vrfReadDataPorts_13_valid_0 = otherTryReadVrf[13] | _storeUnit_vrfReadDataPorts_13_valid;
  wire [4:0]        vrfReadDataPorts_13_bits_vs_0 = otherTryReadVrf[13] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_13_bits_vs;
  wire [2:0]        vrfReadDataPorts_13_bits_instructionIndex_0 = otherTryReadVrf[13] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_13_bits_instructionIndex;
  assign otherUnitDataQueueVec_13_enq_valid = vrfReadResults_13_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_13_deq_ready = dataDeqFire[13];
  wire              vrfReadDataPorts_14_valid_0 = otherTryReadVrf[14] | _storeUnit_vrfReadDataPorts_14_valid;
  wire [4:0]        vrfReadDataPorts_14_bits_vs_0 = otherTryReadVrf[14] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_14_bits_vs;
  wire [2:0]        vrfReadDataPorts_14_bits_instructionIndex_0 = otherTryReadVrf[14] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_14_bits_instructionIndex;
  assign otherUnitDataQueueVec_14_enq_valid = vrfReadResults_14_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_14_deq_ready = dataDeqFire[14];
  wire              vrfReadDataPorts_15_valid_0 = otherTryReadVrf[15] | _storeUnit_vrfReadDataPorts_15_valid;
  wire [4:0]        vrfReadDataPorts_15_bits_vs_0 = otherTryReadVrf[15] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_15_bits_vs;
  wire [2:0]        vrfReadDataPorts_15_bits_instructionIndex_0 = otherTryReadVrf[15] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_15_bits_instructionIndex;
  assign otherUnitDataQueueVec_15_enq_valid = vrfReadResults_15_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_15_deq_ready = dataDeqFire[15];
  wire              vrfReadDataPorts_16_valid_0 = otherTryReadVrf[16] | _storeUnit_vrfReadDataPorts_16_valid;
  wire [4:0]        vrfReadDataPorts_16_bits_vs_0 = otherTryReadVrf[16] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_16_bits_vs;
  wire [2:0]        vrfReadDataPorts_16_bits_instructionIndex_0 = otherTryReadVrf[16] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_16_bits_instructionIndex;
  assign otherUnitDataQueueVec_16_enq_valid = vrfReadResults_16_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_16_deq_ready = dataDeqFire[16];
  wire              vrfReadDataPorts_17_valid_0 = otherTryReadVrf[17] | _storeUnit_vrfReadDataPorts_17_valid;
  wire [4:0]        vrfReadDataPorts_17_bits_vs_0 = otherTryReadVrf[17] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_17_bits_vs;
  wire [2:0]        vrfReadDataPorts_17_bits_instructionIndex_0 = otherTryReadVrf[17] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_17_bits_instructionIndex;
  assign otherUnitDataQueueVec_17_enq_valid = vrfReadResults_17_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_17_deq_ready = dataDeqFire[17];
  wire              vrfReadDataPorts_18_valid_0 = otherTryReadVrf[18] | _storeUnit_vrfReadDataPorts_18_valid;
  wire [4:0]        vrfReadDataPorts_18_bits_vs_0 = otherTryReadVrf[18] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_18_bits_vs;
  wire [2:0]        vrfReadDataPorts_18_bits_instructionIndex_0 = otherTryReadVrf[18] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_18_bits_instructionIndex;
  assign otherUnitDataQueueVec_18_enq_valid = vrfReadResults_18_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_18_deq_ready = dataDeqFire[18];
  wire              vrfReadDataPorts_19_valid_0 = otherTryReadVrf[19] | _storeUnit_vrfReadDataPorts_19_valid;
  wire [4:0]        vrfReadDataPorts_19_bits_vs_0 = otherTryReadVrf[19] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_19_bits_vs;
  wire [2:0]        vrfReadDataPorts_19_bits_instructionIndex_0 = otherTryReadVrf[19] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_19_bits_instructionIndex;
  assign otherUnitDataQueueVec_19_enq_valid = vrfReadResults_19_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_19_deq_ready = dataDeqFire[19];
  wire              vrfReadDataPorts_20_valid_0 = otherTryReadVrf[20] | _storeUnit_vrfReadDataPorts_20_valid;
  wire [4:0]        vrfReadDataPorts_20_bits_vs_0 = otherTryReadVrf[20] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_20_bits_vs;
  wire [2:0]        vrfReadDataPorts_20_bits_instructionIndex_0 = otherTryReadVrf[20] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_20_bits_instructionIndex;
  assign otherUnitDataQueueVec_20_enq_valid = vrfReadResults_20_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_20_deq_ready = dataDeqFire[20];
  wire              vrfReadDataPorts_21_valid_0 = otherTryReadVrf[21] | _storeUnit_vrfReadDataPorts_21_valid;
  wire [4:0]        vrfReadDataPorts_21_bits_vs_0 = otherTryReadVrf[21] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_21_bits_vs;
  wire [2:0]        vrfReadDataPorts_21_bits_instructionIndex_0 = otherTryReadVrf[21] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_21_bits_instructionIndex;
  assign otherUnitDataQueueVec_21_enq_valid = vrfReadResults_21_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_21_deq_ready = dataDeqFire[21];
  wire              vrfReadDataPorts_22_valid_0 = otherTryReadVrf[22] | _storeUnit_vrfReadDataPorts_22_valid;
  wire [4:0]        vrfReadDataPorts_22_bits_vs_0 = otherTryReadVrf[22] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_22_bits_vs;
  wire [2:0]        vrfReadDataPorts_22_bits_instructionIndex_0 = otherTryReadVrf[22] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_22_bits_instructionIndex;
  assign otherUnitDataQueueVec_22_enq_valid = vrfReadResults_22_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_22_deq_ready = dataDeqFire[22];
  wire              vrfReadDataPorts_23_valid_0 = otherTryReadVrf[23] | _storeUnit_vrfReadDataPorts_23_valid;
  wire [4:0]        vrfReadDataPorts_23_bits_vs_0 = otherTryReadVrf[23] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_23_bits_vs;
  wire [2:0]        vrfReadDataPorts_23_bits_instructionIndex_0 = otherTryReadVrf[23] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_23_bits_instructionIndex;
  assign otherUnitDataQueueVec_23_enq_valid = vrfReadResults_23_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_23_deq_ready = dataDeqFire[23];
  wire              vrfReadDataPorts_24_valid_0 = otherTryReadVrf[24] | _storeUnit_vrfReadDataPorts_24_valid;
  wire [4:0]        vrfReadDataPorts_24_bits_vs_0 = otherTryReadVrf[24] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_24_bits_vs;
  wire [2:0]        vrfReadDataPorts_24_bits_instructionIndex_0 = otherTryReadVrf[24] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_24_bits_instructionIndex;
  assign otherUnitDataQueueVec_24_enq_valid = vrfReadResults_24_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_24_deq_ready = dataDeqFire[24];
  wire              vrfReadDataPorts_25_valid_0 = otherTryReadVrf[25] | _storeUnit_vrfReadDataPorts_25_valid;
  wire [4:0]        vrfReadDataPorts_25_bits_vs_0 = otherTryReadVrf[25] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_25_bits_vs;
  wire [2:0]        vrfReadDataPorts_25_bits_instructionIndex_0 = otherTryReadVrf[25] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_25_bits_instructionIndex;
  assign otherUnitDataQueueVec_25_enq_valid = vrfReadResults_25_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_25_deq_ready = dataDeqFire[25];
  wire              vrfReadDataPorts_26_valid_0 = otherTryReadVrf[26] | _storeUnit_vrfReadDataPorts_26_valid;
  wire [4:0]        vrfReadDataPorts_26_bits_vs_0 = otherTryReadVrf[26] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_26_bits_vs;
  wire [2:0]        vrfReadDataPorts_26_bits_instructionIndex_0 = otherTryReadVrf[26] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_26_bits_instructionIndex;
  assign otherUnitDataQueueVec_26_enq_valid = vrfReadResults_26_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_26_deq_ready = dataDeqFire[26];
  wire              vrfReadDataPorts_27_valid_0 = otherTryReadVrf[27] | _storeUnit_vrfReadDataPorts_27_valid;
  wire [4:0]        vrfReadDataPorts_27_bits_vs_0 = otherTryReadVrf[27] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_27_bits_vs;
  wire [2:0]        vrfReadDataPorts_27_bits_instructionIndex_0 = otherTryReadVrf[27] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_27_bits_instructionIndex;
  assign otherUnitDataQueueVec_27_enq_valid = vrfReadResults_27_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_27_deq_ready = dataDeqFire[27];
  wire              vrfReadDataPorts_28_valid_0 = otherTryReadVrf[28] | _storeUnit_vrfReadDataPorts_28_valid;
  wire [4:0]        vrfReadDataPorts_28_bits_vs_0 = otherTryReadVrf[28] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_28_bits_vs;
  wire [2:0]        vrfReadDataPorts_28_bits_instructionIndex_0 = otherTryReadVrf[28] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_28_bits_instructionIndex;
  assign otherUnitDataQueueVec_28_enq_valid = vrfReadResults_28_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_28_deq_ready = dataDeqFire[28];
  wire              vrfReadDataPorts_29_valid_0 = otherTryReadVrf[29] | _storeUnit_vrfReadDataPorts_29_valid;
  wire [4:0]        vrfReadDataPorts_29_bits_vs_0 = otherTryReadVrf[29] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_29_bits_vs;
  wire [2:0]        vrfReadDataPorts_29_bits_instructionIndex_0 = otherTryReadVrf[29] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_29_bits_instructionIndex;
  assign otherUnitDataQueueVec_29_enq_valid = vrfReadResults_29_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_29_deq_ready = dataDeqFire[29];
  wire              vrfReadDataPorts_30_valid_0 = otherTryReadVrf[30] | _storeUnit_vrfReadDataPorts_30_valid;
  wire [4:0]        vrfReadDataPorts_30_bits_vs_0 = otherTryReadVrf[30] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_30_bits_vs;
  wire [2:0]        vrfReadDataPorts_30_bits_instructionIndex_0 = otherTryReadVrf[30] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_30_bits_instructionIndex;
  assign otherUnitDataQueueVec_30_enq_valid = vrfReadResults_30_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_30_deq_ready = dataDeqFire[30];
  wire              vrfReadDataPorts_31_valid_0 = otherTryReadVrf[31] | _storeUnit_vrfReadDataPorts_31_valid;
  wire [4:0]        vrfReadDataPorts_31_bits_vs_0 = otherTryReadVrf[31] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_31_bits_vs;
  wire [2:0]        vrfReadDataPorts_31_bits_instructionIndex_0 = otherTryReadVrf[31] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_31_bits_instructionIndex;
  assign otherUnitDataQueueVec_31_enq_valid = vrfReadResults_31_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_31_deq_ready = dataDeqFire[31];
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_lo_lo_lo_lo = {vrfReadDataPorts_1_ready_0, vrfReadDataPorts_0_ready_0};
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_lo_lo_lo_hi = {vrfReadDataPorts_3_ready_0, vrfReadDataPorts_2_ready_0};
  wire [3:0]        otherUnit_vrfReadDataPorts_ready_lo_lo_lo = {otherUnit_vrfReadDataPorts_ready_lo_lo_lo_hi, otherUnit_vrfReadDataPorts_ready_lo_lo_lo_lo};
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_lo_lo_hi_lo = {vrfReadDataPorts_5_ready_0, vrfReadDataPorts_4_ready_0};
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_lo_lo_hi_hi = {vrfReadDataPorts_7_ready_0, vrfReadDataPorts_6_ready_0};
  wire [3:0]        otherUnit_vrfReadDataPorts_ready_lo_lo_hi = {otherUnit_vrfReadDataPorts_ready_lo_lo_hi_hi, otherUnit_vrfReadDataPorts_ready_lo_lo_hi_lo};
  wire [7:0]        otherUnit_vrfReadDataPorts_ready_lo_lo = {otherUnit_vrfReadDataPorts_ready_lo_lo_hi, otherUnit_vrfReadDataPorts_ready_lo_lo_lo};
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_lo_hi_lo_lo = {vrfReadDataPorts_9_ready_0, vrfReadDataPorts_8_ready_0};
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_lo_hi_lo_hi = {vrfReadDataPorts_11_ready_0, vrfReadDataPorts_10_ready_0};
  wire [3:0]        otherUnit_vrfReadDataPorts_ready_lo_hi_lo = {otherUnit_vrfReadDataPorts_ready_lo_hi_lo_hi, otherUnit_vrfReadDataPorts_ready_lo_hi_lo_lo};
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_lo_hi_hi_lo = {vrfReadDataPorts_13_ready_0, vrfReadDataPorts_12_ready_0};
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_lo_hi_hi_hi = {vrfReadDataPorts_15_ready_0, vrfReadDataPorts_14_ready_0};
  wire [3:0]        otherUnit_vrfReadDataPorts_ready_lo_hi_hi = {otherUnit_vrfReadDataPorts_ready_lo_hi_hi_hi, otherUnit_vrfReadDataPorts_ready_lo_hi_hi_lo};
  wire [7:0]        otherUnit_vrfReadDataPorts_ready_lo_hi = {otherUnit_vrfReadDataPorts_ready_lo_hi_hi, otherUnit_vrfReadDataPorts_ready_lo_hi_lo};
  wire [15:0]       otherUnit_vrfReadDataPorts_ready_lo = {otherUnit_vrfReadDataPorts_ready_lo_hi, otherUnit_vrfReadDataPorts_ready_lo_lo};
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_hi_lo_lo_lo = {vrfReadDataPorts_17_ready_0, vrfReadDataPorts_16_ready_0};
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_hi_lo_lo_hi = {vrfReadDataPorts_19_ready_0, vrfReadDataPorts_18_ready_0};
  wire [3:0]        otherUnit_vrfReadDataPorts_ready_hi_lo_lo = {otherUnit_vrfReadDataPorts_ready_hi_lo_lo_hi, otherUnit_vrfReadDataPorts_ready_hi_lo_lo_lo};
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_hi_lo_hi_lo = {vrfReadDataPorts_21_ready_0, vrfReadDataPorts_20_ready_0};
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_hi_lo_hi_hi = {vrfReadDataPorts_23_ready_0, vrfReadDataPorts_22_ready_0};
  wire [3:0]        otherUnit_vrfReadDataPorts_ready_hi_lo_hi = {otherUnit_vrfReadDataPorts_ready_hi_lo_hi_hi, otherUnit_vrfReadDataPorts_ready_hi_lo_hi_lo};
  wire [7:0]        otherUnit_vrfReadDataPorts_ready_hi_lo = {otherUnit_vrfReadDataPorts_ready_hi_lo_hi, otherUnit_vrfReadDataPorts_ready_hi_lo_lo};
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_hi_hi_lo_lo = {vrfReadDataPorts_25_ready_0, vrfReadDataPorts_24_ready_0};
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_hi_hi_lo_hi = {vrfReadDataPorts_27_ready_0, vrfReadDataPorts_26_ready_0};
  wire [3:0]        otherUnit_vrfReadDataPorts_ready_hi_hi_lo = {otherUnit_vrfReadDataPorts_ready_hi_hi_lo_hi, otherUnit_vrfReadDataPorts_ready_hi_hi_lo_lo};
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_hi_hi_hi_lo = {vrfReadDataPorts_29_ready_0, vrfReadDataPorts_28_ready_0};
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_hi_hi_hi_hi = {vrfReadDataPorts_31_ready_0, vrfReadDataPorts_30_ready_0};
  wire [3:0]        otherUnit_vrfReadDataPorts_ready_hi_hi_hi = {otherUnit_vrfReadDataPorts_ready_hi_hi_hi_hi, otherUnit_vrfReadDataPorts_ready_hi_hi_hi_lo};
  wire [7:0]        otherUnit_vrfReadDataPorts_ready_hi_hi = {otherUnit_vrfReadDataPorts_ready_hi_hi_hi, otherUnit_vrfReadDataPorts_ready_hi_hi_lo};
  wire [15:0]       otherUnit_vrfReadDataPorts_ready_hi = {otherUnit_vrfReadDataPorts_ready_hi_hi, otherUnit_vrfReadDataPorts_ready_hi_lo};
  wire              otherUnit_vrfReadDataPorts_ready = (|(otherTryReadVrf & {otherUnit_vrfReadDataPorts_ready_hi, otherUnit_vrfReadDataPorts_ready_lo})) & otherUnitTargetQueue_enq_ready;
  assign otherUnitTargetQueue_enq_valid = otherUnit_vrfReadDataPorts_ready & _otherUnit_vrfReadDataPorts_valid;
  wire [31:0]       otherUnitTargetQueue_deq_bits;
  wire [1:0]        otherUnit_vrfReadResults_valid_lo_lo_lo_lo = {otherUnitDataQueueVec_1_deq_valid, otherUnitDataQueueVec_0_deq_valid};
  wire [1:0]        otherUnit_vrfReadResults_valid_lo_lo_lo_hi = {otherUnitDataQueueVec_3_deq_valid, otherUnitDataQueueVec_2_deq_valid};
  wire [3:0]        otherUnit_vrfReadResults_valid_lo_lo_lo = {otherUnit_vrfReadResults_valid_lo_lo_lo_hi, otherUnit_vrfReadResults_valid_lo_lo_lo_lo};
  wire [1:0]        otherUnit_vrfReadResults_valid_lo_lo_hi_lo = {otherUnitDataQueueVec_5_deq_valid, otherUnitDataQueueVec_4_deq_valid};
  wire [1:0]        otherUnit_vrfReadResults_valid_lo_lo_hi_hi = {otherUnitDataQueueVec_7_deq_valid, otherUnitDataQueueVec_6_deq_valid};
  wire [3:0]        otherUnit_vrfReadResults_valid_lo_lo_hi = {otherUnit_vrfReadResults_valid_lo_lo_hi_hi, otherUnit_vrfReadResults_valid_lo_lo_hi_lo};
  wire [7:0]        otherUnit_vrfReadResults_valid_lo_lo = {otherUnit_vrfReadResults_valid_lo_lo_hi, otherUnit_vrfReadResults_valid_lo_lo_lo};
  wire [1:0]        otherUnit_vrfReadResults_valid_lo_hi_lo_lo = {otherUnitDataQueueVec_9_deq_valid, otherUnitDataQueueVec_8_deq_valid};
  wire [1:0]        otherUnit_vrfReadResults_valid_lo_hi_lo_hi = {otherUnitDataQueueVec_11_deq_valid, otherUnitDataQueueVec_10_deq_valid};
  wire [3:0]        otherUnit_vrfReadResults_valid_lo_hi_lo = {otherUnit_vrfReadResults_valid_lo_hi_lo_hi, otherUnit_vrfReadResults_valid_lo_hi_lo_lo};
  wire [1:0]        otherUnit_vrfReadResults_valid_lo_hi_hi_lo = {otherUnitDataQueueVec_13_deq_valid, otherUnitDataQueueVec_12_deq_valid};
  wire [1:0]        otherUnit_vrfReadResults_valid_lo_hi_hi_hi = {otherUnitDataQueueVec_15_deq_valid, otherUnitDataQueueVec_14_deq_valid};
  wire [3:0]        otherUnit_vrfReadResults_valid_lo_hi_hi = {otherUnit_vrfReadResults_valid_lo_hi_hi_hi, otherUnit_vrfReadResults_valid_lo_hi_hi_lo};
  wire [7:0]        otherUnit_vrfReadResults_valid_lo_hi = {otherUnit_vrfReadResults_valid_lo_hi_hi, otherUnit_vrfReadResults_valid_lo_hi_lo};
  wire [15:0]       otherUnit_vrfReadResults_valid_lo = {otherUnit_vrfReadResults_valid_lo_hi, otherUnit_vrfReadResults_valid_lo_lo};
  wire [1:0]        otherUnit_vrfReadResults_valid_hi_lo_lo_lo = {otherUnitDataQueueVec_17_deq_valid, otherUnitDataQueueVec_16_deq_valid};
  wire [1:0]        otherUnit_vrfReadResults_valid_hi_lo_lo_hi = {otherUnitDataQueueVec_19_deq_valid, otherUnitDataQueueVec_18_deq_valid};
  wire [3:0]        otherUnit_vrfReadResults_valid_hi_lo_lo = {otherUnit_vrfReadResults_valid_hi_lo_lo_hi, otherUnit_vrfReadResults_valid_hi_lo_lo_lo};
  wire [1:0]        otherUnit_vrfReadResults_valid_hi_lo_hi_lo = {otherUnitDataQueueVec_21_deq_valid, otherUnitDataQueueVec_20_deq_valid};
  wire [1:0]        otherUnit_vrfReadResults_valid_hi_lo_hi_hi = {otherUnitDataQueueVec_23_deq_valid, otherUnitDataQueueVec_22_deq_valid};
  wire [3:0]        otherUnit_vrfReadResults_valid_hi_lo_hi = {otherUnit_vrfReadResults_valid_hi_lo_hi_hi, otherUnit_vrfReadResults_valid_hi_lo_hi_lo};
  wire [7:0]        otherUnit_vrfReadResults_valid_hi_lo = {otherUnit_vrfReadResults_valid_hi_lo_hi, otherUnit_vrfReadResults_valid_hi_lo_lo};
  wire [1:0]        otherUnit_vrfReadResults_valid_hi_hi_lo_lo = {otherUnitDataQueueVec_25_deq_valid, otherUnitDataQueueVec_24_deq_valid};
  wire [1:0]        otherUnit_vrfReadResults_valid_hi_hi_lo_hi = {otherUnitDataQueueVec_27_deq_valid, otherUnitDataQueueVec_26_deq_valid};
  wire [3:0]        otherUnit_vrfReadResults_valid_hi_hi_lo = {otherUnit_vrfReadResults_valid_hi_hi_lo_hi, otherUnit_vrfReadResults_valid_hi_hi_lo_lo};
  wire [1:0]        otherUnit_vrfReadResults_valid_hi_hi_hi_lo = {otherUnitDataQueueVec_29_deq_valid, otherUnitDataQueueVec_28_deq_valid};
  wire [1:0]        otherUnit_vrfReadResults_valid_hi_hi_hi_hi = {otherUnitDataQueueVec_31_deq_valid, otherUnitDataQueueVec_30_deq_valid};
  wire [3:0]        otherUnit_vrfReadResults_valid_hi_hi_hi = {otherUnit_vrfReadResults_valid_hi_hi_hi_hi, otherUnit_vrfReadResults_valid_hi_hi_hi_lo};
  wire [7:0]        otherUnit_vrfReadResults_valid_hi_hi = {otherUnit_vrfReadResults_valid_hi_hi_hi, otherUnit_vrfReadResults_valid_hi_hi_lo};
  wire [15:0]       otherUnit_vrfReadResults_valid_hi = {otherUnit_vrfReadResults_valid_hi_hi, otherUnit_vrfReadResults_valid_hi_lo};
  assign otherUnitTargetQueue_deq_ready = otherUnitTargetQueue_deq_valid & (|(otherUnitTargetQueue_deq_bits & {otherUnit_vrfReadResults_valid_hi, otherUnit_vrfReadResults_valid_lo}));
  assign dataDeqFire = otherUnitTargetQueue_deq_ready ? otherUnitTargetQueue_deq_bits : 32'h0;
  wire [31:0]       otherTryToWrite = _otherUnit_vrfWritePort_valid ? _otherUnit_status_targetLane : 32'h0;
  wire [1:0]        otherUnit_vrfWritePort_ready_lo_lo_lo_lo = {writeQueueVec_1_enq_ready, writeQueueVec_0_enq_ready};
  wire [1:0]        otherUnit_vrfWritePort_ready_lo_lo_lo_hi = {writeQueueVec_3_enq_ready, writeQueueVec_2_enq_ready};
  wire [3:0]        otherUnit_vrfWritePort_ready_lo_lo_lo = {otherUnit_vrfWritePort_ready_lo_lo_lo_hi, otherUnit_vrfWritePort_ready_lo_lo_lo_lo};
  wire [1:0]        otherUnit_vrfWritePort_ready_lo_lo_hi_lo = {writeQueueVec_5_enq_ready, writeQueueVec_4_enq_ready};
  wire [1:0]        otherUnit_vrfWritePort_ready_lo_lo_hi_hi = {writeQueueVec_7_enq_ready, writeQueueVec_6_enq_ready};
  wire [3:0]        otherUnit_vrfWritePort_ready_lo_lo_hi = {otherUnit_vrfWritePort_ready_lo_lo_hi_hi, otherUnit_vrfWritePort_ready_lo_lo_hi_lo};
  wire [7:0]        otherUnit_vrfWritePort_ready_lo_lo = {otherUnit_vrfWritePort_ready_lo_lo_hi, otherUnit_vrfWritePort_ready_lo_lo_lo};
  wire [1:0]        otherUnit_vrfWritePort_ready_lo_hi_lo_lo = {writeQueueVec_9_enq_ready, writeQueueVec_8_enq_ready};
  wire [1:0]        otherUnit_vrfWritePort_ready_lo_hi_lo_hi = {writeQueueVec_11_enq_ready, writeQueueVec_10_enq_ready};
  wire [3:0]        otherUnit_vrfWritePort_ready_lo_hi_lo = {otherUnit_vrfWritePort_ready_lo_hi_lo_hi, otherUnit_vrfWritePort_ready_lo_hi_lo_lo};
  wire [1:0]        otherUnit_vrfWritePort_ready_lo_hi_hi_lo = {writeQueueVec_13_enq_ready, writeQueueVec_12_enq_ready};
  wire [1:0]        otherUnit_vrfWritePort_ready_lo_hi_hi_hi = {writeQueueVec_15_enq_ready, writeQueueVec_14_enq_ready};
  wire [3:0]        otherUnit_vrfWritePort_ready_lo_hi_hi = {otherUnit_vrfWritePort_ready_lo_hi_hi_hi, otherUnit_vrfWritePort_ready_lo_hi_hi_lo};
  wire [7:0]        otherUnit_vrfWritePort_ready_lo_hi = {otherUnit_vrfWritePort_ready_lo_hi_hi, otherUnit_vrfWritePort_ready_lo_hi_lo};
  wire [15:0]       otherUnit_vrfWritePort_ready_lo = {otherUnit_vrfWritePort_ready_lo_hi, otherUnit_vrfWritePort_ready_lo_lo};
  wire [1:0]        otherUnit_vrfWritePort_ready_hi_lo_lo_lo = {writeQueueVec_17_enq_ready, writeQueueVec_16_enq_ready};
  wire [1:0]        otherUnit_vrfWritePort_ready_hi_lo_lo_hi = {writeQueueVec_19_enq_ready, writeQueueVec_18_enq_ready};
  wire [3:0]        otherUnit_vrfWritePort_ready_hi_lo_lo = {otherUnit_vrfWritePort_ready_hi_lo_lo_hi, otherUnit_vrfWritePort_ready_hi_lo_lo_lo};
  wire [1:0]        otherUnit_vrfWritePort_ready_hi_lo_hi_lo = {writeQueueVec_21_enq_ready, writeQueueVec_20_enq_ready};
  wire [1:0]        otherUnit_vrfWritePort_ready_hi_lo_hi_hi = {writeQueueVec_23_enq_ready, writeQueueVec_22_enq_ready};
  wire [3:0]        otherUnit_vrfWritePort_ready_hi_lo_hi = {otherUnit_vrfWritePort_ready_hi_lo_hi_hi, otherUnit_vrfWritePort_ready_hi_lo_hi_lo};
  wire [7:0]        otherUnit_vrfWritePort_ready_hi_lo = {otherUnit_vrfWritePort_ready_hi_lo_hi, otherUnit_vrfWritePort_ready_hi_lo_lo};
  wire [1:0]        otherUnit_vrfWritePort_ready_hi_hi_lo_lo = {writeQueueVec_25_enq_ready, writeQueueVec_24_enq_ready};
  wire [1:0]        otherUnit_vrfWritePort_ready_hi_hi_lo_hi = {writeQueueVec_27_enq_ready, writeQueueVec_26_enq_ready};
  wire [3:0]        otherUnit_vrfWritePort_ready_hi_hi_lo = {otherUnit_vrfWritePort_ready_hi_hi_lo_hi, otherUnit_vrfWritePort_ready_hi_hi_lo_lo};
  wire [1:0]        otherUnit_vrfWritePort_ready_hi_hi_hi_lo = {writeQueueVec_29_enq_ready, writeQueueVec_28_enq_ready};
  wire [1:0]        otherUnit_vrfWritePort_ready_hi_hi_hi_hi = {writeQueueVec_31_enq_ready, writeQueueVec_30_enq_ready};
  wire [3:0]        otherUnit_vrfWritePort_ready_hi_hi_hi = {otherUnit_vrfWritePort_ready_hi_hi_hi_hi, otherUnit_vrfWritePort_ready_hi_hi_hi_lo};
  wire [7:0]        otherUnit_vrfWritePort_ready_hi_hi = {otherUnit_vrfWritePort_ready_hi_hi_hi, otherUnit_vrfWritePort_ready_hi_hi_lo};
  wire [15:0]       otherUnit_vrfWritePort_ready_hi = {otherUnit_vrfWritePort_ready_hi_hi, otherUnit_vrfWritePort_ready_hi_lo};
  assign writeQueueVec_0_enq_valid = otherTryToWrite[0] | _loadUnit_vrfWritePort_0_valid;
  assign writeQueueVec_0_enq_bits_data_vd = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_0_bits_vd;
  assign writeQueueVec_0_enq_bits_data_mask = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_0_bits_mask;
  assign writeQueueVec_0_enq_bits_data_data = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_0_bits_data;
  assign writeQueueVec_0_enq_bits_data_last = otherTryToWrite[0] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_0_enq_bits_data_instructionIndex = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_0_bits_instructionIndex;
  assign writeQueueVec_1_enq_valid = otherTryToWrite[1] | _loadUnit_vrfWritePort_1_valid;
  assign writeQueueVec_1_enq_bits_data_vd = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_1_bits_vd;
  assign writeQueueVec_1_enq_bits_data_mask = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_1_bits_mask;
  assign writeQueueVec_1_enq_bits_data_data = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_1_bits_data;
  assign writeQueueVec_1_enq_bits_data_last = otherTryToWrite[1] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_1_enq_bits_data_instructionIndex = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_1_bits_instructionIndex;
  assign writeQueueVec_2_enq_valid = otherTryToWrite[2] | _loadUnit_vrfWritePort_2_valid;
  assign writeQueueVec_2_enq_bits_data_vd = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_2_bits_vd;
  assign writeQueueVec_2_enq_bits_data_mask = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_2_bits_mask;
  assign writeQueueVec_2_enq_bits_data_data = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_2_bits_data;
  assign writeQueueVec_2_enq_bits_data_last = otherTryToWrite[2] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_2_enq_bits_data_instructionIndex = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_2_bits_instructionIndex;
  assign writeQueueVec_3_enq_valid = otherTryToWrite[3] | _loadUnit_vrfWritePort_3_valid;
  assign writeQueueVec_3_enq_bits_data_vd = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_3_bits_vd;
  assign writeQueueVec_3_enq_bits_data_mask = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_3_bits_mask;
  assign writeQueueVec_3_enq_bits_data_data = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_3_bits_data;
  assign writeQueueVec_3_enq_bits_data_last = otherTryToWrite[3] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_3_enq_bits_data_instructionIndex = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_3_bits_instructionIndex;
  assign writeQueueVec_4_enq_valid = otherTryToWrite[4] | _loadUnit_vrfWritePort_4_valid;
  assign writeQueueVec_4_enq_bits_data_vd = otherTryToWrite[4] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_4_bits_vd;
  assign writeQueueVec_4_enq_bits_data_mask = otherTryToWrite[4] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_4_bits_mask;
  assign writeQueueVec_4_enq_bits_data_data = otherTryToWrite[4] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_4_bits_data;
  assign writeQueueVec_4_enq_bits_data_last = otherTryToWrite[4] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_4_enq_bits_data_instructionIndex = otherTryToWrite[4] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_4_bits_instructionIndex;
  assign writeQueueVec_5_enq_valid = otherTryToWrite[5] | _loadUnit_vrfWritePort_5_valid;
  assign writeQueueVec_5_enq_bits_data_vd = otherTryToWrite[5] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_5_bits_vd;
  assign writeQueueVec_5_enq_bits_data_mask = otherTryToWrite[5] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_5_bits_mask;
  assign writeQueueVec_5_enq_bits_data_data = otherTryToWrite[5] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_5_bits_data;
  assign writeQueueVec_5_enq_bits_data_last = otherTryToWrite[5] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_5_enq_bits_data_instructionIndex = otherTryToWrite[5] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_5_bits_instructionIndex;
  assign writeQueueVec_6_enq_valid = otherTryToWrite[6] | _loadUnit_vrfWritePort_6_valid;
  assign writeQueueVec_6_enq_bits_data_vd = otherTryToWrite[6] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_6_bits_vd;
  assign writeQueueVec_6_enq_bits_data_mask = otherTryToWrite[6] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_6_bits_mask;
  assign writeQueueVec_6_enq_bits_data_data = otherTryToWrite[6] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_6_bits_data;
  assign writeQueueVec_6_enq_bits_data_last = otherTryToWrite[6] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_6_enq_bits_data_instructionIndex = otherTryToWrite[6] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_6_bits_instructionIndex;
  assign writeQueueVec_7_enq_valid = otherTryToWrite[7] | _loadUnit_vrfWritePort_7_valid;
  assign writeQueueVec_7_enq_bits_data_vd = otherTryToWrite[7] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_7_bits_vd;
  assign writeQueueVec_7_enq_bits_data_mask = otherTryToWrite[7] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_7_bits_mask;
  assign writeQueueVec_7_enq_bits_data_data = otherTryToWrite[7] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_7_bits_data;
  assign writeQueueVec_7_enq_bits_data_last = otherTryToWrite[7] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_7_enq_bits_data_instructionIndex = otherTryToWrite[7] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_7_bits_instructionIndex;
  assign writeQueueVec_8_enq_valid = otherTryToWrite[8] | _loadUnit_vrfWritePort_8_valid;
  assign writeQueueVec_8_enq_bits_data_vd = otherTryToWrite[8] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_8_bits_vd;
  assign writeQueueVec_8_enq_bits_data_mask = otherTryToWrite[8] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_8_bits_mask;
  assign writeQueueVec_8_enq_bits_data_data = otherTryToWrite[8] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_8_bits_data;
  assign writeQueueVec_8_enq_bits_data_last = otherTryToWrite[8] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_8_enq_bits_data_instructionIndex = otherTryToWrite[8] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_8_bits_instructionIndex;
  assign writeQueueVec_9_enq_valid = otherTryToWrite[9] | _loadUnit_vrfWritePort_9_valid;
  assign writeQueueVec_9_enq_bits_data_vd = otherTryToWrite[9] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_9_bits_vd;
  assign writeQueueVec_9_enq_bits_data_mask = otherTryToWrite[9] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_9_bits_mask;
  assign writeQueueVec_9_enq_bits_data_data = otherTryToWrite[9] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_9_bits_data;
  assign writeQueueVec_9_enq_bits_data_last = otherTryToWrite[9] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_9_enq_bits_data_instructionIndex = otherTryToWrite[9] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_9_bits_instructionIndex;
  assign writeQueueVec_10_enq_valid = otherTryToWrite[10] | _loadUnit_vrfWritePort_10_valid;
  assign writeQueueVec_10_enq_bits_data_vd = otherTryToWrite[10] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_10_bits_vd;
  assign writeQueueVec_10_enq_bits_data_mask = otherTryToWrite[10] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_10_bits_mask;
  assign writeQueueVec_10_enq_bits_data_data = otherTryToWrite[10] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_10_bits_data;
  assign writeQueueVec_10_enq_bits_data_last = otherTryToWrite[10] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_10_enq_bits_data_instructionIndex = otherTryToWrite[10] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_10_bits_instructionIndex;
  assign writeQueueVec_11_enq_valid = otherTryToWrite[11] | _loadUnit_vrfWritePort_11_valid;
  assign writeQueueVec_11_enq_bits_data_vd = otherTryToWrite[11] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_11_bits_vd;
  assign writeQueueVec_11_enq_bits_data_mask = otherTryToWrite[11] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_11_bits_mask;
  assign writeQueueVec_11_enq_bits_data_data = otherTryToWrite[11] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_11_bits_data;
  assign writeQueueVec_11_enq_bits_data_last = otherTryToWrite[11] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_11_enq_bits_data_instructionIndex = otherTryToWrite[11] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_11_bits_instructionIndex;
  assign writeQueueVec_12_enq_valid = otherTryToWrite[12] | _loadUnit_vrfWritePort_12_valid;
  assign writeQueueVec_12_enq_bits_data_vd = otherTryToWrite[12] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_12_bits_vd;
  assign writeQueueVec_12_enq_bits_data_mask = otherTryToWrite[12] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_12_bits_mask;
  assign writeQueueVec_12_enq_bits_data_data = otherTryToWrite[12] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_12_bits_data;
  assign writeQueueVec_12_enq_bits_data_last = otherTryToWrite[12] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_12_enq_bits_data_instructionIndex = otherTryToWrite[12] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_12_bits_instructionIndex;
  assign writeQueueVec_13_enq_valid = otherTryToWrite[13] | _loadUnit_vrfWritePort_13_valid;
  assign writeQueueVec_13_enq_bits_data_vd = otherTryToWrite[13] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_13_bits_vd;
  assign writeQueueVec_13_enq_bits_data_mask = otherTryToWrite[13] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_13_bits_mask;
  assign writeQueueVec_13_enq_bits_data_data = otherTryToWrite[13] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_13_bits_data;
  assign writeQueueVec_13_enq_bits_data_last = otherTryToWrite[13] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_13_enq_bits_data_instructionIndex = otherTryToWrite[13] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_13_bits_instructionIndex;
  assign writeQueueVec_14_enq_valid = otherTryToWrite[14] | _loadUnit_vrfWritePort_14_valid;
  assign writeQueueVec_14_enq_bits_data_vd = otherTryToWrite[14] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_14_bits_vd;
  assign writeQueueVec_14_enq_bits_data_mask = otherTryToWrite[14] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_14_bits_mask;
  assign writeQueueVec_14_enq_bits_data_data = otherTryToWrite[14] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_14_bits_data;
  assign writeQueueVec_14_enq_bits_data_last = otherTryToWrite[14] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_14_enq_bits_data_instructionIndex = otherTryToWrite[14] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_14_bits_instructionIndex;
  assign writeQueueVec_15_enq_valid = otherTryToWrite[15] | _loadUnit_vrfWritePort_15_valid;
  assign writeQueueVec_15_enq_bits_data_vd = otherTryToWrite[15] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_15_bits_vd;
  assign writeQueueVec_15_enq_bits_data_mask = otherTryToWrite[15] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_15_bits_mask;
  assign writeQueueVec_15_enq_bits_data_data = otherTryToWrite[15] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_15_bits_data;
  assign writeQueueVec_15_enq_bits_data_last = otherTryToWrite[15] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_15_enq_bits_data_instructionIndex = otherTryToWrite[15] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_15_bits_instructionIndex;
  assign writeQueueVec_16_enq_valid = otherTryToWrite[16] | _loadUnit_vrfWritePort_16_valid;
  assign writeQueueVec_16_enq_bits_data_vd = otherTryToWrite[16] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_16_bits_vd;
  assign writeQueueVec_16_enq_bits_data_mask = otherTryToWrite[16] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_16_bits_mask;
  assign writeQueueVec_16_enq_bits_data_data = otherTryToWrite[16] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_16_bits_data;
  assign writeQueueVec_16_enq_bits_data_last = otherTryToWrite[16] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_16_enq_bits_data_instructionIndex = otherTryToWrite[16] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_16_bits_instructionIndex;
  assign writeQueueVec_17_enq_valid = otherTryToWrite[17] | _loadUnit_vrfWritePort_17_valid;
  assign writeQueueVec_17_enq_bits_data_vd = otherTryToWrite[17] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_17_bits_vd;
  assign writeQueueVec_17_enq_bits_data_mask = otherTryToWrite[17] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_17_bits_mask;
  assign writeQueueVec_17_enq_bits_data_data = otherTryToWrite[17] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_17_bits_data;
  assign writeQueueVec_17_enq_bits_data_last = otherTryToWrite[17] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_17_enq_bits_data_instructionIndex = otherTryToWrite[17] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_17_bits_instructionIndex;
  assign writeQueueVec_18_enq_valid = otherTryToWrite[18] | _loadUnit_vrfWritePort_18_valid;
  assign writeQueueVec_18_enq_bits_data_vd = otherTryToWrite[18] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_18_bits_vd;
  assign writeQueueVec_18_enq_bits_data_mask = otherTryToWrite[18] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_18_bits_mask;
  assign writeQueueVec_18_enq_bits_data_data = otherTryToWrite[18] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_18_bits_data;
  assign writeQueueVec_18_enq_bits_data_last = otherTryToWrite[18] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_18_enq_bits_data_instructionIndex = otherTryToWrite[18] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_18_bits_instructionIndex;
  assign writeQueueVec_19_enq_valid = otherTryToWrite[19] | _loadUnit_vrfWritePort_19_valid;
  assign writeQueueVec_19_enq_bits_data_vd = otherTryToWrite[19] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_19_bits_vd;
  assign writeQueueVec_19_enq_bits_data_mask = otherTryToWrite[19] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_19_bits_mask;
  assign writeQueueVec_19_enq_bits_data_data = otherTryToWrite[19] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_19_bits_data;
  assign writeQueueVec_19_enq_bits_data_last = otherTryToWrite[19] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_19_enq_bits_data_instructionIndex = otherTryToWrite[19] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_19_bits_instructionIndex;
  assign writeQueueVec_20_enq_valid = otherTryToWrite[20] | _loadUnit_vrfWritePort_20_valid;
  assign writeQueueVec_20_enq_bits_data_vd = otherTryToWrite[20] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_20_bits_vd;
  assign writeQueueVec_20_enq_bits_data_mask = otherTryToWrite[20] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_20_bits_mask;
  assign writeQueueVec_20_enq_bits_data_data = otherTryToWrite[20] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_20_bits_data;
  assign writeQueueVec_20_enq_bits_data_last = otherTryToWrite[20] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_20_enq_bits_data_instructionIndex = otherTryToWrite[20] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_20_bits_instructionIndex;
  assign writeQueueVec_21_enq_valid = otherTryToWrite[21] | _loadUnit_vrfWritePort_21_valid;
  assign writeQueueVec_21_enq_bits_data_vd = otherTryToWrite[21] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_21_bits_vd;
  assign writeQueueVec_21_enq_bits_data_mask = otherTryToWrite[21] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_21_bits_mask;
  assign writeQueueVec_21_enq_bits_data_data = otherTryToWrite[21] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_21_bits_data;
  assign writeQueueVec_21_enq_bits_data_last = otherTryToWrite[21] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_21_enq_bits_data_instructionIndex = otherTryToWrite[21] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_21_bits_instructionIndex;
  assign writeQueueVec_22_enq_valid = otherTryToWrite[22] | _loadUnit_vrfWritePort_22_valid;
  assign writeQueueVec_22_enq_bits_data_vd = otherTryToWrite[22] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_22_bits_vd;
  assign writeQueueVec_22_enq_bits_data_mask = otherTryToWrite[22] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_22_bits_mask;
  assign writeQueueVec_22_enq_bits_data_data = otherTryToWrite[22] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_22_bits_data;
  assign writeQueueVec_22_enq_bits_data_last = otherTryToWrite[22] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_22_enq_bits_data_instructionIndex = otherTryToWrite[22] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_22_bits_instructionIndex;
  assign writeQueueVec_23_enq_valid = otherTryToWrite[23] | _loadUnit_vrfWritePort_23_valid;
  assign writeQueueVec_23_enq_bits_data_vd = otherTryToWrite[23] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_23_bits_vd;
  assign writeQueueVec_23_enq_bits_data_mask = otherTryToWrite[23] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_23_bits_mask;
  assign writeQueueVec_23_enq_bits_data_data = otherTryToWrite[23] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_23_bits_data;
  assign writeQueueVec_23_enq_bits_data_last = otherTryToWrite[23] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_23_enq_bits_data_instructionIndex = otherTryToWrite[23] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_23_bits_instructionIndex;
  assign writeQueueVec_24_enq_valid = otherTryToWrite[24] | _loadUnit_vrfWritePort_24_valid;
  assign writeQueueVec_24_enq_bits_data_vd = otherTryToWrite[24] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_24_bits_vd;
  assign writeQueueVec_24_enq_bits_data_mask = otherTryToWrite[24] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_24_bits_mask;
  assign writeQueueVec_24_enq_bits_data_data = otherTryToWrite[24] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_24_bits_data;
  assign writeQueueVec_24_enq_bits_data_last = otherTryToWrite[24] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_24_enq_bits_data_instructionIndex = otherTryToWrite[24] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_24_bits_instructionIndex;
  assign writeQueueVec_25_enq_valid = otherTryToWrite[25] | _loadUnit_vrfWritePort_25_valid;
  assign writeQueueVec_25_enq_bits_data_vd = otherTryToWrite[25] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_25_bits_vd;
  assign writeQueueVec_25_enq_bits_data_mask = otherTryToWrite[25] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_25_bits_mask;
  assign writeQueueVec_25_enq_bits_data_data = otherTryToWrite[25] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_25_bits_data;
  assign writeQueueVec_25_enq_bits_data_last = otherTryToWrite[25] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_25_enq_bits_data_instructionIndex = otherTryToWrite[25] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_25_bits_instructionIndex;
  assign writeQueueVec_26_enq_valid = otherTryToWrite[26] | _loadUnit_vrfWritePort_26_valid;
  assign writeQueueVec_26_enq_bits_data_vd = otherTryToWrite[26] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_26_bits_vd;
  assign writeQueueVec_26_enq_bits_data_mask = otherTryToWrite[26] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_26_bits_mask;
  assign writeQueueVec_26_enq_bits_data_data = otherTryToWrite[26] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_26_bits_data;
  assign writeQueueVec_26_enq_bits_data_last = otherTryToWrite[26] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_26_enq_bits_data_instructionIndex = otherTryToWrite[26] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_26_bits_instructionIndex;
  assign writeQueueVec_27_enq_valid = otherTryToWrite[27] | _loadUnit_vrfWritePort_27_valid;
  assign writeQueueVec_27_enq_bits_data_vd = otherTryToWrite[27] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_27_bits_vd;
  assign writeQueueVec_27_enq_bits_data_mask = otherTryToWrite[27] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_27_bits_mask;
  assign writeQueueVec_27_enq_bits_data_data = otherTryToWrite[27] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_27_bits_data;
  assign writeQueueVec_27_enq_bits_data_last = otherTryToWrite[27] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_27_enq_bits_data_instructionIndex = otherTryToWrite[27] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_27_bits_instructionIndex;
  assign writeQueueVec_28_enq_valid = otherTryToWrite[28] | _loadUnit_vrfWritePort_28_valid;
  assign writeQueueVec_28_enq_bits_data_vd = otherTryToWrite[28] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_28_bits_vd;
  assign writeQueueVec_28_enq_bits_data_mask = otherTryToWrite[28] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_28_bits_mask;
  assign writeQueueVec_28_enq_bits_data_data = otherTryToWrite[28] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_28_bits_data;
  assign writeQueueVec_28_enq_bits_data_last = otherTryToWrite[28] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_28_enq_bits_data_instructionIndex = otherTryToWrite[28] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_28_bits_instructionIndex;
  assign writeQueueVec_29_enq_valid = otherTryToWrite[29] | _loadUnit_vrfWritePort_29_valid;
  assign writeQueueVec_29_enq_bits_data_vd = otherTryToWrite[29] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_29_bits_vd;
  assign writeQueueVec_29_enq_bits_data_mask = otherTryToWrite[29] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_29_bits_mask;
  assign writeQueueVec_29_enq_bits_data_data = otherTryToWrite[29] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_29_bits_data;
  assign writeQueueVec_29_enq_bits_data_last = otherTryToWrite[29] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_29_enq_bits_data_instructionIndex = otherTryToWrite[29] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_29_bits_instructionIndex;
  assign writeQueueVec_30_enq_valid = otherTryToWrite[30] | _loadUnit_vrfWritePort_30_valid;
  assign writeQueueVec_30_enq_bits_data_vd = otherTryToWrite[30] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_30_bits_vd;
  assign writeQueueVec_30_enq_bits_data_mask = otherTryToWrite[30] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_30_bits_mask;
  assign writeQueueVec_30_enq_bits_data_data = otherTryToWrite[30] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_30_bits_data;
  assign writeQueueVec_30_enq_bits_data_last = otherTryToWrite[30] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_30_enq_bits_data_instructionIndex = otherTryToWrite[30] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_30_bits_instructionIndex;
  assign writeQueueVec_31_enq_valid = otherTryToWrite[31] | _loadUnit_vrfWritePort_31_valid;
  assign writeQueueVec_31_enq_bits_data_vd = otherTryToWrite[31] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_31_bits_vd;
  assign writeQueueVec_31_enq_bits_data_mask = otherTryToWrite[31] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_31_bits_mask;
  assign writeQueueVec_31_enq_bits_data_data = otherTryToWrite[31] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_31_bits_data;
  assign writeQueueVec_31_enq_bits_data_last = otherTryToWrite[31] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_31_enq_bits_data_instructionIndex = otherTryToWrite[31] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_31_bits_instructionIndex;
  wire [7:0]        _GEN_18 = {5'h0, _loadUnit_status_instructionIndex};
  wire [7:0]        _GEN_19 = {5'h0, _otherUnit_status_instructionIndex};
  wire [7:0]        dataInMSHR = (_loadUnit_status_idle ? 8'h0 : 8'h1 << _GEN_18) | (_otherUnit_status_idle | _otherUnit_status_isStore ? 8'h0 : 8'h1 << _GEN_19);
  reg  [6:0]        queueCount_0;
  reg  [6:0]        queueCount_1;
  reg  [6:0]        queueCount_2;
  reg  [6:0]        queueCount_3;
  reg  [6:0]        queueCount_4;
  reg  [6:0]        queueCount_5;
  reg  [6:0]        queueCount_6;
  reg  [6:0]        queueCount_7;
  wire [7:0]        enqOH = 8'h1 << writeQueueVec_0_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq = _probeWire_slots_0_writeValid_T ? enqOH : 8'h0;
  wire              writeIndexQueue_deq_valid;
  assign writeIndexQueue_deq_valid = ~_writeIndexQueue_fifo_empty;
  wire              writeIndexQueue_enq_ready = ~_writeIndexQueue_fifo_full;
  wire              writeIndexQueue_enq_valid;
  assign writeIndexQueue_enq_valid = writeQueueVec_0_deq_ready & writeQueueVec_0_deq_valid;
  wire [2:0]        writeIndexQueue_deq_bits;
  wire [7:0]        queueDeq = writeIndexQueue_deq_ready & writeIndexQueue_deq_valid ? 8'h1 << writeIndexQueue_deq_bits : 8'h0;
  wire [6:0]        counterUpdate = queueEnq[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_1 = queueEnq[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_2 = queueEnq[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_3 = queueEnq[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_4 = queueEnq[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_5 = queueEnq[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_6 = queueEnq[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_7 = queueEnq[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_0_lo_lo = {|queueCount_1, |queueCount_0};
  wire [1:0]        dataInWriteQueue_0_lo_hi = {|queueCount_3, |queueCount_2};
  wire [3:0]        dataInWriteQueue_0_lo = {dataInWriteQueue_0_lo_hi, dataInWriteQueue_0_lo_lo};
  wire [1:0]        dataInWriteQueue_0_hi_lo = {|queueCount_5, |queueCount_4};
  wire [1:0]        dataInWriteQueue_0_hi_hi = {|queueCount_7, |queueCount_6};
  wire [3:0]        dataInWriteQueue_0_hi = {dataInWriteQueue_0_hi_hi, dataInWriteQueue_0_hi_lo};
  reg  [6:0]        queueCount_0_1;
  reg  [6:0]        queueCount_1_1;
  reg  [6:0]        queueCount_2_1;
  reg  [6:0]        queueCount_3_1;
  reg  [6:0]        queueCount_4_1;
  reg  [6:0]        queueCount_5_1;
  reg  [6:0]        queueCount_6_1;
  reg  [6:0]        queueCount_7_1;
  wire [7:0]        enqOH_1 = 8'h1 << writeQueueVec_1_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_1 = _probeWire_slots_1_writeValid_T ? enqOH_1 : 8'h0;
  wire              writeIndexQueue_1_deq_valid;
  assign writeIndexQueue_1_deq_valid = ~_writeIndexQueue_fifo_1_empty;
  wire              writeIndexQueue_1_enq_ready = ~_writeIndexQueue_fifo_1_full;
  wire              writeIndexQueue_1_enq_valid;
  assign writeIndexQueue_1_enq_valid = writeQueueVec_1_deq_ready & writeQueueVec_1_deq_valid;
  wire [2:0]        writeIndexQueue_1_deq_bits;
  wire [7:0]        queueDeq_1 = writeIndexQueue_1_deq_ready & writeIndexQueue_1_deq_valid ? 8'h1 << writeIndexQueue_1_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_8 = queueEnq_1[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_9 = queueEnq_1[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_10 = queueEnq_1[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_11 = queueEnq_1[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_12 = queueEnq_1[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_13 = queueEnq_1[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_14 = queueEnq_1[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_15 = queueEnq_1[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_1_lo_lo = {|queueCount_1_1, |queueCount_0_1};
  wire [1:0]        dataInWriteQueue_1_lo_hi = {|queueCount_3_1, |queueCount_2_1};
  wire [3:0]        dataInWriteQueue_1_lo = {dataInWriteQueue_1_lo_hi, dataInWriteQueue_1_lo_lo};
  wire [1:0]        dataInWriteQueue_1_hi_lo = {|queueCount_5_1, |queueCount_4_1};
  wire [1:0]        dataInWriteQueue_1_hi_hi = {|queueCount_7_1, |queueCount_6_1};
  wire [3:0]        dataInWriteQueue_1_hi = {dataInWriteQueue_1_hi_hi, dataInWriteQueue_1_hi_lo};
  reg  [6:0]        queueCount_0_2;
  reg  [6:0]        queueCount_1_2;
  reg  [6:0]        queueCount_2_2;
  reg  [6:0]        queueCount_3_2;
  reg  [6:0]        queueCount_4_2;
  reg  [6:0]        queueCount_5_2;
  reg  [6:0]        queueCount_6_2;
  reg  [6:0]        queueCount_7_2;
  wire [7:0]        enqOH_2 = 8'h1 << writeQueueVec_2_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_2 = _probeWire_slots_2_writeValid_T ? enqOH_2 : 8'h0;
  wire              writeIndexQueue_2_deq_valid;
  assign writeIndexQueue_2_deq_valid = ~_writeIndexQueue_fifo_2_empty;
  wire              writeIndexQueue_2_enq_ready = ~_writeIndexQueue_fifo_2_full;
  wire              writeIndexQueue_2_enq_valid;
  assign writeIndexQueue_2_enq_valid = writeQueueVec_2_deq_ready & writeQueueVec_2_deq_valid;
  wire [2:0]        writeIndexQueue_2_deq_bits;
  wire [7:0]        queueDeq_2 = writeIndexQueue_2_deq_ready & writeIndexQueue_2_deq_valid ? 8'h1 << writeIndexQueue_2_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_16 = queueEnq_2[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_17 = queueEnq_2[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_18 = queueEnq_2[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_19 = queueEnq_2[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_20 = queueEnq_2[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_21 = queueEnq_2[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_22 = queueEnq_2[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_23 = queueEnq_2[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_2_lo_lo = {|queueCount_1_2, |queueCount_0_2};
  wire [1:0]        dataInWriteQueue_2_lo_hi = {|queueCount_3_2, |queueCount_2_2};
  wire [3:0]        dataInWriteQueue_2_lo = {dataInWriteQueue_2_lo_hi, dataInWriteQueue_2_lo_lo};
  wire [1:0]        dataInWriteQueue_2_hi_lo = {|queueCount_5_2, |queueCount_4_2};
  wire [1:0]        dataInWriteQueue_2_hi_hi = {|queueCount_7_2, |queueCount_6_2};
  wire [3:0]        dataInWriteQueue_2_hi = {dataInWriteQueue_2_hi_hi, dataInWriteQueue_2_hi_lo};
  reg  [6:0]        queueCount_0_3;
  reg  [6:0]        queueCount_1_3;
  reg  [6:0]        queueCount_2_3;
  reg  [6:0]        queueCount_3_3;
  reg  [6:0]        queueCount_4_3;
  reg  [6:0]        queueCount_5_3;
  reg  [6:0]        queueCount_6_3;
  reg  [6:0]        queueCount_7_3;
  wire [7:0]        enqOH_3 = 8'h1 << writeQueueVec_3_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_3 = _probeWire_slots_3_writeValid_T ? enqOH_3 : 8'h0;
  wire              writeIndexQueue_3_deq_valid;
  assign writeIndexQueue_3_deq_valid = ~_writeIndexQueue_fifo_3_empty;
  wire              writeIndexQueue_3_enq_ready = ~_writeIndexQueue_fifo_3_full;
  wire              writeIndexQueue_3_enq_valid;
  assign writeIndexQueue_3_enq_valid = writeQueueVec_3_deq_ready & writeQueueVec_3_deq_valid;
  wire [2:0]        writeIndexQueue_3_deq_bits;
  wire [7:0]        queueDeq_3 = writeIndexQueue_3_deq_ready & writeIndexQueue_3_deq_valid ? 8'h1 << writeIndexQueue_3_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_24 = queueEnq_3[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_25 = queueEnq_3[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_26 = queueEnq_3[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_27 = queueEnq_3[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_28 = queueEnq_3[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_29 = queueEnq_3[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_30 = queueEnq_3[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_31 = queueEnq_3[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_3_lo_lo = {|queueCount_1_3, |queueCount_0_3};
  wire [1:0]        dataInWriteQueue_3_lo_hi = {|queueCount_3_3, |queueCount_2_3};
  wire [3:0]        dataInWriteQueue_3_lo = {dataInWriteQueue_3_lo_hi, dataInWriteQueue_3_lo_lo};
  wire [1:0]        dataInWriteQueue_3_hi_lo = {|queueCount_5_3, |queueCount_4_3};
  wire [1:0]        dataInWriteQueue_3_hi_hi = {|queueCount_7_3, |queueCount_6_3};
  wire [3:0]        dataInWriteQueue_3_hi = {dataInWriteQueue_3_hi_hi, dataInWriteQueue_3_hi_lo};
  reg  [6:0]        queueCount_0_4;
  reg  [6:0]        queueCount_1_4;
  reg  [6:0]        queueCount_2_4;
  reg  [6:0]        queueCount_3_4;
  reg  [6:0]        queueCount_4_4;
  reg  [6:0]        queueCount_5_4;
  reg  [6:0]        queueCount_6_4;
  reg  [6:0]        queueCount_7_4;
  wire [7:0]        enqOH_4 = 8'h1 << writeQueueVec_4_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_4 = _probeWire_slots_4_writeValid_T ? enqOH_4 : 8'h0;
  wire              writeIndexQueue_4_deq_valid;
  assign writeIndexQueue_4_deq_valid = ~_writeIndexQueue_fifo_4_empty;
  wire              writeIndexQueue_4_enq_ready = ~_writeIndexQueue_fifo_4_full;
  wire              writeIndexQueue_4_enq_valid;
  assign writeIndexQueue_4_enq_valid = writeQueueVec_4_deq_ready & writeQueueVec_4_deq_valid;
  wire [2:0]        writeIndexQueue_4_deq_bits;
  wire [7:0]        queueDeq_4 = writeIndexQueue_4_deq_ready & writeIndexQueue_4_deq_valid ? 8'h1 << writeIndexQueue_4_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_32 = queueEnq_4[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_33 = queueEnq_4[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_34 = queueEnq_4[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_35 = queueEnq_4[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_36 = queueEnq_4[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_37 = queueEnq_4[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_38 = queueEnq_4[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_39 = queueEnq_4[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_4_lo_lo = {|queueCount_1_4, |queueCount_0_4};
  wire [1:0]        dataInWriteQueue_4_lo_hi = {|queueCount_3_4, |queueCount_2_4};
  wire [3:0]        dataInWriteQueue_4_lo = {dataInWriteQueue_4_lo_hi, dataInWriteQueue_4_lo_lo};
  wire [1:0]        dataInWriteQueue_4_hi_lo = {|queueCount_5_4, |queueCount_4_4};
  wire [1:0]        dataInWriteQueue_4_hi_hi = {|queueCount_7_4, |queueCount_6_4};
  wire [3:0]        dataInWriteQueue_4_hi = {dataInWriteQueue_4_hi_hi, dataInWriteQueue_4_hi_lo};
  reg  [6:0]        queueCount_0_5;
  reg  [6:0]        queueCount_1_5;
  reg  [6:0]        queueCount_2_5;
  reg  [6:0]        queueCount_3_5;
  reg  [6:0]        queueCount_4_5;
  reg  [6:0]        queueCount_5_5;
  reg  [6:0]        queueCount_6_5;
  reg  [6:0]        queueCount_7_5;
  wire [7:0]        enqOH_5 = 8'h1 << writeQueueVec_5_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_5 = _probeWire_slots_5_writeValid_T ? enqOH_5 : 8'h0;
  wire              writeIndexQueue_5_deq_valid;
  assign writeIndexQueue_5_deq_valid = ~_writeIndexQueue_fifo_5_empty;
  wire              writeIndexQueue_5_enq_ready = ~_writeIndexQueue_fifo_5_full;
  wire              writeIndexQueue_5_enq_valid;
  assign writeIndexQueue_5_enq_valid = writeQueueVec_5_deq_ready & writeQueueVec_5_deq_valid;
  wire [2:0]        writeIndexQueue_5_deq_bits;
  wire [7:0]        queueDeq_5 = writeIndexQueue_5_deq_ready & writeIndexQueue_5_deq_valid ? 8'h1 << writeIndexQueue_5_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_40 = queueEnq_5[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_41 = queueEnq_5[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_42 = queueEnq_5[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_43 = queueEnq_5[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_44 = queueEnq_5[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_45 = queueEnq_5[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_46 = queueEnq_5[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_47 = queueEnq_5[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_5_lo_lo = {|queueCount_1_5, |queueCount_0_5};
  wire [1:0]        dataInWriteQueue_5_lo_hi = {|queueCount_3_5, |queueCount_2_5};
  wire [3:0]        dataInWriteQueue_5_lo = {dataInWriteQueue_5_lo_hi, dataInWriteQueue_5_lo_lo};
  wire [1:0]        dataInWriteQueue_5_hi_lo = {|queueCount_5_5, |queueCount_4_5};
  wire [1:0]        dataInWriteQueue_5_hi_hi = {|queueCount_7_5, |queueCount_6_5};
  wire [3:0]        dataInWriteQueue_5_hi = {dataInWriteQueue_5_hi_hi, dataInWriteQueue_5_hi_lo};
  reg  [6:0]        queueCount_0_6;
  reg  [6:0]        queueCount_1_6;
  reg  [6:0]        queueCount_2_6;
  reg  [6:0]        queueCount_3_6;
  reg  [6:0]        queueCount_4_6;
  reg  [6:0]        queueCount_5_6;
  reg  [6:0]        queueCount_6_6;
  reg  [6:0]        queueCount_7_6;
  wire [7:0]        enqOH_6 = 8'h1 << writeQueueVec_6_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_6 = _probeWire_slots_6_writeValid_T ? enqOH_6 : 8'h0;
  wire              writeIndexQueue_6_deq_valid;
  assign writeIndexQueue_6_deq_valid = ~_writeIndexQueue_fifo_6_empty;
  wire              writeIndexQueue_6_enq_ready = ~_writeIndexQueue_fifo_6_full;
  wire              writeIndexQueue_6_enq_valid;
  assign writeIndexQueue_6_enq_valid = writeQueueVec_6_deq_ready & writeQueueVec_6_deq_valid;
  wire [2:0]        writeIndexQueue_6_deq_bits;
  wire [7:0]        queueDeq_6 = writeIndexQueue_6_deq_ready & writeIndexQueue_6_deq_valid ? 8'h1 << writeIndexQueue_6_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_48 = queueEnq_6[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_49 = queueEnq_6[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_50 = queueEnq_6[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_51 = queueEnq_6[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_52 = queueEnq_6[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_53 = queueEnq_6[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_54 = queueEnq_6[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_55 = queueEnq_6[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_6_lo_lo = {|queueCount_1_6, |queueCount_0_6};
  wire [1:0]        dataInWriteQueue_6_lo_hi = {|queueCount_3_6, |queueCount_2_6};
  wire [3:0]        dataInWriteQueue_6_lo = {dataInWriteQueue_6_lo_hi, dataInWriteQueue_6_lo_lo};
  wire [1:0]        dataInWriteQueue_6_hi_lo = {|queueCount_5_6, |queueCount_4_6};
  wire [1:0]        dataInWriteQueue_6_hi_hi = {|queueCount_7_6, |queueCount_6_6};
  wire [3:0]        dataInWriteQueue_6_hi = {dataInWriteQueue_6_hi_hi, dataInWriteQueue_6_hi_lo};
  reg  [6:0]        queueCount_0_7;
  reg  [6:0]        queueCount_1_7;
  reg  [6:0]        queueCount_2_7;
  reg  [6:0]        queueCount_3_7;
  reg  [6:0]        queueCount_4_7;
  reg  [6:0]        queueCount_5_7;
  reg  [6:0]        queueCount_6_7;
  reg  [6:0]        queueCount_7_7;
  wire [7:0]        enqOH_7 = 8'h1 << writeQueueVec_7_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_7 = _probeWire_slots_7_writeValid_T ? enqOH_7 : 8'h0;
  wire              writeIndexQueue_7_deq_valid;
  assign writeIndexQueue_7_deq_valid = ~_writeIndexQueue_fifo_7_empty;
  wire              writeIndexQueue_7_enq_ready = ~_writeIndexQueue_fifo_7_full;
  wire              writeIndexQueue_7_enq_valid;
  assign writeIndexQueue_7_enq_valid = writeQueueVec_7_deq_ready & writeQueueVec_7_deq_valid;
  wire [2:0]        writeIndexQueue_7_deq_bits;
  wire [7:0]        queueDeq_7 = writeIndexQueue_7_deq_ready & writeIndexQueue_7_deq_valid ? 8'h1 << writeIndexQueue_7_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_56 = queueEnq_7[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_57 = queueEnq_7[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_58 = queueEnq_7[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_59 = queueEnq_7[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_60 = queueEnq_7[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_61 = queueEnq_7[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_62 = queueEnq_7[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_63 = queueEnq_7[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_7_lo_lo = {|queueCount_1_7, |queueCount_0_7};
  wire [1:0]        dataInWriteQueue_7_lo_hi = {|queueCount_3_7, |queueCount_2_7};
  wire [3:0]        dataInWriteQueue_7_lo = {dataInWriteQueue_7_lo_hi, dataInWriteQueue_7_lo_lo};
  wire [1:0]        dataInWriteQueue_7_hi_lo = {|queueCount_5_7, |queueCount_4_7};
  wire [1:0]        dataInWriteQueue_7_hi_hi = {|queueCount_7_7, |queueCount_6_7};
  wire [3:0]        dataInWriteQueue_7_hi = {dataInWriteQueue_7_hi_hi, dataInWriteQueue_7_hi_lo};
  reg  [6:0]        queueCount_0_8;
  reg  [6:0]        queueCount_1_8;
  reg  [6:0]        queueCount_2_8;
  reg  [6:0]        queueCount_3_8;
  reg  [6:0]        queueCount_4_8;
  reg  [6:0]        queueCount_5_8;
  reg  [6:0]        queueCount_6_8;
  reg  [6:0]        queueCount_7_8;
  wire [7:0]        enqOH_8 = 8'h1 << writeQueueVec_8_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_8 = _probeWire_slots_8_writeValid_T ? enqOH_8 : 8'h0;
  wire              writeIndexQueue_8_deq_valid;
  assign writeIndexQueue_8_deq_valid = ~_writeIndexQueue_fifo_8_empty;
  wire              writeIndexQueue_8_enq_ready = ~_writeIndexQueue_fifo_8_full;
  wire              writeIndexQueue_8_enq_valid;
  assign writeIndexQueue_8_enq_valid = writeQueueVec_8_deq_ready & writeQueueVec_8_deq_valid;
  wire [2:0]        writeIndexQueue_8_deq_bits;
  wire [7:0]        queueDeq_8 = writeIndexQueue_8_deq_ready & writeIndexQueue_8_deq_valid ? 8'h1 << writeIndexQueue_8_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_64 = queueEnq_8[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_65 = queueEnq_8[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_66 = queueEnq_8[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_67 = queueEnq_8[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_68 = queueEnq_8[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_69 = queueEnq_8[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_70 = queueEnq_8[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_71 = queueEnq_8[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_8_lo_lo = {|queueCount_1_8, |queueCount_0_8};
  wire [1:0]        dataInWriteQueue_8_lo_hi = {|queueCount_3_8, |queueCount_2_8};
  wire [3:0]        dataInWriteQueue_8_lo = {dataInWriteQueue_8_lo_hi, dataInWriteQueue_8_lo_lo};
  wire [1:0]        dataInWriteQueue_8_hi_lo = {|queueCount_5_8, |queueCount_4_8};
  wire [1:0]        dataInWriteQueue_8_hi_hi = {|queueCount_7_8, |queueCount_6_8};
  wire [3:0]        dataInWriteQueue_8_hi = {dataInWriteQueue_8_hi_hi, dataInWriteQueue_8_hi_lo};
  reg  [6:0]        queueCount_0_9;
  reg  [6:0]        queueCount_1_9;
  reg  [6:0]        queueCount_2_9;
  reg  [6:0]        queueCount_3_9;
  reg  [6:0]        queueCount_4_9;
  reg  [6:0]        queueCount_5_9;
  reg  [6:0]        queueCount_6_9;
  reg  [6:0]        queueCount_7_9;
  wire [7:0]        enqOH_9 = 8'h1 << writeQueueVec_9_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_9 = _probeWire_slots_9_writeValid_T ? enqOH_9 : 8'h0;
  wire              writeIndexQueue_9_deq_valid;
  assign writeIndexQueue_9_deq_valid = ~_writeIndexQueue_fifo_9_empty;
  wire              writeIndexQueue_9_enq_ready = ~_writeIndexQueue_fifo_9_full;
  wire              writeIndexQueue_9_enq_valid;
  assign writeIndexQueue_9_enq_valid = writeQueueVec_9_deq_ready & writeQueueVec_9_deq_valid;
  wire [2:0]        writeIndexQueue_9_deq_bits;
  wire [7:0]        queueDeq_9 = writeIndexQueue_9_deq_ready & writeIndexQueue_9_deq_valid ? 8'h1 << writeIndexQueue_9_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_72 = queueEnq_9[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_73 = queueEnq_9[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_74 = queueEnq_9[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_75 = queueEnq_9[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_76 = queueEnq_9[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_77 = queueEnq_9[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_78 = queueEnq_9[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_79 = queueEnq_9[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_9_lo_lo = {|queueCount_1_9, |queueCount_0_9};
  wire [1:0]        dataInWriteQueue_9_lo_hi = {|queueCount_3_9, |queueCount_2_9};
  wire [3:0]        dataInWriteQueue_9_lo = {dataInWriteQueue_9_lo_hi, dataInWriteQueue_9_lo_lo};
  wire [1:0]        dataInWriteQueue_9_hi_lo = {|queueCount_5_9, |queueCount_4_9};
  wire [1:0]        dataInWriteQueue_9_hi_hi = {|queueCount_7_9, |queueCount_6_9};
  wire [3:0]        dataInWriteQueue_9_hi = {dataInWriteQueue_9_hi_hi, dataInWriteQueue_9_hi_lo};
  reg  [6:0]        queueCount_0_10;
  reg  [6:0]        queueCount_1_10;
  reg  [6:0]        queueCount_2_10;
  reg  [6:0]        queueCount_3_10;
  reg  [6:0]        queueCount_4_10;
  reg  [6:0]        queueCount_5_10;
  reg  [6:0]        queueCount_6_10;
  reg  [6:0]        queueCount_7_10;
  wire [7:0]        enqOH_10 = 8'h1 << writeQueueVec_10_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_10 = _probeWire_slots_10_writeValid_T ? enqOH_10 : 8'h0;
  wire              writeIndexQueue_10_deq_valid;
  assign writeIndexQueue_10_deq_valid = ~_writeIndexQueue_fifo_10_empty;
  wire              writeIndexQueue_10_enq_ready = ~_writeIndexQueue_fifo_10_full;
  wire              writeIndexQueue_10_enq_valid;
  assign writeIndexQueue_10_enq_valid = writeQueueVec_10_deq_ready & writeQueueVec_10_deq_valid;
  wire [2:0]        writeIndexQueue_10_deq_bits;
  wire [7:0]        queueDeq_10 = writeIndexQueue_10_deq_ready & writeIndexQueue_10_deq_valid ? 8'h1 << writeIndexQueue_10_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_80 = queueEnq_10[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_81 = queueEnq_10[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_82 = queueEnq_10[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_83 = queueEnq_10[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_84 = queueEnq_10[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_85 = queueEnq_10[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_86 = queueEnq_10[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_87 = queueEnq_10[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_10_lo_lo = {|queueCount_1_10, |queueCount_0_10};
  wire [1:0]        dataInWriteQueue_10_lo_hi = {|queueCount_3_10, |queueCount_2_10};
  wire [3:0]        dataInWriteQueue_10_lo = {dataInWriteQueue_10_lo_hi, dataInWriteQueue_10_lo_lo};
  wire [1:0]        dataInWriteQueue_10_hi_lo = {|queueCount_5_10, |queueCount_4_10};
  wire [1:0]        dataInWriteQueue_10_hi_hi = {|queueCount_7_10, |queueCount_6_10};
  wire [3:0]        dataInWriteQueue_10_hi = {dataInWriteQueue_10_hi_hi, dataInWriteQueue_10_hi_lo};
  reg  [6:0]        queueCount_0_11;
  reg  [6:0]        queueCount_1_11;
  reg  [6:0]        queueCount_2_11;
  reg  [6:0]        queueCount_3_11;
  reg  [6:0]        queueCount_4_11;
  reg  [6:0]        queueCount_5_11;
  reg  [6:0]        queueCount_6_11;
  reg  [6:0]        queueCount_7_11;
  wire [7:0]        enqOH_11 = 8'h1 << writeQueueVec_11_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_11 = _probeWire_slots_11_writeValid_T ? enqOH_11 : 8'h0;
  wire              writeIndexQueue_11_deq_valid;
  assign writeIndexQueue_11_deq_valid = ~_writeIndexQueue_fifo_11_empty;
  wire              writeIndexQueue_11_enq_ready = ~_writeIndexQueue_fifo_11_full;
  wire              writeIndexQueue_11_enq_valid;
  assign writeIndexQueue_11_enq_valid = writeQueueVec_11_deq_ready & writeQueueVec_11_deq_valid;
  wire [2:0]        writeIndexQueue_11_deq_bits;
  wire [7:0]        queueDeq_11 = writeIndexQueue_11_deq_ready & writeIndexQueue_11_deq_valid ? 8'h1 << writeIndexQueue_11_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_88 = queueEnq_11[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_89 = queueEnq_11[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_90 = queueEnq_11[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_91 = queueEnq_11[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_92 = queueEnq_11[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_93 = queueEnq_11[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_94 = queueEnq_11[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_95 = queueEnq_11[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_11_lo_lo = {|queueCount_1_11, |queueCount_0_11};
  wire [1:0]        dataInWriteQueue_11_lo_hi = {|queueCount_3_11, |queueCount_2_11};
  wire [3:0]        dataInWriteQueue_11_lo = {dataInWriteQueue_11_lo_hi, dataInWriteQueue_11_lo_lo};
  wire [1:0]        dataInWriteQueue_11_hi_lo = {|queueCount_5_11, |queueCount_4_11};
  wire [1:0]        dataInWriteQueue_11_hi_hi = {|queueCount_7_11, |queueCount_6_11};
  wire [3:0]        dataInWriteQueue_11_hi = {dataInWriteQueue_11_hi_hi, dataInWriteQueue_11_hi_lo};
  reg  [6:0]        queueCount_0_12;
  reg  [6:0]        queueCount_1_12;
  reg  [6:0]        queueCount_2_12;
  reg  [6:0]        queueCount_3_12;
  reg  [6:0]        queueCount_4_12;
  reg  [6:0]        queueCount_5_12;
  reg  [6:0]        queueCount_6_12;
  reg  [6:0]        queueCount_7_12;
  wire [7:0]        enqOH_12 = 8'h1 << writeQueueVec_12_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_12 = _probeWire_slots_12_writeValid_T ? enqOH_12 : 8'h0;
  wire              writeIndexQueue_12_deq_valid;
  assign writeIndexQueue_12_deq_valid = ~_writeIndexQueue_fifo_12_empty;
  wire              writeIndexQueue_12_enq_ready = ~_writeIndexQueue_fifo_12_full;
  wire              writeIndexQueue_12_enq_valid;
  assign writeIndexQueue_12_enq_valid = writeQueueVec_12_deq_ready & writeQueueVec_12_deq_valid;
  wire [2:0]        writeIndexQueue_12_deq_bits;
  wire [7:0]        queueDeq_12 = writeIndexQueue_12_deq_ready & writeIndexQueue_12_deq_valid ? 8'h1 << writeIndexQueue_12_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_96 = queueEnq_12[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_97 = queueEnq_12[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_98 = queueEnq_12[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_99 = queueEnq_12[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_100 = queueEnq_12[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_101 = queueEnq_12[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_102 = queueEnq_12[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_103 = queueEnq_12[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_12_lo_lo = {|queueCount_1_12, |queueCount_0_12};
  wire [1:0]        dataInWriteQueue_12_lo_hi = {|queueCount_3_12, |queueCount_2_12};
  wire [3:0]        dataInWriteQueue_12_lo = {dataInWriteQueue_12_lo_hi, dataInWriteQueue_12_lo_lo};
  wire [1:0]        dataInWriteQueue_12_hi_lo = {|queueCount_5_12, |queueCount_4_12};
  wire [1:0]        dataInWriteQueue_12_hi_hi = {|queueCount_7_12, |queueCount_6_12};
  wire [3:0]        dataInWriteQueue_12_hi = {dataInWriteQueue_12_hi_hi, dataInWriteQueue_12_hi_lo};
  reg  [6:0]        queueCount_0_13;
  reg  [6:0]        queueCount_1_13;
  reg  [6:0]        queueCount_2_13;
  reg  [6:0]        queueCount_3_13;
  reg  [6:0]        queueCount_4_13;
  reg  [6:0]        queueCount_5_13;
  reg  [6:0]        queueCount_6_13;
  reg  [6:0]        queueCount_7_13;
  wire [7:0]        enqOH_13 = 8'h1 << writeQueueVec_13_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_13 = _probeWire_slots_13_writeValid_T ? enqOH_13 : 8'h0;
  wire              writeIndexQueue_13_deq_valid;
  assign writeIndexQueue_13_deq_valid = ~_writeIndexQueue_fifo_13_empty;
  wire              writeIndexQueue_13_enq_ready = ~_writeIndexQueue_fifo_13_full;
  wire              writeIndexQueue_13_enq_valid;
  assign writeIndexQueue_13_enq_valid = writeQueueVec_13_deq_ready & writeQueueVec_13_deq_valid;
  wire [2:0]        writeIndexQueue_13_deq_bits;
  wire [7:0]        queueDeq_13 = writeIndexQueue_13_deq_ready & writeIndexQueue_13_deq_valid ? 8'h1 << writeIndexQueue_13_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_104 = queueEnq_13[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_105 = queueEnq_13[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_106 = queueEnq_13[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_107 = queueEnq_13[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_108 = queueEnq_13[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_109 = queueEnq_13[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_110 = queueEnq_13[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_111 = queueEnq_13[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_13_lo_lo = {|queueCount_1_13, |queueCount_0_13};
  wire [1:0]        dataInWriteQueue_13_lo_hi = {|queueCount_3_13, |queueCount_2_13};
  wire [3:0]        dataInWriteQueue_13_lo = {dataInWriteQueue_13_lo_hi, dataInWriteQueue_13_lo_lo};
  wire [1:0]        dataInWriteQueue_13_hi_lo = {|queueCount_5_13, |queueCount_4_13};
  wire [1:0]        dataInWriteQueue_13_hi_hi = {|queueCount_7_13, |queueCount_6_13};
  wire [3:0]        dataInWriteQueue_13_hi = {dataInWriteQueue_13_hi_hi, dataInWriteQueue_13_hi_lo};
  reg  [6:0]        queueCount_0_14;
  reg  [6:0]        queueCount_1_14;
  reg  [6:0]        queueCount_2_14;
  reg  [6:0]        queueCount_3_14;
  reg  [6:0]        queueCount_4_14;
  reg  [6:0]        queueCount_5_14;
  reg  [6:0]        queueCount_6_14;
  reg  [6:0]        queueCount_7_14;
  wire [7:0]        enqOH_14 = 8'h1 << writeQueueVec_14_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_14 = _probeWire_slots_14_writeValid_T ? enqOH_14 : 8'h0;
  wire              writeIndexQueue_14_deq_valid;
  assign writeIndexQueue_14_deq_valid = ~_writeIndexQueue_fifo_14_empty;
  wire              writeIndexQueue_14_enq_ready = ~_writeIndexQueue_fifo_14_full;
  wire              writeIndexQueue_14_enq_valid;
  assign writeIndexQueue_14_enq_valid = writeQueueVec_14_deq_ready & writeQueueVec_14_deq_valid;
  wire [2:0]        writeIndexQueue_14_deq_bits;
  wire [7:0]        queueDeq_14 = writeIndexQueue_14_deq_ready & writeIndexQueue_14_deq_valid ? 8'h1 << writeIndexQueue_14_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_112 = queueEnq_14[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_113 = queueEnq_14[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_114 = queueEnq_14[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_115 = queueEnq_14[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_116 = queueEnq_14[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_117 = queueEnq_14[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_118 = queueEnq_14[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_119 = queueEnq_14[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_14_lo_lo = {|queueCount_1_14, |queueCount_0_14};
  wire [1:0]        dataInWriteQueue_14_lo_hi = {|queueCount_3_14, |queueCount_2_14};
  wire [3:0]        dataInWriteQueue_14_lo = {dataInWriteQueue_14_lo_hi, dataInWriteQueue_14_lo_lo};
  wire [1:0]        dataInWriteQueue_14_hi_lo = {|queueCount_5_14, |queueCount_4_14};
  wire [1:0]        dataInWriteQueue_14_hi_hi = {|queueCount_7_14, |queueCount_6_14};
  wire [3:0]        dataInWriteQueue_14_hi = {dataInWriteQueue_14_hi_hi, dataInWriteQueue_14_hi_lo};
  reg  [6:0]        queueCount_0_15;
  reg  [6:0]        queueCount_1_15;
  reg  [6:0]        queueCount_2_15;
  reg  [6:0]        queueCount_3_15;
  reg  [6:0]        queueCount_4_15;
  reg  [6:0]        queueCount_5_15;
  reg  [6:0]        queueCount_6_15;
  reg  [6:0]        queueCount_7_15;
  wire [7:0]        enqOH_15 = 8'h1 << writeQueueVec_15_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_15 = _probeWire_slots_15_writeValid_T ? enqOH_15 : 8'h0;
  wire              writeIndexQueue_15_deq_valid;
  assign writeIndexQueue_15_deq_valid = ~_writeIndexQueue_fifo_15_empty;
  wire              writeIndexQueue_15_enq_ready = ~_writeIndexQueue_fifo_15_full;
  wire              writeIndexQueue_15_enq_valid;
  assign writeIndexQueue_15_enq_valid = writeQueueVec_15_deq_ready & writeQueueVec_15_deq_valid;
  wire [2:0]        writeIndexQueue_15_deq_bits;
  wire [7:0]        queueDeq_15 = writeIndexQueue_15_deq_ready & writeIndexQueue_15_deq_valid ? 8'h1 << writeIndexQueue_15_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_120 = queueEnq_15[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_121 = queueEnq_15[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_122 = queueEnq_15[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_123 = queueEnq_15[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_124 = queueEnq_15[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_125 = queueEnq_15[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_126 = queueEnq_15[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_127 = queueEnq_15[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_15_lo_lo = {|queueCount_1_15, |queueCount_0_15};
  wire [1:0]        dataInWriteQueue_15_lo_hi = {|queueCount_3_15, |queueCount_2_15};
  wire [3:0]        dataInWriteQueue_15_lo = {dataInWriteQueue_15_lo_hi, dataInWriteQueue_15_lo_lo};
  wire [1:0]        dataInWriteQueue_15_hi_lo = {|queueCount_5_15, |queueCount_4_15};
  wire [1:0]        dataInWriteQueue_15_hi_hi = {|queueCount_7_15, |queueCount_6_15};
  wire [3:0]        dataInWriteQueue_15_hi = {dataInWriteQueue_15_hi_hi, dataInWriteQueue_15_hi_lo};
  reg  [6:0]        queueCount_0_16;
  reg  [6:0]        queueCount_1_16;
  reg  [6:0]        queueCount_2_16;
  reg  [6:0]        queueCount_3_16;
  reg  [6:0]        queueCount_4_16;
  reg  [6:0]        queueCount_5_16;
  reg  [6:0]        queueCount_6_16;
  reg  [6:0]        queueCount_7_16;
  wire [7:0]        enqOH_16 = 8'h1 << writeQueueVec_16_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_16 = _probeWire_slots_16_writeValid_T ? enqOH_16 : 8'h0;
  wire              writeIndexQueue_16_deq_valid;
  assign writeIndexQueue_16_deq_valid = ~_writeIndexQueue_fifo_16_empty;
  wire              writeIndexQueue_16_enq_ready = ~_writeIndexQueue_fifo_16_full;
  wire              writeIndexQueue_16_enq_valid;
  assign writeIndexQueue_16_enq_valid = writeQueueVec_16_deq_ready & writeQueueVec_16_deq_valid;
  wire [2:0]        writeIndexQueue_16_deq_bits;
  wire [7:0]        queueDeq_16 = writeIndexQueue_16_deq_ready & writeIndexQueue_16_deq_valid ? 8'h1 << writeIndexQueue_16_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_128 = queueEnq_16[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_129 = queueEnq_16[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_130 = queueEnq_16[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_131 = queueEnq_16[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_132 = queueEnq_16[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_133 = queueEnq_16[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_134 = queueEnq_16[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_135 = queueEnq_16[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_16_lo_lo = {|queueCount_1_16, |queueCount_0_16};
  wire [1:0]        dataInWriteQueue_16_lo_hi = {|queueCount_3_16, |queueCount_2_16};
  wire [3:0]        dataInWriteQueue_16_lo = {dataInWriteQueue_16_lo_hi, dataInWriteQueue_16_lo_lo};
  wire [1:0]        dataInWriteQueue_16_hi_lo = {|queueCount_5_16, |queueCount_4_16};
  wire [1:0]        dataInWriteQueue_16_hi_hi = {|queueCount_7_16, |queueCount_6_16};
  wire [3:0]        dataInWriteQueue_16_hi = {dataInWriteQueue_16_hi_hi, dataInWriteQueue_16_hi_lo};
  reg  [6:0]        queueCount_0_17;
  reg  [6:0]        queueCount_1_17;
  reg  [6:0]        queueCount_2_17;
  reg  [6:0]        queueCount_3_17;
  reg  [6:0]        queueCount_4_17;
  reg  [6:0]        queueCount_5_17;
  reg  [6:0]        queueCount_6_17;
  reg  [6:0]        queueCount_7_17;
  wire [7:0]        enqOH_17 = 8'h1 << writeQueueVec_17_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_17 = _probeWire_slots_17_writeValid_T ? enqOH_17 : 8'h0;
  wire              writeIndexQueue_17_deq_valid;
  assign writeIndexQueue_17_deq_valid = ~_writeIndexQueue_fifo_17_empty;
  wire              writeIndexQueue_17_enq_ready = ~_writeIndexQueue_fifo_17_full;
  wire              writeIndexQueue_17_enq_valid;
  assign writeIndexQueue_17_enq_valid = writeQueueVec_17_deq_ready & writeQueueVec_17_deq_valid;
  wire [2:0]        writeIndexQueue_17_deq_bits;
  wire [7:0]        queueDeq_17 = writeIndexQueue_17_deq_ready & writeIndexQueue_17_deq_valid ? 8'h1 << writeIndexQueue_17_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_136 = queueEnq_17[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_137 = queueEnq_17[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_138 = queueEnq_17[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_139 = queueEnq_17[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_140 = queueEnq_17[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_141 = queueEnq_17[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_142 = queueEnq_17[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_143 = queueEnq_17[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_17_lo_lo = {|queueCount_1_17, |queueCount_0_17};
  wire [1:0]        dataInWriteQueue_17_lo_hi = {|queueCount_3_17, |queueCount_2_17};
  wire [3:0]        dataInWriteQueue_17_lo = {dataInWriteQueue_17_lo_hi, dataInWriteQueue_17_lo_lo};
  wire [1:0]        dataInWriteQueue_17_hi_lo = {|queueCount_5_17, |queueCount_4_17};
  wire [1:0]        dataInWriteQueue_17_hi_hi = {|queueCount_7_17, |queueCount_6_17};
  wire [3:0]        dataInWriteQueue_17_hi = {dataInWriteQueue_17_hi_hi, dataInWriteQueue_17_hi_lo};
  reg  [6:0]        queueCount_0_18;
  reg  [6:0]        queueCount_1_18;
  reg  [6:0]        queueCount_2_18;
  reg  [6:0]        queueCount_3_18;
  reg  [6:0]        queueCount_4_18;
  reg  [6:0]        queueCount_5_18;
  reg  [6:0]        queueCount_6_18;
  reg  [6:0]        queueCount_7_18;
  wire [7:0]        enqOH_18 = 8'h1 << writeQueueVec_18_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_18 = _probeWire_slots_18_writeValid_T ? enqOH_18 : 8'h0;
  wire              writeIndexQueue_18_deq_valid;
  assign writeIndexQueue_18_deq_valid = ~_writeIndexQueue_fifo_18_empty;
  wire              writeIndexQueue_18_enq_ready = ~_writeIndexQueue_fifo_18_full;
  wire              writeIndexQueue_18_enq_valid;
  assign writeIndexQueue_18_enq_valid = writeQueueVec_18_deq_ready & writeQueueVec_18_deq_valid;
  wire [2:0]        writeIndexQueue_18_deq_bits;
  wire [7:0]        queueDeq_18 = writeIndexQueue_18_deq_ready & writeIndexQueue_18_deq_valid ? 8'h1 << writeIndexQueue_18_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_144 = queueEnq_18[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_145 = queueEnq_18[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_146 = queueEnq_18[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_147 = queueEnq_18[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_148 = queueEnq_18[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_149 = queueEnq_18[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_150 = queueEnq_18[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_151 = queueEnq_18[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_18_lo_lo = {|queueCount_1_18, |queueCount_0_18};
  wire [1:0]        dataInWriteQueue_18_lo_hi = {|queueCount_3_18, |queueCount_2_18};
  wire [3:0]        dataInWriteQueue_18_lo = {dataInWriteQueue_18_lo_hi, dataInWriteQueue_18_lo_lo};
  wire [1:0]        dataInWriteQueue_18_hi_lo = {|queueCount_5_18, |queueCount_4_18};
  wire [1:0]        dataInWriteQueue_18_hi_hi = {|queueCount_7_18, |queueCount_6_18};
  wire [3:0]        dataInWriteQueue_18_hi = {dataInWriteQueue_18_hi_hi, dataInWriteQueue_18_hi_lo};
  reg  [6:0]        queueCount_0_19;
  reg  [6:0]        queueCount_1_19;
  reg  [6:0]        queueCount_2_19;
  reg  [6:0]        queueCount_3_19;
  reg  [6:0]        queueCount_4_19;
  reg  [6:0]        queueCount_5_19;
  reg  [6:0]        queueCount_6_19;
  reg  [6:0]        queueCount_7_19;
  wire [7:0]        enqOH_19 = 8'h1 << writeQueueVec_19_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_19 = _probeWire_slots_19_writeValid_T ? enqOH_19 : 8'h0;
  wire              writeIndexQueue_19_deq_valid;
  assign writeIndexQueue_19_deq_valid = ~_writeIndexQueue_fifo_19_empty;
  wire              writeIndexQueue_19_enq_ready = ~_writeIndexQueue_fifo_19_full;
  wire              writeIndexQueue_19_enq_valid;
  assign writeIndexQueue_19_enq_valid = writeQueueVec_19_deq_ready & writeQueueVec_19_deq_valid;
  wire [2:0]        writeIndexQueue_19_deq_bits;
  wire [7:0]        queueDeq_19 = writeIndexQueue_19_deq_ready & writeIndexQueue_19_deq_valid ? 8'h1 << writeIndexQueue_19_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_152 = queueEnq_19[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_153 = queueEnq_19[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_154 = queueEnq_19[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_155 = queueEnq_19[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_156 = queueEnq_19[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_157 = queueEnq_19[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_158 = queueEnq_19[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_159 = queueEnq_19[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_19_lo_lo = {|queueCount_1_19, |queueCount_0_19};
  wire [1:0]        dataInWriteQueue_19_lo_hi = {|queueCount_3_19, |queueCount_2_19};
  wire [3:0]        dataInWriteQueue_19_lo = {dataInWriteQueue_19_lo_hi, dataInWriteQueue_19_lo_lo};
  wire [1:0]        dataInWriteQueue_19_hi_lo = {|queueCount_5_19, |queueCount_4_19};
  wire [1:0]        dataInWriteQueue_19_hi_hi = {|queueCount_7_19, |queueCount_6_19};
  wire [3:0]        dataInWriteQueue_19_hi = {dataInWriteQueue_19_hi_hi, dataInWriteQueue_19_hi_lo};
  reg  [6:0]        queueCount_0_20;
  reg  [6:0]        queueCount_1_20;
  reg  [6:0]        queueCount_2_20;
  reg  [6:0]        queueCount_3_20;
  reg  [6:0]        queueCount_4_20;
  reg  [6:0]        queueCount_5_20;
  reg  [6:0]        queueCount_6_20;
  reg  [6:0]        queueCount_7_20;
  wire [7:0]        enqOH_20 = 8'h1 << writeQueueVec_20_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_20 = _probeWire_slots_20_writeValid_T ? enqOH_20 : 8'h0;
  wire              writeIndexQueue_20_deq_valid;
  assign writeIndexQueue_20_deq_valid = ~_writeIndexQueue_fifo_20_empty;
  wire              writeIndexQueue_20_enq_ready = ~_writeIndexQueue_fifo_20_full;
  wire              writeIndexQueue_20_enq_valid;
  assign writeIndexQueue_20_enq_valid = writeQueueVec_20_deq_ready & writeQueueVec_20_deq_valid;
  wire [2:0]        writeIndexQueue_20_deq_bits;
  wire [7:0]        queueDeq_20 = writeIndexQueue_20_deq_ready & writeIndexQueue_20_deq_valid ? 8'h1 << writeIndexQueue_20_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_160 = queueEnq_20[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_161 = queueEnq_20[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_162 = queueEnq_20[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_163 = queueEnq_20[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_164 = queueEnq_20[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_165 = queueEnq_20[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_166 = queueEnq_20[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_167 = queueEnq_20[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_20_lo_lo = {|queueCount_1_20, |queueCount_0_20};
  wire [1:0]        dataInWriteQueue_20_lo_hi = {|queueCount_3_20, |queueCount_2_20};
  wire [3:0]        dataInWriteQueue_20_lo = {dataInWriteQueue_20_lo_hi, dataInWriteQueue_20_lo_lo};
  wire [1:0]        dataInWriteQueue_20_hi_lo = {|queueCount_5_20, |queueCount_4_20};
  wire [1:0]        dataInWriteQueue_20_hi_hi = {|queueCount_7_20, |queueCount_6_20};
  wire [3:0]        dataInWriteQueue_20_hi = {dataInWriteQueue_20_hi_hi, dataInWriteQueue_20_hi_lo};
  reg  [6:0]        queueCount_0_21;
  reg  [6:0]        queueCount_1_21;
  reg  [6:0]        queueCount_2_21;
  reg  [6:0]        queueCount_3_21;
  reg  [6:0]        queueCount_4_21;
  reg  [6:0]        queueCount_5_21;
  reg  [6:0]        queueCount_6_21;
  reg  [6:0]        queueCount_7_21;
  wire [7:0]        enqOH_21 = 8'h1 << writeQueueVec_21_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_21 = _probeWire_slots_21_writeValid_T ? enqOH_21 : 8'h0;
  wire              writeIndexQueue_21_deq_valid;
  assign writeIndexQueue_21_deq_valid = ~_writeIndexQueue_fifo_21_empty;
  wire              writeIndexQueue_21_enq_ready = ~_writeIndexQueue_fifo_21_full;
  wire              writeIndexQueue_21_enq_valid;
  assign writeIndexQueue_21_enq_valid = writeQueueVec_21_deq_ready & writeQueueVec_21_deq_valid;
  wire [2:0]        writeIndexQueue_21_deq_bits;
  wire [7:0]        queueDeq_21 = writeIndexQueue_21_deq_ready & writeIndexQueue_21_deq_valid ? 8'h1 << writeIndexQueue_21_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_168 = queueEnq_21[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_169 = queueEnq_21[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_170 = queueEnq_21[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_171 = queueEnq_21[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_172 = queueEnq_21[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_173 = queueEnq_21[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_174 = queueEnq_21[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_175 = queueEnq_21[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_21_lo_lo = {|queueCount_1_21, |queueCount_0_21};
  wire [1:0]        dataInWriteQueue_21_lo_hi = {|queueCount_3_21, |queueCount_2_21};
  wire [3:0]        dataInWriteQueue_21_lo = {dataInWriteQueue_21_lo_hi, dataInWriteQueue_21_lo_lo};
  wire [1:0]        dataInWriteQueue_21_hi_lo = {|queueCount_5_21, |queueCount_4_21};
  wire [1:0]        dataInWriteQueue_21_hi_hi = {|queueCount_7_21, |queueCount_6_21};
  wire [3:0]        dataInWriteQueue_21_hi = {dataInWriteQueue_21_hi_hi, dataInWriteQueue_21_hi_lo};
  reg  [6:0]        queueCount_0_22;
  reg  [6:0]        queueCount_1_22;
  reg  [6:0]        queueCount_2_22;
  reg  [6:0]        queueCount_3_22;
  reg  [6:0]        queueCount_4_22;
  reg  [6:0]        queueCount_5_22;
  reg  [6:0]        queueCount_6_22;
  reg  [6:0]        queueCount_7_22;
  wire [7:0]        enqOH_22 = 8'h1 << writeQueueVec_22_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_22 = _probeWire_slots_22_writeValid_T ? enqOH_22 : 8'h0;
  wire              writeIndexQueue_22_deq_valid;
  assign writeIndexQueue_22_deq_valid = ~_writeIndexQueue_fifo_22_empty;
  wire              writeIndexQueue_22_enq_ready = ~_writeIndexQueue_fifo_22_full;
  wire              writeIndexQueue_22_enq_valid;
  assign writeIndexQueue_22_enq_valid = writeQueueVec_22_deq_ready & writeQueueVec_22_deq_valid;
  wire [2:0]        writeIndexQueue_22_deq_bits;
  wire [7:0]        queueDeq_22 = writeIndexQueue_22_deq_ready & writeIndexQueue_22_deq_valid ? 8'h1 << writeIndexQueue_22_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_176 = queueEnq_22[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_177 = queueEnq_22[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_178 = queueEnq_22[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_179 = queueEnq_22[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_180 = queueEnq_22[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_181 = queueEnq_22[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_182 = queueEnq_22[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_183 = queueEnq_22[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_22_lo_lo = {|queueCount_1_22, |queueCount_0_22};
  wire [1:0]        dataInWriteQueue_22_lo_hi = {|queueCount_3_22, |queueCount_2_22};
  wire [3:0]        dataInWriteQueue_22_lo = {dataInWriteQueue_22_lo_hi, dataInWriteQueue_22_lo_lo};
  wire [1:0]        dataInWriteQueue_22_hi_lo = {|queueCount_5_22, |queueCount_4_22};
  wire [1:0]        dataInWriteQueue_22_hi_hi = {|queueCount_7_22, |queueCount_6_22};
  wire [3:0]        dataInWriteQueue_22_hi = {dataInWriteQueue_22_hi_hi, dataInWriteQueue_22_hi_lo};
  reg  [6:0]        queueCount_0_23;
  reg  [6:0]        queueCount_1_23;
  reg  [6:0]        queueCount_2_23;
  reg  [6:0]        queueCount_3_23;
  reg  [6:0]        queueCount_4_23;
  reg  [6:0]        queueCount_5_23;
  reg  [6:0]        queueCount_6_23;
  reg  [6:0]        queueCount_7_23;
  wire [7:0]        enqOH_23 = 8'h1 << writeQueueVec_23_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_23 = _probeWire_slots_23_writeValid_T ? enqOH_23 : 8'h0;
  wire              writeIndexQueue_23_deq_valid;
  assign writeIndexQueue_23_deq_valid = ~_writeIndexQueue_fifo_23_empty;
  wire              writeIndexQueue_23_enq_ready = ~_writeIndexQueue_fifo_23_full;
  wire              writeIndexQueue_23_enq_valid;
  assign writeIndexQueue_23_enq_valid = writeQueueVec_23_deq_ready & writeQueueVec_23_deq_valid;
  wire [2:0]        writeIndexQueue_23_deq_bits;
  wire [7:0]        queueDeq_23 = writeIndexQueue_23_deq_ready & writeIndexQueue_23_deq_valid ? 8'h1 << writeIndexQueue_23_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_184 = queueEnq_23[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_185 = queueEnq_23[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_186 = queueEnq_23[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_187 = queueEnq_23[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_188 = queueEnq_23[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_189 = queueEnq_23[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_190 = queueEnq_23[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_191 = queueEnq_23[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_23_lo_lo = {|queueCount_1_23, |queueCount_0_23};
  wire [1:0]        dataInWriteQueue_23_lo_hi = {|queueCount_3_23, |queueCount_2_23};
  wire [3:0]        dataInWriteQueue_23_lo = {dataInWriteQueue_23_lo_hi, dataInWriteQueue_23_lo_lo};
  wire [1:0]        dataInWriteQueue_23_hi_lo = {|queueCount_5_23, |queueCount_4_23};
  wire [1:0]        dataInWriteQueue_23_hi_hi = {|queueCount_7_23, |queueCount_6_23};
  wire [3:0]        dataInWriteQueue_23_hi = {dataInWriteQueue_23_hi_hi, dataInWriteQueue_23_hi_lo};
  reg  [6:0]        queueCount_0_24;
  reg  [6:0]        queueCount_1_24;
  reg  [6:0]        queueCount_2_24;
  reg  [6:0]        queueCount_3_24;
  reg  [6:0]        queueCount_4_24;
  reg  [6:0]        queueCount_5_24;
  reg  [6:0]        queueCount_6_24;
  reg  [6:0]        queueCount_7_24;
  wire [7:0]        enqOH_24 = 8'h1 << writeQueueVec_24_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_24 = _probeWire_slots_24_writeValid_T ? enqOH_24 : 8'h0;
  wire              writeIndexQueue_24_deq_valid;
  assign writeIndexQueue_24_deq_valid = ~_writeIndexQueue_fifo_24_empty;
  wire              writeIndexQueue_24_enq_ready = ~_writeIndexQueue_fifo_24_full;
  wire              writeIndexQueue_24_enq_valid;
  assign writeIndexQueue_24_enq_valid = writeQueueVec_24_deq_ready & writeQueueVec_24_deq_valid;
  wire [2:0]        writeIndexQueue_24_deq_bits;
  wire [7:0]        queueDeq_24 = writeIndexQueue_24_deq_ready & writeIndexQueue_24_deq_valid ? 8'h1 << writeIndexQueue_24_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_192 = queueEnq_24[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_193 = queueEnq_24[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_194 = queueEnq_24[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_195 = queueEnq_24[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_196 = queueEnq_24[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_197 = queueEnq_24[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_198 = queueEnq_24[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_199 = queueEnq_24[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_24_lo_lo = {|queueCount_1_24, |queueCount_0_24};
  wire [1:0]        dataInWriteQueue_24_lo_hi = {|queueCount_3_24, |queueCount_2_24};
  wire [3:0]        dataInWriteQueue_24_lo = {dataInWriteQueue_24_lo_hi, dataInWriteQueue_24_lo_lo};
  wire [1:0]        dataInWriteQueue_24_hi_lo = {|queueCount_5_24, |queueCount_4_24};
  wire [1:0]        dataInWriteQueue_24_hi_hi = {|queueCount_7_24, |queueCount_6_24};
  wire [3:0]        dataInWriteQueue_24_hi = {dataInWriteQueue_24_hi_hi, dataInWriteQueue_24_hi_lo};
  reg  [6:0]        queueCount_0_25;
  reg  [6:0]        queueCount_1_25;
  reg  [6:0]        queueCount_2_25;
  reg  [6:0]        queueCount_3_25;
  reg  [6:0]        queueCount_4_25;
  reg  [6:0]        queueCount_5_25;
  reg  [6:0]        queueCount_6_25;
  reg  [6:0]        queueCount_7_25;
  wire [7:0]        enqOH_25 = 8'h1 << writeQueueVec_25_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_25 = _probeWire_slots_25_writeValid_T ? enqOH_25 : 8'h0;
  wire              writeIndexQueue_25_deq_valid;
  assign writeIndexQueue_25_deq_valid = ~_writeIndexQueue_fifo_25_empty;
  wire              writeIndexQueue_25_enq_ready = ~_writeIndexQueue_fifo_25_full;
  wire              writeIndexQueue_25_enq_valid;
  assign writeIndexQueue_25_enq_valid = writeQueueVec_25_deq_ready & writeQueueVec_25_deq_valid;
  wire [2:0]        writeIndexQueue_25_deq_bits;
  wire [7:0]        queueDeq_25 = writeIndexQueue_25_deq_ready & writeIndexQueue_25_deq_valid ? 8'h1 << writeIndexQueue_25_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_200 = queueEnq_25[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_201 = queueEnq_25[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_202 = queueEnq_25[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_203 = queueEnq_25[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_204 = queueEnq_25[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_205 = queueEnq_25[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_206 = queueEnq_25[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_207 = queueEnq_25[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_25_lo_lo = {|queueCount_1_25, |queueCount_0_25};
  wire [1:0]        dataInWriteQueue_25_lo_hi = {|queueCount_3_25, |queueCount_2_25};
  wire [3:0]        dataInWriteQueue_25_lo = {dataInWriteQueue_25_lo_hi, dataInWriteQueue_25_lo_lo};
  wire [1:0]        dataInWriteQueue_25_hi_lo = {|queueCount_5_25, |queueCount_4_25};
  wire [1:0]        dataInWriteQueue_25_hi_hi = {|queueCount_7_25, |queueCount_6_25};
  wire [3:0]        dataInWriteQueue_25_hi = {dataInWriteQueue_25_hi_hi, dataInWriteQueue_25_hi_lo};
  reg  [6:0]        queueCount_0_26;
  reg  [6:0]        queueCount_1_26;
  reg  [6:0]        queueCount_2_26;
  reg  [6:0]        queueCount_3_26;
  reg  [6:0]        queueCount_4_26;
  reg  [6:0]        queueCount_5_26;
  reg  [6:0]        queueCount_6_26;
  reg  [6:0]        queueCount_7_26;
  wire [7:0]        enqOH_26 = 8'h1 << writeQueueVec_26_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_26 = _probeWire_slots_26_writeValid_T ? enqOH_26 : 8'h0;
  wire              writeIndexQueue_26_deq_valid;
  assign writeIndexQueue_26_deq_valid = ~_writeIndexQueue_fifo_26_empty;
  wire              writeIndexQueue_26_enq_ready = ~_writeIndexQueue_fifo_26_full;
  wire              writeIndexQueue_26_enq_valid;
  assign writeIndexQueue_26_enq_valid = writeQueueVec_26_deq_ready & writeQueueVec_26_deq_valid;
  wire [2:0]        writeIndexQueue_26_deq_bits;
  wire [7:0]        queueDeq_26 = writeIndexQueue_26_deq_ready & writeIndexQueue_26_deq_valid ? 8'h1 << writeIndexQueue_26_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_208 = queueEnq_26[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_209 = queueEnq_26[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_210 = queueEnq_26[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_211 = queueEnq_26[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_212 = queueEnq_26[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_213 = queueEnq_26[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_214 = queueEnq_26[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_215 = queueEnq_26[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_26_lo_lo = {|queueCount_1_26, |queueCount_0_26};
  wire [1:0]        dataInWriteQueue_26_lo_hi = {|queueCount_3_26, |queueCount_2_26};
  wire [3:0]        dataInWriteQueue_26_lo = {dataInWriteQueue_26_lo_hi, dataInWriteQueue_26_lo_lo};
  wire [1:0]        dataInWriteQueue_26_hi_lo = {|queueCount_5_26, |queueCount_4_26};
  wire [1:0]        dataInWriteQueue_26_hi_hi = {|queueCount_7_26, |queueCount_6_26};
  wire [3:0]        dataInWriteQueue_26_hi = {dataInWriteQueue_26_hi_hi, dataInWriteQueue_26_hi_lo};
  reg  [6:0]        queueCount_0_27;
  reg  [6:0]        queueCount_1_27;
  reg  [6:0]        queueCount_2_27;
  reg  [6:0]        queueCount_3_27;
  reg  [6:0]        queueCount_4_27;
  reg  [6:0]        queueCount_5_27;
  reg  [6:0]        queueCount_6_27;
  reg  [6:0]        queueCount_7_27;
  wire [7:0]        enqOH_27 = 8'h1 << writeQueueVec_27_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_27 = _probeWire_slots_27_writeValid_T ? enqOH_27 : 8'h0;
  wire              writeIndexQueue_27_deq_valid;
  assign writeIndexQueue_27_deq_valid = ~_writeIndexQueue_fifo_27_empty;
  wire              writeIndexQueue_27_enq_ready = ~_writeIndexQueue_fifo_27_full;
  wire              writeIndexQueue_27_enq_valid;
  assign writeIndexQueue_27_enq_valid = writeQueueVec_27_deq_ready & writeQueueVec_27_deq_valid;
  wire [2:0]        writeIndexQueue_27_deq_bits;
  wire [7:0]        queueDeq_27 = writeIndexQueue_27_deq_ready & writeIndexQueue_27_deq_valid ? 8'h1 << writeIndexQueue_27_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_216 = queueEnq_27[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_217 = queueEnq_27[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_218 = queueEnq_27[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_219 = queueEnq_27[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_220 = queueEnq_27[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_221 = queueEnq_27[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_222 = queueEnq_27[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_223 = queueEnq_27[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_27_lo_lo = {|queueCount_1_27, |queueCount_0_27};
  wire [1:0]        dataInWriteQueue_27_lo_hi = {|queueCount_3_27, |queueCount_2_27};
  wire [3:0]        dataInWriteQueue_27_lo = {dataInWriteQueue_27_lo_hi, dataInWriteQueue_27_lo_lo};
  wire [1:0]        dataInWriteQueue_27_hi_lo = {|queueCount_5_27, |queueCount_4_27};
  wire [1:0]        dataInWriteQueue_27_hi_hi = {|queueCount_7_27, |queueCount_6_27};
  wire [3:0]        dataInWriteQueue_27_hi = {dataInWriteQueue_27_hi_hi, dataInWriteQueue_27_hi_lo};
  reg  [6:0]        queueCount_0_28;
  reg  [6:0]        queueCount_1_28;
  reg  [6:0]        queueCount_2_28;
  reg  [6:0]        queueCount_3_28;
  reg  [6:0]        queueCount_4_28;
  reg  [6:0]        queueCount_5_28;
  reg  [6:0]        queueCount_6_28;
  reg  [6:0]        queueCount_7_28;
  wire [7:0]        enqOH_28 = 8'h1 << writeQueueVec_28_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_28 = _probeWire_slots_28_writeValid_T ? enqOH_28 : 8'h0;
  wire              writeIndexQueue_28_deq_valid;
  assign writeIndexQueue_28_deq_valid = ~_writeIndexQueue_fifo_28_empty;
  wire              writeIndexQueue_28_enq_ready = ~_writeIndexQueue_fifo_28_full;
  wire              writeIndexQueue_28_enq_valid;
  assign writeIndexQueue_28_enq_valid = writeQueueVec_28_deq_ready & writeQueueVec_28_deq_valid;
  wire [2:0]        writeIndexQueue_28_deq_bits;
  wire [7:0]        queueDeq_28 = writeIndexQueue_28_deq_ready & writeIndexQueue_28_deq_valid ? 8'h1 << writeIndexQueue_28_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_224 = queueEnq_28[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_225 = queueEnq_28[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_226 = queueEnq_28[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_227 = queueEnq_28[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_228 = queueEnq_28[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_229 = queueEnq_28[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_230 = queueEnq_28[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_231 = queueEnq_28[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_28_lo_lo = {|queueCount_1_28, |queueCount_0_28};
  wire [1:0]        dataInWriteQueue_28_lo_hi = {|queueCount_3_28, |queueCount_2_28};
  wire [3:0]        dataInWriteQueue_28_lo = {dataInWriteQueue_28_lo_hi, dataInWriteQueue_28_lo_lo};
  wire [1:0]        dataInWriteQueue_28_hi_lo = {|queueCount_5_28, |queueCount_4_28};
  wire [1:0]        dataInWriteQueue_28_hi_hi = {|queueCount_7_28, |queueCount_6_28};
  wire [3:0]        dataInWriteQueue_28_hi = {dataInWriteQueue_28_hi_hi, dataInWriteQueue_28_hi_lo};
  reg  [6:0]        queueCount_0_29;
  reg  [6:0]        queueCount_1_29;
  reg  [6:0]        queueCount_2_29;
  reg  [6:0]        queueCount_3_29;
  reg  [6:0]        queueCount_4_29;
  reg  [6:0]        queueCount_5_29;
  reg  [6:0]        queueCount_6_29;
  reg  [6:0]        queueCount_7_29;
  wire [7:0]        enqOH_29 = 8'h1 << writeQueueVec_29_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_29 = _probeWire_slots_29_writeValid_T ? enqOH_29 : 8'h0;
  wire              writeIndexQueue_29_deq_valid;
  assign writeIndexQueue_29_deq_valid = ~_writeIndexQueue_fifo_29_empty;
  wire              writeIndexQueue_29_enq_ready = ~_writeIndexQueue_fifo_29_full;
  wire              writeIndexQueue_29_enq_valid;
  assign writeIndexQueue_29_enq_valid = writeQueueVec_29_deq_ready & writeQueueVec_29_deq_valid;
  wire [2:0]        writeIndexQueue_29_deq_bits;
  wire [7:0]        queueDeq_29 = writeIndexQueue_29_deq_ready & writeIndexQueue_29_deq_valid ? 8'h1 << writeIndexQueue_29_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_232 = queueEnq_29[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_233 = queueEnq_29[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_234 = queueEnq_29[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_235 = queueEnq_29[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_236 = queueEnq_29[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_237 = queueEnq_29[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_238 = queueEnq_29[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_239 = queueEnq_29[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_29_lo_lo = {|queueCount_1_29, |queueCount_0_29};
  wire [1:0]        dataInWriteQueue_29_lo_hi = {|queueCount_3_29, |queueCount_2_29};
  wire [3:0]        dataInWriteQueue_29_lo = {dataInWriteQueue_29_lo_hi, dataInWriteQueue_29_lo_lo};
  wire [1:0]        dataInWriteQueue_29_hi_lo = {|queueCount_5_29, |queueCount_4_29};
  wire [1:0]        dataInWriteQueue_29_hi_hi = {|queueCount_7_29, |queueCount_6_29};
  wire [3:0]        dataInWriteQueue_29_hi = {dataInWriteQueue_29_hi_hi, dataInWriteQueue_29_hi_lo};
  reg  [6:0]        queueCount_0_30;
  reg  [6:0]        queueCount_1_30;
  reg  [6:0]        queueCount_2_30;
  reg  [6:0]        queueCount_3_30;
  reg  [6:0]        queueCount_4_30;
  reg  [6:0]        queueCount_5_30;
  reg  [6:0]        queueCount_6_30;
  reg  [6:0]        queueCount_7_30;
  wire [7:0]        enqOH_30 = 8'h1 << writeQueueVec_30_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_30 = _probeWire_slots_30_writeValid_T ? enqOH_30 : 8'h0;
  wire              writeIndexQueue_30_deq_valid;
  assign writeIndexQueue_30_deq_valid = ~_writeIndexQueue_fifo_30_empty;
  wire              writeIndexQueue_30_enq_ready = ~_writeIndexQueue_fifo_30_full;
  wire              writeIndexQueue_30_enq_valid;
  assign writeIndexQueue_30_enq_valid = writeQueueVec_30_deq_ready & writeQueueVec_30_deq_valid;
  wire [2:0]        writeIndexQueue_30_deq_bits;
  wire [7:0]        queueDeq_30 = writeIndexQueue_30_deq_ready & writeIndexQueue_30_deq_valid ? 8'h1 << writeIndexQueue_30_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_240 = queueEnq_30[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_241 = queueEnq_30[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_242 = queueEnq_30[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_243 = queueEnq_30[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_244 = queueEnq_30[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_245 = queueEnq_30[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_246 = queueEnq_30[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_247 = queueEnq_30[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_30_lo_lo = {|queueCount_1_30, |queueCount_0_30};
  wire [1:0]        dataInWriteQueue_30_lo_hi = {|queueCount_3_30, |queueCount_2_30};
  wire [3:0]        dataInWriteQueue_30_lo = {dataInWriteQueue_30_lo_hi, dataInWriteQueue_30_lo_lo};
  wire [1:0]        dataInWriteQueue_30_hi_lo = {|queueCount_5_30, |queueCount_4_30};
  wire [1:0]        dataInWriteQueue_30_hi_hi = {|queueCount_7_30, |queueCount_6_30};
  wire [3:0]        dataInWriteQueue_30_hi = {dataInWriteQueue_30_hi_hi, dataInWriteQueue_30_hi_lo};
  reg  [6:0]        queueCount_0_31;
  reg  [6:0]        queueCount_1_31;
  reg  [6:0]        queueCount_2_31;
  reg  [6:0]        queueCount_3_31;
  reg  [6:0]        queueCount_4_31;
  reg  [6:0]        queueCount_5_31;
  reg  [6:0]        queueCount_6_31;
  reg  [6:0]        queueCount_7_31;
  wire [7:0]        enqOH_31 = 8'h1 << writeQueueVec_31_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_31 = _probeWire_slots_31_writeValid_T ? enqOH_31 : 8'h0;
  wire              writeIndexQueue_31_deq_valid;
  assign writeIndexQueue_31_deq_valid = ~_writeIndexQueue_fifo_31_empty;
  wire              writeIndexQueue_31_enq_ready = ~_writeIndexQueue_fifo_31_full;
  wire              writeIndexQueue_31_enq_valid;
  assign writeIndexQueue_31_enq_valid = writeQueueVec_31_deq_ready & writeQueueVec_31_deq_valid;
  wire [2:0]        writeIndexQueue_31_deq_bits;
  wire [7:0]        queueDeq_31 = writeIndexQueue_31_deq_ready & writeIndexQueue_31_deq_valid ? 8'h1 << writeIndexQueue_31_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_248 = queueEnq_31[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_249 = queueEnq_31[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_250 = queueEnq_31[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_251 = queueEnq_31[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_252 = queueEnq_31[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_253 = queueEnq_31[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_254 = queueEnq_31[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_255 = queueEnq_31[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_31_lo_lo = {|queueCount_1_31, |queueCount_0_31};
  wire [1:0]        dataInWriteQueue_31_lo_hi = {|queueCount_3_31, |queueCount_2_31};
  wire [3:0]        dataInWriteQueue_31_lo = {dataInWriteQueue_31_lo_hi, dataInWriteQueue_31_lo_lo};
  wire [1:0]        dataInWriteQueue_31_hi_lo = {|queueCount_5_31, |queueCount_4_31};
  wire [1:0]        dataInWriteQueue_31_hi_hi = {|queueCount_7_31, |queueCount_6_31};
  wire [3:0]        dataInWriteQueue_31_hi = {dataInWriteQueue_31_hi_hi, dataInWriteQueue_31_hi_lo};
  wire              sourceQueue_deq_valid;
  assign sourceQueue_deq_valid = ~_sourceQueue_fifo_empty;
  wire              sourceQueue_enq_ready = ~_sourceQueue_fifo_full;
  wire              sourceQueue_enq_valid;
  wire              sourceQueue_deq_ready;
  wire              axi4Port_ar_valid_0 = _loadUnit_memRequest_valid & sourceQueue_enq_ready;
  wire              axi4Port_r_ready_0;
  assign sourceQueue_enq_valid = _loadUnit_memRequest_valid & axi4Port_ar_ready_0;
  assign sourceQueue_deq_ready = axi4Port_r_ready_0 & axi4Port_r_valid_0;
  assign dataQueue_deq_valid = ~_dataQueue_fifo_empty;
  wire              axi4Port_w_valid_0 = dataQueue_deq_valid;
  wire [1023:0]     dataQueue_dataOut_data;
  wire [1023:0]     axi4Port_w_bits_data_0 = dataQueue_deq_bits_data;
  wire [127:0]      dataQueue_dataOut_mask;
  wire [127:0]      axi4Port_w_bits_strb_0 = dataQueue_deq_bits_mask;
  wire [3:0]        dataQueue_dataOut_index;
  wire [31:0]       dataQueue_dataOut_address;
  wire [3:0]        dataQueue_enq_bits_index;
  wire [31:0]       dataQueue_enq_bits_address;
  wire [35:0]       dataQueue_dataIn_lo = {dataQueue_enq_bits_index, dataQueue_enq_bits_address};
  wire [1023:0]     dataQueue_enq_bits_data;
  wire [127:0]      dataQueue_enq_bits_mask;
  wire [1151:0]     dataQueue_dataIn_hi = {dataQueue_enq_bits_data, dataQueue_enq_bits_mask};
  wire [1187:0]     dataQueue_dataIn = {dataQueue_dataIn_hi, dataQueue_dataIn_lo};
  assign dataQueue_dataOut_address = _dataQueue_fifo_data_out[31:0];
  assign dataQueue_dataOut_index = _dataQueue_fifo_data_out[35:32];
  assign dataQueue_dataOut_mask = _dataQueue_fifo_data_out[163:36];
  assign dataQueue_dataOut_data = _dataQueue_fifo_data_out[1187:164];
  assign dataQueue_deq_bits_data = dataQueue_dataOut_data;
  assign dataQueue_deq_bits_mask = dataQueue_dataOut_mask;
  wire [3:0]        dataQueue_deq_bits_index = dataQueue_dataOut_index;
  wire [31:0]       dataQueue_deq_bits_address = dataQueue_dataOut_address;
  wire              dataQueue_enq_ready = ~_dataQueue_fifo_full;
  wire              dataQueue_enq_valid;
  wire              axi4Port_aw_valid_0 = _storeUnit_memRequest_valid & dataQueue_enq_ready;
  wire [1:0]        axi4Port_aw_bits_id_0 = _storeUnit_memRequest_bits_index[1:0];
  assign dataQueue_enq_valid = _storeUnit_memRequest_valid & axi4Port_aw_ready_0;
  wire              simpleSourceQueue_deq_valid;
  assign simpleSourceQueue_deq_valid = ~_simpleSourceQueue_fifo_empty;
  wire              simpleSourceQueue_enq_ready = ~_simpleSourceQueue_fifo_full;
  wire              simpleSourceQueue_enq_valid;
  wire              simpleSourceQueue_deq_ready;
  wire              simpleAccessPorts_ar_valid_0 = _otherUnit_memReadRequest_valid & simpleSourceQueue_enq_ready;
  wire              simpleAccessPorts_r_ready_0;
  assign simpleSourceQueue_enq_valid = _otherUnit_memReadRequest_valid & simpleAccessPorts_ar_ready_0;
  assign simpleSourceQueue_deq_ready = simpleAccessPorts_r_ready_0 & simpleAccessPorts_r_valid_0;
  assign simpleDataQueue_deq_valid = ~_simpleDataQueue_fifo_empty;
  wire              simpleAccessPorts_w_valid_0 = simpleDataQueue_deq_valid;
  wire [31:0]       simpleDataQueue_dataOut_data;
  wire [31:0]       simpleAccessPorts_w_bits_data_0 = simpleDataQueue_deq_bits_data;
  wire [3:0]        simpleDataQueue_dataOut_mask;
  wire [3:0]        simpleAccessPorts_w_bits_strb_0 = simpleDataQueue_deq_bits_mask;
  wire [7:0]        simpleDataQueue_dataOut_source;
  wire [31:0]       simpleDataQueue_dataOut_address;
  wire [1:0]        simpleDataQueue_dataOut_size;
  wire [31:0]       simpleDataQueue_enq_bits_address;
  wire [1:0]        simpleDataQueue_enq_bits_size;
  wire [33:0]       simpleDataQueue_dataIn_lo = {simpleDataQueue_enq_bits_address, simpleDataQueue_enq_bits_size};
  wire [31:0]       simpleDataQueue_enq_bits_data;
  wire [3:0]        simpleDataQueue_enq_bits_mask;
  wire [35:0]       simpleDataQueue_dataIn_hi_hi = {simpleDataQueue_enq_bits_data, simpleDataQueue_enq_bits_mask};
  wire [7:0]        simpleDataQueue_enq_bits_source;
  wire [43:0]       simpleDataQueue_dataIn_hi = {simpleDataQueue_dataIn_hi_hi, simpleDataQueue_enq_bits_source};
  wire [77:0]       simpleDataQueue_dataIn = {simpleDataQueue_dataIn_hi, simpleDataQueue_dataIn_lo};
  assign simpleDataQueue_dataOut_size = _simpleDataQueue_fifo_data_out[1:0];
  assign simpleDataQueue_dataOut_address = _simpleDataQueue_fifo_data_out[33:2];
  assign simpleDataQueue_dataOut_source = _simpleDataQueue_fifo_data_out[41:34];
  assign simpleDataQueue_dataOut_mask = _simpleDataQueue_fifo_data_out[45:42];
  assign simpleDataQueue_dataOut_data = _simpleDataQueue_fifo_data_out[77:46];
  assign simpleDataQueue_deq_bits_data = simpleDataQueue_dataOut_data;
  assign simpleDataQueue_deq_bits_mask = simpleDataQueue_dataOut_mask;
  wire [7:0]        simpleDataQueue_deq_bits_source = simpleDataQueue_dataOut_source;
  wire [31:0]       simpleDataQueue_deq_bits_address = simpleDataQueue_dataOut_address;
  wire [1:0]        simpleDataQueue_deq_bits_size = simpleDataQueue_dataOut_size;
  wire              simpleDataQueue_enq_ready = ~_simpleDataQueue_fifo_full;
  wire              simpleDataQueue_enq_valid;
  wire              simpleAccessPorts_aw_valid_0 = _otherUnit_memWriteRequest_valid & dataQueue_enq_ready;
  wire [2:0]        simpleAccessPorts_aw_bits_size_0 = {1'h0, _otherUnit_memWriteRequest_bits_size};
  wire [1:0]        simpleAccessPorts_aw_bits_id_0 = _otherUnit_memWriteRequest_bits_source[1:0];
  assign simpleDataQueue_enq_valid = _otherUnit_memWriteRequest_valid & simpleAccessPorts_aw_ready_0;
  wire [1:0]        tokenIO_offsetGroupRelease_lo_lo_lo_lo = {_otherUnit_offsetRelease_1, _otherUnit_offsetRelease_0};
  wire [1:0]        tokenIO_offsetGroupRelease_lo_lo_lo_hi = {_otherUnit_offsetRelease_3, _otherUnit_offsetRelease_2};
  wire [3:0]        tokenIO_offsetGroupRelease_lo_lo_lo = {tokenIO_offsetGroupRelease_lo_lo_lo_hi, tokenIO_offsetGroupRelease_lo_lo_lo_lo};
  wire [1:0]        tokenIO_offsetGroupRelease_lo_lo_hi_lo = {_otherUnit_offsetRelease_5, _otherUnit_offsetRelease_4};
  wire [1:0]        tokenIO_offsetGroupRelease_lo_lo_hi_hi = {_otherUnit_offsetRelease_7, _otherUnit_offsetRelease_6};
  wire [3:0]        tokenIO_offsetGroupRelease_lo_lo_hi = {tokenIO_offsetGroupRelease_lo_lo_hi_hi, tokenIO_offsetGroupRelease_lo_lo_hi_lo};
  wire [7:0]        tokenIO_offsetGroupRelease_lo_lo = {tokenIO_offsetGroupRelease_lo_lo_hi, tokenIO_offsetGroupRelease_lo_lo_lo};
  wire [1:0]        tokenIO_offsetGroupRelease_lo_hi_lo_lo = {_otherUnit_offsetRelease_9, _otherUnit_offsetRelease_8};
  wire [1:0]        tokenIO_offsetGroupRelease_lo_hi_lo_hi = {_otherUnit_offsetRelease_11, _otherUnit_offsetRelease_10};
  wire [3:0]        tokenIO_offsetGroupRelease_lo_hi_lo = {tokenIO_offsetGroupRelease_lo_hi_lo_hi, tokenIO_offsetGroupRelease_lo_hi_lo_lo};
  wire [1:0]        tokenIO_offsetGroupRelease_lo_hi_hi_lo = {_otherUnit_offsetRelease_13, _otherUnit_offsetRelease_12};
  wire [1:0]        tokenIO_offsetGroupRelease_lo_hi_hi_hi = {_otherUnit_offsetRelease_15, _otherUnit_offsetRelease_14};
  wire [3:0]        tokenIO_offsetGroupRelease_lo_hi_hi = {tokenIO_offsetGroupRelease_lo_hi_hi_hi, tokenIO_offsetGroupRelease_lo_hi_hi_lo};
  wire [7:0]        tokenIO_offsetGroupRelease_lo_hi = {tokenIO_offsetGroupRelease_lo_hi_hi, tokenIO_offsetGroupRelease_lo_hi_lo};
  wire [15:0]       tokenIO_offsetGroupRelease_lo = {tokenIO_offsetGroupRelease_lo_hi, tokenIO_offsetGroupRelease_lo_lo};
  wire [1:0]        tokenIO_offsetGroupRelease_hi_lo_lo_lo = {_otherUnit_offsetRelease_17, _otherUnit_offsetRelease_16};
  wire [1:0]        tokenIO_offsetGroupRelease_hi_lo_lo_hi = {_otherUnit_offsetRelease_19, _otherUnit_offsetRelease_18};
  wire [3:0]        tokenIO_offsetGroupRelease_hi_lo_lo = {tokenIO_offsetGroupRelease_hi_lo_lo_hi, tokenIO_offsetGroupRelease_hi_lo_lo_lo};
  wire [1:0]        tokenIO_offsetGroupRelease_hi_lo_hi_lo = {_otherUnit_offsetRelease_21, _otherUnit_offsetRelease_20};
  wire [1:0]        tokenIO_offsetGroupRelease_hi_lo_hi_hi = {_otherUnit_offsetRelease_23, _otherUnit_offsetRelease_22};
  wire [3:0]        tokenIO_offsetGroupRelease_hi_lo_hi = {tokenIO_offsetGroupRelease_hi_lo_hi_hi, tokenIO_offsetGroupRelease_hi_lo_hi_lo};
  wire [7:0]        tokenIO_offsetGroupRelease_hi_lo = {tokenIO_offsetGroupRelease_hi_lo_hi, tokenIO_offsetGroupRelease_hi_lo_lo};
  wire [1:0]        tokenIO_offsetGroupRelease_hi_hi_lo_lo = {_otherUnit_offsetRelease_25, _otherUnit_offsetRelease_24};
  wire [1:0]        tokenIO_offsetGroupRelease_hi_hi_lo_hi = {_otherUnit_offsetRelease_27, _otherUnit_offsetRelease_26};
  wire [3:0]        tokenIO_offsetGroupRelease_hi_hi_lo = {tokenIO_offsetGroupRelease_hi_hi_lo_hi, tokenIO_offsetGroupRelease_hi_hi_lo_lo};
  wire [1:0]        tokenIO_offsetGroupRelease_hi_hi_hi_lo = {_otherUnit_offsetRelease_29, _otherUnit_offsetRelease_28};
  wire [1:0]        tokenIO_offsetGroupRelease_hi_hi_hi_hi = {_otherUnit_offsetRelease_31, _otherUnit_offsetRelease_30};
  wire [3:0]        tokenIO_offsetGroupRelease_hi_hi_hi = {tokenIO_offsetGroupRelease_hi_hi_hi_hi, tokenIO_offsetGroupRelease_hi_hi_hi_lo};
  wire [7:0]        tokenIO_offsetGroupRelease_hi_hi = {tokenIO_offsetGroupRelease_hi_hi_hi, tokenIO_offsetGroupRelease_hi_hi_lo};
  wire [15:0]       tokenIO_offsetGroupRelease_hi = {tokenIO_offsetGroupRelease_hi_hi, tokenIO_offsetGroupRelease_hi_lo};
  wire              unitOrder =
    _loadUnit_status_instructionIndex == _storeUnit_status_instructionIndex | _loadUnit_status_instructionIndex[1:0] < _storeUnit_status_instructionIndex[1:0] ^ _loadUnit_status_instructionIndex[2] ^ _storeUnit_status_instructionIndex[2];
  wire              loadAddressConflict = _loadUnit_status_startAddress >= _storeUnit_status_startAddress & _loadUnit_status_startAddress <= _storeUnit_status_endAddress;
  wire              storeAddressConflict = _storeUnit_status_startAddress >= _loadUnit_status_startAddress & _storeUnit_status_startAddress <= _loadUnit_status_endAddress;
  wire              stallLoad = ~unitOrder & loadAddressConflict & ~_storeUnit_status_idle;
  wire              stallStore = unitOrder & storeAddressConflict & ~_loadUnit_status_idle;
  always @(posedge clock) begin
    if (reset) begin
      v0_0 <= 32'h0;
      v0_1 <= 32'h0;
      v0_2 <= 32'h0;
      v0_3 <= 32'h0;
      v0_4 <= 32'h0;
      v0_5 <= 32'h0;
      v0_6 <= 32'h0;
      v0_7 <= 32'h0;
      v0_8 <= 32'h0;
      v0_9 <= 32'h0;
      v0_10 <= 32'h0;
      v0_11 <= 32'h0;
      v0_12 <= 32'h0;
      v0_13 <= 32'h0;
      v0_14 <= 32'h0;
      v0_15 <= 32'h0;
      v0_16 <= 32'h0;
      v0_17 <= 32'h0;
      v0_18 <= 32'h0;
      v0_19 <= 32'h0;
      v0_20 <= 32'h0;
      v0_21 <= 32'h0;
      v0_22 <= 32'h0;
      v0_23 <= 32'h0;
      v0_24 <= 32'h0;
      v0_25 <= 32'h0;
      v0_26 <= 32'h0;
      v0_27 <= 32'h0;
      v0_28 <= 32'h0;
      v0_29 <= 32'h0;
      v0_30 <= 32'h0;
      v0_31 <= 32'h0;
      queueCount_0 <= 7'h0;
      queueCount_1 <= 7'h0;
      queueCount_2 <= 7'h0;
      queueCount_3 <= 7'h0;
      queueCount_4 <= 7'h0;
      queueCount_5 <= 7'h0;
      queueCount_6 <= 7'h0;
      queueCount_7 <= 7'h0;
      queueCount_0_1 <= 7'h0;
      queueCount_1_1 <= 7'h0;
      queueCount_2_1 <= 7'h0;
      queueCount_3_1 <= 7'h0;
      queueCount_4_1 <= 7'h0;
      queueCount_5_1 <= 7'h0;
      queueCount_6_1 <= 7'h0;
      queueCount_7_1 <= 7'h0;
      queueCount_0_2 <= 7'h0;
      queueCount_1_2 <= 7'h0;
      queueCount_2_2 <= 7'h0;
      queueCount_3_2 <= 7'h0;
      queueCount_4_2 <= 7'h0;
      queueCount_5_2 <= 7'h0;
      queueCount_6_2 <= 7'h0;
      queueCount_7_2 <= 7'h0;
      queueCount_0_3 <= 7'h0;
      queueCount_1_3 <= 7'h0;
      queueCount_2_3 <= 7'h0;
      queueCount_3_3 <= 7'h0;
      queueCount_4_3 <= 7'h0;
      queueCount_5_3 <= 7'h0;
      queueCount_6_3 <= 7'h0;
      queueCount_7_3 <= 7'h0;
      queueCount_0_4 <= 7'h0;
      queueCount_1_4 <= 7'h0;
      queueCount_2_4 <= 7'h0;
      queueCount_3_4 <= 7'h0;
      queueCount_4_4 <= 7'h0;
      queueCount_5_4 <= 7'h0;
      queueCount_6_4 <= 7'h0;
      queueCount_7_4 <= 7'h0;
      queueCount_0_5 <= 7'h0;
      queueCount_1_5 <= 7'h0;
      queueCount_2_5 <= 7'h0;
      queueCount_3_5 <= 7'h0;
      queueCount_4_5 <= 7'h0;
      queueCount_5_5 <= 7'h0;
      queueCount_6_5 <= 7'h0;
      queueCount_7_5 <= 7'h0;
      queueCount_0_6 <= 7'h0;
      queueCount_1_6 <= 7'h0;
      queueCount_2_6 <= 7'h0;
      queueCount_3_6 <= 7'h0;
      queueCount_4_6 <= 7'h0;
      queueCount_5_6 <= 7'h0;
      queueCount_6_6 <= 7'h0;
      queueCount_7_6 <= 7'h0;
      queueCount_0_7 <= 7'h0;
      queueCount_1_7 <= 7'h0;
      queueCount_2_7 <= 7'h0;
      queueCount_3_7 <= 7'h0;
      queueCount_4_7 <= 7'h0;
      queueCount_5_7 <= 7'h0;
      queueCount_6_7 <= 7'h0;
      queueCount_7_7 <= 7'h0;
      queueCount_0_8 <= 7'h0;
      queueCount_1_8 <= 7'h0;
      queueCount_2_8 <= 7'h0;
      queueCount_3_8 <= 7'h0;
      queueCount_4_8 <= 7'h0;
      queueCount_5_8 <= 7'h0;
      queueCount_6_8 <= 7'h0;
      queueCount_7_8 <= 7'h0;
      queueCount_0_9 <= 7'h0;
      queueCount_1_9 <= 7'h0;
      queueCount_2_9 <= 7'h0;
      queueCount_3_9 <= 7'h0;
      queueCount_4_9 <= 7'h0;
      queueCount_5_9 <= 7'h0;
      queueCount_6_9 <= 7'h0;
      queueCount_7_9 <= 7'h0;
      queueCount_0_10 <= 7'h0;
      queueCount_1_10 <= 7'h0;
      queueCount_2_10 <= 7'h0;
      queueCount_3_10 <= 7'h0;
      queueCount_4_10 <= 7'h0;
      queueCount_5_10 <= 7'h0;
      queueCount_6_10 <= 7'h0;
      queueCount_7_10 <= 7'h0;
      queueCount_0_11 <= 7'h0;
      queueCount_1_11 <= 7'h0;
      queueCount_2_11 <= 7'h0;
      queueCount_3_11 <= 7'h0;
      queueCount_4_11 <= 7'h0;
      queueCount_5_11 <= 7'h0;
      queueCount_6_11 <= 7'h0;
      queueCount_7_11 <= 7'h0;
      queueCount_0_12 <= 7'h0;
      queueCount_1_12 <= 7'h0;
      queueCount_2_12 <= 7'h0;
      queueCount_3_12 <= 7'h0;
      queueCount_4_12 <= 7'h0;
      queueCount_5_12 <= 7'h0;
      queueCount_6_12 <= 7'h0;
      queueCount_7_12 <= 7'h0;
      queueCount_0_13 <= 7'h0;
      queueCount_1_13 <= 7'h0;
      queueCount_2_13 <= 7'h0;
      queueCount_3_13 <= 7'h0;
      queueCount_4_13 <= 7'h0;
      queueCount_5_13 <= 7'h0;
      queueCount_6_13 <= 7'h0;
      queueCount_7_13 <= 7'h0;
      queueCount_0_14 <= 7'h0;
      queueCount_1_14 <= 7'h0;
      queueCount_2_14 <= 7'h0;
      queueCount_3_14 <= 7'h0;
      queueCount_4_14 <= 7'h0;
      queueCount_5_14 <= 7'h0;
      queueCount_6_14 <= 7'h0;
      queueCount_7_14 <= 7'h0;
      queueCount_0_15 <= 7'h0;
      queueCount_1_15 <= 7'h0;
      queueCount_2_15 <= 7'h0;
      queueCount_3_15 <= 7'h0;
      queueCount_4_15 <= 7'h0;
      queueCount_5_15 <= 7'h0;
      queueCount_6_15 <= 7'h0;
      queueCount_7_15 <= 7'h0;
      queueCount_0_16 <= 7'h0;
      queueCount_1_16 <= 7'h0;
      queueCount_2_16 <= 7'h0;
      queueCount_3_16 <= 7'h0;
      queueCount_4_16 <= 7'h0;
      queueCount_5_16 <= 7'h0;
      queueCount_6_16 <= 7'h0;
      queueCount_7_16 <= 7'h0;
      queueCount_0_17 <= 7'h0;
      queueCount_1_17 <= 7'h0;
      queueCount_2_17 <= 7'h0;
      queueCount_3_17 <= 7'h0;
      queueCount_4_17 <= 7'h0;
      queueCount_5_17 <= 7'h0;
      queueCount_6_17 <= 7'h0;
      queueCount_7_17 <= 7'h0;
      queueCount_0_18 <= 7'h0;
      queueCount_1_18 <= 7'h0;
      queueCount_2_18 <= 7'h0;
      queueCount_3_18 <= 7'h0;
      queueCount_4_18 <= 7'h0;
      queueCount_5_18 <= 7'h0;
      queueCount_6_18 <= 7'h0;
      queueCount_7_18 <= 7'h0;
      queueCount_0_19 <= 7'h0;
      queueCount_1_19 <= 7'h0;
      queueCount_2_19 <= 7'h0;
      queueCount_3_19 <= 7'h0;
      queueCount_4_19 <= 7'h0;
      queueCount_5_19 <= 7'h0;
      queueCount_6_19 <= 7'h0;
      queueCount_7_19 <= 7'h0;
      queueCount_0_20 <= 7'h0;
      queueCount_1_20 <= 7'h0;
      queueCount_2_20 <= 7'h0;
      queueCount_3_20 <= 7'h0;
      queueCount_4_20 <= 7'h0;
      queueCount_5_20 <= 7'h0;
      queueCount_6_20 <= 7'h0;
      queueCount_7_20 <= 7'h0;
      queueCount_0_21 <= 7'h0;
      queueCount_1_21 <= 7'h0;
      queueCount_2_21 <= 7'h0;
      queueCount_3_21 <= 7'h0;
      queueCount_4_21 <= 7'h0;
      queueCount_5_21 <= 7'h0;
      queueCount_6_21 <= 7'h0;
      queueCount_7_21 <= 7'h0;
      queueCount_0_22 <= 7'h0;
      queueCount_1_22 <= 7'h0;
      queueCount_2_22 <= 7'h0;
      queueCount_3_22 <= 7'h0;
      queueCount_4_22 <= 7'h0;
      queueCount_5_22 <= 7'h0;
      queueCount_6_22 <= 7'h0;
      queueCount_7_22 <= 7'h0;
      queueCount_0_23 <= 7'h0;
      queueCount_1_23 <= 7'h0;
      queueCount_2_23 <= 7'h0;
      queueCount_3_23 <= 7'h0;
      queueCount_4_23 <= 7'h0;
      queueCount_5_23 <= 7'h0;
      queueCount_6_23 <= 7'h0;
      queueCount_7_23 <= 7'h0;
      queueCount_0_24 <= 7'h0;
      queueCount_1_24 <= 7'h0;
      queueCount_2_24 <= 7'h0;
      queueCount_3_24 <= 7'h0;
      queueCount_4_24 <= 7'h0;
      queueCount_5_24 <= 7'h0;
      queueCount_6_24 <= 7'h0;
      queueCount_7_24 <= 7'h0;
      queueCount_0_25 <= 7'h0;
      queueCount_1_25 <= 7'h0;
      queueCount_2_25 <= 7'h0;
      queueCount_3_25 <= 7'h0;
      queueCount_4_25 <= 7'h0;
      queueCount_5_25 <= 7'h0;
      queueCount_6_25 <= 7'h0;
      queueCount_7_25 <= 7'h0;
      queueCount_0_26 <= 7'h0;
      queueCount_1_26 <= 7'h0;
      queueCount_2_26 <= 7'h0;
      queueCount_3_26 <= 7'h0;
      queueCount_4_26 <= 7'h0;
      queueCount_5_26 <= 7'h0;
      queueCount_6_26 <= 7'h0;
      queueCount_7_26 <= 7'h0;
      queueCount_0_27 <= 7'h0;
      queueCount_1_27 <= 7'h0;
      queueCount_2_27 <= 7'h0;
      queueCount_3_27 <= 7'h0;
      queueCount_4_27 <= 7'h0;
      queueCount_5_27 <= 7'h0;
      queueCount_6_27 <= 7'h0;
      queueCount_7_27 <= 7'h0;
      queueCount_0_28 <= 7'h0;
      queueCount_1_28 <= 7'h0;
      queueCount_2_28 <= 7'h0;
      queueCount_3_28 <= 7'h0;
      queueCount_4_28 <= 7'h0;
      queueCount_5_28 <= 7'h0;
      queueCount_6_28 <= 7'h0;
      queueCount_7_28 <= 7'h0;
      queueCount_0_29 <= 7'h0;
      queueCount_1_29 <= 7'h0;
      queueCount_2_29 <= 7'h0;
      queueCount_3_29 <= 7'h0;
      queueCount_4_29 <= 7'h0;
      queueCount_5_29 <= 7'h0;
      queueCount_6_29 <= 7'h0;
      queueCount_7_29 <= 7'h0;
      queueCount_0_30 <= 7'h0;
      queueCount_1_30 <= 7'h0;
      queueCount_2_30 <= 7'h0;
      queueCount_3_30 <= 7'h0;
      queueCount_4_30 <= 7'h0;
      queueCount_5_30 <= 7'h0;
      queueCount_6_30 <= 7'h0;
      queueCount_7_30 <= 7'h0;
      queueCount_0_31 <= 7'h0;
      queueCount_1_31 <= 7'h0;
      queueCount_2_31 <= 7'h0;
      queueCount_3_31 <= 7'h0;
      queueCount_4_31 <= 7'h0;
      queueCount_5_31 <= 7'h0;
      queueCount_6_31 <= 7'h0;
      queueCount_7_31 <= 7'h0;
    end
    else begin
      if (v0UpdateVec_0_valid)
        v0_0 <= v0_0 & ~maskExt | maskExt & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid)
        v0_1 <= v0_1 & ~maskExt_1 | maskExt_1 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid)
        v0_2 <= v0_2 & ~maskExt_2 | maskExt_2 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid)
        v0_3 <= v0_3 & ~maskExt_3 | maskExt_3 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_4_valid)
        v0_4 <= v0_4 & ~maskExt_4 | maskExt_4 & v0UpdateVec_4_bits_data;
      if (v0UpdateVec_5_valid)
        v0_5 <= v0_5 & ~maskExt_5 | maskExt_5 & v0UpdateVec_5_bits_data;
      if (v0UpdateVec_6_valid)
        v0_6 <= v0_6 & ~maskExt_6 | maskExt_6 & v0UpdateVec_6_bits_data;
      if (v0UpdateVec_7_valid)
        v0_7 <= v0_7 & ~maskExt_7 | maskExt_7 & v0UpdateVec_7_bits_data;
      if (v0UpdateVec_8_valid)
        v0_8 <= v0_8 & ~maskExt_8 | maskExt_8 & v0UpdateVec_8_bits_data;
      if (v0UpdateVec_9_valid)
        v0_9 <= v0_9 & ~maskExt_9 | maskExt_9 & v0UpdateVec_9_bits_data;
      if (v0UpdateVec_10_valid)
        v0_10 <= v0_10 & ~maskExt_10 | maskExt_10 & v0UpdateVec_10_bits_data;
      if (v0UpdateVec_11_valid)
        v0_11 <= v0_11 & ~maskExt_11 | maskExt_11 & v0UpdateVec_11_bits_data;
      if (v0UpdateVec_12_valid)
        v0_12 <= v0_12 & ~maskExt_12 | maskExt_12 & v0UpdateVec_12_bits_data;
      if (v0UpdateVec_13_valid)
        v0_13 <= v0_13 & ~maskExt_13 | maskExt_13 & v0UpdateVec_13_bits_data;
      if (v0UpdateVec_14_valid)
        v0_14 <= v0_14 & ~maskExt_14 | maskExt_14 & v0UpdateVec_14_bits_data;
      if (v0UpdateVec_15_valid)
        v0_15 <= v0_15 & ~maskExt_15 | maskExt_15 & v0UpdateVec_15_bits_data;
      if (v0UpdateVec_16_valid)
        v0_16 <= v0_16 & ~maskExt_16 | maskExt_16 & v0UpdateVec_16_bits_data;
      if (v0UpdateVec_17_valid)
        v0_17 <= v0_17 & ~maskExt_17 | maskExt_17 & v0UpdateVec_17_bits_data;
      if (v0UpdateVec_18_valid)
        v0_18 <= v0_18 & ~maskExt_18 | maskExt_18 & v0UpdateVec_18_bits_data;
      if (v0UpdateVec_19_valid)
        v0_19 <= v0_19 & ~maskExt_19 | maskExt_19 & v0UpdateVec_19_bits_data;
      if (v0UpdateVec_20_valid)
        v0_20 <= v0_20 & ~maskExt_20 | maskExt_20 & v0UpdateVec_20_bits_data;
      if (v0UpdateVec_21_valid)
        v0_21 <= v0_21 & ~maskExt_21 | maskExt_21 & v0UpdateVec_21_bits_data;
      if (v0UpdateVec_22_valid)
        v0_22 <= v0_22 & ~maskExt_22 | maskExt_22 & v0UpdateVec_22_bits_data;
      if (v0UpdateVec_23_valid)
        v0_23 <= v0_23 & ~maskExt_23 | maskExt_23 & v0UpdateVec_23_bits_data;
      if (v0UpdateVec_24_valid)
        v0_24 <= v0_24 & ~maskExt_24 | maskExt_24 & v0UpdateVec_24_bits_data;
      if (v0UpdateVec_25_valid)
        v0_25 <= v0_25 & ~maskExt_25 | maskExt_25 & v0UpdateVec_25_bits_data;
      if (v0UpdateVec_26_valid)
        v0_26 <= v0_26 & ~maskExt_26 | maskExt_26 & v0UpdateVec_26_bits_data;
      if (v0UpdateVec_27_valid)
        v0_27 <= v0_27 & ~maskExt_27 | maskExt_27 & v0UpdateVec_27_bits_data;
      if (v0UpdateVec_28_valid)
        v0_28 <= v0_28 & ~maskExt_28 | maskExt_28 & v0UpdateVec_28_bits_data;
      if (v0UpdateVec_29_valid)
        v0_29 <= v0_29 & ~maskExt_29 | maskExt_29 & v0UpdateVec_29_bits_data;
      if (v0UpdateVec_30_valid)
        v0_30 <= v0_30 & ~maskExt_30 | maskExt_30 & v0UpdateVec_30_bits_data;
      if (v0UpdateVec_31_valid)
        v0_31 <= v0_31 & ~maskExt_31 | maskExt_31 & v0UpdateVec_31_bits_data;
      if (queueEnq[0] ^ queueDeq[0])
        queueCount_0 <= queueCount_0 + counterUpdate;
      if (queueEnq[1] ^ queueDeq[1])
        queueCount_1 <= queueCount_1 + counterUpdate_1;
      if (queueEnq[2] ^ queueDeq[2])
        queueCount_2 <= queueCount_2 + counterUpdate_2;
      if (queueEnq[3] ^ queueDeq[3])
        queueCount_3 <= queueCount_3 + counterUpdate_3;
      if (queueEnq[4] ^ queueDeq[4])
        queueCount_4 <= queueCount_4 + counterUpdate_4;
      if (queueEnq[5] ^ queueDeq[5])
        queueCount_5 <= queueCount_5 + counterUpdate_5;
      if (queueEnq[6] ^ queueDeq[6])
        queueCount_6 <= queueCount_6 + counterUpdate_6;
      if (queueEnq[7] ^ queueDeq[7])
        queueCount_7 <= queueCount_7 + counterUpdate_7;
      if (queueEnq_1[0] ^ queueDeq_1[0])
        queueCount_0_1 <= queueCount_0_1 + counterUpdate_8;
      if (queueEnq_1[1] ^ queueDeq_1[1])
        queueCount_1_1 <= queueCount_1_1 + counterUpdate_9;
      if (queueEnq_1[2] ^ queueDeq_1[2])
        queueCount_2_1 <= queueCount_2_1 + counterUpdate_10;
      if (queueEnq_1[3] ^ queueDeq_1[3])
        queueCount_3_1 <= queueCount_3_1 + counterUpdate_11;
      if (queueEnq_1[4] ^ queueDeq_1[4])
        queueCount_4_1 <= queueCount_4_1 + counterUpdate_12;
      if (queueEnq_1[5] ^ queueDeq_1[5])
        queueCount_5_1 <= queueCount_5_1 + counterUpdate_13;
      if (queueEnq_1[6] ^ queueDeq_1[6])
        queueCount_6_1 <= queueCount_6_1 + counterUpdate_14;
      if (queueEnq_1[7] ^ queueDeq_1[7])
        queueCount_7_1 <= queueCount_7_1 + counterUpdate_15;
      if (queueEnq_2[0] ^ queueDeq_2[0])
        queueCount_0_2 <= queueCount_0_2 + counterUpdate_16;
      if (queueEnq_2[1] ^ queueDeq_2[1])
        queueCount_1_2 <= queueCount_1_2 + counterUpdate_17;
      if (queueEnq_2[2] ^ queueDeq_2[2])
        queueCount_2_2 <= queueCount_2_2 + counterUpdate_18;
      if (queueEnq_2[3] ^ queueDeq_2[3])
        queueCount_3_2 <= queueCount_3_2 + counterUpdate_19;
      if (queueEnq_2[4] ^ queueDeq_2[4])
        queueCount_4_2 <= queueCount_4_2 + counterUpdate_20;
      if (queueEnq_2[5] ^ queueDeq_2[5])
        queueCount_5_2 <= queueCount_5_2 + counterUpdate_21;
      if (queueEnq_2[6] ^ queueDeq_2[6])
        queueCount_6_2 <= queueCount_6_2 + counterUpdate_22;
      if (queueEnq_2[7] ^ queueDeq_2[7])
        queueCount_7_2 <= queueCount_7_2 + counterUpdate_23;
      if (queueEnq_3[0] ^ queueDeq_3[0])
        queueCount_0_3 <= queueCount_0_3 + counterUpdate_24;
      if (queueEnq_3[1] ^ queueDeq_3[1])
        queueCount_1_3 <= queueCount_1_3 + counterUpdate_25;
      if (queueEnq_3[2] ^ queueDeq_3[2])
        queueCount_2_3 <= queueCount_2_3 + counterUpdate_26;
      if (queueEnq_3[3] ^ queueDeq_3[3])
        queueCount_3_3 <= queueCount_3_3 + counterUpdate_27;
      if (queueEnq_3[4] ^ queueDeq_3[4])
        queueCount_4_3 <= queueCount_4_3 + counterUpdate_28;
      if (queueEnq_3[5] ^ queueDeq_3[5])
        queueCount_5_3 <= queueCount_5_3 + counterUpdate_29;
      if (queueEnq_3[6] ^ queueDeq_3[6])
        queueCount_6_3 <= queueCount_6_3 + counterUpdate_30;
      if (queueEnq_3[7] ^ queueDeq_3[7])
        queueCount_7_3 <= queueCount_7_3 + counterUpdate_31;
      if (queueEnq_4[0] ^ queueDeq_4[0])
        queueCount_0_4 <= queueCount_0_4 + counterUpdate_32;
      if (queueEnq_4[1] ^ queueDeq_4[1])
        queueCount_1_4 <= queueCount_1_4 + counterUpdate_33;
      if (queueEnq_4[2] ^ queueDeq_4[2])
        queueCount_2_4 <= queueCount_2_4 + counterUpdate_34;
      if (queueEnq_4[3] ^ queueDeq_4[3])
        queueCount_3_4 <= queueCount_3_4 + counterUpdate_35;
      if (queueEnq_4[4] ^ queueDeq_4[4])
        queueCount_4_4 <= queueCount_4_4 + counterUpdate_36;
      if (queueEnq_4[5] ^ queueDeq_4[5])
        queueCount_5_4 <= queueCount_5_4 + counterUpdate_37;
      if (queueEnq_4[6] ^ queueDeq_4[6])
        queueCount_6_4 <= queueCount_6_4 + counterUpdate_38;
      if (queueEnq_4[7] ^ queueDeq_4[7])
        queueCount_7_4 <= queueCount_7_4 + counterUpdate_39;
      if (queueEnq_5[0] ^ queueDeq_5[0])
        queueCount_0_5 <= queueCount_0_5 + counterUpdate_40;
      if (queueEnq_5[1] ^ queueDeq_5[1])
        queueCount_1_5 <= queueCount_1_5 + counterUpdate_41;
      if (queueEnq_5[2] ^ queueDeq_5[2])
        queueCount_2_5 <= queueCount_2_5 + counterUpdate_42;
      if (queueEnq_5[3] ^ queueDeq_5[3])
        queueCount_3_5 <= queueCount_3_5 + counterUpdate_43;
      if (queueEnq_5[4] ^ queueDeq_5[4])
        queueCount_4_5 <= queueCount_4_5 + counterUpdate_44;
      if (queueEnq_5[5] ^ queueDeq_5[5])
        queueCount_5_5 <= queueCount_5_5 + counterUpdate_45;
      if (queueEnq_5[6] ^ queueDeq_5[6])
        queueCount_6_5 <= queueCount_6_5 + counterUpdate_46;
      if (queueEnq_5[7] ^ queueDeq_5[7])
        queueCount_7_5 <= queueCount_7_5 + counterUpdate_47;
      if (queueEnq_6[0] ^ queueDeq_6[0])
        queueCount_0_6 <= queueCount_0_6 + counterUpdate_48;
      if (queueEnq_6[1] ^ queueDeq_6[1])
        queueCount_1_6 <= queueCount_1_6 + counterUpdate_49;
      if (queueEnq_6[2] ^ queueDeq_6[2])
        queueCount_2_6 <= queueCount_2_6 + counterUpdate_50;
      if (queueEnq_6[3] ^ queueDeq_6[3])
        queueCount_3_6 <= queueCount_3_6 + counterUpdate_51;
      if (queueEnq_6[4] ^ queueDeq_6[4])
        queueCount_4_6 <= queueCount_4_6 + counterUpdate_52;
      if (queueEnq_6[5] ^ queueDeq_6[5])
        queueCount_5_6 <= queueCount_5_6 + counterUpdate_53;
      if (queueEnq_6[6] ^ queueDeq_6[6])
        queueCount_6_6 <= queueCount_6_6 + counterUpdate_54;
      if (queueEnq_6[7] ^ queueDeq_6[7])
        queueCount_7_6 <= queueCount_7_6 + counterUpdate_55;
      if (queueEnq_7[0] ^ queueDeq_7[0])
        queueCount_0_7 <= queueCount_0_7 + counterUpdate_56;
      if (queueEnq_7[1] ^ queueDeq_7[1])
        queueCount_1_7 <= queueCount_1_7 + counterUpdate_57;
      if (queueEnq_7[2] ^ queueDeq_7[2])
        queueCount_2_7 <= queueCount_2_7 + counterUpdate_58;
      if (queueEnq_7[3] ^ queueDeq_7[3])
        queueCount_3_7 <= queueCount_3_7 + counterUpdate_59;
      if (queueEnq_7[4] ^ queueDeq_7[4])
        queueCount_4_7 <= queueCount_4_7 + counterUpdate_60;
      if (queueEnq_7[5] ^ queueDeq_7[5])
        queueCount_5_7 <= queueCount_5_7 + counterUpdate_61;
      if (queueEnq_7[6] ^ queueDeq_7[6])
        queueCount_6_7 <= queueCount_6_7 + counterUpdate_62;
      if (queueEnq_7[7] ^ queueDeq_7[7])
        queueCount_7_7 <= queueCount_7_7 + counterUpdate_63;
      if (queueEnq_8[0] ^ queueDeq_8[0])
        queueCount_0_8 <= queueCount_0_8 + counterUpdate_64;
      if (queueEnq_8[1] ^ queueDeq_8[1])
        queueCount_1_8 <= queueCount_1_8 + counterUpdate_65;
      if (queueEnq_8[2] ^ queueDeq_8[2])
        queueCount_2_8 <= queueCount_2_8 + counterUpdate_66;
      if (queueEnq_8[3] ^ queueDeq_8[3])
        queueCount_3_8 <= queueCount_3_8 + counterUpdate_67;
      if (queueEnq_8[4] ^ queueDeq_8[4])
        queueCount_4_8 <= queueCount_4_8 + counterUpdate_68;
      if (queueEnq_8[5] ^ queueDeq_8[5])
        queueCount_5_8 <= queueCount_5_8 + counterUpdate_69;
      if (queueEnq_8[6] ^ queueDeq_8[6])
        queueCount_6_8 <= queueCount_6_8 + counterUpdate_70;
      if (queueEnq_8[7] ^ queueDeq_8[7])
        queueCount_7_8 <= queueCount_7_8 + counterUpdate_71;
      if (queueEnq_9[0] ^ queueDeq_9[0])
        queueCount_0_9 <= queueCount_0_9 + counterUpdate_72;
      if (queueEnq_9[1] ^ queueDeq_9[1])
        queueCount_1_9 <= queueCount_1_9 + counterUpdate_73;
      if (queueEnq_9[2] ^ queueDeq_9[2])
        queueCount_2_9 <= queueCount_2_9 + counterUpdate_74;
      if (queueEnq_9[3] ^ queueDeq_9[3])
        queueCount_3_9 <= queueCount_3_9 + counterUpdate_75;
      if (queueEnq_9[4] ^ queueDeq_9[4])
        queueCount_4_9 <= queueCount_4_9 + counterUpdate_76;
      if (queueEnq_9[5] ^ queueDeq_9[5])
        queueCount_5_9 <= queueCount_5_9 + counterUpdate_77;
      if (queueEnq_9[6] ^ queueDeq_9[6])
        queueCount_6_9 <= queueCount_6_9 + counterUpdate_78;
      if (queueEnq_9[7] ^ queueDeq_9[7])
        queueCount_7_9 <= queueCount_7_9 + counterUpdate_79;
      if (queueEnq_10[0] ^ queueDeq_10[0])
        queueCount_0_10 <= queueCount_0_10 + counterUpdate_80;
      if (queueEnq_10[1] ^ queueDeq_10[1])
        queueCount_1_10 <= queueCount_1_10 + counterUpdate_81;
      if (queueEnq_10[2] ^ queueDeq_10[2])
        queueCount_2_10 <= queueCount_2_10 + counterUpdate_82;
      if (queueEnq_10[3] ^ queueDeq_10[3])
        queueCount_3_10 <= queueCount_3_10 + counterUpdate_83;
      if (queueEnq_10[4] ^ queueDeq_10[4])
        queueCount_4_10 <= queueCount_4_10 + counterUpdate_84;
      if (queueEnq_10[5] ^ queueDeq_10[5])
        queueCount_5_10 <= queueCount_5_10 + counterUpdate_85;
      if (queueEnq_10[6] ^ queueDeq_10[6])
        queueCount_6_10 <= queueCount_6_10 + counterUpdate_86;
      if (queueEnq_10[7] ^ queueDeq_10[7])
        queueCount_7_10 <= queueCount_7_10 + counterUpdate_87;
      if (queueEnq_11[0] ^ queueDeq_11[0])
        queueCount_0_11 <= queueCount_0_11 + counterUpdate_88;
      if (queueEnq_11[1] ^ queueDeq_11[1])
        queueCount_1_11 <= queueCount_1_11 + counterUpdate_89;
      if (queueEnq_11[2] ^ queueDeq_11[2])
        queueCount_2_11 <= queueCount_2_11 + counterUpdate_90;
      if (queueEnq_11[3] ^ queueDeq_11[3])
        queueCount_3_11 <= queueCount_3_11 + counterUpdate_91;
      if (queueEnq_11[4] ^ queueDeq_11[4])
        queueCount_4_11 <= queueCount_4_11 + counterUpdate_92;
      if (queueEnq_11[5] ^ queueDeq_11[5])
        queueCount_5_11 <= queueCount_5_11 + counterUpdate_93;
      if (queueEnq_11[6] ^ queueDeq_11[6])
        queueCount_6_11 <= queueCount_6_11 + counterUpdate_94;
      if (queueEnq_11[7] ^ queueDeq_11[7])
        queueCount_7_11 <= queueCount_7_11 + counterUpdate_95;
      if (queueEnq_12[0] ^ queueDeq_12[0])
        queueCount_0_12 <= queueCount_0_12 + counterUpdate_96;
      if (queueEnq_12[1] ^ queueDeq_12[1])
        queueCount_1_12 <= queueCount_1_12 + counterUpdate_97;
      if (queueEnq_12[2] ^ queueDeq_12[2])
        queueCount_2_12 <= queueCount_2_12 + counterUpdate_98;
      if (queueEnq_12[3] ^ queueDeq_12[3])
        queueCount_3_12 <= queueCount_3_12 + counterUpdate_99;
      if (queueEnq_12[4] ^ queueDeq_12[4])
        queueCount_4_12 <= queueCount_4_12 + counterUpdate_100;
      if (queueEnq_12[5] ^ queueDeq_12[5])
        queueCount_5_12 <= queueCount_5_12 + counterUpdate_101;
      if (queueEnq_12[6] ^ queueDeq_12[6])
        queueCount_6_12 <= queueCount_6_12 + counterUpdate_102;
      if (queueEnq_12[7] ^ queueDeq_12[7])
        queueCount_7_12 <= queueCount_7_12 + counterUpdate_103;
      if (queueEnq_13[0] ^ queueDeq_13[0])
        queueCount_0_13 <= queueCount_0_13 + counterUpdate_104;
      if (queueEnq_13[1] ^ queueDeq_13[1])
        queueCount_1_13 <= queueCount_1_13 + counterUpdate_105;
      if (queueEnq_13[2] ^ queueDeq_13[2])
        queueCount_2_13 <= queueCount_2_13 + counterUpdate_106;
      if (queueEnq_13[3] ^ queueDeq_13[3])
        queueCount_3_13 <= queueCount_3_13 + counterUpdate_107;
      if (queueEnq_13[4] ^ queueDeq_13[4])
        queueCount_4_13 <= queueCount_4_13 + counterUpdate_108;
      if (queueEnq_13[5] ^ queueDeq_13[5])
        queueCount_5_13 <= queueCount_5_13 + counterUpdate_109;
      if (queueEnq_13[6] ^ queueDeq_13[6])
        queueCount_6_13 <= queueCount_6_13 + counterUpdate_110;
      if (queueEnq_13[7] ^ queueDeq_13[7])
        queueCount_7_13 <= queueCount_7_13 + counterUpdate_111;
      if (queueEnq_14[0] ^ queueDeq_14[0])
        queueCount_0_14 <= queueCount_0_14 + counterUpdate_112;
      if (queueEnq_14[1] ^ queueDeq_14[1])
        queueCount_1_14 <= queueCount_1_14 + counterUpdate_113;
      if (queueEnq_14[2] ^ queueDeq_14[2])
        queueCount_2_14 <= queueCount_2_14 + counterUpdate_114;
      if (queueEnq_14[3] ^ queueDeq_14[3])
        queueCount_3_14 <= queueCount_3_14 + counterUpdate_115;
      if (queueEnq_14[4] ^ queueDeq_14[4])
        queueCount_4_14 <= queueCount_4_14 + counterUpdate_116;
      if (queueEnq_14[5] ^ queueDeq_14[5])
        queueCount_5_14 <= queueCount_5_14 + counterUpdate_117;
      if (queueEnq_14[6] ^ queueDeq_14[6])
        queueCount_6_14 <= queueCount_6_14 + counterUpdate_118;
      if (queueEnq_14[7] ^ queueDeq_14[7])
        queueCount_7_14 <= queueCount_7_14 + counterUpdate_119;
      if (queueEnq_15[0] ^ queueDeq_15[0])
        queueCount_0_15 <= queueCount_0_15 + counterUpdate_120;
      if (queueEnq_15[1] ^ queueDeq_15[1])
        queueCount_1_15 <= queueCount_1_15 + counterUpdate_121;
      if (queueEnq_15[2] ^ queueDeq_15[2])
        queueCount_2_15 <= queueCount_2_15 + counterUpdate_122;
      if (queueEnq_15[3] ^ queueDeq_15[3])
        queueCount_3_15 <= queueCount_3_15 + counterUpdate_123;
      if (queueEnq_15[4] ^ queueDeq_15[4])
        queueCount_4_15 <= queueCount_4_15 + counterUpdate_124;
      if (queueEnq_15[5] ^ queueDeq_15[5])
        queueCount_5_15 <= queueCount_5_15 + counterUpdate_125;
      if (queueEnq_15[6] ^ queueDeq_15[6])
        queueCount_6_15 <= queueCount_6_15 + counterUpdate_126;
      if (queueEnq_15[7] ^ queueDeq_15[7])
        queueCount_7_15 <= queueCount_7_15 + counterUpdate_127;
      if (queueEnq_16[0] ^ queueDeq_16[0])
        queueCount_0_16 <= queueCount_0_16 + counterUpdate_128;
      if (queueEnq_16[1] ^ queueDeq_16[1])
        queueCount_1_16 <= queueCount_1_16 + counterUpdate_129;
      if (queueEnq_16[2] ^ queueDeq_16[2])
        queueCount_2_16 <= queueCount_2_16 + counterUpdate_130;
      if (queueEnq_16[3] ^ queueDeq_16[3])
        queueCount_3_16 <= queueCount_3_16 + counterUpdate_131;
      if (queueEnq_16[4] ^ queueDeq_16[4])
        queueCount_4_16 <= queueCount_4_16 + counterUpdate_132;
      if (queueEnq_16[5] ^ queueDeq_16[5])
        queueCount_5_16 <= queueCount_5_16 + counterUpdate_133;
      if (queueEnq_16[6] ^ queueDeq_16[6])
        queueCount_6_16 <= queueCount_6_16 + counterUpdate_134;
      if (queueEnq_16[7] ^ queueDeq_16[7])
        queueCount_7_16 <= queueCount_7_16 + counterUpdate_135;
      if (queueEnq_17[0] ^ queueDeq_17[0])
        queueCount_0_17 <= queueCount_0_17 + counterUpdate_136;
      if (queueEnq_17[1] ^ queueDeq_17[1])
        queueCount_1_17 <= queueCount_1_17 + counterUpdate_137;
      if (queueEnq_17[2] ^ queueDeq_17[2])
        queueCount_2_17 <= queueCount_2_17 + counterUpdate_138;
      if (queueEnq_17[3] ^ queueDeq_17[3])
        queueCount_3_17 <= queueCount_3_17 + counterUpdate_139;
      if (queueEnq_17[4] ^ queueDeq_17[4])
        queueCount_4_17 <= queueCount_4_17 + counterUpdate_140;
      if (queueEnq_17[5] ^ queueDeq_17[5])
        queueCount_5_17 <= queueCount_5_17 + counterUpdate_141;
      if (queueEnq_17[6] ^ queueDeq_17[6])
        queueCount_6_17 <= queueCount_6_17 + counterUpdate_142;
      if (queueEnq_17[7] ^ queueDeq_17[7])
        queueCount_7_17 <= queueCount_7_17 + counterUpdate_143;
      if (queueEnq_18[0] ^ queueDeq_18[0])
        queueCount_0_18 <= queueCount_0_18 + counterUpdate_144;
      if (queueEnq_18[1] ^ queueDeq_18[1])
        queueCount_1_18 <= queueCount_1_18 + counterUpdate_145;
      if (queueEnq_18[2] ^ queueDeq_18[2])
        queueCount_2_18 <= queueCount_2_18 + counterUpdate_146;
      if (queueEnq_18[3] ^ queueDeq_18[3])
        queueCount_3_18 <= queueCount_3_18 + counterUpdate_147;
      if (queueEnq_18[4] ^ queueDeq_18[4])
        queueCount_4_18 <= queueCount_4_18 + counterUpdate_148;
      if (queueEnq_18[5] ^ queueDeq_18[5])
        queueCount_5_18 <= queueCount_5_18 + counterUpdate_149;
      if (queueEnq_18[6] ^ queueDeq_18[6])
        queueCount_6_18 <= queueCount_6_18 + counterUpdate_150;
      if (queueEnq_18[7] ^ queueDeq_18[7])
        queueCount_7_18 <= queueCount_7_18 + counterUpdate_151;
      if (queueEnq_19[0] ^ queueDeq_19[0])
        queueCount_0_19 <= queueCount_0_19 + counterUpdate_152;
      if (queueEnq_19[1] ^ queueDeq_19[1])
        queueCount_1_19 <= queueCount_1_19 + counterUpdate_153;
      if (queueEnq_19[2] ^ queueDeq_19[2])
        queueCount_2_19 <= queueCount_2_19 + counterUpdate_154;
      if (queueEnq_19[3] ^ queueDeq_19[3])
        queueCount_3_19 <= queueCount_3_19 + counterUpdate_155;
      if (queueEnq_19[4] ^ queueDeq_19[4])
        queueCount_4_19 <= queueCount_4_19 + counterUpdate_156;
      if (queueEnq_19[5] ^ queueDeq_19[5])
        queueCount_5_19 <= queueCount_5_19 + counterUpdate_157;
      if (queueEnq_19[6] ^ queueDeq_19[6])
        queueCount_6_19 <= queueCount_6_19 + counterUpdate_158;
      if (queueEnq_19[7] ^ queueDeq_19[7])
        queueCount_7_19 <= queueCount_7_19 + counterUpdate_159;
      if (queueEnq_20[0] ^ queueDeq_20[0])
        queueCount_0_20 <= queueCount_0_20 + counterUpdate_160;
      if (queueEnq_20[1] ^ queueDeq_20[1])
        queueCount_1_20 <= queueCount_1_20 + counterUpdate_161;
      if (queueEnq_20[2] ^ queueDeq_20[2])
        queueCount_2_20 <= queueCount_2_20 + counterUpdate_162;
      if (queueEnq_20[3] ^ queueDeq_20[3])
        queueCount_3_20 <= queueCount_3_20 + counterUpdate_163;
      if (queueEnq_20[4] ^ queueDeq_20[4])
        queueCount_4_20 <= queueCount_4_20 + counterUpdate_164;
      if (queueEnq_20[5] ^ queueDeq_20[5])
        queueCount_5_20 <= queueCount_5_20 + counterUpdate_165;
      if (queueEnq_20[6] ^ queueDeq_20[6])
        queueCount_6_20 <= queueCount_6_20 + counterUpdate_166;
      if (queueEnq_20[7] ^ queueDeq_20[7])
        queueCount_7_20 <= queueCount_7_20 + counterUpdate_167;
      if (queueEnq_21[0] ^ queueDeq_21[0])
        queueCount_0_21 <= queueCount_0_21 + counterUpdate_168;
      if (queueEnq_21[1] ^ queueDeq_21[1])
        queueCount_1_21 <= queueCount_1_21 + counterUpdate_169;
      if (queueEnq_21[2] ^ queueDeq_21[2])
        queueCount_2_21 <= queueCount_2_21 + counterUpdate_170;
      if (queueEnq_21[3] ^ queueDeq_21[3])
        queueCount_3_21 <= queueCount_3_21 + counterUpdate_171;
      if (queueEnq_21[4] ^ queueDeq_21[4])
        queueCount_4_21 <= queueCount_4_21 + counterUpdate_172;
      if (queueEnq_21[5] ^ queueDeq_21[5])
        queueCount_5_21 <= queueCount_5_21 + counterUpdate_173;
      if (queueEnq_21[6] ^ queueDeq_21[6])
        queueCount_6_21 <= queueCount_6_21 + counterUpdate_174;
      if (queueEnq_21[7] ^ queueDeq_21[7])
        queueCount_7_21 <= queueCount_7_21 + counterUpdate_175;
      if (queueEnq_22[0] ^ queueDeq_22[0])
        queueCount_0_22 <= queueCount_0_22 + counterUpdate_176;
      if (queueEnq_22[1] ^ queueDeq_22[1])
        queueCount_1_22 <= queueCount_1_22 + counterUpdate_177;
      if (queueEnq_22[2] ^ queueDeq_22[2])
        queueCount_2_22 <= queueCount_2_22 + counterUpdate_178;
      if (queueEnq_22[3] ^ queueDeq_22[3])
        queueCount_3_22 <= queueCount_3_22 + counterUpdate_179;
      if (queueEnq_22[4] ^ queueDeq_22[4])
        queueCount_4_22 <= queueCount_4_22 + counterUpdate_180;
      if (queueEnq_22[5] ^ queueDeq_22[5])
        queueCount_5_22 <= queueCount_5_22 + counterUpdate_181;
      if (queueEnq_22[6] ^ queueDeq_22[6])
        queueCount_6_22 <= queueCount_6_22 + counterUpdate_182;
      if (queueEnq_22[7] ^ queueDeq_22[7])
        queueCount_7_22 <= queueCount_7_22 + counterUpdate_183;
      if (queueEnq_23[0] ^ queueDeq_23[0])
        queueCount_0_23 <= queueCount_0_23 + counterUpdate_184;
      if (queueEnq_23[1] ^ queueDeq_23[1])
        queueCount_1_23 <= queueCount_1_23 + counterUpdate_185;
      if (queueEnq_23[2] ^ queueDeq_23[2])
        queueCount_2_23 <= queueCount_2_23 + counterUpdate_186;
      if (queueEnq_23[3] ^ queueDeq_23[3])
        queueCount_3_23 <= queueCount_3_23 + counterUpdate_187;
      if (queueEnq_23[4] ^ queueDeq_23[4])
        queueCount_4_23 <= queueCount_4_23 + counterUpdate_188;
      if (queueEnq_23[5] ^ queueDeq_23[5])
        queueCount_5_23 <= queueCount_5_23 + counterUpdate_189;
      if (queueEnq_23[6] ^ queueDeq_23[6])
        queueCount_6_23 <= queueCount_6_23 + counterUpdate_190;
      if (queueEnq_23[7] ^ queueDeq_23[7])
        queueCount_7_23 <= queueCount_7_23 + counterUpdate_191;
      if (queueEnq_24[0] ^ queueDeq_24[0])
        queueCount_0_24 <= queueCount_0_24 + counterUpdate_192;
      if (queueEnq_24[1] ^ queueDeq_24[1])
        queueCount_1_24 <= queueCount_1_24 + counterUpdate_193;
      if (queueEnq_24[2] ^ queueDeq_24[2])
        queueCount_2_24 <= queueCount_2_24 + counterUpdate_194;
      if (queueEnq_24[3] ^ queueDeq_24[3])
        queueCount_3_24 <= queueCount_3_24 + counterUpdate_195;
      if (queueEnq_24[4] ^ queueDeq_24[4])
        queueCount_4_24 <= queueCount_4_24 + counterUpdate_196;
      if (queueEnq_24[5] ^ queueDeq_24[5])
        queueCount_5_24 <= queueCount_5_24 + counterUpdate_197;
      if (queueEnq_24[6] ^ queueDeq_24[6])
        queueCount_6_24 <= queueCount_6_24 + counterUpdate_198;
      if (queueEnq_24[7] ^ queueDeq_24[7])
        queueCount_7_24 <= queueCount_7_24 + counterUpdate_199;
      if (queueEnq_25[0] ^ queueDeq_25[0])
        queueCount_0_25 <= queueCount_0_25 + counterUpdate_200;
      if (queueEnq_25[1] ^ queueDeq_25[1])
        queueCount_1_25 <= queueCount_1_25 + counterUpdate_201;
      if (queueEnq_25[2] ^ queueDeq_25[2])
        queueCount_2_25 <= queueCount_2_25 + counterUpdate_202;
      if (queueEnq_25[3] ^ queueDeq_25[3])
        queueCount_3_25 <= queueCount_3_25 + counterUpdate_203;
      if (queueEnq_25[4] ^ queueDeq_25[4])
        queueCount_4_25 <= queueCount_4_25 + counterUpdate_204;
      if (queueEnq_25[5] ^ queueDeq_25[5])
        queueCount_5_25 <= queueCount_5_25 + counterUpdate_205;
      if (queueEnq_25[6] ^ queueDeq_25[6])
        queueCount_6_25 <= queueCount_6_25 + counterUpdate_206;
      if (queueEnq_25[7] ^ queueDeq_25[7])
        queueCount_7_25 <= queueCount_7_25 + counterUpdate_207;
      if (queueEnq_26[0] ^ queueDeq_26[0])
        queueCount_0_26 <= queueCount_0_26 + counterUpdate_208;
      if (queueEnq_26[1] ^ queueDeq_26[1])
        queueCount_1_26 <= queueCount_1_26 + counterUpdate_209;
      if (queueEnq_26[2] ^ queueDeq_26[2])
        queueCount_2_26 <= queueCount_2_26 + counterUpdate_210;
      if (queueEnq_26[3] ^ queueDeq_26[3])
        queueCount_3_26 <= queueCount_3_26 + counterUpdate_211;
      if (queueEnq_26[4] ^ queueDeq_26[4])
        queueCount_4_26 <= queueCount_4_26 + counterUpdate_212;
      if (queueEnq_26[5] ^ queueDeq_26[5])
        queueCount_5_26 <= queueCount_5_26 + counterUpdate_213;
      if (queueEnq_26[6] ^ queueDeq_26[6])
        queueCount_6_26 <= queueCount_6_26 + counterUpdate_214;
      if (queueEnq_26[7] ^ queueDeq_26[7])
        queueCount_7_26 <= queueCount_7_26 + counterUpdate_215;
      if (queueEnq_27[0] ^ queueDeq_27[0])
        queueCount_0_27 <= queueCount_0_27 + counterUpdate_216;
      if (queueEnq_27[1] ^ queueDeq_27[1])
        queueCount_1_27 <= queueCount_1_27 + counterUpdate_217;
      if (queueEnq_27[2] ^ queueDeq_27[2])
        queueCount_2_27 <= queueCount_2_27 + counterUpdate_218;
      if (queueEnq_27[3] ^ queueDeq_27[3])
        queueCount_3_27 <= queueCount_3_27 + counterUpdate_219;
      if (queueEnq_27[4] ^ queueDeq_27[4])
        queueCount_4_27 <= queueCount_4_27 + counterUpdate_220;
      if (queueEnq_27[5] ^ queueDeq_27[5])
        queueCount_5_27 <= queueCount_5_27 + counterUpdate_221;
      if (queueEnq_27[6] ^ queueDeq_27[6])
        queueCount_6_27 <= queueCount_6_27 + counterUpdate_222;
      if (queueEnq_27[7] ^ queueDeq_27[7])
        queueCount_7_27 <= queueCount_7_27 + counterUpdate_223;
      if (queueEnq_28[0] ^ queueDeq_28[0])
        queueCount_0_28 <= queueCount_0_28 + counterUpdate_224;
      if (queueEnq_28[1] ^ queueDeq_28[1])
        queueCount_1_28 <= queueCount_1_28 + counterUpdate_225;
      if (queueEnq_28[2] ^ queueDeq_28[2])
        queueCount_2_28 <= queueCount_2_28 + counterUpdate_226;
      if (queueEnq_28[3] ^ queueDeq_28[3])
        queueCount_3_28 <= queueCount_3_28 + counterUpdate_227;
      if (queueEnq_28[4] ^ queueDeq_28[4])
        queueCount_4_28 <= queueCount_4_28 + counterUpdate_228;
      if (queueEnq_28[5] ^ queueDeq_28[5])
        queueCount_5_28 <= queueCount_5_28 + counterUpdate_229;
      if (queueEnq_28[6] ^ queueDeq_28[6])
        queueCount_6_28 <= queueCount_6_28 + counterUpdate_230;
      if (queueEnq_28[7] ^ queueDeq_28[7])
        queueCount_7_28 <= queueCount_7_28 + counterUpdate_231;
      if (queueEnq_29[0] ^ queueDeq_29[0])
        queueCount_0_29 <= queueCount_0_29 + counterUpdate_232;
      if (queueEnq_29[1] ^ queueDeq_29[1])
        queueCount_1_29 <= queueCount_1_29 + counterUpdate_233;
      if (queueEnq_29[2] ^ queueDeq_29[2])
        queueCount_2_29 <= queueCount_2_29 + counterUpdate_234;
      if (queueEnq_29[3] ^ queueDeq_29[3])
        queueCount_3_29 <= queueCount_3_29 + counterUpdate_235;
      if (queueEnq_29[4] ^ queueDeq_29[4])
        queueCount_4_29 <= queueCount_4_29 + counterUpdate_236;
      if (queueEnq_29[5] ^ queueDeq_29[5])
        queueCount_5_29 <= queueCount_5_29 + counterUpdate_237;
      if (queueEnq_29[6] ^ queueDeq_29[6])
        queueCount_6_29 <= queueCount_6_29 + counterUpdate_238;
      if (queueEnq_29[7] ^ queueDeq_29[7])
        queueCount_7_29 <= queueCount_7_29 + counterUpdate_239;
      if (queueEnq_30[0] ^ queueDeq_30[0])
        queueCount_0_30 <= queueCount_0_30 + counterUpdate_240;
      if (queueEnq_30[1] ^ queueDeq_30[1])
        queueCount_1_30 <= queueCount_1_30 + counterUpdate_241;
      if (queueEnq_30[2] ^ queueDeq_30[2])
        queueCount_2_30 <= queueCount_2_30 + counterUpdate_242;
      if (queueEnq_30[3] ^ queueDeq_30[3])
        queueCount_3_30 <= queueCount_3_30 + counterUpdate_243;
      if (queueEnq_30[4] ^ queueDeq_30[4])
        queueCount_4_30 <= queueCount_4_30 + counterUpdate_244;
      if (queueEnq_30[5] ^ queueDeq_30[5])
        queueCount_5_30 <= queueCount_5_30 + counterUpdate_245;
      if (queueEnq_30[6] ^ queueDeq_30[6])
        queueCount_6_30 <= queueCount_6_30 + counterUpdate_246;
      if (queueEnq_30[7] ^ queueDeq_30[7])
        queueCount_7_30 <= queueCount_7_30 + counterUpdate_247;
      if (queueEnq_31[0] ^ queueDeq_31[0])
        queueCount_0_31 <= queueCount_0_31 + counterUpdate_248;
      if (queueEnq_31[1] ^ queueDeq_31[1])
        queueCount_1_31 <= queueCount_1_31 + counterUpdate_249;
      if (queueEnq_31[2] ^ queueDeq_31[2])
        queueCount_2_31 <= queueCount_2_31 + counterUpdate_250;
      if (queueEnq_31[3] ^ queueDeq_31[3])
        queueCount_3_31 <= queueCount_3_31 + counterUpdate_251;
      if (queueEnq_31[4] ^ queueDeq_31[4])
        queueCount_4_31 <= queueCount_4_31 + counterUpdate_252;
      if (queueEnq_31[5] ^ queueDeq_31[5])
        queueCount_5_31 <= queueCount_5_31 + counterUpdate_253;
      if (queueEnq_31[6] ^ queueDeq_31[6])
        queueCount_6_31 <= queueCount_6_31 + counterUpdate_254;
      if (queueEnq_31[7] ^ queueDeq_31[7])
        queueCount_7_31 <= queueCount_7_31 + counterUpdate_255;
    end
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:87];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [6:0] i = 7'h0; i < 7'h58; i += 7'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        v0_0 = _RANDOM[7'h0];
        v0_1 = _RANDOM[7'h1];
        v0_2 = _RANDOM[7'h2];
        v0_3 = _RANDOM[7'h3];
        v0_4 = _RANDOM[7'h4];
        v0_5 = _RANDOM[7'h5];
        v0_6 = _RANDOM[7'h6];
        v0_7 = _RANDOM[7'h7];
        v0_8 = _RANDOM[7'h8];
        v0_9 = _RANDOM[7'h9];
        v0_10 = _RANDOM[7'hA];
        v0_11 = _RANDOM[7'hB];
        v0_12 = _RANDOM[7'hC];
        v0_13 = _RANDOM[7'hD];
        v0_14 = _RANDOM[7'hE];
        v0_15 = _RANDOM[7'hF];
        v0_16 = _RANDOM[7'h10];
        v0_17 = _RANDOM[7'h11];
        v0_18 = _RANDOM[7'h12];
        v0_19 = _RANDOM[7'h13];
        v0_20 = _RANDOM[7'h14];
        v0_21 = _RANDOM[7'h15];
        v0_22 = _RANDOM[7'h16];
        v0_23 = _RANDOM[7'h17];
        v0_24 = _RANDOM[7'h18];
        v0_25 = _RANDOM[7'h19];
        v0_26 = _RANDOM[7'h1A];
        v0_27 = _RANDOM[7'h1B];
        v0_28 = _RANDOM[7'h1C];
        v0_29 = _RANDOM[7'h1D];
        v0_30 = _RANDOM[7'h1E];
        v0_31 = _RANDOM[7'h1F];
        queueCount_0 = _RANDOM[7'h20][6:0];
        queueCount_1 = _RANDOM[7'h20][13:7];
        queueCount_2 = _RANDOM[7'h20][20:14];
        queueCount_3 = _RANDOM[7'h20][27:21];
        queueCount_4 = {_RANDOM[7'h20][31:28], _RANDOM[7'h21][2:0]};
        queueCount_5 = _RANDOM[7'h21][9:3];
        queueCount_6 = _RANDOM[7'h21][16:10];
        queueCount_7 = _RANDOM[7'h21][23:17];
        queueCount_0_1 = _RANDOM[7'h21][30:24];
        queueCount_1_1 = {_RANDOM[7'h21][31], _RANDOM[7'h22][5:0]};
        queueCount_2_1 = _RANDOM[7'h22][12:6];
        queueCount_3_1 = _RANDOM[7'h22][19:13];
        queueCount_4_1 = _RANDOM[7'h22][26:20];
        queueCount_5_1 = {_RANDOM[7'h22][31:27], _RANDOM[7'h23][1:0]};
        queueCount_6_1 = _RANDOM[7'h23][8:2];
        queueCount_7_1 = _RANDOM[7'h23][15:9];
        queueCount_0_2 = _RANDOM[7'h23][22:16];
        queueCount_1_2 = _RANDOM[7'h23][29:23];
        queueCount_2_2 = {_RANDOM[7'h23][31:30], _RANDOM[7'h24][4:0]};
        queueCount_3_2 = _RANDOM[7'h24][11:5];
        queueCount_4_2 = _RANDOM[7'h24][18:12];
        queueCount_5_2 = _RANDOM[7'h24][25:19];
        queueCount_6_2 = {_RANDOM[7'h24][31:26], _RANDOM[7'h25][0]};
        queueCount_7_2 = _RANDOM[7'h25][7:1];
        queueCount_0_3 = _RANDOM[7'h25][14:8];
        queueCount_1_3 = _RANDOM[7'h25][21:15];
        queueCount_2_3 = _RANDOM[7'h25][28:22];
        queueCount_3_3 = {_RANDOM[7'h25][31:29], _RANDOM[7'h26][3:0]};
        queueCount_4_3 = _RANDOM[7'h26][10:4];
        queueCount_5_3 = _RANDOM[7'h26][17:11];
        queueCount_6_3 = _RANDOM[7'h26][24:18];
        queueCount_7_3 = _RANDOM[7'h26][31:25];
        queueCount_0_4 = _RANDOM[7'h27][6:0];
        queueCount_1_4 = _RANDOM[7'h27][13:7];
        queueCount_2_4 = _RANDOM[7'h27][20:14];
        queueCount_3_4 = _RANDOM[7'h27][27:21];
        queueCount_4_4 = {_RANDOM[7'h27][31:28], _RANDOM[7'h28][2:0]};
        queueCount_5_4 = _RANDOM[7'h28][9:3];
        queueCount_6_4 = _RANDOM[7'h28][16:10];
        queueCount_7_4 = _RANDOM[7'h28][23:17];
        queueCount_0_5 = _RANDOM[7'h28][30:24];
        queueCount_1_5 = {_RANDOM[7'h28][31], _RANDOM[7'h29][5:0]};
        queueCount_2_5 = _RANDOM[7'h29][12:6];
        queueCount_3_5 = _RANDOM[7'h29][19:13];
        queueCount_4_5 = _RANDOM[7'h29][26:20];
        queueCount_5_5 = {_RANDOM[7'h29][31:27], _RANDOM[7'h2A][1:0]};
        queueCount_6_5 = _RANDOM[7'h2A][8:2];
        queueCount_7_5 = _RANDOM[7'h2A][15:9];
        queueCount_0_6 = _RANDOM[7'h2A][22:16];
        queueCount_1_6 = _RANDOM[7'h2A][29:23];
        queueCount_2_6 = {_RANDOM[7'h2A][31:30], _RANDOM[7'h2B][4:0]};
        queueCount_3_6 = _RANDOM[7'h2B][11:5];
        queueCount_4_6 = _RANDOM[7'h2B][18:12];
        queueCount_5_6 = _RANDOM[7'h2B][25:19];
        queueCount_6_6 = {_RANDOM[7'h2B][31:26], _RANDOM[7'h2C][0]};
        queueCount_7_6 = _RANDOM[7'h2C][7:1];
        queueCount_0_7 = _RANDOM[7'h2C][14:8];
        queueCount_1_7 = _RANDOM[7'h2C][21:15];
        queueCount_2_7 = _RANDOM[7'h2C][28:22];
        queueCount_3_7 = {_RANDOM[7'h2C][31:29], _RANDOM[7'h2D][3:0]};
        queueCount_4_7 = _RANDOM[7'h2D][10:4];
        queueCount_5_7 = _RANDOM[7'h2D][17:11];
        queueCount_6_7 = _RANDOM[7'h2D][24:18];
        queueCount_7_7 = _RANDOM[7'h2D][31:25];
        queueCount_0_8 = _RANDOM[7'h2E][6:0];
        queueCount_1_8 = _RANDOM[7'h2E][13:7];
        queueCount_2_8 = _RANDOM[7'h2E][20:14];
        queueCount_3_8 = _RANDOM[7'h2E][27:21];
        queueCount_4_8 = {_RANDOM[7'h2E][31:28], _RANDOM[7'h2F][2:0]};
        queueCount_5_8 = _RANDOM[7'h2F][9:3];
        queueCount_6_8 = _RANDOM[7'h2F][16:10];
        queueCount_7_8 = _RANDOM[7'h2F][23:17];
        queueCount_0_9 = _RANDOM[7'h2F][30:24];
        queueCount_1_9 = {_RANDOM[7'h2F][31], _RANDOM[7'h30][5:0]};
        queueCount_2_9 = _RANDOM[7'h30][12:6];
        queueCount_3_9 = _RANDOM[7'h30][19:13];
        queueCount_4_9 = _RANDOM[7'h30][26:20];
        queueCount_5_9 = {_RANDOM[7'h30][31:27], _RANDOM[7'h31][1:0]};
        queueCount_6_9 = _RANDOM[7'h31][8:2];
        queueCount_7_9 = _RANDOM[7'h31][15:9];
        queueCount_0_10 = _RANDOM[7'h31][22:16];
        queueCount_1_10 = _RANDOM[7'h31][29:23];
        queueCount_2_10 = {_RANDOM[7'h31][31:30], _RANDOM[7'h32][4:0]};
        queueCount_3_10 = _RANDOM[7'h32][11:5];
        queueCount_4_10 = _RANDOM[7'h32][18:12];
        queueCount_5_10 = _RANDOM[7'h32][25:19];
        queueCount_6_10 = {_RANDOM[7'h32][31:26], _RANDOM[7'h33][0]};
        queueCount_7_10 = _RANDOM[7'h33][7:1];
        queueCount_0_11 = _RANDOM[7'h33][14:8];
        queueCount_1_11 = _RANDOM[7'h33][21:15];
        queueCount_2_11 = _RANDOM[7'h33][28:22];
        queueCount_3_11 = {_RANDOM[7'h33][31:29], _RANDOM[7'h34][3:0]};
        queueCount_4_11 = _RANDOM[7'h34][10:4];
        queueCount_5_11 = _RANDOM[7'h34][17:11];
        queueCount_6_11 = _RANDOM[7'h34][24:18];
        queueCount_7_11 = _RANDOM[7'h34][31:25];
        queueCount_0_12 = _RANDOM[7'h35][6:0];
        queueCount_1_12 = _RANDOM[7'h35][13:7];
        queueCount_2_12 = _RANDOM[7'h35][20:14];
        queueCount_3_12 = _RANDOM[7'h35][27:21];
        queueCount_4_12 = {_RANDOM[7'h35][31:28], _RANDOM[7'h36][2:0]};
        queueCount_5_12 = _RANDOM[7'h36][9:3];
        queueCount_6_12 = _RANDOM[7'h36][16:10];
        queueCount_7_12 = _RANDOM[7'h36][23:17];
        queueCount_0_13 = _RANDOM[7'h36][30:24];
        queueCount_1_13 = {_RANDOM[7'h36][31], _RANDOM[7'h37][5:0]};
        queueCount_2_13 = _RANDOM[7'h37][12:6];
        queueCount_3_13 = _RANDOM[7'h37][19:13];
        queueCount_4_13 = _RANDOM[7'h37][26:20];
        queueCount_5_13 = {_RANDOM[7'h37][31:27], _RANDOM[7'h38][1:0]};
        queueCount_6_13 = _RANDOM[7'h38][8:2];
        queueCount_7_13 = _RANDOM[7'h38][15:9];
        queueCount_0_14 = _RANDOM[7'h38][22:16];
        queueCount_1_14 = _RANDOM[7'h38][29:23];
        queueCount_2_14 = {_RANDOM[7'h38][31:30], _RANDOM[7'h39][4:0]};
        queueCount_3_14 = _RANDOM[7'h39][11:5];
        queueCount_4_14 = _RANDOM[7'h39][18:12];
        queueCount_5_14 = _RANDOM[7'h39][25:19];
        queueCount_6_14 = {_RANDOM[7'h39][31:26], _RANDOM[7'h3A][0]};
        queueCount_7_14 = _RANDOM[7'h3A][7:1];
        queueCount_0_15 = _RANDOM[7'h3A][14:8];
        queueCount_1_15 = _RANDOM[7'h3A][21:15];
        queueCount_2_15 = _RANDOM[7'h3A][28:22];
        queueCount_3_15 = {_RANDOM[7'h3A][31:29], _RANDOM[7'h3B][3:0]};
        queueCount_4_15 = _RANDOM[7'h3B][10:4];
        queueCount_5_15 = _RANDOM[7'h3B][17:11];
        queueCount_6_15 = _RANDOM[7'h3B][24:18];
        queueCount_7_15 = _RANDOM[7'h3B][31:25];
        queueCount_0_16 = _RANDOM[7'h3C][6:0];
        queueCount_1_16 = _RANDOM[7'h3C][13:7];
        queueCount_2_16 = _RANDOM[7'h3C][20:14];
        queueCount_3_16 = _RANDOM[7'h3C][27:21];
        queueCount_4_16 = {_RANDOM[7'h3C][31:28], _RANDOM[7'h3D][2:0]};
        queueCount_5_16 = _RANDOM[7'h3D][9:3];
        queueCount_6_16 = _RANDOM[7'h3D][16:10];
        queueCount_7_16 = _RANDOM[7'h3D][23:17];
        queueCount_0_17 = _RANDOM[7'h3D][30:24];
        queueCount_1_17 = {_RANDOM[7'h3D][31], _RANDOM[7'h3E][5:0]};
        queueCount_2_17 = _RANDOM[7'h3E][12:6];
        queueCount_3_17 = _RANDOM[7'h3E][19:13];
        queueCount_4_17 = _RANDOM[7'h3E][26:20];
        queueCount_5_17 = {_RANDOM[7'h3E][31:27], _RANDOM[7'h3F][1:0]};
        queueCount_6_17 = _RANDOM[7'h3F][8:2];
        queueCount_7_17 = _RANDOM[7'h3F][15:9];
        queueCount_0_18 = _RANDOM[7'h3F][22:16];
        queueCount_1_18 = _RANDOM[7'h3F][29:23];
        queueCount_2_18 = {_RANDOM[7'h3F][31:30], _RANDOM[7'h40][4:0]};
        queueCount_3_18 = _RANDOM[7'h40][11:5];
        queueCount_4_18 = _RANDOM[7'h40][18:12];
        queueCount_5_18 = _RANDOM[7'h40][25:19];
        queueCount_6_18 = {_RANDOM[7'h40][31:26], _RANDOM[7'h41][0]};
        queueCount_7_18 = _RANDOM[7'h41][7:1];
        queueCount_0_19 = _RANDOM[7'h41][14:8];
        queueCount_1_19 = _RANDOM[7'h41][21:15];
        queueCount_2_19 = _RANDOM[7'h41][28:22];
        queueCount_3_19 = {_RANDOM[7'h41][31:29], _RANDOM[7'h42][3:0]};
        queueCount_4_19 = _RANDOM[7'h42][10:4];
        queueCount_5_19 = _RANDOM[7'h42][17:11];
        queueCount_6_19 = _RANDOM[7'h42][24:18];
        queueCount_7_19 = _RANDOM[7'h42][31:25];
        queueCount_0_20 = _RANDOM[7'h43][6:0];
        queueCount_1_20 = _RANDOM[7'h43][13:7];
        queueCount_2_20 = _RANDOM[7'h43][20:14];
        queueCount_3_20 = _RANDOM[7'h43][27:21];
        queueCount_4_20 = {_RANDOM[7'h43][31:28], _RANDOM[7'h44][2:0]};
        queueCount_5_20 = _RANDOM[7'h44][9:3];
        queueCount_6_20 = _RANDOM[7'h44][16:10];
        queueCount_7_20 = _RANDOM[7'h44][23:17];
        queueCount_0_21 = _RANDOM[7'h44][30:24];
        queueCount_1_21 = {_RANDOM[7'h44][31], _RANDOM[7'h45][5:0]};
        queueCount_2_21 = _RANDOM[7'h45][12:6];
        queueCount_3_21 = _RANDOM[7'h45][19:13];
        queueCount_4_21 = _RANDOM[7'h45][26:20];
        queueCount_5_21 = {_RANDOM[7'h45][31:27], _RANDOM[7'h46][1:0]};
        queueCount_6_21 = _RANDOM[7'h46][8:2];
        queueCount_7_21 = _RANDOM[7'h46][15:9];
        queueCount_0_22 = _RANDOM[7'h46][22:16];
        queueCount_1_22 = _RANDOM[7'h46][29:23];
        queueCount_2_22 = {_RANDOM[7'h46][31:30], _RANDOM[7'h47][4:0]};
        queueCount_3_22 = _RANDOM[7'h47][11:5];
        queueCount_4_22 = _RANDOM[7'h47][18:12];
        queueCount_5_22 = _RANDOM[7'h47][25:19];
        queueCount_6_22 = {_RANDOM[7'h47][31:26], _RANDOM[7'h48][0]};
        queueCount_7_22 = _RANDOM[7'h48][7:1];
        queueCount_0_23 = _RANDOM[7'h48][14:8];
        queueCount_1_23 = _RANDOM[7'h48][21:15];
        queueCount_2_23 = _RANDOM[7'h48][28:22];
        queueCount_3_23 = {_RANDOM[7'h48][31:29], _RANDOM[7'h49][3:0]};
        queueCount_4_23 = _RANDOM[7'h49][10:4];
        queueCount_5_23 = _RANDOM[7'h49][17:11];
        queueCount_6_23 = _RANDOM[7'h49][24:18];
        queueCount_7_23 = _RANDOM[7'h49][31:25];
        queueCount_0_24 = _RANDOM[7'h4A][6:0];
        queueCount_1_24 = _RANDOM[7'h4A][13:7];
        queueCount_2_24 = _RANDOM[7'h4A][20:14];
        queueCount_3_24 = _RANDOM[7'h4A][27:21];
        queueCount_4_24 = {_RANDOM[7'h4A][31:28], _RANDOM[7'h4B][2:0]};
        queueCount_5_24 = _RANDOM[7'h4B][9:3];
        queueCount_6_24 = _RANDOM[7'h4B][16:10];
        queueCount_7_24 = _RANDOM[7'h4B][23:17];
        queueCount_0_25 = _RANDOM[7'h4B][30:24];
        queueCount_1_25 = {_RANDOM[7'h4B][31], _RANDOM[7'h4C][5:0]};
        queueCount_2_25 = _RANDOM[7'h4C][12:6];
        queueCount_3_25 = _RANDOM[7'h4C][19:13];
        queueCount_4_25 = _RANDOM[7'h4C][26:20];
        queueCount_5_25 = {_RANDOM[7'h4C][31:27], _RANDOM[7'h4D][1:0]};
        queueCount_6_25 = _RANDOM[7'h4D][8:2];
        queueCount_7_25 = _RANDOM[7'h4D][15:9];
        queueCount_0_26 = _RANDOM[7'h4D][22:16];
        queueCount_1_26 = _RANDOM[7'h4D][29:23];
        queueCount_2_26 = {_RANDOM[7'h4D][31:30], _RANDOM[7'h4E][4:0]};
        queueCount_3_26 = _RANDOM[7'h4E][11:5];
        queueCount_4_26 = _RANDOM[7'h4E][18:12];
        queueCount_5_26 = _RANDOM[7'h4E][25:19];
        queueCount_6_26 = {_RANDOM[7'h4E][31:26], _RANDOM[7'h4F][0]};
        queueCount_7_26 = _RANDOM[7'h4F][7:1];
        queueCount_0_27 = _RANDOM[7'h4F][14:8];
        queueCount_1_27 = _RANDOM[7'h4F][21:15];
        queueCount_2_27 = _RANDOM[7'h4F][28:22];
        queueCount_3_27 = {_RANDOM[7'h4F][31:29], _RANDOM[7'h50][3:0]};
        queueCount_4_27 = _RANDOM[7'h50][10:4];
        queueCount_5_27 = _RANDOM[7'h50][17:11];
        queueCount_6_27 = _RANDOM[7'h50][24:18];
        queueCount_7_27 = _RANDOM[7'h50][31:25];
        queueCount_0_28 = _RANDOM[7'h51][6:0];
        queueCount_1_28 = _RANDOM[7'h51][13:7];
        queueCount_2_28 = _RANDOM[7'h51][20:14];
        queueCount_3_28 = _RANDOM[7'h51][27:21];
        queueCount_4_28 = {_RANDOM[7'h51][31:28], _RANDOM[7'h52][2:0]};
        queueCount_5_28 = _RANDOM[7'h52][9:3];
        queueCount_6_28 = _RANDOM[7'h52][16:10];
        queueCount_7_28 = _RANDOM[7'h52][23:17];
        queueCount_0_29 = _RANDOM[7'h52][30:24];
        queueCount_1_29 = {_RANDOM[7'h52][31], _RANDOM[7'h53][5:0]};
        queueCount_2_29 = _RANDOM[7'h53][12:6];
        queueCount_3_29 = _RANDOM[7'h53][19:13];
        queueCount_4_29 = _RANDOM[7'h53][26:20];
        queueCount_5_29 = {_RANDOM[7'h53][31:27], _RANDOM[7'h54][1:0]};
        queueCount_6_29 = _RANDOM[7'h54][8:2];
        queueCount_7_29 = _RANDOM[7'h54][15:9];
        queueCount_0_30 = _RANDOM[7'h54][22:16];
        queueCount_1_30 = _RANDOM[7'h54][29:23];
        queueCount_2_30 = {_RANDOM[7'h54][31:30], _RANDOM[7'h55][4:0]};
        queueCount_3_30 = _RANDOM[7'h55][11:5];
        queueCount_4_30 = _RANDOM[7'h55][18:12];
        queueCount_5_30 = _RANDOM[7'h55][25:19];
        queueCount_6_30 = {_RANDOM[7'h55][31:26], _RANDOM[7'h56][0]};
        queueCount_7_30 = _RANDOM[7'h56][7:1];
        queueCount_0_31 = _RANDOM[7'h56][14:8];
        queueCount_1_31 = _RANDOM[7'h56][21:15];
        queueCount_2_31 = _RANDOM[7'h56][28:22];
        queueCount_3_31 = {_RANDOM[7'h56][31:29], _RANDOM[7'h57][3:0]};
        queueCount_4_31 = _RANDOM[7'h57][10:4];
        queueCount_5_31 = _RANDOM[7'h57][17:11];
        queueCount_6_31 = _RANDOM[7'h57][24:18];
        queueCount_7_31 = _RANDOM[7'h57][31:25];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  wire [3:0]        sourceQueue_deq_bits;
  wire [31:0]       axi4Port_aw_bits_addr_0;
  assign axi4Port_aw_bits_addr_0 = _storeUnit_memRequest_bits_address;
  assign dataQueue_enq_bits_index = _storeUnit_memRequest_bits_index;
  assign dataQueue_enq_bits_address = _storeUnit_memRequest_bits_address;
  wire [9:0]        simpleSourceQueue_deq_bits;
  wire [31:0]       simpleAccessPorts_aw_bits_addr_0;
  assign simpleAccessPorts_aw_bits_addr_0 = _otherUnit_memWriteRequest_bits_address;
  wire [31:0]       otherUnitTargetQueue_enq_bits;
  assign otherUnitTargetQueue_enq_bits = _otherUnit_status_targetLane;
  assign simpleDataQueue_enq_bits_source = _otherUnit_memWriteRequest_bits_source;
  assign simpleDataQueue_enq_bits_address = _otherUnit_memWriteRequest_bits_address;
  assign simpleDataQueue_enq_bits_size = _otherUnit_memWriteRequest_bits_size;
  wire              writeQueueVec_0_empty;
  assign writeQueueVec_0_empty = _writeQueueVec_fifo_empty;
  wire              writeQueueVec_0_full;
  assign writeQueueVec_0_full = _writeQueueVec_fifo_full;
  wire              writeQueueVec_1_empty;
  assign writeQueueVec_1_empty = _writeQueueVec_fifo_1_empty;
  wire              writeQueueVec_1_full;
  assign writeQueueVec_1_full = _writeQueueVec_fifo_1_full;
  wire              writeQueueVec_2_empty;
  assign writeQueueVec_2_empty = _writeQueueVec_fifo_2_empty;
  wire              writeQueueVec_2_full;
  assign writeQueueVec_2_full = _writeQueueVec_fifo_2_full;
  wire              writeQueueVec_3_empty;
  assign writeQueueVec_3_empty = _writeQueueVec_fifo_3_empty;
  wire              writeQueueVec_3_full;
  assign writeQueueVec_3_full = _writeQueueVec_fifo_3_full;
  wire              writeQueueVec_4_empty;
  assign writeQueueVec_4_empty = _writeQueueVec_fifo_4_empty;
  wire              writeQueueVec_4_full;
  assign writeQueueVec_4_full = _writeQueueVec_fifo_4_full;
  wire              writeQueueVec_5_empty;
  assign writeQueueVec_5_empty = _writeQueueVec_fifo_5_empty;
  wire              writeQueueVec_5_full;
  assign writeQueueVec_5_full = _writeQueueVec_fifo_5_full;
  wire              writeQueueVec_6_empty;
  assign writeQueueVec_6_empty = _writeQueueVec_fifo_6_empty;
  wire              writeQueueVec_6_full;
  assign writeQueueVec_6_full = _writeQueueVec_fifo_6_full;
  wire              writeQueueVec_7_empty;
  assign writeQueueVec_7_empty = _writeQueueVec_fifo_7_empty;
  wire              writeQueueVec_7_full;
  assign writeQueueVec_7_full = _writeQueueVec_fifo_7_full;
  wire              writeQueueVec_8_empty;
  assign writeQueueVec_8_empty = _writeQueueVec_fifo_8_empty;
  wire              writeQueueVec_8_full;
  assign writeQueueVec_8_full = _writeQueueVec_fifo_8_full;
  wire              writeQueueVec_9_empty;
  assign writeQueueVec_9_empty = _writeQueueVec_fifo_9_empty;
  wire              writeQueueVec_9_full;
  assign writeQueueVec_9_full = _writeQueueVec_fifo_9_full;
  wire              writeQueueVec_10_empty;
  assign writeQueueVec_10_empty = _writeQueueVec_fifo_10_empty;
  wire              writeQueueVec_10_full;
  assign writeQueueVec_10_full = _writeQueueVec_fifo_10_full;
  wire              writeQueueVec_11_empty;
  assign writeQueueVec_11_empty = _writeQueueVec_fifo_11_empty;
  wire              writeQueueVec_11_full;
  assign writeQueueVec_11_full = _writeQueueVec_fifo_11_full;
  wire              writeQueueVec_12_empty;
  assign writeQueueVec_12_empty = _writeQueueVec_fifo_12_empty;
  wire              writeQueueVec_12_full;
  assign writeQueueVec_12_full = _writeQueueVec_fifo_12_full;
  wire              writeQueueVec_13_empty;
  assign writeQueueVec_13_empty = _writeQueueVec_fifo_13_empty;
  wire              writeQueueVec_13_full;
  assign writeQueueVec_13_full = _writeQueueVec_fifo_13_full;
  wire              writeQueueVec_14_empty;
  assign writeQueueVec_14_empty = _writeQueueVec_fifo_14_empty;
  wire              writeQueueVec_14_full;
  assign writeQueueVec_14_full = _writeQueueVec_fifo_14_full;
  wire              writeQueueVec_15_empty;
  assign writeQueueVec_15_empty = _writeQueueVec_fifo_15_empty;
  wire              writeQueueVec_15_full;
  assign writeQueueVec_15_full = _writeQueueVec_fifo_15_full;
  wire              writeQueueVec_16_empty;
  assign writeQueueVec_16_empty = _writeQueueVec_fifo_16_empty;
  wire              writeQueueVec_16_full;
  assign writeQueueVec_16_full = _writeQueueVec_fifo_16_full;
  wire              writeQueueVec_17_empty;
  assign writeQueueVec_17_empty = _writeQueueVec_fifo_17_empty;
  wire              writeQueueVec_17_full;
  assign writeQueueVec_17_full = _writeQueueVec_fifo_17_full;
  wire              writeQueueVec_18_empty;
  assign writeQueueVec_18_empty = _writeQueueVec_fifo_18_empty;
  wire              writeQueueVec_18_full;
  assign writeQueueVec_18_full = _writeQueueVec_fifo_18_full;
  wire              writeQueueVec_19_empty;
  assign writeQueueVec_19_empty = _writeQueueVec_fifo_19_empty;
  wire              writeQueueVec_19_full;
  assign writeQueueVec_19_full = _writeQueueVec_fifo_19_full;
  wire              writeQueueVec_20_empty;
  assign writeQueueVec_20_empty = _writeQueueVec_fifo_20_empty;
  wire              writeQueueVec_20_full;
  assign writeQueueVec_20_full = _writeQueueVec_fifo_20_full;
  wire              writeQueueVec_21_empty;
  assign writeQueueVec_21_empty = _writeQueueVec_fifo_21_empty;
  wire              writeQueueVec_21_full;
  assign writeQueueVec_21_full = _writeQueueVec_fifo_21_full;
  wire              writeQueueVec_22_empty;
  assign writeQueueVec_22_empty = _writeQueueVec_fifo_22_empty;
  wire              writeQueueVec_22_full;
  assign writeQueueVec_22_full = _writeQueueVec_fifo_22_full;
  wire              writeQueueVec_23_empty;
  assign writeQueueVec_23_empty = _writeQueueVec_fifo_23_empty;
  wire              writeQueueVec_23_full;
  assign writeQueueVec_23_full = _writeQueueVec_fifo_23_full;
  wire              writeQueueVec_24_empty;
  assign writeQueueVec_24_empty = _writeQueueVec_fifo_24_empty;
  wire              writeQueueVec_24_full;
  assign writeQueueVec_24_full = _writeQueueVec_fifo_24_full;
  wire              writeQueueVec_25_empty;
  assign writeQueueVec_25_empty = _writeQueueVec_fifo_25_empty;
  wire              writeQueueVec_25_full;
  assign writeQueueVec_25_full = _writeQueueVec_fifo_25_full;
  wire              writeQueueVec_26_empty;
  assign writeQueueVec_26_empty = _writeQueueVec_fifo_26_empty;
  wire              writeQueueVec_26_full;
  assign writeQueueVec_26_full = _writeQueueVec_fifo_26_full;
  wire              writeQueueVec_27_empty;
  assign writeQueueVec_27_empty = _writeQueueVec_fifo_27_empty;
  wire              writeQueueVec_27_full;
  assign writeQueueVec_27_full = _writeQueueVec_fifo_27_full;
  wire              writeQueueVec_28_empty;
  assign writeQueueVec_28_empty = _writeQueueVec_fifo_28_empty;
  wire              writeQueueVec_28_full;
  assign writeQueueVec_28_full = _writeQueueVec_fifo_28_full;
  wire              writeQueueVec_29_empty;
  assign writeQueueVec_29_empty = _writeQueueVec_fifo_29_empty;
  wire              writeQueueVec_29_full;
  assign writeQueueVec_29_full = _writeQueueVec_fifo_29_full;
  wire              writeQueueVec_30_empty;
  assign writeQueueVec_30_empty = _writeQueueVec_fifo_30_empty;
  wire              writeQueueVec_30_full;
  assign writeQueueVec_30_full = _writeQueueVec_fifo_30_full;
  wire              writeQueueVec_31_empty;
  assign writeQueueVec_31_empty = _writeQueueVec_fifo_31_empty;
  wire              writeQueueVec_31_full;
  assign writeQueueVec_31_full = _writeQueueVec_fifo_31_full;
  assign otherUnitTargetQueue_empty = _otherUnitTargetQueue_fifo_empty;
  wire              otherUnitTargetQueue_full;
  assign otherUnitTargetQueue_full = _otherUnitTargetQueue_fifo_full;
  wire              otherUnitDataQueueVec_0_empty;
  assign otherUnitDataQueueVec_0_empty = _otherUnitDataQueueVec_fifo_empty;
  wire              otherUnitDataQueueVec_0_full;
  assign otherUnitDataQueueVec_0_full = _otherUnitDataQueueVec_fifo_full;
  wire              otherUnitDataQueueVec_1_empty;
  assign otherUnitDataQueueVec_1_empty = _otherUnitDataQueueVec_fifo_1_empty;
  wire              otherUnitDataQueueVec_1_full;
  assign otherUnitDataQueueVec_1_full = _otherUnitDataQueueVec_fifo_1_full;
  wire              otherUnitDataQueueVec_2_empty;
  assign otherUnitDataQueueVec_2_empty = _otherUnitDataQueueVec_fifo_2_empty;
  wire              otherUnitDataQueueVec_2_full;
  assign otherUnitDataQueueVec_2_full = _otherUnitDataQueueVec_fifo_2_full;
  wire              otherUnitDataQueueVec_3_empty;
  assign otherUnitDataQueueVec_3_empty = _otherUnitDataQueueVec_fifo_3_empty;
  wire              otherUnitDataQueueVec_3_full;
  assign otherUnitDataQueueVec_3_full = _otherUnitDataQueueVec_fifo_3_full;
  wire              otherUnitDataQueueVec_4_empty;
  assign otherUnitDataQueueVec_4_empty = _otherUnitDataQueueVec_fifo_4_empty;
  wire              otherUnitDataQueueVec_4_full;
  assign otherUnitDataQueueVec_4_full = _otherUnitDataQueueVec_fifo_4_full;
  wire              otherUnitDataQueueVec_5_empty;
  assign otherUnitDataQueueVec_5_empty = _otherUnitDataQueueVec_fifo_5_empty;
  wire              otherUnitDataQueueVec_5_full;
  assign otherUnitDataQueueVec_5_full = _otherUnitDataQueueVec_fifo_5_full;
  wire              otherUnitDataQueueVec_6_empty;
  assign otherUnitDataQueueVec_6_empty = _otherUnitDataQueueVec_fifo_6_empty;
  wire              otherUnitDataQueueVec_6_full;
  assign otherUnitDataQueueVec_6_full = _otherUnitDataQueueVec_fifo_6_full;
  wire              otherUnitDataQueueVec_7_empty;
  assign otherUnitDataQueueVec_7_empty = _otherUnitDataQueueVec_fifo_7_empty;
  wire              otherUnitDataQueueVec_7_full;
  assign otherUnitDataQueueVec_7_full = _otherUnitDataQueueVec_fifo_7_full;
  wire              otherUnitDataQueueVec_8_empty;
  assign otherUnitDataQueueVec_8_empty = _otherUnitDataQueueVec_fifo_8_empty;
  wire              otherUnitDataQueueVec_8_full;
  assign otherUnitDataQueueVec_8_full = _otherUnitDataQueueVec_fifo_8_full;
  wire              otherUnitDataQueueVec_9_empty;
  assign otherUnitDataQueueVec_9_empty = _otherUnitDataQueueVec_fifo_9_empty;
  wire              otherUnitDataQueueVec_9_full;
  assign otherUnitDataQueueVec_9_full = _otherUnitDataQueueVec_fifo_9_full;
  wire              otherUnitDataQueueVec_10_empty;
  assign otherUnitDataQueueVec_10_empty = _otherUnitDataQueueVec_fifo_10_empty;
  wire              otherUnitDataQueueVec_10_full;
  assign otherUnitDataQueueVec_10_full = _otherUnitDataQueueVec_fifo_10_full;
  wire              otherUnitDataQueueVec_11_empty;
  assign otherUnitDataQueueVec_11_empty = _otherUnitDataQueueVec_fifo_11_empty;
  wire              otherUnitDataQueueVec_11_full;
  assign otherUnitDataQueueVec_11_full = _otherUnitDataQueueVec_fifo_11_full;
  wire              otherUnitDataQueueVec_12_empty;
  assign otherUnitDataQueueVec_12_empty = _otherUnitDataQueueVec_fifo_12_empty;
  wire              otherUnitDataQueueVec_12_full;
  assign otherUnitDataQueueVec_12_full = _otherUnitDataQueueVec_fifo_12_full;
  wire              otherUnitDataQueueVec_13_empty;
  assign otherUnitDataQueueVec_13_empty = _otherUnitDataQueueVec_fifo_13_empty;
  wire              otherUnitDataQueueVec_13_full;
  assign otherUnitDataQueueVec_13_full = _otherUnitDataQueueVec_fifo_13_full;
  wire              otherUnitDataQueueVec_14_empty;
  assign otherUnitDataQueueVec_14_empty = _otherUnitDataQueueVec_fifo_14_empty;
  wire              otherUnitDataQueueVec_14_full;
  assign otherUnitDataQueueVec_14_full = _otherUnitDataQueueVec_fifo_14_full;
  wire              otherUnitDataQueueVec_15_empty;
  assign otherUnitDataQueueVec_15_empty = _otherUnitDataQueueVec_fifo_15_empty;
  wire              otherUnitDataQueueVec_15_full;
  assign otherUnitDataQueueVec_15_full = _otherUnitDataQueueVec_fifo_15_full;
  wire              otherUnitDataQueueVec_16_empty;
  assign otherUnitDataQueueVec_16_empty = _otherUnitDataQueueVec_fifo_16_empty;
  wire              otherUnitDataQueueVec_16_full;
  assign otherUnitDataQueueVec_16_full = _otherUnitDataQueueVec_fifo_16_full;
  wire              otherUnitDataQueueVec_17_empty;
  assign otherUnitDataQueueVec_17_empty = _otherUnitDataQueueVec_fifo_17_empty;
  wire              otherUnitDataQueueVec_17_full;
  assign otherUnitDataQueueVec_17_full = _otherUnitDataQueueVec_fifo_17_full;
  wire              otherUnitDataQueueVec_18_empty;
  assign otherUnitDataQueueVec_18_empty = _otherUnitDataQueueVec_fifo_18_empty;
  wire              otherUnitDataQueueVec_18_full;
  assign otherUnitDataQueueVec_18_full = _otherUnitDataQueueVec_fifo_18_full;
  wire              otherUnitDataQueueVec_19_empty;
  assign otherUnitDataQueueVec_19_empty = _otherUnitDataQueueVec_fifo_19_empty;
  wire              otherUnitDataQueueVec_19_full;
  assign otherUnitDataQueueVec_19_full = _otherUnitDataQueueVec_fifo_19_full;
  wire              otherUnitDataQueueVec_20_empty;
  assign otherUnitDataQueueVec_20_empty = _otherUnitDataQueueVec_fifo_20_empty;
  wire              otherUnitDataQueueVec_20_full;
  assign otherUnitDataQueueVec_20_full = _otherUnitDataQueueVec_fifo_20_full;
  wire              otherUnitDataQueueVec_21_empty;
  assign otherUnitDataQueueVec_21_empty = _otherUnitDataQueueVec_fifo_21_empty;
  wire              otherUnitDataQueueVec_21_full;
  assign otherUnitDataQueueVec_21_full = _otherUnitDataQueueVec_fifo_21_full;
  wire              otherUnitDataQueueVec_22_empty;
  assign otherUnitDataQueueVec_22_empty = _otherUnitDataQueueVec_fifo_22_empty;
  wire              otherUnitDataQueueVec_22_full;
  assign otherUnitDataQueueVec_22_full = _otherUnitDataQueueVec_fifo_22_full;
  wire              otherUnitDataQueueVec_23_empty;
  assign otherUnitDataQueueVec_23_empty = _otherUnitDataQueueVec_fifo_23_empty;
  wire              otherUnitDataQueueVec_23_full;
  assign otherUnitDataQueueVec_23_full = _otherUnitDataQueueVec_fifo_23_full;
  wire              otherUnitDataQueueVec_24_empty;
  assign otherUnitDataQueueVec_24_empty = _otherUnitDataQueueVec_fifo_24_empty;
  wire              otherUnitDataQueueVec_24_full;
  assign otherUnitDataQueueVec_24_full = _otherUnitDataQueueVec_fifo_24_full;
  wire              otherUnitDataQueueVec_25_empty;
  assign otherUnitDataQueueVec_25_empty = _otherUnitDataQueueVec_fifo_25_empty;
  wire              otherUnitDataQueueVec_25_full;
  assign otherUnitDataQueueVec_25_full = _otherUnitDataQueueVec_fifo_25_full;
  wire              otherUnitDataQueueVec_26_empty;
  assign otherUnitDataQueueVec_26_empty = _otherUnitDataQueueVec_fifo_26_empty;
  wire              otherUnitDataQueueVec_26_full;
  assign otherUnitDataQueueVec_26_full = _otherUnitDataQueueVec_fifo_26_full;
  wire              otherUnitDataQueueVec_27_empty;
  assign otherUnitDataQueueVec_27_empty = _otherUnitDataQueueVec_fifo_27_empty;
  wire              otherUnitDataQueueVec_27_full;
  assign otherUnitDataQueueVec_27_full = _otherUnitDataQueueVec_fifo_27_full;
  wire              otherUnitDataQueueVec_28_empty;
  assign otherUnitDataQueueVec_28_empty = _otherUnitDataQueueVec_fifo_28_empty;
  wire              otherUnitDataQueueVec_28_full;
  assign otherUnitDataQueueVec_28_full = _otherUnitDataQueueVec_fifo_28_full;
  wire              otherUnitDataQueueVec_29_empty;
  assign otherUnitDataQueueVec_29_empty = _otherUnitDataQueueVec_fifo_29_empty;
  wire              otherUnitDataQueueVec_29_full;
  assign otherUnitDataQueueVec_29_full = _otherUnitDataQueueVec_fifo_29_full;
  wire              otherUnitDataQueueVec_30_empty;
  assign otherUnitDataQueueVec_30_empty = _otherUnitDataQueueVec_fifo_30_empty;
  wire              otherUnitDataQueueVec_30_full;
  assign otherUnitDataQueueVec_30_full = _otherUnitDataQueueVec_fifo_30_full;
  wire              otherUnitDataQueueVec_31_empty;
  assign otherUnitDataQueueVec_31_empty = _otherUnitDataQueueVec_fifo_31_empty;
  wire              otherUnitDataQueueVec_31_full;
  assign otherUnitDataQueueVec_31_full = _otherUnitDataQueueVec_fifo_31_full;
  wire              writeIndexQueue_empty;
  assign writeIndexQueue_empty = _writeIndexQueue_fifo_empty;
  wire              writeIndexQueue_full;
  assign writeIndexQueue_full = _writeIndexQueue_fifo_full;
  wire              writeIndexQueue_1_empty;
  assign writeIndexQueue_1_empty = _writeIndexQueue_fifo_1_empty;
  wire              writeIndexQueue_1_full;
  assign writeIndexQueue_1_full = _writeIndexQueue_fifo_1_full;
  wire              writeIndexQueue_2_empty;
  assign writeIndexQueue_2_empty = _writeIndexQueue_fifo_2_empty;
  wire              writeIndexQueue_2_full;
  assign writeIndexQueue_2_full = _writeIndexQueue_fifo_2_full;
  wire              writeIndexQueue_3_empty;
  assign writeIndexQueue_3_empty = _writeIndexQueue_fifo_3_empty;
  wire              writeIndexQueue_3_full;
  assign writeIndexQueue_3_full = _writeIndexQueue_fifo_3_full;
  wire              writeIndexQueue_4_empty;
  assign writeIndexQueue_4_empty = _writeIndexQueue_fifo_4_empty;
  wire              writeIndexQueue_4_full;
  assign writeIndexQueue_4_full = _writeIndexQueue_fifo_4_full;
  wire              writeIndexQueue_5_empty;
  assign writeIndexQueue_5_empty = _writeIndexQueue_fifo_5_empty;
  wire              writeIndexQueue_5_full;
  assign writeIndexQueue_5_full = _writeIndexQueue_fifo_5_full;
  wire              writeIndexQueue_6_empty;
  assign writeIndexQueue_6_empty = _writeIndexQueue_fifo_6_empty;
  wire              writeIndexQueue_6_full;
  assign writeIndexQueue_6_full = _writeIndexQueue_fifo_6_full;
  wire              writeIndexQueue_7_empty;
  assign writeIndexQueue_7_empty = _writeIndexQueue_fifo_7_empty;
  wire              writeIndexQueue_7_full;
  assign writeIndexQueue_7_full = _writeIndexQueue_fifo_7_full;
  wire              writeIndexQueue_8_empty;
  assign writeIndexQueue_8_empty = _writeIndexQueue_fifo_8_empty;
  wire              writeIndexQueue_8_full;
  assign writeIndexQueue_8_full = _writeIndexQueue_fifo_8_full;
  wire              writeIndexQueue_9_empty;
  assign writeIndexQueue_9_empty = _writeIndexQueue_fifo_9_empty;
  wire              writeIndexQueue_9_full;
  assign writeIndexQueue_9_full = _writeIndexQueue_fifo_9_full;
  wire              writeIndexQueue_10_empty;
  assign writeIndexQueue_10_empty = _writeIndexQueue_fifo_10_empty;
  wire              writeIndexQueue_10_full;
  assign writeIndexQueue_10_full = _writeIndexQueue_fifo_10_full;
  wire              writeIndexQueue_11_empty;
  assign writeIndexQueue_11_empty = _writeIndexQueue_fifo_11_empty;
  wire              writeIndexQueue_11_full;
  assign writeIndexQueue_11_full = _writeIndexQueue_fifo_11_full;
  wire              writeIndexQueue_12_empty;
  assign writeIndexQueue_12_empty = _writeIndexQueue_fifo_12_empty;
  wire              writeIndexQueue_12_full;
  assign writeIndexQueue_12_full = _writeIndexQueue_fifo_12_full;
  wire              writeIndexQueue_13_empty;
  assign writeIndexQueue_13_empty = _writeIndexQueue_fifo_13_empty;
  wire              writeIndexQueue_13_full;
  assign writeIndexQueue_13_full = _writeIndexQueue_fifo_13_full;
  wire              writeIndexQueue_14_empty;
  assign writeIndexQueue_14_empty = _writeIndexQueue_fifo_14_empty;
  wire              writeIndexQueue_14_full;
  assign writeIndexQueue_14_full = _writeIndexQueue_fifo_14_full;
  wire              writeIndexQueue_15_empty;
  assign writeIndexQueue_15_empty = _writeIndexQueue_fifo_15_empty;
  wire              writeIndexQueue_15_full;
  assign writeIndexQueue_15_full = _writeIndexQueue_fifo_15_full;
  wire              writeIndexQueue_16_empty;
  assign writeIndexQueue_16_empty = _writeIndexQueue_fifo_16_empty;
  wire              writeIndexQueue_16_full;
  assign writeIndexQueue_16_full = _writeIndexQueue_fifo_16_full;
  wire              writeIndexQueue_17_empty;
  assign writeIndexQueue_17_empty = _writeIndexQueue_fifo_17_empty;
  wire              writeIndexQueue_17_full;
  assign writeIndexQueue_17_full = _writeIndexQueue_fifo_17_full;
  wire              writeIndexQueue_18_empty;
  assign writeIndexQueue_18_empty = _writeIndexQueue_fifo_18_empty;
  wire              writeIndexQueue_18_full;
  assign writeIndexQueue_18_full = _writeIndexQueue_fifo_18_full;
  wire              writeIndexQueue_19_empty;
  assign writeIndexQueue_19_empty = _writeIndexQueue_fifo_19_empty;
  wire              writeIndexQueue_19_full;
  assign writeIndexQueue_19_full = _writeIndexQueue_fifo_19_full;
  wire              writeIndexQueue_20_empty;
  assign writeIndexQueue_20_empty = _writeIndexQueue_fifo_20_empty;
  wire              writeIndexQueue_20_full;
  assign writeIndexQueue_20_full = _writeIndexQueue_fifo_20_full;
  wire              writeIndexQueue_21_empty;
  assign writeIndexQueue_21_empty = _writeIndexQueue_fifo_21_empty;
  wire              writeIndexQueue_21_full;
  assign writeIndexQueue_21_full = _writeIndexQueue_fifo_21_full;
  wire              writeIndexQueue_22_empty;
  assign writeIndexQueue_22_empty = _writeIndexQueue_fifo_22_empty;
  wire              writeIndexQueue_22_full;
  assign writeIndexQueue_22_full = _writeIndexQueue_fifo_22_full;
  wire              writeIndexQueue_23_empty;
  assign writeIndexQueue_23_empty = _writeIndexQueue_fifo_23_empty;
  wire              writeIndexQueue_23_full;
  assign writeIndexQueue_23_full = _writeIndexQueue_fifo_23_full;
  wire              writeIndexQueue_24_empty;
  assign writeIndexQueue_24_empty = _writeIndexQueue_fifo_24_empty;
  wire              writeIndexQueue_24_full;
  assign writeIndexQueue_24_full = _writeIndexQueue_fifo_24_full;
  wire              writeIndexQueue_25_empty;
  assign writeIndexQueue_25_empty = _writeIndexQueue_fifo_25_empty;
  wire              writeIndexQueue_25_full;
  assign writeIndexQueue_25_full = _writeIndexQueue_fifo_25_full;
  wire              writeIndexQueue_26_empty;
  assign writeIndexQueue_26_empty = _writeIndexQueue_fifo_26_empty;
  wire              writeIndexQueue_26_full;
  assign writeIndexQueue_26_full = _writeIndexQueue_fifo_26_full;
  wire              writeIndexQueue_27_empty;
  assign writeIndexQueue_27_empty = _writeIndexQueue_fifo_27_empty;
  wire              writeIndexQueue_27_full;
  assign writeIndexQueue_27_full = _writeIndexQueue_fifo_27_full;
  wire              writeIndexQueue_28_empty;
  assign writeIndexQueue_28_empty = _writeIndexQueue_fifo_28_empty;
  wire              writeIndexQueue_28_full;
  assign writeIndexQueue_28_full = _writeIndexQueue_fifo_28_full;
  wire              writeIndexQueue_29_empty;
  assign writeIndexQueue_29_empty = _writeIndexQueue_fifo_29_empty;
  wire              writeIndexQueue_29_full;
  assign writeIndexQueue_29_full = _writeIndexQueue_fifo_29_full;
  wire              writeIndexQueue_30_empty;
  assign writeIndexQueue_30_empty = _writeIndexQueue_fifo_30_empty;
  wire              writeIndexQueue_30_full;
  assign writeIndexQueue_30_full = _writeIndexQueue_fifo_30_full;
  wire              writeIndexQueue_31_empty;
  assign writeIndexQueue_31_empty = _writeIndexQueue_fifo_31_empty;
  wire              writeIndexQueue_31_full;
  assign writeIndexQueue_31_full = _writeIndexQueue_fifo_31_full;
  wire              sourceQueue_empty;
  assign sourceQueue_empty = _sourceQueue_fifo_empty;
  wire              sourceQueue_full;
  assign sourceQueue_full = _sourceQueue_fifo_full;
  wire              dataQueue_empty;
  assign dataQueue_empty = _dataQueue_fifo_empty;
  wire              dataQueue_full;
  assign dataQueue_full = _dataQueue_fifo_full;
  wire              simpleSourceQueue_empty;
  assign simpleSourceQueue_empty = _simpleSourceQueue_fifo_empty;
  wire              simpleSourceQueue_full;
  assign simpleSourceQueue_full = _simpleSourceQueue_fifo_full;
  wire              simpleDataQueue_empty;
  assign simpleDataQueue_empty = _simpleDataQueue_fifo_empty;
  wire              simpleDataQueue_full;
  assign simpleDataQueue_full = _simpleDataQueue_fifo_full;
  LoadUnit loadUnit (
    .clock                                                  (clock),
    .reset                                                  (reset),
    .lsuRequest_valid                                       (reqEnq_0),
    .lsuRequest_bits_instructionInformation_nf              (request_bits_instructionInformation_nf_0),
    .lsuRequest_bits_instructionInformation_mew             (request_bits_instructionInformation_mew_0),
    .lsuRequest_bits_instructionInformation_mop             (request_bits_instructionInformation_mop_0),
    .lsuRequest_bits_instructionInformation_lumop           (request_bits_instructionInformation_lumop_0),
    .lsuRequest_bits_instructionInformation_eew             (request_bits_instructionInformation_eew_0),
    .lsuRequest_bits_instructionInformation_vs3             (request_bits_instructionInformation_vs3_0),
    .lsuRequest_bits_instructionInformation_isStore         (request_bits_instructionInformation_isStore_0),
    .lsuRequest_bits_instructionInformation_maskedLoadStore (request_bits_instructionInformation_maskedLoadStore_0),
    .lsuRequest_bits_rs1Data                                (request_bits_rs1Data_0),
    .lsuRequest_bits_rs2Data                                (request_bits_rs2Data_0),
    .lsuRequest_bits_instructionIndex                       (request_bits_instructionIndex_0),
    .csrInterface_vl                                        (csrInterface_vl),
    .csrInterface_vStart                                    (csrInterface_vStart),
    .csrInterface_vlmul                                     (csrInterface_vlmul),
    .csrInterface_vSew                                      (csrInterface_vSew),
    .csrInterface_vxrm                                      (csrInterface_vxrm),
    .csrInterface_vta                                       (csrInterface_vta),
    .csrInterface_vma                                       (csrInterface_vma),
    .maskInput                                              (_GEN_15[maskSelect]),
    .maskSelect_valid                                       (_loadUnit_maskSelect_valid),
    .maskSelect_bits                                        (_loadUnit_maskSelect_bits),
    .addressConflict                                        (stallLoad),
    .memRequest_ready                                       (sourceQueue_enq_ready & axi4Port_ar_ready_0),
    .memRequest_valid                                       (_loadUnit_memRequest_valid),
    .memRequest_bits_src                                    (sourceQueue_enq_bits),
    .memRequest_bits_address                                (axi4Port_ar_bits_addr_0),
    .memResponse_ready                                      (axi4Port_r_ready_0),
    .memResponse_valid                                      (axi4Port_r_valid_0),
    .memResponse_bits_data                                  (axi4Port_r_bits_data_0),
    .memResponse_bits_index                                 (sourceQueue_deq_bits),
    .status_idle                                            (_loadUnit_status_idle),
    .status_last                                            (_loadUnit_status_last),
    .status_instructionIndex                                (_loadUnit_status_instructionIndex),
    .status_changeMaskGroup                                 (/* unused */),
    .status_startAddress                                    (_loadUnit_status_startAddress),
    .status_endAddress                                      (_loadUnit_status_endAddress),
    .vrfWritePort_0_ready                                   (writeQueueVec_0_enq_ready & ~(otherTryToWrite[0])),
    .vrfWritePort_0_valid                                   (_loadUnit_vrfWritePort_0_valid),
    .vrfWritePort_0_bits_vd                                 (_loadUnit_vrfWritePort_0_bits_vd),
    .vrfWritePort_0_bits_mask                               (_loadUnit_vrfWritePort_0_bits_mask),
    .vrfWritePort_0_bits_data                               (_loadUnit_vrfWritePort_0_bits_data),
    .vrfWritePort_0_bits_instructionIndex                   (_loadUnit_vrfWritePort_0_bits_instructionIndex),
    .vrfWritePort_1_ready                                   (writeQueueVec_1_enq_ready & ~(otherTryToWrite[1])),
    .vrfWritePort_1_valid                                   (_loadUnit_vrfWritePort_1_valid),
    .vrfWritePort_1_bits_vd                                 (_loadUnit_vrfWritePort_1_bits_vd),
    .vrfWritePort_1_bits_mask                               (_loadUnit_vrfWritePort_1_bits_mask),
    .vrfWritePort_1_bits_data                               (_loadUnit_vrfWritePort_1_bits_data),
    .vrfWritePort_1_bits_instructionIndex                   (_loadUnit_vrfWritePort_1_bits_instructionIndex),
    .vrfWritePort_2_ready                                   (writeQueueVec_2_enq_ready & ~(otherTryToWrite[2])),
    .vrfWritePort_2_valid                                   (_loadUnit_vrfWritePort_2_valid),
    .vrfWritePort_2_bits_vd                                 (_loadUnit_vrfWritePort_2_bits_vd),
    .vrfWritePort_2_bits_mask                               (_loadUnit_vrfWritePort_2_bits_mask),
    .vrfWritePort_2_bits_data                               (_loadUnit_vrfWritePort_2_bits_data),
    .vrfWritePort_2_bits_instructionIndex                   (_loadUnit_vrfWritePort_2_bits_instructionIndex),
    .vrfWritePort_3_ready                                   (writeQueueVec_3_enq_ready & ~(otherTryToWrite[3])),
    .vrfWritePort_3_valid                                   (_loadUnit_vrfWritePort_3_valid),
    .vrfWritePort_3_bits_vd                                 (_loadUnit_vrfWritePort_3_bits_vd),
    .vrfWritePort_3_bits_mask                               (_loadUnit_vrfWritePort_3_bits_mask),
    .vrfWritePort_3_bits_data                               (_loadUnit_vrfWritePort_3_bits_data),
    .vrfWritePort_3_bits_instructionIndex                   (_loadUnit_vrfWritePort_3_bits_instructionIndex),
    .vrfWritePort_4_ready                                   (writeQueueVec_4_enq_ready & ~(otherTryToWrite[4])),
    .vrfWritePort_4_valid                                   (_loadUnit_vrfWritePort_4_valid),
    .vrfWritePort_4_bits_vd                                 (_loadUnit_vrfWritePort_4_bits_vd),
    .vrfWritePort_4_bits_mask                               (_loadUnit_vrfWritePort_4_bits_mask),
    .vrfWritePort_4_bits_data                               (_loadUnit_vrfWritePort_4_bits_data),
    .vrfWritePort_4_bits_instructionIndex                   (_loadUnit_vrfWritePort_4_bits_instructionIndex),
    .vrfWritePort_5_ready                                   (writeQueueVec_5_enq_ready & ~(otherTryToWrite[5])),
    .vrfWritePort_5_valid                                   (_loadUnit_vrfWritePort_5_valid),
    .vrfWritePort_5_bits_vd                                 (_loadUnit_vrfWritePort_5_bits_vd),
    .vrfWritePort_5_bits_mask                               (_loadUnit_vrfWritePort_5_bits_mask),
    .vrfWritePort_5_bits_data                               (_loadUnit_vrfWritePort_5_bits_data),
    .vrfWritePort_5_bits_instructionIndex                   (_loadUnit_vrfWritePort_5_bits_instructionIndex),
    .vrfWritePort_6_ready                                   (writeQueueVec_6_enq_ready & ~(otherTryToWrite[6])),
    .vrfWritePort_6_valid                                   (_loadUnit_vrfWritePort_6_valid),
    .vrfWritePort_6_bits_vd                                 (_loadUnit_vrfWritePort_6_bits_vd),
    .vrfWritePort_6_bits_mask                               (_loadUnit_vrfWritePort_6_bits_mask),
    .vrfWritePort_6_bits_data                               (_loadUnit_vrfWritePort_6_bits_data),
    .vrfWritePort_6_bits_instructionIndex                   (_loadUnit_vrfWritePort_6_bits_instructionIndex),
    .vrfWritePort_7_ready                                   (writeQueueVec_7_enq_ready & ~(otherTryToWrite[7])),
    .vrfWritePort_7_valid                                   (_loadUnit_vrfWritePort_7_valid),
    .vrfWritePort_7_bits_vd                                 (_loadUnit_vrfWritePort_7_bits_vd),
    .vrfWritePort_7_bits_mask                               (_loadUnit_vrfWritePort_7_bits_mask),
    .vrfWritePort_7_bits_data                               (_loadUnit_vrfWritePort_7_bits_data),
    .vrfWritePort_7_bits_instructionIndex                   (_loadUnit_vrfWritePort_7_bits_instructionIndex),
    .vrfWritePort_8_ready                                   (writeQueueVec_8_enq_ready & ~(otherTryToWrite[8])),
    .vrfWritePort_8_valid                                   (_loadUnit_vrfWritePort_8_valid),
    .vrfWritePort_8_bits_vd                                 (_loadUnit_vrfWritePort_8_bits_vd),
    .vrfWritePort_8_bits_mask                               (_loadUnit_vrfWritePort_8_bits_mask),
    .vrfWritePort_8_bits_data                               (_loadUnit_vrfWritePort_8_bits_data),
    .vrfWritePort_8_bits_instructionIndex                   (_loadUnit_vrfWritePort_8_bits_instructionIndex),
    .vrfWritePort_9_ready                                   (writeQueueVec_9_enq_ready & ~(otherTryToWrite[9])),
    .vrfWritePort_9_valid                                   (_loadUnit_vrfWritePort_9_valid),
    .vrfWritePort_9_bits_vd                                 (_loadUnit_vrfWritePort_9_bits_vd),
    .vrfWritePort_9_bits_mask                               (_loadUnit_vrfWritePort_9_bits_mask),
    .vrfWritePort_9_bits_data                               (_loadUnit_vrfWritePort_9_bits_data),
    .vrfWritePort_9_bits_instructionIndex                   (_loadUnit_vrfWritePort_9_bits_instructionIndex),
    .vrfWritePort_10_ready                                  (writeQueueVec_10_enq_ready & ~(otherTryToWrite[10])),
    .vrfWritePort_10_valid                                  (_loadUnit_vrfWritePort_10_valid),
    .vrfWritePort_10_bits_vd                                (_loadUnit_vrfWritePort_10_bits_vd),
    .vrfWritePort_10_bits_mask                              (_loadUnit_vrfWritePort_10_bits_mask),
    .vrfWritePort_10_bits_data                              (_loadUnit_vrfWritePort_10_bits_data),
    .vrfWritePort_10_bits_instructionIndex                  (_loadUnit_vrfWritePort_10_bits_instructionIndex),
    .vrfWritePort_11_ready                                  (writeQueueVec_11_enq_ready & ~(otherTryToWrite[11])),
    .vrfWritePort_11_valid                                  (_loadUnit_vrfWritePort_11_valid),
    .vrfWritePort_11_bits_vd                                (_loadUnit_vrfWritePort_11_bits_vd),
    .vrfWritePort_11_bits_mask                              (_loadUnit_vrfWritePort_11_bits_mask),
    .vrfWritePort_11_bits_data                              (_loadUnit_vrfWritePort_11_bits_data),
    .vrfWritePort_11_bits_instructionIndex                  (_loadUnit_vrfWritePort_11_bits_instructionIndex),
    .vrfWritePort_12_ready                                  (writeQueueVec_12_enq_ready & ~(otherTryToWrite[12])),
    .vrfWritePort_12_valid                                  (_loadUnit_vrfWritePort_12_valid),
    .vrfWritePort_12_bits_vd                                (_loadUnit_vrfWritePort_12_bits_vd),
    .vrfWritePort_12_bits_mask                              (_loadUnit_vrfWritePort_12_bits_mask),
    .vrfWritePort_12_bits_data                              (_loadUnit_vrfWritePort_12_bits_data),
    .vrfWritePort_12_bits_instructionIndex                  (_loadUnit_vrfWritePort_12_bits_instructionIndex),
    .vrfWritePort_13_ready                                  (writeQueueVec_13_enq_ready & ~(otherTryToWrite[13])),
    .vrfWritePort_13_valid                                  (_loadUnit_vrfWritePort_13_valid),
    .vrfWritePort_13_bits_vd                                (_loadUnit_vrfWritePort_13_bits_vd),
    .vrfWritePort_13_bits_mask                              (_loadUnit_vrfWritePort_13_bits_mask),
    .vrfWritePort_13_bits_data                              (_loadUnit_vrfWritePort_13_bits_data),
    .vrfWritePort_13_bits_instructionIndex                  (_loadUnit_vrfWritePort_13_bits_instructionIndex),
    .vrfWritePort_14_ready                                  (writeQueueVec_14_enq_ready & ~(otherTryToWrite[14])),
    .vrfWritePort_14_valid                                  (_loadUnit_vrfWritePort_14_valid),
    .vrfWritePort_14_bits_vd                                (_loadUnit_vrfWritePort_14_bits_vd),
    .vrfWritePort_14_bits_mask                              (_loadUnit_vrfWritePort_14_bits_mask),
    .vrfWritePort_14_bits_data                              (_loadUnit_vrfWritePort_14_bits_data),
    .vrfWritePort_14_bits_instructionIndex                  (_loadUnit_vrfWritePort_14_bits_instructionIndex),
    .vrfWritePort_15_ready                                  (writeQueueVec_15_enq_ready & ~(otherTryToWrite[15])),
    .vrfWritePort_15_valid                                  (_loadUnit_vrfWritePort_15_valid),
    .vrfWritePort_15_bits_vd                                (_loadUnit_vrfWritePort_15_bits_vd),
    .vrfWritePort_15_bits_mask                              (_loadUnit_vrfWritePort_15_bits_mask),
    .vrfWritePort_15_bits_data                              (_loadUnit_vrfWritePort_15_bits_data),
    .vrfWritePort_15_bits_instructionIndex                  (_loadUnit_vrfWritePort_15_bits_instructionIndex),
    .vrfWritePort_16_ready                                  (writeQueueVec_16_enq_ready & ~(otherTryToWrite[16])),
    .vrfWritePort_16_valid                                  (_loadUnit_vrfWritePort_16_valid),
    .vrfWritePort_16_bits_vd                                (_loadUnit_vrfWritePort_16_bits_vd),
    .vrfWritePort_16_bits_mask                              (_loadUnit_vrfWritePort_16_bits_mask),
    .vrfWritePort_16_bits_data                              (_loadUnit_vrfWritePort_16_bits_data),
    .vrfWritePort_16_bits_instructionIndex                  (_loadUnit_vrfWritePort_16_bits_instructionIndex),
    .vrfWritePort_17_ready                                  (writeQueueVec_17_enq_ready & ~(otherTryToWrite[17])),
    .vrfWritePort_17_valid                                  (_loadUnit_vrfWritePort_17_valid),
    .vrfWritePort_17_bits_vd                                (_loadUnit_vrfWritePort_17_bits_vd),
    .vrfWritePort_17_bits_mask                              (_loadUnit_vrfWritePort_17_bits_mask),
    .vrfWritePort_17_bits_data                              (_loadUnit_vrfWritePort_17_bits_data),
    .vrfWritePort_17_bits_instructionIndex                  (_loadUnit_vrfWritePort_17_bits_instructionIndex),
    .vrfWritePort_18_ready                                  (writeQueueVec_18_enq_ready & ~(otherTryToWrite[18])),
    .vrfWritePort_18_valid                                  (_loadUnit_vrfWritePort_18_valid),
    .vrfWritePort_18_bits_vd                                (_loadUnit_vrfWritePort_18_bits_vd),
    .vrfWritePort_18_bits_mask                              (_loadUnit_vrfWritePort_18_bits_mask),
    .vrfWritePort_18_bits_data                              (_loadUnit_vrfWritePort_18_bits_data),
    .vrfWritePort_18_bits_instructionIndex                  (_loadUnit_vrfWritePort_18_bits_instructionIndex),
    .vrfWritePort_19_ready                                  (writeQueueVec_19_enq_ready & ~(otherTryToWrite[19])),
    .vrfWritePort_19_valid                                  (_loadUnit_vrfWritePort_19_valid),
    .vrfWritePort_19_bits_vd                                (_loadUnit_vrfWritePort_19_bits_vd),
    .vrfWritePort_19_bits_mask                              (_loadUnit_vrfWritePort_19_bits_mask),
    .vrfWritePort_19_bits_data                              (_loadUnit_vrfWritePort_19_bits_data),
    .vrfWritePort_19_bits_instructionIndex                  (_loadUnit_vrfWritePort_19_bits_instructionIndex),
    .vrfWritePort_20_ready                                  (writeQueueVec_20_enq_ready & ~(otherTryToWrite[20])),
    .vrfWritePort_20_valid                                  (_loadUnit_vrfWritePort_20_valid),
    .vrfWritePort_20_bits_vd                                (_loadUnit_vrfWritePort_20_bits_vd),
    .vrfWritePort_20_bits_mask                              (_loadUnit_vrfWritePort_20_bits_mask),
    .vrfWritePort_20_bits_data                              (_loadUnit_vrfWritePort_20_bits_data),
    .vrfWritePort_20_bits_instructionIndex                  (_loadUnit_vrfWritePort_20_bits_instructionIndex),
    .vrfWritePort_21_ready                                  (writeQueueVec_21_enq_ready & ~(otherTryToWrite[21])),
    .vrfWritePort_21_valid                                  (_loadUnit_vrfWritePort_21_valid),
    .vrfWritePort_21_bits_vd                                (_loadUnit_vrfWritePort_21_bits_vd),
    .vrfWritePort_21_bits_mask                              (_loadUnit_vrfWritePort_21_bits_mask),
    .vrfWritePort_21_bits_data                              (_loadUnit_vrfWritePort_21_bits_data),
    .vrfWritePort_21_bits_instructionIndex                  (_loadUnit_vrfWritePort_21_bits_instructionIndex),
    .vrfWritePort_22_ready                                  (writeQueueVec_22_enq_ready & ~(otherTryToWrite[22])),
    .vrfWritePort_22_valid                                  (_loadUnit_vrfWritePort_22_valid),
    .vrfWritePort_22_bits_vd                                (_loadUnit_vrfWritePort_22_bits_vd),
    .vrfWritePort_22_bits_mask                              (_loadUnit_vrfWritePort_22_bits_mask),
    .vrfWritePort_22_bits_data                              (_loadUnit_vrfWritePort_22_bits_data),
    .vrfWritePort_22_bits_instructionIndex                  (_loadUnit_vrfWritePort_22_bits_instructionIndex),
    .vrfWritePort_23_ready                                  (writeQueueVec_23_enq_ready & ~(otherTryToWrite[23])),
    .vrfWritePort_23_valid                                  (_loadUnit_vrfWritePort_23_valid),
    .vrfWritePort_23_bits_vd                                (_loadUnit_vrfWritePort_23_bits_vd),
    .vrfWritePort_23_bits_mask                              (_loadUnit_vrfWritePort_23_bits_mask),
    .vrfWritePort_23_bits_data                              (_loadUnit_vrfWritePort_23_bits_data),
    .vrfWritePort_23_bits_instructionIndex                  (_loadUnit_vrfWritePort_23_bits_instructionIndex),
    .vrfWritePort_24_ready                                  (writeQueueVec_24_enq_ready & ~(otherTryToWrite[24])),
    .vrfWritePort_24_valid                                  (_loadUnit_vrfWritePort_24_valid),
    .vrfWritePort_24_bits_vd                                (_loadUnit_vrfWritePort_24_bits_vd),
    .vrfWritePort_24_bits_mask                              (_loadUnit_vrfWritePort_24_bits_mask),
    .vrfWritePort_24_bits_data                              (_loadUnit_vrfWritePort_24_bits_data),
    .vrfWritePort_24_bits_instructionIndex                  (_loadUnit_vrfWritePort_24_bits_instructionIndex),
    .vrfWritePort_25_ready                                  (writeQueueVec_25_enq_ready & ~(otherTryToWrite[25])),
    .vrfWritePort_25_valid                                  (_loadUnit_vrfWritePort_25_valid),
    .vrfWritePort_25_bits_vd                                (_loadUnit_vrfWritePort_25_bits_vd),
    .vrfWritePort_25_bits_mask                              (_loadUnit_vrfWritePort_25_bits_mask),
    .vrfWritePort_25_bits_data                              (_loadUnit_vrfWritePort_25_bits_data),
    .vrfWritePort_25_bits_instructionIndex                  (_loadUnit_vrfWritePort_25_bits_instructionIndex),
    .vrfWritePort_26_ready                                  (writeQueueVec_26_enq_ready & ~(otherTryToWrite[26])),
    .vrfWritePort_26_valid                                  (_loadUnit_vrfWritePort_26_valid),
    .vrfWritePort_26_bits_vd                                (_loadUnit_vrfWritePort_26_bits_vd),
    .vrfWritePort_26_bits_mask                              (_loadUnit_vrfWritePort_26_bits_mask),
    .vrfWritePort_26_bits_data                              (_loadUnit_vrfWritePort_26_bits_data),
    .vrfWritePort_26_bits_instructionIndex                  (_loadUnit_vrfWritePort_26_bits_instructionIndex),
    .vrfWritePort_27_ready                                  (writeQueueVec_27_enq_ready & ~(otherTryToWrite[27])),
    .vrfWritePort_27_valid                                  (_loadUnit_vrfWritePort_27_valid),
    .vrfWritePort_27_bits_vd                                (_loadUnit_vrfWritePort_27_bits_vd),
    .vrfWritePort_27_bits_mask                              (_loadUnit_vrfWritePort_27_bits_mask),
    .vrfWritePort_27_bits_data                              (_loadUnit_vrfWritePort_27_bits_data),
    .vrfWritePort_27_bits_instructionIndex                  (_loadUnit_vrfWritePort_27_bits_instructionIndex),
    .vrfWritePort_28_ready                                  (writeQueueVec_28_enq_ready & ~(otherTryToWrite[28])),
    .vrfWritePort_28_valid                                  (_loadUnit_vrfWritePort_28_valid),
    .vrfWritePort_28_bits_vd                                (_loadUnit_vrfWritePort_28_bits_vd),
    .vrfWritePort_28_bits_mask                              (_loadUnit_vrfWritePort_28_bits_mask),
    .vrfWritePort_28_bits_data                              (_loadUnit_vrfWritePort_28_bits_data),
    .vrfWritePort_28_bits_instructionIndex                  (_loadUnit_vrfWritePort_28_bits_instructionIndex),
    .vrfWritePort_29_ready                                  (writeQueueVec_29_enq_ready & ~(otherTryToWrite[29])),
    .vrfWritePort_29_valid                                  (_loadUnit_vrfWritePort_29_valid),
    .vrfWritePort_29_bits_vd                                (_loadUnit_vrfWritePort_29_bits_vd),
    .vrfWritePort_29_bits_mask                              (_loadUnit_vrfWritePort_29_bits_mask),
    .vrfWritePort_29_bits_data                              (_loadUnit_vrfWritePort_29_bits_data),
    .vrfWritePort_29_bits_instructionIndex                  (_loadUnit_vrfWritePort_29_bits_instructionIndex),
    .vrfWritePort_30_ready                                  (writeQueueVec_30_enq_ready & ~(otherTryToWrite[30])),
    .vrfWritePort_30_valid                                  (_loadUnit_vrfWritePort_30_valid),
    .vrfWritePort_30_bits_vd                                (_loadUnit_vrfWritePort_30_bits_vd),
    .vrfWritePort_30_bits_mask                              (_loadUnit_vrfWritePort_30_bits_mask),
    .vrfWritePort_30_bits_data                              (_loadUnit_vrfWritePort_30_bits_data),
    .vrfWritePort_30_bits_instructionIndex                  (_loadUnit_vrfWritePort_30_bits_instructionIndex),
    .vrfWritePort_31_ready                                  (writeQueueVec_31_enq_ready & ~(otherTryToWrite[31])),
    .vrfWritePort_31_valid                                  (_loadUnit_vrfWritePort_31_valid),
    .vrfWritePort_31_bits_vd                                (_loadUnit_vrfWritePort_31_bits_vd),
    .vrfWritePort_31_bits_mask                              (_loadUnit_vrfWritePort_31_bits_mask),
    .vrfWritePort_31_bits_data                              (_loadUnit_vrfWritePort_31_bits_data),
    .vrfWritePort_31_bits_instructionIndex                  (_loadUnit_vrfWritePort_31_bits_instructionIndex)
  );
  StoreUnit storeUnit (
    .clock                                                  (clock),
    .reset                                                  (reset),
    .lsuRequest_valid                                       (reqEnq_1),
    .lsuRequest_bits_instructionInformation_nf              (request_bits_instructionInformation_nf_0),
    .lsuRequest_bits_instructionInformation_mew             (request_bits_instructionInformation_mew_0),
    .lsuRequest_bits_instructionInformation_mop             (request_bits_instructionInformation_mop_0),
    .lsuRequest_bits_instructionInformation_lumop           (request_bits_instructionInformation_lumop_0),
    .lsuRequest_bits_instructionInformation_eew             (request_bits_instructionInformation_eew_0),
    .lsuRequest_bits_instructionInformation_vs3             (request_bits_instructionInformation_vs3_0),
    .lsuRequest_bits_instructionInformation_isStore         (request_bits_instructionInformation_isStore_0),
    .lsuRequest_bits_instructionInformation_maskedLoadStore (request_bits_instructionInformation_maskedLoadStore_0),
    .lsuRequest_bits_rs1Data                                (request_bits_rs1Data_0),
    .lsuRequest_bits_rs2Data                                (request_bits_rs2Data_0),
    .lsuRequest_bits_instructionIndex                       (request_bits_instructionIndex_0),
    .csrInterface_vl                                        (csrInterface_vl),
    .csrInterface_vStart                                    (csrInterface_vStart),
    .csrInterface_vlmul                                     (csrInterface_vlmul),
    .csrInterface_vSew                                      (csrInterface_vSew),
    .csrInterface_vxrm                                      (csrInterface_vxrm),
    .csrInterface_vta                                       (csrInterface_vta),
    .csrInterface_vma                                       (csrInterface_vma),
    .maskInput                                              (_GEN_16[maskSelect_1]),
    .maskSelect_valid                                       (_storeUnit_maskSelect_valid),
    .maskSelect_bits                                        (_storeUnit_maskSelect_bits),
    .memRequest_ready                                       (axi4Port_aw_ready_0 & dataQueue_enq_ready),
    .memRequest_valid                                       (_storeUnit_memRequest_valid),
    .memRequest_bits_data                                   (dataQueue_enq_bits_data),
    .memRequest_bits_mask                                   (dataQueue_enq_bits_mask),
    .memRequest_bits_index                                  (_storeUnit_memRequest_bits_index),
    .memRequest_bits_address                                (_storeUnit_memRequest_bits_address),
    .status_idle                                            (_storeUnit_status_idle),
    .status_last                                            (_storeUnit_status_last),
    .status_instructionIndex                                (_storeUnit_status_instructionIndex),
    .status_changeMaskGroup                                 (/* unused */),
    .status_startAddress                                    (_storeUnit_status_startAddress),
    .status_endAddress                                      (_storeUnit_status_endAddress),
    .vrfReadDataPorts_0_ready                               (vrfReadDataPorts_0_ready_0 & ~(otherTryReadVrf[0])),
    .vrfReadDataPorts_0_valid                               (_storeUnit_vrfReadDataPorts_0_valid),
    .vrfReadDataPorts_0_bits_vs                             (_storeUnit_vrfReadDataPorts_0_bits_vs),
    .vrfReadDataPorts_0_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_0_bits_instructionIndex),
    .vrfReadDataPorts_1_ready                               (vrfReadDataPorts_1_ready_0 & ~(otherTryReadVrf[1])),
    .vrfReadDataPorts_1_valid                               (_storeUnit_vrfReadDataPorts_1_valid),
    .vrfReadDataPorts_1_bits_vs                             (_storeUnit_vrfReadDataPorts_1_bits_vs),
    .vrfReadDataPorts_1_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_1_bits_instructionIndex),
    .vrfReadDataPorts_2_ready                               (vrfReadDataPorts_2_ready_0 & ~(otherTryReadVrf[2])),
    .vrfReadDataPorts_2_valid                               (_storeUnit_vrfReadDataPorts_2_valid),
    .vrfReadDataPorts_2_bits_vs                             (_storeUnit_vrfReadDataPorts_2_bits_vs),
    .vrfReadDataPorts_2_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_2_bits_instructionIndex),
    .vrfReadDataPorts_3_ready                               (vrfReadDataPorts_3_ready_0 & ~(otherTryReadVrf[3])),
    .vrfReadDataPorts_3_valid                               (_storeUnit_vrfReadDataPorts_3_valid),
    .vrfReadDataPorts_3_bits_vs                             (_storeUnit_vrfReadDataPorts_3_bits_vs),
    .vrfReadDataPorts_3_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_3_bits_instructionIndex),
    .vrfReadDataPorts_4_ready                               (vrfReadDataPorts_4_ready_0 & ~(otherTryReadVrf[4])),
    .vrfReadDataPorts_4_valid                               (_storeUnit_vrfReadDataPorts_4_valid),
    .vrfReadDataPorts_4_bits_vs                             (_storeUnit_vrfReadDataPorts_4_bits_vs),
    .vrfReadDataPorts_4_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_4_bits_instructionIndex),
    .vrfReadDataPorts_5_ready                               (vrfReadDataPorts_5_ready_0 & ~(otherTryReadVrf[5])),
    .vrfReadDataPorts_5_valid                               (_storeUnit_vrfReadDataPorts_5_valid),
    .vrfReadDataPorts_5_bits_vs                             (_storeUnit_vrfReadDataPorts_5_bits_vs),
    .vrfReadDataPorts_5_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_5_bits_instructionIndex),
    .vrfReadDataPorts_6_ready                               (vrfReadDataPorts_6_ready_0 & ~(otherTryReadVrf[6])),
    .vrfReadDataPorts_6_valid                               (_storeUnit_vrfReadDataPorts_6_valid),
    .vrfReadDataPorts_6_bits_vs                             (_storeUnit_vrfReadDataPorts_6_bits_vs),
    .vrfReadDataPorts_6_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_6_bits_instructionIndex),
    .vrfReadDataPorts_7_ready                               (vrfReadDataPorts_7_ready_0 & ~(otherTryReadVrf[7])),
    .vrfReadDataPorts_7_valid                               (_storeUnit_vrfReadDataPorts_7_valid),
    .vrfReadDataPorts_7_bits_vs                             (_storeUnit_vrfReadDataPorts_7_bits_vs),
    .vrfReadDataPorts_7_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_7_bits_instructionIndex),
    .vrfReadDataPorts_8_ready                               (vrfReadDataPorts_8_ready_0 & ~(otherTryReadVrf[8])),
    .vrfReadDataPorts_8_valid                               (_storeUnit_vrfReadDataPorts_8_valid),
    .vrfReadDataPorts_8_bits_vs                             (_storeUnit_vrfReadDataPorts_8_bits_vs),
    .vrfReadDataPorts_8_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_8_bits_instructionIndex),
    .vrfReadDataPorts_9_ready                               (vrfReadDataPorts_9_ready_0 & ~(otherTryReadVrf[9])),
    .vrfReadDataPorts_9_valid                               (_storeUnit_vrfReadDataPorts_9_valid),
    .vrfReadDataPorts_9_bits_vs                             (_storeUnit_vrfReadDataPorts_9_bits_vs),
    .vrfReadDataPorts_9_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_9_bits_instructionIndex),
    .vrfReadDataPorts_10_ready                              (vrfReadDataPorts_10_ready_0 & ~(otherTryReadVrf[10])),
    .vrfReadDataPorts_10_valid                              (_storeUnit_vrfReadDataPorts_10_valid),
    .vrfReadDataPorts_10_bits_vs                            (_storeUnit_vrfReadDataPorts_10_bits_vs),
    .vrfReadDataPorts_10_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_10_bits_instructionIndex),
    .vrfReadDataPorts_11_ready                              (vrfReadDataPorts_11_ready_0 & ~(otherTryReadVrf[11])),
    .vrfReadDataPorts_11_valid                              (_storeUnit_vrfReadDataPorts_11_valid),
    .vrfReadDataPorts_11_bits_vs                            (_storeUnit_vrfReadDataPorts_11_bits_vs),
    .vrfReadDataPorts_11_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_11_bits_instructionIndex),
    .vrfReadDataPorts_12_ready                              (vrfReadDataPorts_12_ready_0 & ~(otherTryReadVrf[12])),
    .vrfReadDataPorts_12_valid                              (_storeUnit_vrfReadDataPorts_12_valid),
    .vrfReadDataPorts_12_bits_vs                            (_storeUnit_vrfReadDataPorts_12_bits_vs),
    .vrfReadDataPorts_12_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_12_bits_instructionIndex),
    .vrfReadDataPorts_13_ready                              (vrfReadDataPorts_13_ready_0 & ~(otherTryReadVrf[13])),
    .vrfReadDataPorts_13_valid                              (_storeUnit_vrfReadDataPorts_13_valid),
    .vrfReadDataPorts_13_bits_vs                            (_storeUnit_vrfReadDataPorts_13_bits_vs),
    .vrfReadDataPorts_13_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_13_bits_instructionIndex),
    .vrfReadDataPorts_14_ready                              (vrfReadDataPorts_14_ready_0 & ~(otherTryReadVrf[14])),
    .vrfReadDataPorts_14_valid                              (_storeUnit_vrfReadDataPorts_14_valid),
    .vrfReadDataPorts_14_bits_vs                            (_storeUnit_vrfReadDataPorts_14_bits_vs),
    .vrfReadDataPorts_14_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_14_bits_instructionIndex),
    .vrfReadDataPorts_15_ready                              (vrfReadDataPorts_15_ready_0 & ~(otherTryReadVrf[15])),
    .vrfReadDataPorts_15_valid                              (_storeUnit_vrfReadDataPorts_15_valid),
    .vrfReadDataPorts_15_bits_vs                            (_storeUnit_vrfReadDataPorts_15_bits_vs),
    .vrfReadDataPorts_15_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_15_bits_instructionIndex),
    .vrfReadDataPorts_16_ready                              (vrfReadDataPorts_16_ready_0 & ~(otherTryReadVrf[16])),
    .vrfReadDataPorts_16_valid                              (_storeUnit_vrfReadDataPorts_16_valid),
    .vrfReadDataPorts_16_bits_vs                            (_storeUnit_vrfReadDataPorts_16_bits_vs),
    .vrfReadDataPorts_16_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_16_bits_instructionIndex),
    .vrfReadDataPorts_17_ready                              (vrfReadDataPorts_17_ready_0 & ~(otherTryReadVrf[17])),
    .vrfReadDataPorts_17_valid                              (_storeUnit_vrfReadDataPorts_17_valid),
    .vrfReadDataPorts_17_bits_vs                            (_storeUnit_vrfReadDataPorts_17_bits_vs),
    .vrfReadDataPorts_17_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_17_bits_instructionIndex),
    .vrfReadDataPorts_18_ready                              (vrfReadDataPorts_18_ready_0 & ~(otherTryReadVrf[18])),
    .vrfReadDataPorts_18_valid                              (_storeUnit_vrfReadDataPorts_18_valid),
    .vrfReadDataPorts_18_bits_vs                            (_storeUnit_vrfReadDataPorts_18_bits_vs),
    .vrfReadDataPorts_18_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_18_bits_instructionIndex),
    .vrfReadDataPorts_19_ready                              (vrfReadDataPorts_19_ready_0 & ~(otherTryReadVrf[19])),
    .vrfReadDataPorts_19_valid                              (_storeUnit_vrfReadDataPorts_19_valid),
    .vrfReadDataPorts_19_bits_vs                            (_storeUnit_vrfReadDataPorts_19_bits_vs),
    .vrfReadDataPorts_19_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_19_bits_instructionIndex),
    .vrfReadDataPorts_20_ready                              (vrfReadDataPorts_20_ready_0 & ~(otherTryReadVrf[20])),
    .vrfReadDataPorts_20_valid                              (_storeUnit_vrfReadDataPorts_20_valid),
    .vrfReadDataPorts_20_bits_vs                            (_storeUnit_vrfReadDataPorts_20_bits_vs),
    .vrfReadDataPorts_20_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_20_bits_instructionIndex),
    .vrfReadDataPorts_21_ready                              (vrfReadDataPorts_21_ready_0 & ~(otherTryReadVrf[21])),
    .vrfReadDataPorts_21_valid                              (_storeUnit_vrfReadDataPorts_21_valid),
    .vrfReadDataPorts_21_bits_vs                            (_storeUnit_vrfReadDataPorts_21_bits_vs),
    .vrfReadDataPorts_21_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_21_bits_instructionIndex),
    .vrfReadDataPorts_22_ready                              (vrfReadDataPorts_22_ready_0 & ~(otherTryReadVrf[22])),
    .vrfReadDataPorts_22_valid                              (_storeUnit_vrfReadDataPorts_22_valid),
    .vrfReadDataPorts_22_bits_vs                            (_storeUnit_vrfReadDataPorts_22_bits_vs),
    .vrfReadDataPorts_22_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_22_bits_instructionIndex),
    .vrfReadDataPorts_23_ready                              (vrfReadDataPorts_23_ready_0 & ~(otherTryReadVrf[23])),
    .vrfReadDataPorts_23_valid                              (_storeUnit_vrfReadDataPorts_23_valid),
    .vrfReadDataPorts_23_bits_vs                            (_storeUnit_vrfReadDataPorts_23_bits_vs),
    .vrfReadDataPorts_23_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_23_bits_instructionIndex),
    .vrfReadDataPorts_24_ready                              (vrfReadDataPorts_24_ready_0 & ~(otherTryReadVrf[24])),
    .vrfReadDataPorts_24_valid                              (_storeUnit_vrfReadDataPorts_24_valid),
    .vrfReadDataPorts_24_bits_vs                            (_storeUnit_vrfReadDataPorts_24_bits_vs),
    .vrfReadDataPorts_24_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_24_bits_instructionIndex),
    .vrfReadDataPorts_25_ready                              (vrfReadDataPorts_25_ready_0 & ~(otherTryReadVrf[25])),
    .vrfReadDataPorts_25_valid                              (_storeUnit_vrfReadDataPorts_25_valid),
    .vrfReadDataPorts_25_bits_vs                            (_storeUnit_vrfReadDataPorts_25_bits_vs),
    .vrfReadDataPorts_25_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_25_bits_instructionIndex),
    .vrfReadDataPorts_26_ready                              (vrfReadDataPorts_26_ready_0 & ~(otherTryReadVrf[26])),
    .vrfReadDataPorts_26_valid                              (_storeUnit_vrfReadDataPorts_26_valid),
    .vrfReadDataPorts_26_bits_vs                            (_storeUnit_vrfReadDataPorts_26_bits_vs),
    .vrfReadDataPorts_26_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_26_bits_instructionIndex),
    .vrfReadDataPorts_27_ready                              (vrfReadDataPorts_27_ready_0 & ~(otherTryReadVrf[27])),
    .vrfReadDataPorts_27_valid                              (_storeUnit_vrfReadDataPorts_27_valid),
    .vrfReadDataPorts_27_bits_vs                            (_storeUnit_vrfReadDataPorts_27_bits_vs),
    .vrfReadDataPorts_27_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_27_bits_instructionIndex),
    .vrfReadDataPorts_28_ready                              (vrfReadDataPorts_28_ready_0 & ~(otherTryReadVrf[28])),
    .vrfReadDataPorts_28_valid                              (_storeUnit_vrfReadDataPorts_28_valid),
    .vrfReadDataPorts_28_bits_vs                            (_storeUnit_vrfReadDataPorts_28_bits_vs),
    .vrfReadDataPorts_28_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_28_bits_instructionIndex),
    .vrfReadDataPorts_29_ready                              (vrfReadDataPorts_29_ready_0 & ~(otherTryReadVrf[29])),
    .vrfReadDataPorts_29_valid                              (_storeUnit_vrfReadDataPorts_29_valid),
    .vrfReadDataPorts_29_bits_vs                            (_storeUnit_vrfReadDataPorts_29_bits_vs),
    .vrfReadDataPorts_29_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_29_bits_instructionIndex),
    .vrfReadDataPorts_30_ready                              (vrfReadDataPorts_30_ready_0 & ~(otherTryReadVrf[30])),
    .vrfReadDataPorts_30_valid                              (_storeUnit_vrfReadDataPorts_30_valid),
    .vrfReadDataPorts_30_bits_vs                            (_storeUnit_vrfReadDataPorts_30_bits_vs),
    .vrfReadDataPorts_30_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_30_bits_instructionIndex),
    .vrfReadDataPorts_31_ready                              (vrfReadDataPorts_31_ready_0 & ~(otherTryReadVrf[31])),
    .vrfReadDataPorts_31_valid                              (_storeUnit_vrfReadDataPorts_31_valid),
    .vrfReadDataPorts_31_bits_vs                            (_storeUnit_vrfReadDataPorts_31_bits_vs),
    .vrfReadDataPorts_31_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_31_bits_instructionIndex),
    .vrfReadResults_0_valid                                 (vrfReadResults_0_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_0_bits                                  (vrfReadResults_0_bits),
    .vrfReadResults_1_valid                                 (vrfReadResults_1_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_1_bits                                  (vrfReadResults_1_bits),
    .vrfReadResults_2_valid                                 (vrfReadResults_2_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_2_bits                                  (vrfReadResults_2_bits),
    .vrfReadResults_3_valid                                 (vrfReadResults_3_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_3_bits                                  (vrfReadResults_3_bits),
    .vrfReadResults_4_valid                                 (vrfReadResults_4_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_4_bits                                  (vrfReadResults_4_bits),
    .vrfReadResults_5_valid                                 (vrfReadResults_5_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_5_bits                                  (vrfReadResults_5_bits),
    .vrfReadResults_6_valid                                 (vrfReadResults_6_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_6_bits                                  (vrfReadResults_6_bits),
    .vrfReadResults_7_valid                                 (vrfReadResults_7_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_7_bits                                  (vrfReadResults_7_bits),
    .vrfReadResults_8_valid                                 (vrfReadResults_8_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_8_bits                                  (vrfReadResults_8_bits),
    .vrfReadResults_9_valid                                 (vrfReadResults_9_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_9_bits                                  (vrfReadResults_9_bits),
    .vrfReadResults_10_valid                                (vrfReadResults_10_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_10_bits                                 (vrfReadResults_10_bits),
    .vrfReadResults_11_valid                                (vrfReadResults_11_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_11_bits                                 (vrfReadResults_11_bits),
    .vrfReadResults_12_valid                                (vrfReadResults_12_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_12_bits                                 (vrfReadResults_12_bits),
    .vrfReadResults_13_valid                                (vrfReadResults_13_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_13_bits                                 (vrfReadResults_13_bits),
    .vrfReadResults_14_valid                                (vrfReadResults_14_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_14_bits                                 (vrfReadResults_14_bits),
    .vrfReadResults_15_valid                                (vrfReadResults_15_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_15_bits                                 (vrfReadResults_15_bits),
    .vrfReadResults_16_valid                                (vrfReadResults_16_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_16_bits                                 (vrfReadResults_16_bits),
    .vrfReadResults_17_valid                                (vrfReadResults_17_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_17_bits                                 (vrfReadResults_17_bits),
    .vrfReadResults_18_valid                                (vrfReadResults_18_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_18_bits                                 (vrfReadResults_18_bits),
    .vrfReadResults_19_valid                                (vrfReadResults_19_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_19_bits                                 (vrfReadResults_19_bits),
    .vrfReadResults_20_valid                                (vrfReadResults_20_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_20_bits                                 (vrfReadResults_20_bits),
    .vrfReadResults_21_valid                                (vrfReadResults_21_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_21_bits                                 (vrfReadResults_21_bits),
    .vrfReadResults_22_valid                                (vrfReadResults_22_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_22_bits                                 (vrfReadResults_22_bits),
    .vrfReadResults_23_valid                                (vrfReadResults_23_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_23_bits                                 (vrfReadResults_23_bits),
    .vrfReadResults_24_valid                                (vrfReadResults_24_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_24_bits                                 (vrfReadResults_24_bits),
    .vrfReadResults_25_valid                                (vrfReadResults_25_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_25_bits                                 (vrfReadResults_25_bits),
    .vrfReadResults_26_valid                                (vrfReadResults_26_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_26_bits                                 (vrfReadResults_26_bits),
    .vrfReadResults_27_valid                                (vrfReadResults_27_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_27_bits                                 (vrfReadResults_27_bits),
    .vrfReadResults_28_valid                                (vrfReadResults_28_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_28_bits                                 (vrfReadResults_28_bits),
    .vrfReadResults_29_valid                                (vrfReadResults_29_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_29_bits                                 (vrfReadResults_29_bits),
    .vrfReadResults_30_valid                                (vrfReadResults_30_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_30_bits                                 (vrfReadResults_30_bits),
    .vrfReadResults_31_valid                                (vrfReadResults_31_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_31_bits                                 (vrfReadResults_31_bits),
    .storeResponse                                          (axi4Port_b_valid_0)
  );
  SimpleAccessUnit otherUnit (
    .clock                                                  (clock),
    .reset                                                  (reset),
    .lsuRequest_valid                                       (reqEnq_2),
    .lsuRequest_bits_instructionInformation_nf              (request_bits_instructionInformation_nf_0),
    .lsuRequest_bits_instructionInformation_mew             (request_bits_instructionInformation_mew_0),
    .lsuRequest_bits_instructionInformation_mop             (request_bits_instructionInformation_mop_0),
    .lsuRequest_bits_instructionInformation_lumop           (request_bits_instructionInformation_lumop_0),
    .lsuRequest_bits_instructionInformation_eew             (request_bits_instructionInformation_eew_0),
    .lsuRequest_bits_instructionInformation_vs3             (request_bits_instructionInformation_vs3_0),
    .lsuRequest_bits_instructionInformation_isStore         (request_bits_instructionInformation_isStore_0),
    .lsuRequest_bits_instructionInformation_maskedLoadStore (request_bits_instructionInformation_maskedLoadStore_0),
    .lsuRequest_bits_rs1Data                                (request_bits_rs1Data_0),
    .lsuRequest_bits_rs2Data                                (request_bits_rs2Data_0),
    .lsuRequest_bits_instructionIndex                       (request_bits_instructionIndex_0),
    .vrfReadDataPorts_ready                                 (otherUnit_vrfReadDataPorts_ready),
    .vrfReadDataPorts_valid                                 (_otherUnit_vrfReadDataPorts_valid),
    .vrfReadDataPorts_bits_vs                               (_otherUnit_vrfReadDataPorts_bits_vs),
    .vrfReadDataPorts_bits_instructionIndex                 (_otherUnit_vrfReadDataPorts_bits_instructionIndex),
    .vrfReadResults_valid                                   (otherUnitTargetQueue_deq_ready),
    .vrfReadResults_bits
      ((otherUnitTargetQueue_deq_bits[0] ? otherUnitDataQueueVec_0_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[1] ? otherUnitDataQueueVec_1_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[2] ? otherUnitDataQueueVec_2_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[3] ? otherUnitDataQueueVec_3_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[4] ? otherUnitDataQueueVec_4_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[5] ? otherUnitDataQueueVec_5_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[6] ? otherUnitDataQueueVec_6_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[7] ? otherUnitDataQueueVec_7_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[8] ? otherUnitDataQueueVec_8_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[9] ? otherUnitDataQueueVec_9_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[10] ? otherUnitDataQueueVec_10_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[11] ? otherUnitDataQueueVec_11_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[12] ? otherUnitDataQueueVec_12_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[13] ? otherUnitDataQueueVec_13_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[14] ? otherUnitDataQueueVec_14_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[15] ? otherUnitDataQueueVec_15_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[16] ? otherUnitDataQueueVec_16_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[17] ? otherUnitDataQueueVec_17_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[18] ? otherUnitDataQueueVec_18_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[19] ? otherUnitDataQueueVec_19_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[20] ? otherUnitDataQueueVec_20_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[21] ? otherUnitDataQueueVec_21_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[22] ? otherUnitDataQueueVec_22_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[23] ? otherUnitDataQueueVec_23_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[24] ? otherUnitDataQueueVec_24_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[25] ? otherUnitDataQueueVec_25_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[26] ? otherUnitDataQueueVec_26_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[27] ? otherUnitDataQueueVec_27_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[28] ? otherUnitDataQueueVec_28_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[29] ? otherUnitDataQueueVec_29_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[30] ? otherUnitDataQueueVec_30_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[31] ? otherUnitDataQueueVec_31_deq_bits : 32'h0)),
    .offsetReadResult_0_valid                               (offsetReadResult_0_valid),
    .offsetReadResult_0_bits                                (offsetReadResult_0_bits),
    .offsetReadResult_1_valid                               (offsetReadResult_1_valid),
    .offsetReadResult_1_bits                                (offsetReadResult_1_bits),
    .offsetReadResult_2_valid                               (offsetReadResult_2_valid),
    .offsetReadResult_2_bits                                (offsetReadResult_2_bits),
    .offsetReadResult_3_valid                               (offsetReadResult_3_valid),
    .offsetReadResult_3_bits                                (offsetReadResult_3_bits),
    .offsetReadResult_4_valid                               (offsetReadResult_4_valid),
    .offsetReadResult_4_bits                                (offsetReadResult_4_bits),
    .offsetReadResult_5_valid                               (offsetReadResult_5_valid),
    .offsetReadResult_5_bits                                (offsetReadResult_5_bits),
    .offsetReadResult_6_valid                               (offsetReadResult_6_valid),
    .offsetReadResult_6_bits                                (offsetReadResult_6_bits),
    .offsetReadResult_7_valid                               (offsetReadResult_7_valid),
    .offsetReadResult_7_bits                                (offsetReadResult_7_bits),
    .offsetReadResult_8_valid                               (offsetReadResult_8_valid),
    .offsetReadResult_8_bits                                (offsetReadResult_8_bits),
    .offsetReadResult_9_valid                               (offsetReadResult_9_valid),
    .offsetReadResult_9_bits                                (offsetReadResult_9_bits),
    .offsetReadResult_10_valid                              (offsetReadResult_10_valid),
    .offsetReadResult_10_bits                               (offsetReadResult_10_bits),
    .offsetReadResult_11_valid                              (offsetReadResult_11_valid),
    .offsetReadResult_11_bits                               (offsetReadResult_11_bits),
    .offsetReadResult_12_valid                              (offsetReadResult_12_valid),
    .offsetReadResult_12_bits                               (offsetReadResult_12_bits),
    .offsetReadResult_13_valid                              (offsetReadResult_13_valid),
    .offsetReadResult_13_bits                               (offsetReadResult_13_bits),
    .offsetReadResult_14_valid                              (offsetReadResult_14_valid),
    .offsetReadResult_14_bits                               (offsetReadResult_14_bits),
    .offsetReadResult_15_valid                              (offsetReadResult_15_valid),
    .offsetReadResult_15_bits                               (offsetReadResult_15_bits),
    .offsetReadResult_16_valid                              (offsetReadResult_16_valid),
    .offsetReadResult_16_bits                               (offsetReadResult_16_bits),
    .offsetReadResult_17_valid                              (offsetReadResult_17_valid),
    .offsetReadResult_17_bits                               (offsetReadResult_17_bits),
    .offsetReadResult_18_valid                              (offsetReadResult_18_valid),
    .offsetReadResult_18_bits                               (offsetReadResult_18_bits),
    .offsetReadResult_19_valid                              (offsetReadResult_19_valid),
    .offsetReadResult_19_bits                               (offsetReadResult_19_bits),
    .offsetReadResult_20_valid                              (offsetReadResult_20_valid),
    .offsetReadResult_20_bits                               (offsetReadResult_20_bits),
    .offsetReadResult_21_valid                              (offsetReadResult_21_valid),
    .offsetReadResult_21_bits                               (offsetReadResult_21_bits),
    .offsetReadResult_22_valid                              (offsetReadResult_22_valid),
    .offsetReadResult_22_bits                               (offsetReadResult_22_bits),
    .offsetReadResult_23_valid                              (offsetReadResult_23_valid),
    .offsetReadResult_23_bits                               (offsetReadResult_23_bits),
    .offsetReadResult_24_valid                              (offsetReadResult_24_valid),
    .offsetReadResult_24_bits                               (offsetReadResult_24_bits),
    .offsetReadResult_25_valid                              (offsetReadResult_25_valid),
    .offsetReadResult_25_bits                               (offsetReadResult_25_bits),
    .offsetReadResult_26_valid                              (offsetReadResult_26_valid),
    .offsetReadResult_26_bits                               (offsetReadResult_26_bits),
    .offsetReadResult_27_valid                              (offsetReadResult_27_valid),
    .offsetReadResult_27_bits                               (offsetReadResult_27_bits),
    .offsetReadResult_28_valid                              (offsetReadResult_28_valid),
    .offsetReadResult_28_bits                               (offsetReadResult_28_bits),
    .offsetReadResult_29_valid                              (offsetReadResult_29_valid),
    .offsetReadResult_29_bits                               (offsetReadResult_29_bits),
    .offsetReadResult_30_valid                              (offsetReadResult_30_valid),
    .offsetReadResult_30_bits                               (offsetReadResult_30_bits),
    .offsetReadResult_31_valid                              (offsetReadResult_31_valid),
    .offsetReadResult_31_bits                               (offsetReadResult_31_bits),
    .maskInput                                              (_GEN_17[maskSelect_2]),
    .maskSelect_valid                                       (_otherUnit_maskSelect_valid),
    .maskSelect_bits                                        (_otherUnit_maskSelect_bits),
    .memReadRequest_ready                                   (simpleSourceQueue_enq_ready & simpleAccessPorts_ar_ready_0),
    .memReadRequest_valid                                   (_otherUnit_memReadRequest_valid),
    .memReadRequest_bits_address                            (simpleAccessPorts_ar_bits_addr_0),
    .memReadRequest_bits_source                             (simpleSourceQueue_enq_bits),
    .memReadResponse_ready                                  (simpleAccessPorts_r_ready_0),
    .memReadResponse_valid                                  (simpleAccessPorts_r_valid_0),
    .memReadResponse_bits_data                              (simpleAccessPorts_r_bits_data_0),
    .memReadResponse_bits_source                            (simpleSourceQueue_deq_bits),
    .memWriteRequest_ready                                  (simpleAccessPorts_aw_ready_0 & simpleDataQueue_enq_ready),
    .memWriteRequest_valid                                  (_otherUnit_memWriteRequest_valid),
    .memWriteRequest_bits_data                              (simpleDataQueue_enq_bits_data),
    .memWriteRequest_bits_mask                              (simpleDataQueue_enq_bits_mask),
    .memWriteRequest_bits_source                            (_otherUnit_memWriteRequest_bits_source),
    .memWriteRequest_bits_address                           (_otherUnit_memWriteRequest_bits_address),
    .memWriteRequest_bits_size                              (_otherUnit_memWriteRequest_bits_size),
    .vrfWritePort_ready                                     (|(_otherUnit_status_targetLane & {otherUnit_vrfWritePort_ready_hi, otherUnit_vrfWritePort_ready_lo})),
    .vrfWritePort_valid                                     (_otherUnit_vrfWritePort_valid),
    .vrfWritePort_bits_vd                                   (_otherUnit_vrfWritePort_bits_vd),
    .vrfWritePort_bits_mask                                 (_otherUnit_vrfWritePort_bits_mask),
    .vrfWritePort_bits_data                                 (_otherUnit_vrfWritePort_bits_data),
    .vrfWritePort_bits_last                                 (_otherUnit_vrfWritePort_bits_last),
    .vrfWritePort_bits_instructionIndex                     (_otherUnit_vrfWritePort_bits_instructionIndex),
    .csrInterface_vl                                        (csrInterface_vl),
    .csrInterface_vStart                                    (csrInterface_vStart),
    .csrInterface_vlmul                                     (csrInterface_vlmul),
    .csrInterface_vSew                                      (csrInterface_vSew),
    .csrInterface_vxrm                                      (csrInterface_vxrm),
    .csrInterface_vta                                       (csrInterface_vta),
    .csrInterface_vma                                       (csrInterface_vma),
    .status_idle                                            (_otherUnit_status_idle),
    .status_last                                            (_otherUnit_status_last),
    .status_instructionIndex                                (_otherUnit_status_instructionIndex),
    .status_targetLane                                      (_otherUnit_status_targetLane),
    .status_isStore                                         (_otherUnit_status_isStore),
    .offsetRelease_0                                        (_otherUnit_offsetRelease_0),
    .offsetRelease_1                                        (_otherUnit_offsetRelease_1),
    .offsetRelease_2                                        (_otherUnit_offsetRelease_2),
    .offsetRelease_3                                        (_otherUnit_offsetRelease_3),
    .offsetRelease_4                                        (_otherUnit_offsetRelease_4),
    .offsetRelease_5                                        (_otherUnit_offsetRelease_5),
    .offsetRelease_6                                        (_otherUnit_offsetRelease_6),
    .offsetRelease_7                                        (_otherUnit_offsetRelease_7),
    .offsetRelease_8                                        (_otherUnit_offsetRelease_8),
    .offsetRelease_9                                        (_otherUnit_offsetRelease_9),
    .offsetRelease_10                                       (_otherUnit_offsetRelease_10),
    .offsetRelease_11                                       (_otherUnit_offsetRelease_11),
    .offsetRelease_12                                       (_otherUnit_offsetRelease_12),
    .offsetRelease_13                                       (_otherUnit_offsetRelease_13),
    .offsetRelease_14                                       (_otherUnit_offsetRelease_14),
    .offsetRelease_15                                       (_otherUnit_offsetRelease_15),
    .offsetRelease_16                                       (_otherUnit_offsetRelease_16),
    .offsetRelease_17                                       (_otherUnit_offsetRelease_17),
    .offsetRelease_18                                       (_otherUnit_offsetRelease_18),
    .offsetRelease_19                                       (_otherUnit_offsetRelease_19),
    .offsetRelease_20                                       (_otherUnit_offsetRelease_20),
    .offsetRelease_21                                       (_otherUnit_offsetRelease_21),
    .offsetRelease_22                                       (_otherUnit_offsetRelease_22),
    .offsetRelease_23                                       (_otherUnit_offsetRelease_23),
    .offsetRelease_24                                       (_otherUnit_offsetRelease_24),
    .offsetRelease_25                                       (_otherUnit_offsetRelease_25),
    .offsetRelease_26                                       (_otherUnit_offsetRelease_26),
    .offsetRelease_27                                       (_otherUnit_offsetRelease_27),
    .offsetRelease_28                                       (_otherUnit_offsetRelease_28),
    .offsetRelease_29                                       (_otherUnit_offsetRelease_29),
    .offsetRelease_30                                       (_otherUnit_offsetRelease_30),
    .offsetRelease_31                                       (_otherUnit_offsetRelease_31)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_0_writeValid_T & ~(_writeQueueVec_fifo_empty & writeQueueVec_0_deq_ready))),
    .pop_req_n    (~(writeQueueVec_0_deq_ready & ~_writeQueueVec_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn),
    .empty        (_writeQueueVec_fifo_empty),
    .almost_empty (writeQueueVec_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_0_almostFull),
    .full         (_writeQueueVec_fifo_full),
    .error        (_writeQueueVec_fifo_error),
    .data_out     (_writeQueueVec_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_1_writeValid_T & ~(_writeQueueVec_fifo_1_empty & writeQueueVec_1_deq_ready))),
    .pop_req_n    (~(writeQueueVec_1_deq_ready & ~_writeQueueVec_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_1),
    .empty        (_writeQueueVec_fifo_1_empty),
    .almost_empty (writeQueueVec_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_1_almostFull),
    .full         (_writeQueueVec_fifo_1_full),
    .error        (_writeQueueVec_fifo_1_error),
    .data_out     (_writeQueueVec_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_2_writeValid_T & ~(_writeQueueVec_fifo_2_empty & writeQueueVec_2_deq_ready))),
    .pop_req_n    (~(writeQueueVec_2_deq_ready & ~_writeQueueVec_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_2),
    .empty        (_writeQueueVec_fifo_2_empty),
    .almost_empty (writeQueueVec_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_2_almostFull),
    .full         (_writeQueueVec_fifo_2_full),
    .error        (_writeQueueVec_fifo_2_error),
    .data_out     (_writeQueueVec_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_3_writeValid_T & ~(_writeQueueVec_fifo_3_empty & writeQueueVec_3_deq_ready))),
    .pop_req_n    (~(writeQueueVec_3_deq_ready & ~_writeQueueVec_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_3),
    .empty        (_writeQueueVec_fifo_3_empty),
    .almost_empty (writeQueueVec_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_3_almostFull),
    .full         (_writeQueueVec_fifo_3_full),
    .error        (_writeQueueVec_fifo_3_error),
    .data_out     (_writeQueueVec_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_4_writeValid_T & ~(_writeQueueVec_fifo_4_empty & writeQueueVec_4_deq_ready))),
    .pop_req_n    (~(writeQueueVec_4_deq_ready & ~_writeQueueVec_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_4),
    .empty        (_writeQueueVec_fifo_4_empty),
    .almost_empty (writeQueueVec_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_4_almostFull),
    .full         (_writeQueueVec_fifo_4_full),
    .error        (_writeQueueVec_fifo_4_error),
    .data_out     (_writeQueueVec_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_5_writeValid_T & ~(_writeQueueVec_fifo_5_empty & writeQueueVec_5_deq_ready))),
    .pop_req_n    (~(writeQueueVec_5_deq_ready & ~_writeQueueVec_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_5),
    .empty        (_writeQueueVec_fifo_5_empty),
    .almost_empty (writeQueueVec_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_5_almostFull),
    .full         (_writeQueueVec_fifo_5_full),
    .error        (_writeQueueVec_fifo_5_error),
    .data_out     (_writeQueueVec_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_6_writeValid_T & ~(_writeQueueVec_fifo_6_empty & writeQueueVec_6_deq_ready))),
    .pop_req_n    (~(writeQueueVec_6_deq_ready & ~_writeQueueVec_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_6),
    .empty        (_writeQueueVec_fifo_6_empty),
    .almost_empty (writeQueueVec_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_6_almostFull),
    .full         (_writeQueueVec_fifo_6_full),
    .error        (_writeQueueVec_fifo_6_error),
    .data_out     (_writeQueueVec_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_7_writeValid_T & ~(_writeQueueVec_fifo_7_empty & writeQueueVec_7_deq_ready))),
    .pop_req_n    (~(writeQueueVec_7_deq_ready & ~_writeQueueVec_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_7),
    .empty        (_writeQueueVec_fifo_7_empty),
    .almost_empty (writeQueueVec_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_7_almostFull),
    .full         (_writeQueueVec_fifo_7_full),
    .error        (_writeQueueVec_fifo_7_error),
    .data_out     (_writeQueueVec_fifo_7_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_8_writeValid_T & ~(_writeQueueVec_fifo_8_empty & writeQueueVec_8_deq_ready))),
    .pop_req_n    (~(writeQueueVec_8_deq_ready & ~_writeQueueVec_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_8),
    .empty        (_writeQueueVec_fifo_8_empty),
    .almost_empty (writeQueueVec_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_8_almostFull),
    .full         (_writeQueueVec_fifo_8_full),
    .error        (_writeQueueVec_fifo_8_error),
    .data_out     (_writeQueueVec_fifo_8_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_9_writeValid_T & ~(_writeQueueVec_fifo_9_empty & writeQueueVec_9_deq_ready))),
    .pop_req_n    (~(writeQueueVec_9_deq_ready & ~_writeQueueVec_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_9),
    .empty        (_writeQueueVec_fifo_9_empty),
    .almost_empty (writeQueueVec_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_9_almostFull),
    .full         (_writeQueueVec_fifo_9_full),
    .error        (_writeQueueVec_fifo_9_error),
    .data_out     (_writeQueueVec_fifo_9_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_10_writeValid_T & ~(_writeQueueVec_fifo_10_empty & writeQueueVec_10_deq_ready))),
    .pop_req_n    (~(writeQueueVec_10_deq_ready & ~_writeQueueVec_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_10),
    .empty        (_writeQueueVec_fifo_10_empty),
    .almost_empty (writeQueueVec_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_10_almostFull),
    .full         (_writeQueueVec_fifo_10_full),
    .error        (_writeQueueVec_fifo_10_error),
    .data_out     (_writeQueueVec_fifo_10_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_11_writeValid_T & ~(_writeQueueVec_fifo_11_empty & writeQueueVec_11_deq_ready))),
    .pop_req_n    (~(writeQueueVec_11_deq_ready & ~_writeQueueVec_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_11),
    .empty        (_writeQueueVec_fifo_11_empty),
    .almost_empty (writeQueueVec_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_11_almostFull),
    .full         (_writeQueueVec_fifo_11_full),
    .error        (_writeQueueVec_fifo_11_error),
    .data_out     (_writeQueueVec_fifo_11_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_12_writeValid_T & ~(_writeQueueVec_fifo_12_empty & writeQueueVec_12_deq_ready))),
    .pop_req_n    (~(writeQueueVec_12_deq_ready & ~_writeQueueVec_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_12),
    .empty        (_writeQueueVec_fifo_12_empty),
    .almost_empty (writeQueueVec_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_12_almostFull),
    .full         (_writeQueueVec_fifo_12_full),
    .error        (_writeQueueVec_fifo_12_error),
    .data_out     (_writeQueueVec_fifo_12_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_13_writeValid_T & ~(_writeQueueVec_fifo_13_empty & writeQueueVec_13_deq_ready))),
    .pop_req_n    (~(writeQueueVec_13_deq_ready & ~_writeQueueVec_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_13),
    .empty        (_writeQueueVec_fifo_13_empty),
    .almost_empty (writeQueueVec_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_13_almostFull),
    .full         (_writeQueueVec_fifo_13_full),
    .error        (_writeQueueVec_fifo_13_error),
    .data_out     (_writeQueueVec_fifo_13_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_14_writeValid_T & ~(_writeQueueVec_fifo_14_empty & writeQueueVec_14_deq_ready))),
    .pop_req_n    (~(writeQueueVec_14_deq_ready & ~_writeQueueVec_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_14),
    .empty        (_writeQueueVec_fifo_14_empty),
    .almost_empty (writeQueueVec_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_14_almostFull),
    .full         (_writeQueueVec_fifo_14_full),
    .error        (_writeQueueVec_fifo_14_error),
    .data_out     (_writeQueueVec_fifo_14_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_15_writeValid_T & ~(_writeQueueVec_fifo_15_empty & writeQueueVec_15_deq_ready))),
    .pop_req_n    (~(writeQueueVec_15_deq_ready & ~_writeQueueVec_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_15),
    .empty        (_writeQueueVec_fifo_15_empty),
    .almost_empty (writeQueueVec_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_15_almostFull),
    .full         (_writeQueueVec_fifo_15_full),
    .error        (_writeQueueVec_fifo_15_error),
    .data_out     (_writeQueueVec_fifo_15_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_16 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_16_writeValid_T & ~(_writeQueueVec_fifo_16_empty & writeQueueVec_16_deq_ready))),
    .pop_req_n    (~(writeQueueVec_16_deq_ready & ~_writeQueueVec_fifo_16_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_16),
    .empty        (_writeQueueVec_fifo_16_empty),
    .almost_empty (writeQueueVec_16_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_16_almostFull),
    .full         (_writeQueueVec_fifo_16_full),
    .error        (_writeQueueVec_fifo_16_error),
    .data_out     (_writeQueueVec_fifo_16_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_17 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_17_writeValid_T & ~(_writeQueueVec_fifo_17_empty & writeQueueVec_17_deq_ready))),
    .pop_req_n    (~(writeQueueVec_17_deq_ready & ~_writeQueueVec_fifo_17_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_17),
    .empty        (_writeQueueVec_fifo_17_empty),
    .almost_empty (writeQueueVec_17_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_17_almostFull),
    .full         (_writeQueueVec_fifo_17_full),
    .error        (_writeQueueVec_fifo_17_error),
    .data_out     (_writeQueueVec_fifo_17_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_18 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_18_writeValid_T & ~(_writeQueueVec_fifo_18_empty & writeQueueVec_18_deq_ready))),
    .pop_req_n    (~(writeQueueVec_18_deq_ready & ~_writeQueueVec_fifo_18_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_18),
    .empty        (_writeQueueVec_fifo_18_empty),
    .almost_empty (writeQueueVec_18_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_18_almostFull),
    .full         (_writeQueueVec_fifo_18_full),
    .error        (_writeQueueVec_fifo_18_error),
    .data_out     (_writeQueueVec_fifo_18_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_19 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_19_writeValid_T & ~(_writeQueueVec_fifo_19_empty & writeQueueVec_19_deq_ready))),
    .pop_req_n    (~(writeQueueVec_19_deq_ready & ~_writeQueueVec_fifo_19_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_19),
    .empty        (_writeQueueVec_fifo_19_empty),
    .almost_empty (writeQueueVec_19_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_19_almostFull),
    .full         (_writeQueueVec_fifo_19_full),
    .error        (_writeQueueVec_fifo_19_error),
    .data_out     (_writeQueueVec_fifo_19_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_20 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_20_writeValid_T & ~(_writeQueueVec_fifo_20_empty & writeQueueVec_20_deq_ready))),
    .pop_req_n    (~(writeQueueVec_20_deq_ready & ~_writeQueueVec_fifo_20_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_20),
    .empty        (_writeQueueVec_fifo_20_empty),
    .almost_empty (writeQueueVec_20_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_20_almostFull),
    .full         (_writeQueueVec_fifo_20_full),
    .error        (_writeQueueVec_fifo_20_error),
    .data_out     (_writeQueueVec_fifo_20_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_21 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_21_writeValid_T & ~(_writeQueueVec_fifo_21_empty & writeQueueVec_21_deq_ready))),
    .pop_req_n    (~(writeQueueVec_21_deq_ready & ~_writeQueueVec_fifo_21_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_21),
    .empty        (_writeQueueVec_fifo_21_empty),
    .almost_empty (writeQueueVec_21_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_21_almostFull),
    .full         (_writeQueueVec_fifo_21_full),
    .error        (_writeQueueVec_fifo_21_error),
    .data_out     (_writeQueueVec_fifo_21_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_22 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_22_writeValid_T & ~(_writeQueueVec_fifo_22_empty & writeQueueVec_22_deq_ready))),
    .pop_req_n    (~(writeQueueVec_22_deq_ready & ~_writeQueueVec_fifo_22_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_22),
    .empty        (_writeQueueVec_fifo_22_empty),
    .almost_empty (writeQueueVec_22_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_22_almostFull),
    .full         (_writeQueueVec_fifo_22_full),
    .error        (_writeQueueVec_fifo_22_error),
    .data_out     (_writeQueueVec_fifo_22_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_23 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_23_writeValid_T & ~(_writeQueueVec_fifo_23_empty & writeQueueVec_23_deq_ready))),
    .pop_req_n    (~(writeQueueVec_23_deq_ready & ~_writeQueueVec_fifo_23_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_23),
    .empty        (_writeQueueVec_fifo_23_empty),
    .almost_empty (writeQueueVec_23_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_23_almostFull),
    .full         (_writeQueueVec_fifo_23_full),
    .error        (_writeQueueVec_fifo_23_error),
    .data_out     (_writeQueueVec_fifo_23_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_24 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_24_writeValid_T & ~(_writeQueueVec_fifo_24_empty & writeQueueVec_24_deq_ready))),
    .pop_req_n    (~(writeQueueVec_24_deq_ready & ~_writeQueueVec_fifo_24_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_24),
    .empty        (_writeQueueVec_fifo_24_empty),
    .almost_empty (writeQueueVec_24_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_24_almostFull),
    .full         (_writeQueueVec_fifo_24_full),
    .error        (_writeQueueVec_fifo_24_error),
    .data_out     (_writeQueueVec_fifo_24_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_25 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_25_writeValid_T & ~(_writeQueueVec_fifo_25_empty & writeQueueVec_25_deq_ready))),
    .pop_req_n    (~(writeQueueVec_25_deq_ready & ~_writeQueueVec_fifo_25_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_25),
    .empty        (_writeQueueVec_fifo_25_empty),
    .almost_empty (writeQueueVec_25_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_25_almostFull),
    .full         (_writeQueueVec_fifo_25_full),
    .error        (_writeQueueVec_fifo_25_error),
    .data_out     (_writeQueueVec_fifo_25_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_26 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_26_writeValid_T & ~(_writeQueueVec_fifo_26_empty & writeQueueVec_26_deq_ready))),
    .pop_req_n    (~(writeQueueVec_26_deq_ready & ~_writeQueueVec_fifo_26_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_26),
    .empty        (_writeQueueVec_fifo_26_empty),
    .almost_empty (writeQueueVec_26_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_26_almostFull),
    .full         (_writeQueueVec_fifo_26_full),
    .error        (_writeQueueVec_fifo_26_error),
    .data_out     (_writeQueueVec_fifo_26_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_27 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_27_writeValid_T & ~(_writeQueueVec_fifo_27_empty & writeQueueVec_27_deq_ready))),
    .pop_req_n    (~(writeQueueVec_27_deq_ready & ~_writeQueueVec_fifo_27_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_27),
    .empty        (_writeQueueVec_fifo_27_empty),
    .almost_empty (writeQueueVec_27_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_27_almostFull),
    .full         (_writeQueueVec_fifo_27_full),
    .error        (_writeQueueVec_fifo_27_error),
    .data_out     (_writeQueueVec_fifo_27_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_28 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_28_writeValid_T & ~(_writeQueueVec_fifo_28_empty & writeQueueVec_28_deq_ready))),
    .pop_req_n    (~(writeQueueVec_28_deq_ready & ~_writeQueueVec_fifo_28_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_28),
    .empty        (_writeQueueVec_fifo_28_empty),
    .almost_empty (writeQueueVec_28_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_28_almostFull),
    .full         (_writeQueueVec_fifo_28_full),
    .error        (_writeQueueVec_fifo_28_error),
    .data_out     (_writeQueueVec_fifo_28_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_29 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_29_writeValid_T & ~(_writeQueueVec_fifo_29_empty & writeQueueVec_29_deq_ready))),
    .pop_req_n    (~(writeQueueVec_29_deq_ready & ~_writeQueueVec_fifo_29_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_29),
    .empty        (_writeQueueVec_fifo_29_empty),
    .almost_empty (writeQueueVec_29_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_29_almostFull),
    .full         (_writeQueueVec_fifo_29_full),
    .error        (_writeQueueVec_fifo_29_error),
    .data_out     (_writeQueueVec_fifo_29_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_30 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_30_writeValid_T & ~(_writeQueueVec_fifo_30_empty & writeQueueVec_30_deq_ready))),
    .pop_req_n    (~(writeQueueVec_30_deq_ready & ~_writeQueueVec_fifo_30_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_30),
    .empty        (_writeQueueVec_fifo_30_empty),
    .almost_empty (writeQueueVec_30_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_30_almostFull),
    .full         (_writeQueueVec_fifo_30_full),
    .error        (_writeQueueVec_fifo_30_error),
    .data_out     (_writeQueueVec_fifo_30_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(77)
  ) writeQueueVec_fifo_31 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_31_writeValid_T & ~(_writeQueueVec_fifo_31_empty & writeQueueVec_31_deq_ready))),
    .pop_req_n    (~(writeQueueVec_31_deq_ready & ~_writeQueueVec_fifo_31_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_31),
    .empty        (_writeQueueVec_fifo_31_empty),
    .almost_empty (writeQueueVec_31_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_31_almostFull),
    .full         (_writeQueueVec_fifo_31_full),
    .error        (_writeQueueVec_fifo_31_error),
    .data_out     (_writeQueueVec_fifo_31_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitTargetQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitTargetQueue_enq_ready & otherUnitTargetQueue_enq_valid)),
    .pop_req_n    (~(otherUnitTargetQueue_deq_ready & ~_otherUnitTargetQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitTargetQueue_enq_bits),
    .empty        (_otherUnitTargetQueue_fifo_empty),
    .almost_empty (otherUnitTargetQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitTargetQueue_almostFull),
    .full         (_otherUnitTargetQueue_fifo_full),
    .error        (_otherUnitTargetQueue_fifo_error),
    .data_out     (otherUnitTargetQueue_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_0_enq_ready & otherUnitDataQueueVec_0_enq_valid & ~(_otherUnitDataQueueVec_fifo_empty & otherUnitDataQueueVec_0_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_0_deq_ready & ~_otherUnitDataQueueVec_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_0_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_empty),
    .almost_empty (otherUnitDataQueueVec_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_0_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_full),
    .error        (_otherUnitDataQueueVec_fifo_error),
    .data_out     (_otherUnitDataQueueVec_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_1_enq_ready & otherUnitDataQueueVec_1_enq_valid & ~(_otherUnitDataQueueVec_fifo_1_empty & otherUnitDataQueueVec_1_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_1_deq_ready & ~_otherUnitDataQueueVec_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_1_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_1_empty),
    .almost_empty (otherUnitDataQueueVec_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_1_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_1_full),
    .error        (_otherUnitDataQueueVec_fifo_1_error),
    .data_out     (_otherUnitDataQueueVec_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_2_enq_ready & otherUnitDataQueueVec_2_enq_valid & ~(_otherUnitDataQueueVec_fifo_2_empty & otherUnitDataQueueVec_2_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_2_deq_ready & ~_otherUnitDataQueueVec_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_2_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_2_empty),
    .almost_empty (otherUnitDataQueueVec_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_2_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_2_full),
    .error        (_otherUnitDataQueueVec_fifo_2_error),
    .data_out     (_otherUnitDataQueueVec_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_3_enq_ready & otherUnitDataQueueVec_3_enq_valid & ~(_otherUnitDataQueueVec_fifo_3_empty & otherUnitDataQueueVec_3_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_3_deq_ready & ~_otherUnitDataQueueVec_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_3_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_3_empty),
    .almost_empty (otherUnitDataQueueVec_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_3_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_3_full),
    .error        (_otherUnitDataQueueVec_fifo_3_error),
    .data_out     (_otherUnitDataQueueVec_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_4_enq_ready & otherUnitDataQueueVec_4_enq_valid & ~(_otherUnitDataQueueVec_fifo_4_empty & otherUnitDataQueueVec_4_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_4_deq_ready & ~_otherUnitDataQueueVec_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_4_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_4_empty),
    .almost_empty (otherUnitDataQueueVec_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_4_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_4_full),
    .error        (_otherUnitDataQueueVec_fifo_4_error),
    .data_out     (_otherUnitDataQueueVec_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_5_enq_ready & otherUnitDataQueueVec_5_enq_valid & ~(_otherUnitDataQueueVec_fifo_5_empty & otherUnitDataQueueVec_5_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_5_deq_ready & ~_otherUnitDataQueueVec_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_5_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_5_empty),
    .almost_empty (otherUnitDataQueueVec_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_5_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_5_full),
    .error        (_otherUnitDataQueueVec_fifo_5_error),
    .data_out     (_otherUnitDataQueueVec_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_6_enq_ready & otherUnitDataQueueVec_6_enq_valid & ~(_otherUnitDataQueueVec_fifo_6_empty & otherUnitDataQueueVec_6_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_6_deq_ready & ~_otherUnitDataQueueVec_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_6_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_6_empty),
    .almost_empty (otherUnitDataQueueVec_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_6_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_6_full),
    .error        (_otherUnitDataQueueVec_fifo_6_error),
    .data_out     (_otherUnitDataQueueVec_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_7_enq_ready & otherUnitDataQueueVec_7_enq_valid & ~(_otherUnitDataQueueVec_fifo_7_empty & otherUnitDataQueueVec_7_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_7_deq_ready & ~_otherUnitDataQueueVec_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_7_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_7_empty),
    .almost_empty (otherUnitDataQueueVec_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_7_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_7_full),
    .error        (_otherUnitDataQueueVec_fifo_7_error),
    .data_out     (_otherUnitDataQueueVec_fifo_7_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_8_enq_ready & otherUnitDataQueueVec_8_enq_valid & ~(_otherUnitDataQueueVec_fifo_8_empty & otherUnitDataQueueVec_8_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_8_deq_ready & ~_otherUnitDataQueueVec_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_8_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_8_empty),
    .almost_empty (otherUnitDataQueueVec_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_8_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_8_full),
    .error        (_otherUnitDataQueueVec_fifo_8_error),
    .data_out     (_otherUnitDataQueueVec_fifo_8_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_9_enq_ready & otherUnitDataQueueVec_9_enq_valid & ~(_otherUnitDataQueueVec_fifo_9_empty & otherUnitDataQueueVec_9_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_9_deq_ready & ~_otherUnitDataQueueVec_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_9_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_9_empty),
    .almost_empty (otherUnitDataQueueVec_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_9_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_9_full),
    .error        (_otherUnitDataQueueVec_fifo_9_error),
    .data_out     (_otherUnitDataQueueVec_fifo_9_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_10_enq_ready & otherUnitDataQueueVec_10_enq_valid & ~(_otherUnitDataQueueVec_fifo_10_empty & otherUnitDataQueueVec_10_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_10_deq_ready & ~_otherUnitDataQueueVec_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_10_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_10_empty),
    .almost_empty (otherUnitDataQueueVec_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_10_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_10_full),
    .error        (_otherUnitDataQueueVec_fifo_10_error),
    .data_out     (_otherUnitDataQueueVec_fifo_10_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_11_enq_ready & otherUnitDataQueueVec_11_enq_valid & ~(_otherUnitDataQueueVec_fifo_11_empty & otherUnitDataQueueVec_11_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_11_deq_ready & ~_otherUnitDataQueueVec_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_11_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_11_empty),
    .almost_empty (otherUnitDataQueueVec_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_11_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_11_full),
    .error        (_otherUnitDataQueueVec_fifo_11_error),
    .data_out     (_otherUnitDataQueueVec_fifo_11_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_12_enq_ready & otherUnitDataQueueVec_12_enq_valid & ~(_otherUnitDataQueueVec_fifo_12_empty & otherUnitDataQueueVec_12_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_12_deq_ready & ~_otherUnitDataQueueVec_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_12_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_12_empty),
    .almost_empty (otherUnitDataQueueVec_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_12_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_12_full),
    .error        (_otherUnitDataQueueVec_fifo_12_error),
    .data_out     (_otherUnitDataQueueVec_fifo_12_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_13_enq_ready & otherUnitDataQueueVec_13_enq_valid & ~(_otherUnitDataQueueVec_fifo_13_empty & otherUnitDataQueueVec_13_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_13_deq_ready & ~_otherUnitDataQueueVec_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_13_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_13_empty),
    .almost_empty (otherUnitDataQueueVec_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_13_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_13_full),
    .error        (_otherUnitDataQueueVec_fifo_13_error),
    .data_out     (_otherUnitDataQueueVec_fifo_13_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_14_enq_ready & otherUnitDataQueueVec_14_enq_valid & ~(_otherUnitDataQueueVec_fifo_14_empty & otherUnitDataQueueVec_14_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_14_deq_ready & ~_otherUnitDataQueueVec_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_14_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_14_empty),
    .almost_empty (otherUnitDataQueueVec_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_14_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_14_full),
    .error        (_otherUnitDataQueueVec_fifo_14_error),
    .data_out     (_otherUnitDataQueueVec_fifo_14_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_15_enq_ready & otherUnitDataQueueVec_15_enq_valid & ~(_otherUnitDataQueueVec_fifo_15_empty & otherUnitDataQueueVec_15_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_15_deq_ready & ~_otherUnitDataQueueVec_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_15_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_15_empty),
    .almost_empty (otherUnitDataQueueVec_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_15_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_15_full),
    .error        (_otherUnitDataQueueVec_fifo_15_error),
    .data_out     (_otherUnitDataQueueVec_fifo_15_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_16 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_16_enq_ready & otherUnitDataQueueVec_16_enq_valid & ~(_otherUnitDataQueueVec_fifo_16_empty & otherUnitDataQueueVec_16_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_16_deq_ready & ~_otherUnitDataQueueVec_fifo_16_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_16_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_16_empty),
    .almost_empty (otherUnitDataQueueVec_16_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_16_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_16_full),
    .error        (_otherUnitDataQueueVec_fifo_16_error),
    .data_out     (_otherUnitDataQueueVec_fifo_16_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_17 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_17_enq_ready & otherUnitDataQueueVec_17_enq_valid & ~(_otherUnitDataQueueVec_fifo_17_empty & otherUnitDataQueueVec_17_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_17_deq_ready & ~_otherUnitDataQueueVec_fifo_17_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_17_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_17_empty),
    .almost_empty (otherUnitDataQueueVec_17_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_17_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_17_full),
    .error        (_otherUnitDataQueueVec_fifo_17_error),
    .data_out     (_otherUnitDataQueueVec_fifo_17_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_18 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_18_enq_ready & otherUnitDataQueueVec_18_enq_valid & ~(_otherUnitDataQueueVec_fifo_18_empty & otherUnitDataQueueVec_18_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_18_deq_ready & ~_otherUnitDataQueueVec_fifo_18_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_18_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_18_empty),
    .almost_empty (otherUnitDataQueueVec_18_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_18_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_18_full),
    .error        (_otherUnitDataQueueVec_fifo_18_error),
    .data_out     (_otherUnitDataQueueVec_fifo_18_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_19 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_19_enq_ready & otherUnitDataQueueVec_19_enq_valid & ~(_otherUnitDataQueueVec_fifo_19_empty & otherUnitDataQueueVec_19_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_19_deq_ready & ~_otherUnitDataQueueVec_fifo_19_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_19_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_19_empty),
    .almost_empty (otherUnitDataQueueVec_19_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_19_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_19_full),
    .error        (_otherUnitDataQueueVec_fifo_19_error),
    .data_out     (_otherUnitDataQueueVec_fifo_19_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_20 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_20_enq_ready & otherUnitDataQueueVec_20_enq_valid & ~(_otherUnitDataQueueVec_fifo_20_empty & otherUnitDataQueueVec_20_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_20_deq_ready & ~_otherUnitDataQueueVec_fifo_20_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_20_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_20_empty),
    .almost_empty (otherUnitDataQueueVec_20_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_20_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_20_full),
    .error        (_otherUnitDataQueueVec_fifo_20_error),
    .data_out     (_otherUnitDataQueueVec_fifo_20_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_21 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_21_enq_ready & otherUnitDataQueueVec_21_enq_valid & ~(_otherUnitDataQueueVec_fifo_21_empty & otherUnitDataQueueVec_21_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_21_deq_ready & ~_otherUnitDataQueueVec_fifo_21_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_21_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_21_empty),
    .almost_empty (otherUnitDataQueueVec_21_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_21_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_21_full),
    .error        (_otherUnitDataQueueVec_fifo_21_error),
    .data_out     (_otherUnitDataQueueVec_fifo_21_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_22 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_22_enq_ready & otherUnitDataQueueVec_22_enq_valid & ~(_otherUnitDataQueueVec_fifo_22_empty & otherUnitDataQueueVec_22_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_22_deq_ready & ~_otherUnitDataQueueVec_fifo_22_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_22_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_22_empty),
    .almost_empty (otherUnitDataQueueVec_22_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_22_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_22_full),
    .error        (_otherUnitDataQueueVec_fifo_22_error),
    .data_out     (_otherUnitDataQueueVec_fifo_22_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_23 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_23_enq_ready & otherUnitDataQueueVec_23_enq_valid & ~(_otherUnitDataQueueVec_fifo_23_empty & otherUnitDataQueueVec_23_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_23_deq_ready & ~_otherUnitDataQueueVec_fifo_23_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_23_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_23_empty),
    .almost_empty (otherUnitDataQueueVec_23_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_23_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_23_full),
    .error        (_otherUnitDataQueueVec_fifo_23_error),
    .data_out     (_otherUnitDataQueueVec_fifo_23_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_24 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_24_enq_ready & otherUnitDataQueueVec_24_enq_valid & ~(_otherUnitDataQueueVec_fifo_24_empty & otherUnitDataQueueVec_24_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_24_deq_ready & ~_otherUnitDataQueueVec_fifo_24_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_24_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_24_empty),
    .almost_empty (otherUnitDataQueueVec_24_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_24_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_24_full),
    .error        (_otherUnitDataQueueVec_fifo_24_error),
    .data_out     (_otherUnitDataQueueVec_fifo_24_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_25 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_25_enq_ready & otherUnitDataQueueVec_25_enq_valid & ~(_otherUnitDataQueueVec_fifo_25_empty & otherUnitDataQueueVec_25_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_25_deq_ready & ~_otherUnitDataQueueVec_fifo_25_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_25_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_25_empty),
    .almost_empty (otherUnitDataQueueVec_25_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_25_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_25_full),
    .error        (_otherUnitDataQueueVec_fifo_25_error),
    .data_out     (_otherUnitDataQueueVec_fifo_25_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_26 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_26_enq_ready & otherUnitDataQueueVec_26_enq_valid & ~(_otherUnitDataQueueVec_fifo_26_empty & otherUnitDataQueueVec_26_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_26_deq_ready & ~_otherUnitDataQueueVec_fifo_26_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_26_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_26_empty),
    .almost_empty (otherUnitDataQueueVec_26_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_26_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_26_full),
    .error        (_otherUnitDataQueueVec_fifo_26_error),
    .data_out     (_otherUnitDataQueueVec_fifo_26_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_27 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_27_enq_ready & otherUnitDataQueueVec_27_enq_valid & ~(_otherUnitDataQueueVec_fifo_27_empty & otherUnitDataQueueVec_27_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_27_deq_ready & ~_otherUnitDataQueueVec_fifo_27_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_27_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_27_empty),
    .almost_empty (otherUnitDataQueueVec_27_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_27_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_27_full),
    .error        (_otherUnitDataQueueVec_fifo_27_error),
    .data_out     (_otherUnitDataQueueVec_fifo_27_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_28 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_28_enq_ready & otherUnitDataQueueVec_28_enq_valid & ~(_otherUnitDataQueueVec_fifo_28_empty & otherUnitDataQueueVec_28_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_28_deq_ready & ~_otherUnitDataQueueVec_fifo_28_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_28_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_28_empty),
    .almost_empty (otherUnitDataQueueVec_28_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_28_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_28_full),
    .error        (_otherUnitDataQueueVec_fifo_28_error),
    .data_out     (_otherUnitDataQueueVec_fifo_28_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_29 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_29_enq_ready & otherUnitDataQueueVec_29_enq_valid & ~(_otherUnitDataQueueVec_fifo_29_empty & otherUnitDataQueueVec_29_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_29_deq_ready & ~_otherUnitDataQueueVec_fifo_29_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_29_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_29_empty),
    .almost_empty (otherUnitDataQueueVec_29_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_29_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_29_full),
    .error        (_otherUnitDataQueueVec_fifo_29_error),
    .data_out     (_otherUnitDataQueueVec_fifo_29_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_30 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_30_enq_ready & otherUnitDataQueueVec_30_enq_valid & ~(_otherUnitDataQueueVec_fifo_30_empty & otherUnitDataQueueVec_30_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_30_deq_ready & ~_otherUnitDataQueueVec_fifo_30_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_30_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_30_empty),
    .almost_empty (otherUnitDataQueueVec_30_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_30_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_30_full),
    .error        (_otherUnitDataQueueVec_fifo_30_error),
    .data_out     (_otherUnitDataQueueVec_fifo_30_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_31 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_31_enq_ready & otherUnitDataQueueVec_31_enq_valid & ~(_otherUnitDataQueueVec_fifo_31_empty & otherUnitDataQueueVec_31_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_31_deq_ready & ~_otherUnitDataQueueVec_fifo_31_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_31_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_31_empty),
    .almost_empty (otherUnitDataQueueVec_31_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_31_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_31_full),
    .error        (_otherUnitDataQueueVec_fifo_31_error),
    .data_out     (_otherUnitDataQueueVec_fifo_31_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_enq_ready & writeIndexQueue_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_deq_ready & ~_writeIndexQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_enq_bits),
    .empty        (_writeIndexQueue_fifo_empty),
    .almost_empty (writeIndexQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_almostFull),
    .full         (_writeIndexQueue_fifo_full),
    .error        (_writeIndexQueue_fifo_error),
    .data_out     (writeIndexQueue_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_1_enq_ready & writeIndexQueue_1_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_1_deq_ready & ~_writeIndexQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_1_enq_bits),
    .empty        (_writeIndexQueue_fifo_1_empty),
    .almost_empty (writeIndexQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_1_almostFull),
    .full         (_writeIndexQueue_fifo_1_full),
    .error        (_writeIndexQueue_fifo_1_error),
    .data_out     (writeIndexQueue_1_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_2_enq_ready & writeIndexQueue_2_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_2_deq_ready & ~_writeIndexQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_2_enq_bits),
    .empty        (_writeIndexQueue_fifo_2_empty),
    .almost_empty (writeIndexQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_2_almostFull),
    .full         (_writeIndexQueue_fifo_2_full),
    .error        (_writeIndexQueue_fifo_2_error),
    .data_out     (writeIndexQueue_2_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_3_enq_ready & writeIndexQueue_3_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_3_deq_ready & ~_writeIndexQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_3_enq_bits),
    .empty        (_writeIndexQueue_fifo_3_empty),
    .almost_empty (writeIndexQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_3_almostFull),
    .full         (_writeIndexQueue_fifo_3_full),
    .error        (_writeIndexQueue_fifo_3_error),
    .data_out     (writeIndexQueue_3_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_4_enq_ready & writeIndexQueue_4_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_4_deq_ready & ~_writeIndexQueue_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_4_enq_bits),
    .empty        (_writeIndexQueue_fifo_4_empty),
    .almost_empty (writeIndexQueue_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_4_almostFull),
    .full         (_writeIndexQueue_fifo_4_full),
    .error        (_writeIndexQueue_fifo_4_error),
    .data_out     (writeIndexQueue_4_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_5_enq_ready & writeIndexQueue_5_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_5_deq_ready & ~_writeIndexQueue_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_5_enq_bits),
    .empty        (_writeIndexQueue_fifo_5_empty),
    .almost_empty (writeIndexQueue_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_5_almostFull),
    .full         (_writeIndexQueue_fifo_5_full),
    .error        (_writeIndexQueue_fifo_5_error),
    .data_out     (writeIndexQueue_5_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_6_enq_ready & writeIndexQueue_6_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_6_deq_ready & ~_writeIndexQueue_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_6_enq_bits),
    .empty        (_writeIndexQueue_fifo_6_empty),
    .almost_empty (writeIndexQueue_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_6_almostFull),
    .full         (_writeIndexQueue_fifo_6_full),
    .error        (_writeIndexQueue_fifo_6_error),
    .data_out     (writeIndexQueue_6_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_7_enq_ready & writeIndexQueue_7_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_7_deq_ready & ~_writeIndexQueue_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_7_enq_bits),
    .empty        (_writeIndexQueue_fifo_7_empty),
    .almost_empty (writeIndexQueue_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_7_almostFull),
    .full         (_writeIndexQueue_fifo_7_full),
    .error        (_writeIndexQueue_fifo_7_error),
    .data_out     (writeIndexQueue_7_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_8_enq_ready & writeIndexQueue_8_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_8_deq_ready & ~_writeIndexQueue_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_8_enq_bits),
    .empty        (_writeIndexQueue_fifo_8_empty),
    .almost_empty (writeIndexQueue_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_8_almostFull),
    .full         (_writeIndexQueue_fifo_8_full),
    .error        (_writeIndexQueue_fifo_8_error),
    .data_out     (writeIndexQueue_8_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_9_enq_ready & writeIndexQueue_9_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_9_deq_ready & ~_writeIndexQueue_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_9_enq_bits),
    .empty        (_writeIndexQueue_fifo_9_empty),
    .almost_empty (writeIndexQueue_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_9_almostFull),
    .full         (_writeIndexQueue_fifo_9_full),
    .error        (_writeIndexQueue_fifo_9_error),
    .data_out     (writeIndexQueue_9_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_10_enq_ready & writeIndexQueue_10_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_10_deq_ready & ~_writeIndexQueue_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_10_enq_bits),
    .empty        (_writeIndexQueue_fifo_10_empty),
    .almost_empty (writeIndexQueue_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_10_almostFull),
    .full         (_writeIndexQueue_fifo_10_full),
    .error        (_writeIndexQueue_fifo_10_error),
    .data_out     (writeIndexQueue_10_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_11_enq_ready & writeIndexQueue_11_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_11_deq_ready & ~_writeIndexQueue_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_11_enq_bits),
    .empty        (_writeIndexQueue_fifo_11_empty),
    .almost_empty (writeIndexQueue_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_11_almostFull),
    .full         (_writeIndexQueue_fifo_11_full),
    .error        (_writeIndexQueue_fifo_11_error),
    .data_out     (writeIndexQueue_11_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_12_enq_ready & writeIndexQueue_12_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_12_deq_ready & ~_writeIndexQueue_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_12_enq_bits),
    .empty        (_writeIndexQueue_fifo_12_empty),
    .almost_empty (writeIndexQueue_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_12_almostFull),
    .full         (_writeIndexQueue_fifo_12_full),
    .error        (_writeIndexQueue_fifo_12_error),
    .data_out     (writeIndexQueue_12_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_13_enq_ready & writeIndexQueue_13_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_13_deq_ready & ~_writeIndexQueue_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_13_enq_bits),
    .empty        (_writeIndexQueue_fifo_13_empty),
    .almost_empty (writeIndexQueue_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_13_almostFull),
    .full         (_writeIndexQueue_fifo_13_full),
    .error        (_writeIndexQueue_fifo_13_error),
    .data_out     (writeIndexQueue_13_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_14_enq_ready & writeIndexQueue_14_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_14_deq_ready & ~_writeIndexQueue_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_14_enq_bits),
    .empty        (_writeIndexQueue_fifo_14_empty),
    .almost_empty (writeIndexQueue_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_14_almostFull),
    .full         (_writeIndexQueue_fifo_14_full),
    .error        (_writeIndexQueue_fifo_14_error),
    .data_out     (writeIndexQueue_14_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_15_enq_ready & writeIndexQueue_15_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_15_deq_ready & ~_writeIndexQueue_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_15_enq_bits),
    .empty        (_writeIndexQueue_fifo_15_empty),
    .almost_empty (writeIndexQueue_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_15_almostFull),
    .full         (_writeIndexQueue_fifo_15_full),
    .error        (_writeIndexQueue_fifo_15_error),
    .data_out     (writeIndexQueue_15_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_16 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_16_enq_ready & writeIndexQueue_16_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_16_deq_ready & ~_writeIndexQueue_fifo_16_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_16_enq_bits),
    .empty        (_writeIndexQueue_fifo_16_empty),
    .almost_empty (writeIndexQueue_16_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_16_almostFull),
    .full         (_writeIndexQueue_fifo_16_full),
    .error        (_writeIndexQueue_fifo_16_error),
    .data_out     (writeIndexQueue_16_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_17 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_17_enq_ready & writeIndexQueue_17_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_17_deq_ready & ~_writeIndexQueue_fifo_17_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_17_enq_bits),
    .empty        (_writeIndexQueue_fifo_17_empty),
    .almost_empty (writeIndexQueue_17_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_17_almostFull),
    .full         (_writeIndexQueue_fifo_17_full),
    .error        (_writeIndexQueue_fifo_17_error),
    .data_out     (writeIndexQueue_17_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_18 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_18_enq_ready & writeIndexQueue_18_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_18_deq_ready & ~_writeIndexQueue_fifo_18_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_18_enq_bits),
    .empty        (_writeIndexQueue_fifo_18_empty),
    .almost_empty (writeIndexQueue_18_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_18_almostFull),
    .full         (_writeIndexQueue_fifo_18_full),
    .error        (_writeIndexQueue_fifo_18_error),
    .data_out     (writeIndexQueue_18_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_19 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_19_enq_ready & writeIndexQueue_19_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_19_deq_ready & ~_writeIndexQueue_fifo_19_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_19_enq_bits),
    .empty        (_writeIndexQueue_fifo_19_empty),
    .almost_empty (writeIndexQueue_19_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_19_almostFull),
    .full         (_writeIndexQueue_fifo_19_full),
    .error        (_writeIndexQueue_fifo_19_error),
    .data_out     (writeIndexQueue_19_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_20 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_20_enq_ready & writeIndexQueue_20_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_20_deq_ready & ~_writeIndexQueue_fifo_20_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_20_enq_bits),
    .empty        (_writeIndexQueue_fifo_20_empty),
    .almost_empty (writeIndexQueue_20_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_20_almostFull),
    .full         (_writeIndexQueue_fifo_20_full),
    .error        (_writeIndexQueue_fifo_20_error),
    .data_out     (writeIndexQueue_20_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_21 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_21_enq_ready & writeIndexQueue_21_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_21_deq_ready & ~_writeIndexQueue_fifo_21_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_21_enq_bits),
    .empty        (_writeIndexQueue_fifo_21_empty),
    .almost_empty (writeIndexQueue_21_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_21_almostFull),
    .full         (_writeIndexQueue_fifo_21_full),
    .error        (_writeIndexQueue_fifo_21_error),
    .data_out     (writeIndexQueue_21_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_22 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_22_enq_ready & writeIndexQueue_22_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_22_deq_ready & ~_writeIndexQueue_fifo_22_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_22_enq_bits),
    .empty        (_writeIndexQueue_fifo_22_empty),
    .almost_empty (writeIndexQueue_22_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_22_almostFull),
    .full         (_writeIndexQueue_fifo_22_full),
    .error        (_writeIndexQueue_fifo_22_error),
    .data_out     (writeIndexQueue_22_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_23 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_23_enq_ready & writeIndexQueue_23_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_23_deq_ready & ~_writeIndexQueue_fifo_23_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_23_enq_bits),
    .empty        (_writeIndexQueue_fifo_23_empty),
    .almost_empty (writeIndexQueue_23_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_23_almostFull),
    .full         (_writeIndexQueue_fifo_23_full),
    .error        (_writeIndexQueue_fifo_23_error),
    .data_out     (writeIndexQueue_23_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_24 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_24_enq_ready & writeIndexQueue_24_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_24_deq_ready & ~_writeIndexQueue_fifo_24_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_24_enq_bits),
    .empty        (_writeIndexQueue_fifo_24_empty),
    .almost_empty (writeIndexQueue_24_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_24_almostFull),
    .full         (_writeIndexQueue_fifo_24_full),
    .error        (_writeIndexQueue_fifo_24_error),
    .data_out     (writeIndexQueue_24_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_25 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_25_enq_ready & writeIndexQueue_25_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_25_deq_ready & ~_writeIndexQueue_fifo_25_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_25_enq_bits),
    .empty        (_writeIndexQueue_fifo_25_empty),
    .almost_empty (writeIndexQueue_25_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_25_almostFull),
    .full         (_writeIndexQueue_fifo_25_full),
    .error        (_writeIndexQueue_fifo_25_error),
    .data_out     (writeIndexQueue_25_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_26 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_26_enq_ready & writeIndexQueue_26_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_26_deq_ready & ~_writeIndexQueue_fifo_26_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_26_enq_bits),
    .empty        (_writeIndexQueue_fifo_26_empty),
    .almost_empty (writeIndexQueue_26_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_26_almostFull),
    .full         (_writeIndexQueue_fifo_26_full),
    .error        (_writeIndexQueue_fifo_26_error),
    .data_out     (writeIndexQueue_26_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_27 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_27_enq_ready & writeIndexQueue_27_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_27_deq_ready & ~_writeIndexQueue_fifo_27_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_27_enq_bits),
    .empty        (_writeIndexQueue_fifo_27_empty),
    .almost_empty (writeIndexQueue_27_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_27_almostFull),
    .full         (_writeIndexQueue_fifo_27_full),
    .error        (_writeIndexQueue_fifo_27_error),
    .data_out     (writeIndexQueue_27_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_28 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_28_enq_ready & writeIndexQueue_28_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_28_deq_ready & ~_writeIndexQueue_fifo_28_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_28_enq_bits),
    .empty        (_writeIndexQueue_fifo_28_empty),
    .almost_empty (writeIndexQueue_28_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_28_almostFull),
    .full         (_writeIndexQueue_fifo_28_full),
    .error        (_writeIndexQueue_fifo_28_error),
    .data_out     (writeIndexQueue_28_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_29 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_29_enq_ready & writeIndexQueue_29_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_29_deq_ready & ~_writeIndexQueue_fifo_29_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_29_enq_bits),
    .empty        (_writeIndexQueue_fifo_29_empty),
    .almost_empty (writeIndexQueue_29_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_29_almostFull),
    .full         (_writeIndexQueue_fifo_29_full),
    .error        (_writeIndexQueue_fifo_29_error),
    .data_out     (writeIndexQueue_29_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_30 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_30_enq_ready & writeIndexQueue_30_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_30_deq_ready & ~_writeIndexQueue_fifo_30_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_30_enq_bits),
    .empty        (_writeIndexQueue_fifo_30_empty),
    .almost_empty (writeIndexQueue_30_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_30_almostFull),
    .full         (_writeIndexQueue_fifo_30_full),
    .error        (_writeIndexQueue_fifo_30_error),
    .data_out     (writeIndexQueue_30_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_31 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_31_enq_ready & writeIndexQueue_31_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_31_deq_ready & ~_writeIndexQueue_fifo_31_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_31_enq_bits),
    .empty        (_writeIndexQueue_fifo_31_empty),
    .almost_empty (writeIndexQueue_31_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_31_almostFull),
    .full         (_writeIndexQueue_fifo_31_full),
    .error        (_writeIndexQueue_fifo_31_error),
    .data_out     (writeIndexQueue_31_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(4)
  ) sourceQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sourceQueue_enq_ready & sourceQueue_enq_valid)),
    .pop_req_n    (~(sourceQueue_deq_ready & ~_sourceQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (sourceQueue_enq_bits),
    .empty        (_sourceQueue_fifo_empty),
    .almost_empty (sourceQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sourceQueue_almostFull),
    .full         (_sourceQueue_fifo_full),
    .error        (_sourceQueue_fifo_error),
    .data_out     (sourceQueue_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(2),
    .err_mode(2),
    .rst_mode(3),
    .width(1188)
  ) dataQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(dataQueue_enq_ready & dataQueue_enq_valid)),
    .pop_req_n    (~(dataQueue_deq_ready & ~_dataQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (dataQueue_dataIn),
    .empty        (_dataQueue_fifo_empty),
    .almost_empty (dataQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (dataQueue_almostFull),
    .full         (_dataQueue_fifo_full),
    .error        (_dataQueue_fifo_error),
    .data_out     (_dataQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(10)
  ) simpleSourceQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(simpleSourceQueue_enq_ready & simpleSourceQueue_enq_valid)),
    .pop_req_n    (~(simpleSourceQueue_deq_ready & ~_simpleSourceQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (simpleSourceQueue_enq_bits),
    .empty        (_simpleSourceQueue_fifo_empty),
    .almost_empty (simpleSourceQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (simpleSourceQueue_almostFull),
    .full         (_simpleSourceQueue_fifo_full),
    .error        (_simpleSourceQueue_fifo_error),
    .data_out     (simpleSourceQueue_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(2),
    .err_mode(2),
    .rst_mode(3),
    .width(78)
  ) simpleDataQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(simpleDataQueue_enq_ready & simpleDataQueue_enq_valid)),
    .pop_req_n    (~(simpleDataQueue_deq_ready & ~_simpleDataQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (simpleDataQueue_dataIn),
    .empty        (_simpleDataQueue_fifo_empty),
    .almost_empty (simpleDataQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (simpleDataQueue_almostFull),
    .full         (_simpleDataQueue_fifo_full),
    .error        (_simpleDataQueue_fifo_error),
    .data_out     (_simpleDataQueue_fifo_data_out)
  );
  assign request_ready = request_ready_0;
  assign axi4Port_aw_valid = axi4Port_aw_valid_0;
  assign axi4Port_aw_bits_id = axi4Port_aw_bits_id_0;
  assign axi4Port_aw_bits_addr = axi4Port_aw_bits_addr_0;
  assign axi4Port_w_valid = axi4Port_w_valid_0;
  assign axi4Port_w_bits_data = axi4Port_w_bits_data_0;
  assign axi4Port_w_bits_strb = axi4Port_w_bits_strb_0;
  assign axi4Port_ar_valid = axi4Port_ar_valid_0;
  assign axi4Port_ar_bits_addr = axi4Port_ar_bits_addr_0;
  assign axi4Port_r_ready = axi4Port_r_ready_0;
  assign simpleAccessPorts_aw_valid = simpleAccessPorts_aw_valid_0;
  assign simpleAccessPorts_aw_bits_id = simpleAccessPorts_aw_bits_id_0;
  assign simpleAccessPorts_aw_bits_addr = simpleAccessPorts_aw_bits_addr_0;
  assign simpleAccessPorts_aw_bits_size = simpleAccessPorts_aw_bits_size_0;
  assign simpleAccessPorts_w_valid = simpleAccessPorts_w_valid_0;
  assign simpleAccessPorts_w_bits_data = simpleAccessPorts_w_bits_data_0;
  assign simpleAccessPorts_w_bits_strb = simpleAccessPorts_w_bits_strb_0;
  assign simpleAccessPorts_ar_valid = simpleAccessPorts_ar_valid_0;
  assign simpleAccessPorts_ar_bits_addr = simpleAccessPorts_ar_bits_addr_0;
  assign simpleAccessPorts_r_ready = simpleAccessPorts_r_ready_0;
  assign vrfReadDataPorts_0_valid = vrfReadDataPorts_0_valid_0;
  assign vrfReadDataPorts_0_bits_vs = vrfReadDataPorts_0_bits_vs_0;
  assign vrfReadDataPorts_0_bits_instructionIndex = vrfReadDataPorts_0_bits_instructionIndex_0;
  assign vrfReadDataPorts_1_valid = vrfReadDataPorts_1_valid_0;
  assign vrfReadDataPorts_1_bits_vs = vrfReadDataPorts_1_bits_vs_0;
  assign vrfReadDataPorts_1_bits_instructionIndex = vrfReadDataPorts_1_bits_instructionIndex_0;
  assign vrfReadDataPorts_2_valid = vrfReadDataPorts_2_valid_0;
  assign vrfReadDataPorts_2_bits_vs = vrfReadDataPorts_2_bits_vs_0;
  assign vrfReadDataPorts_2_bits_instructionIndex = vrfReadDataPorts_2_bits_instructionIndex_0;
  assign vrfReadDataPorts_3_valid = vrfReadDataPorts_3_valid_0;
  assign vrfReadDataPorts_3_bits_vs = vrfReadDataPorts_3_bits_vs_0;
  assign vrfReadDataPorts_3_bits_instructionIndex = vrfReadDataPorts_3_bits_instructionIndex_0;
  assign vrfReadDataPorts_4_valid = vrfReadDataPorts_4_valid_0;
  assign vrfReadDataPorts_4_bits_vs = vrfReadDataPorts_4_bits_vs_0;
  assign vrfReadDataPorts_4_bits_instructionIndex = vrfReadDataPorts_4_bits_instructionIndex_0;
  assign vrfReadDataPorts_5_valid = vrfReadDataPorts_5_valid_0;
  assign vrfReadDataPorts_5_bits_vs = vrfReadDataPorts_5_bits_vs_0;
  assign vrfReadDataPorts_5_bits_instructionIndex = vrfReadDataPorts_5_bits_instructionIndex_0;
  assign vrfReadDataPorts_6_valid = vrfReadDataPorts_6_valid_0;
  assign vrfReadDataPorts_6_bits_vs = vrfReadDataPorts_6_bits_vs_0;
  assign vrfReadDataPorts_6_bits_instructionIndex = vrfReadDataPorts_6_bits_instructionIndex_0;
  assign vrfReadDataPorts_7_valid = vrfReadDataPorts_7_valid_0;
  assign vrfReadDataPorts_7_bits_vs = vrfReadDataPorts_7_bits_vs_0;
  assign vrfReadDataPorts_7_bits_instructionIndex = vrfReadDataPorts_7_bits_instructionIndex_0;
  assign vrfReadDataPorts_8_valid = vrfReadDataPorts_8_valid_0;
  assign vrfReadDataPorts_8_bits_vs = vrfReadDataPorts_8_bits_vs_0;
  assign vrfReadDataPorts_8_bits_instructionIndex = vrfReadDataPorts_8_bits_instructionIndex_0;
  assign vrfReadDataPorts_9_valid = vrfReadDataPorts_9_valid_0;
  assign vrfReadDataPorts_9_bits_vs = vrfReadDataPorts_9_bits_vs_0;
  assign vrfReadDataPorts_9_bits_instructionIndex = vrfReadDataPorts_9_bits_instructionIndex_0;
  assign vrfReadDataPorts_10_valid = vrfReadDataPorts_10_valid_0;
  assign vrfReadDataPorts_10_bits_vs = vrfReadDataPorts_10_bits_vs_0;
  assign vrfReadDataPorts_10_bits_instructionIndex = vrfReadDataPorts_10_bits_instructionIndex_0;
  assign vrfReadDataPorts_11_valid = vrfReadDataPorts_11_valid_0;
  assign vrfReadDataPorts_11_bits_vs = vrfReadDataPorts_11_bits_vs_0;
  assign vrfReadDataPorts_11_bits_instructionIndex = vrfReadDataPorts_11_bits_instructionIndex_0;
  assign vrfReadDataPorts_12_valid = vrfReadDataPorts_12_valid_0;
  assign vrfReadDataPorts_12_bits_vs = vrfReadDataPorts_12_bits_vs_0;
  assign vrfReadDataPorts_12_bits_instructionIndex = vrfReadDataPorts_12_bits_instructionIndex_0;
  assign vrfReadDataPorts_13_valid = vrfReadDataPorts_13_valid_0;
  assign vrfReadDataPorts_13_bits_vs = vrfReadDataPorts_13_bits_vs_0;
  assign vrfReadDataPorts_13_bits_instructionIndex = vrfReadDataPorts_13_bits_instructionIndex_0;
  assign vrfReadDataPorts_14_valid = vrfReadDataPorts_14_valid_0;
  assign vrfReadDataPorts_14_bits_vs = vrfReadDataPorts_14_bits_vs_0;
  assign vrfReadDataPorts_14_bits_instructionIndex = vrfReadDataPorts_14_bits_instructionIndex_0;
  assign vrfReadDataPorts_15_valid = vrfReadDataPorts_15_valid_0;
  assign vrfReadDataPorts_15_bits_vs = vrfReadDataPorts_15_bits_vs_0;
  assign vrfReadDataPorts_15_bits_instructionIndex = vrfReadDataPorts_15_bits_instructionIndex_0;
  assign vrfReadDataPorts_16_valid = vrfReadDataPorts_16_valid_0;
  assign vrfReadDataPorts_16_bits_vs = vrfReadDataPorts_16_bits_vs_0;
  assign vrfReadDataPorts_16_bits_instructionIndex = vrfReadDataPorts_16_bits_instructionIndex_0;
  assign vrfReadDataPorts_17_valid = vrfReadDataPorts_17_valid_0;
  assign vrfReadDataPorts_17_bits_vs = vrfReadDataPorts_17_bits_vs_0;
  assign vrfReadDataPorts_17_bits_instructionIndex = vrfReadDataPorts_17_bits_instructionIndex_0;
  assign vrfReadDataPorts_18_valid = vrfReadDataPorts_18_valid_0;
  assign vrfReadDataPorts_18_bits_vs = vrfReadDataPorts_18_bits_vs_0;
  assign vrfReadDataPorts_18_bits_instructionIndex = vrfReadDataPorts_18_bits_instructionIndex_0;
  assign vrfReadDataPorts_19_valid = vrfReadDataPorts_19_valid_0;
  assign vrfReadDataPorts_19_bits_vs = vrfReadDataPorts_19_bits_vs_0;
  assign vrfReadDataPorts_19_bits_instructionIndex = vrfReadDataPorts_19_bits_instructionIndex_0;
  assign vrfReadDataPorts_20_valid = vrfReadDataPorts_20_valid_0;
  assign vrfReadDataPorts_20_bits_vs = vrfReadDataPorts_20_bits_vs_0;
  assign vrfReadDataPorts_20_bits_instructionIndex = vrfReadDataPorts_20_bits_instructionIndex_0;
  assign vrfReadDataPorts_21_valid = vrfReadDataPorts_21_valid_0;
  assign vrfReadDataPorts_21_bits_vs = vrfReadDataPorts_21_bits_vs_0;
  assign vrfReadDataPorts_21_bits_instructionIndex = vrfReadDataPorts_21_bits_instructionIndex_0;
  assign vrfReadDataPorts_22_valid = vrfReadDataPorts_22_valid_0;
  assign vrfReadDataPorts_22_bits_vs = vrfReadDataPorts_22_bits_vs_0;
  assign vrfReadDataPorts_22_bits_instructionIndex = vrfReadDataPorts_22_bits_instructionIndex_0;
  assign vrfReadDataPorts_23_valid = vrfReadDataPorts_23_valid_0;
  assign vrfReadDataPorts_23_bits_vs = vrfReadDataPorts_23_bits_vs_0;
  assign vrfReadDataPorts_23_bits_instructionIndex = vrfReadDataPorts_23_bits_instructionIndex_0;
  assign vrfReadDataPorts_24_valid = vrfReadDataPorts_24_valid_0;
  assign vrfReadDataPorts_24_bits_vs = vrfReadDataPorts_24_bits_vs_0;
  assign vrfReadDataPorts_24_bits_instructionIndex = vrfReadDataPorts_24_bits_instructionIndex_0;
  assign vrfReadDataPorts_25_valid = vrfReadDataPorts_25_valid_0;
  assign vrfReadDataPorts_25_bits_vs = vrfReadDataPorts_25_bits_vs_0;
  assign vrfReadDataPorts_25_bits_instructionIndex = vrfReadDataPorts_25_bits_instructionIndex_0;
  assign vrfReadDataPorts_26_valid = vrfReadDataPorts_26_valid_0;
  assign vrfReadDataPorts_26_bits_vs = vrfReadDataPorts_26_bits_vs_0;
  assign vrfReadDataPorts_26_bits_instructionIndex = vrfReadDataPorts_26_bits_instructionIndex_0;
  assign vrfReadDataPorts_27_valid = vrfReadDataPorts_27_valid_0;
  assign vrfReadDataPorts_27_bits_vs = vrfReadDataPorts_27_bits_vs_0;
  assign vrfReadDataPorts_27_bits_instructionIndex = vrfReadDataPorts_27_bits_instructionIndex_0;
  assign vrfReadDataPorts_28_valid = vrfReadDataPorts_28_valid_0;
  assign vrfReadDataPorts_28_bits_vs = vrfReadDataPorts_28_bits_vs_0;
  assign vrfReadDataPorts_28_bits_instructionIndex = vrfReadDataPorts_28_bits_instructionIndex_0;
  assign vrfReadDataPorts_29_valid = vrfReadDataPorts_29_valid_0;
  assign vrfReadDataPorts_29_bits_vs = vrfReadDataPorts_29_bits_vs_0;
  assign vrfReadDataPorts_29_bits_instructionIndex = vrfReadDataPorts_29_bits_instructionIndex_0;
  assign vrfReadDataPorts_30_valid = vrfReadDataPorts_30_valid_0;
  assign vrfReadDataPorts_30_bits_vs = vrfReadDataPorts_30_bits_vs_0;
  assign vrfReadDataPorts_30_bits_instructionIndex = vrfReadDataPorts_30_bits_instructionIndex_0;
  assign vrfReadDataPorts_31_valid = vrfReadDataPorts_31_valid_0;
  assign vrfReadDataPorts_31_bits_vs = vrfReadDataPorts_31_bits_vs_0;
  assign vrfReadDataPorts_31_bits_instructionIndex = vrfReadDataPorts_31_bits_instructionIndex_0;
  assign vrfWritePort_0_valid = vrfWritePort_0_valid_0;
  assign vrfWritePort_0_bits_vd = vrfWritePort_0_bits_vd_0;
  assign vrfWritePort_0_bits_mask = vrfWritePort_0_bits_mask_0;
  assign vrfWritePort_0_bits_data = vrfWritePort_0_bits_data_0;
  assign vrfWritePort_0_bits_last = vrfWritePort_0_bits_last_0;
  assign vrfWritePort_0_bits_instructionIndex = vrfWritePort_0_bits_instructionIndex_0;
  assign vrfWritePort_1_valid = vrfWritePort_1_valid_0;
  assign vrfWritePort_1_bits_vd = vrfWritePort_1_bits_vd_0;
  assign vrfWritePort_1_bits_mask = vrfWritePort_1_bits_mask_0;
  assign vrfWritePort_1_bits_data = vrfWritePort_1_bits_data_0;
  assign vrfWritePort_1_bits_last = vrfWritePort_1_bits_last_0;
  assign vrfWritePort_1_bits_instructionIndex = vrfWritePort_1_bits_instructionIndex_0;
  assign vrfWritePort_2_valid = vrfWritePort_2_valid_0;
  assign vrfWritePort_2_bits_vd = vrfWritePort_2_bits_vd_0;
  assign vrfWritePort_2_bits_mask = vrfWritePort_2_bits_mask_0;
  assign vrfWritePort_2_bits_data = vrfWritePort_2_bits_data_0;
  assign vrfWritePort_2_bits_last = vrfWritePort_2_bits_last_0;
  assign vrfWritePort_2_bits_instructionIndex = vrfWritePort_2_bits_instructionIndex_0;
  assign vrfWritePort_3_valid = vrfWritePort_3_valid_0;
  assign vrfWritePort_3_bits_vd = vrfWritePort_3_bits_vd_0;
  assign vrfWritePort_3_bits_mask = vrfWritePort_3_bits_mask_0;
  assign vrfWritePort_3_bits_data = vrfWritePort_3_bits_data_0;
  assign vrfWritePort_3_bits_last = vrfWritePort_3_bits_last_0;
  assign vrfWritePort_3_bits_instructionIndex = vrfWritePort_3_bits_instructionIndex_0;
  assign vrfWritePort_4_valid = vrfWritePort_4_valid_0;
  assign vrfWritePort_4_bits_vd = vrfWritePort_4_bits_vd_0;
  assign vrfWritePort_4_bits_mask = vrfWritePort_4_bits_mask_0;
  assign vrfWritePort_4_bits_data = vrfWritePort_4_bits_data_0;
  assign vrfWritePort_4_bits_last = vrfWritePort_4_bits_last_0;
  assign vrfWritePort_4_bits_instructionIndex = vrfWritePort_4_bits_instructionIndex_0;
  assign vrfWritePort_5_valid = vrfWritePort_5_valid_0;
  assign vrfWritePort_5_bits_vd = vrfWritePort_5_bits_vd_0;
  assign vrfWritePort_5_bits_mask = vrfWritePort_5_bits_mask_0;
  assign vrfWritePort_5_bits_data = vrfWritePort_5_bits_data_0;
  assign vrfWritePort_5_bits_last = vrfWritePort_5_bits_last_0;
  assign vrfWritePort_5_bits_instructionIndex = vrfWritePort_5_bits_instructionIndex_0;
  assign vrfWritePort_6_valid = vrfWritePort_6_valid_0;
  assign vrfWritePort_6_bits_vd = vrfWritePort_6_bits_vd_0;
  assign vrfWritePort_6_bits_mask = vrfWritePort_6_bits_mask_0;
  assign vrfWritePort_6_bits_data = vrfWritePort_6_bits_data_0;
  assign vrfWritePort_6_bits_last = vrfWritePort_6_bits_last_0;
  assign vrfWritePort_6_bits_instructionIndex = vrfWritePort_6_bits_instructionIndex_0;
  assign vrfWritePort_7_valid = vrfWritePort_7_valid_0;
  assign vrfWritePort_7_bits_vd = vrfWritePort_7_bits_vd_0;
  assign vrfWritePort_7_bits_mask = vrfWritePort_7_bits_mask_0;
  assign vrfWritePort_7_bits_data = vrfWritePort_7_bits_data_0;
  assign vrfWritePort_7_bits_last = vrfWritePort_7_bits_last_0;
  assign vrfWritePort_7_bits_instructionIndex = vrfWritePort_7_bits_instructionIndex_0;
  assign vrfWritePort_8_valid = vrfWritePort_8_valid_0;
  assign vrfWritePort_8_bits_vd = vrfWritePort_8_bits_vd_0;
  assign vrfWritePort_8_bits_mask = vrfWritePort_8_bits_mask_0;
  assign vrfWritePort_8_bits_data = vrfWritePort_8_bits_data_0;
  assign vrfWritePort_8_bits_last = vrfWritePort_8_bits_last_0;
  assign vrfWritePort_8_bits_instructionIndex = vrfWritePort_8_bits_instructionIndex_0;
  assign vrfWritePort_9_valid = vrfWritePort_9_valid_0;
  assign vrfWritePort_9_bits_vd = vrfWritePort_9_bits_vd_0;
  assign vrfWritePort_9_bits_mask = vrfWritePort_9_bits_mask_0;
  assign vrfWritePort_9_bits_data = vrfWritePort_9_bits_data_0;
  assign vrfWritePort_9_bits_last = vrfWritePort_9_bits_last_0;
  assign vrfWritePort_9_bits_instructionIndex = vrfWritePort_9_bits_instructionIndex_0;
  assign vrfWritePort_10_valid = vrfWritePort_10_valid_0;
  assign vrfWritePort_10_bits_vd = vrfWritePort_10_bits_vd_0;
  assign vrfWritePort_10_bits_mask = vrfWritePort_10_bits_mask_0;
  assign vrfWritePort_10_bits_data = vrfWritePort_10_bits_data_0;
  assign vrfWritePort_10_bits_last = vrfWritePort_10_bits_last_0;
  assign vrfWritePort_10_bits_instructionIndex = vrfWritePort_10_bits_instructionIndex_0;
  assign vrfWritePort_11_valid = vrfWritePort_11_valid_0;
  assign vrfWritePort_11_bits_vd = vrfWritePort_11_bits_vd_0;
  assign vrfWritePort_11_bits_mask = vrfWritePort_11_bits_mask_0;
  assign vrfWritePort_11_bits_data = vrfWritePort_11_bits_data_0;
  assign vrfWritePort_11_bits_last = vrfWritePort_11_bits_last_0;
  assign vrfWritePort_11_bits_instructionIndex = vrfWritePort_11_bits_instructionIndex_0;
  assign vrfWritePort_12_valid = vrfWritePort_12_valid_0;
  assign vrfWritePort_12_bits_vd = vrfWritePort_12_bits_vd_0;
  assign vrfWritePort_12_bits_mask = vrfWritePort_12_bits_mask_0;
  assign vrfWritePort_12_bits_data = vrfWritePort_12_bits_data_0;
  assign vrfWritePort_12_bits_last = vrfWritePort_12_bits_last_0;
  assign vrfWritePort_12_bits_instructionIndex = vrfWritePort_12_bits_instructionIndex_0;
  assign vrfWritePort_13_valid = vrfWritePort_13_valid_0;
  assign vrfWritePort_13_bits_vd = vrfWritePort_13_bits_vd_0;
  assign vrfWritePort_13_bits_mask = vrfWritePort_13_bits_mask_0;
  assign vrfWritePort_13_bits_data = vrfWritePort_13_bits_data_0;
  assign vrfWritePort_13_bits_last = vrfWritePort_13_bits_last_0;
  assign vrfWritePort_13_bits_instructionIndex = vrfWritePort_13_bits_instructionIndex_0;
  assign vrfWritePort_14_valid = vrfWritePort_14_valid_0;
  assign vrfWritePort_14_bits_vd = vrfWritePort_14_bits_vd_0;
  assign vrfWritePort_14_bits_mask = vrfWritePort_14_bits_mask_0;
  assign vrfWritePort_14_bits_data = vrfWritePort_14_bits_data_0;
  assign vrfWritePort_14_bits_last = vrfWritePort_14_bits_last_0;
  assign vrfWritePort_14_bits_instructionIndex = vrfWritePort_14_bits_instructionIndex_0;
  assign vrfWritePort_15_valid = vrfWritePort_15_valid_0;
  assign vrfWritePort_15_bits_vd = vrfWritePort_15_bits_vd_0;
  assign vrfWritePort_15_bits_mask = vrfWritePort_15_bits_mask_0;
  assign vrfWritePort_15_bits_data = vrfWritePort_15_bits_data_0;
  assign vrfWritePort_15_bits_last = vrfWritePort_15_bits_last_0;
  assign vrfWritePort_15_bits_instructionIndex = vrfWritePort_15_bits_instructionIndex_0;
  assign vrfWritePort_16_valid = vrfWritePort_16_valid_0;
  assign vrfWritePort_16_bits_vd = vrfWritePort_16_bits_vd_0;
  assign vrfWritePort_16_bits_mask = vrfWritePort_16_bits_mask_0;
  assign vrfWritePort_16_bits_data = vrfWritePort_16_bits_data_0;
  assign vrfWritePort_16_bits_last = vrfWritePort_16_bits_last_0;
  assign vrfWritePort_16_bits_instructionIndex = vrfWritePort_16_bits_instructionIndex_0;
  assign vrfWritePort_17_valid = vrfWritePort_17_valid_0;
  assign vrfWritePort_17_bits_vd = vrfWritePort_17_bits_vd_0;
  assign vrfWritePort_17_bits_mask = vrfWritePort_17_bits_mask_0;
  assign vrfWritePort_17_bits_data = vrfWritePort_17_bits_data_0;
  assign vrfWritePort_17_bits_last = vrfWritePort_17_bits_last_0;
  assign vrfWritePort_17_bits_instructionIndex = vrfWritePort_17_bits_instructionIndex_0;
  assign vrfWritePort_18_valid = vrfWritePort_18_valid_0;
  assign vrfWritePort_18_bits_vd = vrfWritePort_18_bits_vd_0;
  assign vrfWritePort_18_bits_mask = vrfWritePort_18_bits_mask_0;
  assign vrfWritePort_18_bits_data = vrfWritePort_18_bits_data_0;
  assign vrfWritePort_18_bits_last = vrfWritePort_18_bits_last_0;
  assign vrfWritePort_18_bits_instructionIndex = vrfWritePort_18_bits_instructionIndex_0;
  assign vrfWritePort_19_valid = vrfWritePort_19_valid_0;
  assign vrfWritePort_19_bits_vd = vrfWritePort_19_bits_vd_0;
  assign vrfWritePort_19_bits_mask = vrfWritePort_19_bits_mask_0;
  assign vrfWritePort_19_bits_data = vrfWritePort_19_bits_data_0;
  assign vrfWritePort_19_bits_last = vrfWritePort_19_bits_last_0;
  assign vrfWritePort_19_bits_instructionIndex = vrfWritePort_19_bits_instructionIndex_0;
  assign vrfWritePort_20_valid = vrfWritePort_20_valid_0;
  assign vrfWritePort_20_bits_vd = vrfWritePort_20_bits_vd_0;
  assign vrfWritePort_20_bits_mask = vrfWritePort_20_bits_mask_0;
  assign vrfWritePort_20_bits_data = vrfWritePort_20_bits_data_0;
  assign vrfWritePort_20_bits_last = vrfWritePort_20_bits_last_0;
  assign vrfWritePort_20_bits_instructionIndex = vrfWritePort_20_bits_instructionIndex_0;
  assign vrfWritePort_21_valid = vrfWritePort_21_valid_0;
  assign vrfWritePort_21_bits_vd = vrfWritePort_21_bits_vd_0;
  assign vrfWritePort_21_bits_mask = vrfWritePort_21_bits_mask_0;
  assign vrfWritePort_21_bits_data = vrfWritePort_21_bits_data_0;
  assign vrfWritePort_21_bits_last = vrfWritePort_21_bits_last_0;
  assign vrfWritePort_21_bits_instructionIndex = vrfWritePort_21_bits_instructionIndex_0;
  assign vrfWritePort_22_valid = vrfWritePort_22_valid_0;
  assign vrfWritePort_22_bits_vd = vrfWritePort_22_bits_vd_0;
  assign vrfWritePort_22_bits_mask = vrfWritePort_22_bits_mask_0;
  assign vrfWritePort_22_bits_data = vrfWritePort_22_bits_data_0;
  assign vrfWritePort_22_bits_last = vrfWritePort_22_bits_last_0;
  assign vrfWritePort_22_bits_instructionIndex = vrfWritePort_22_bits_instructionIndex_0;
  assign vrfWritePort_23_valid = vrfWritePort_23_valid_0;
  assign vrfWritePort_23_bits_vd = vrfWritePort_23_bits_vd_0;
  assign vrfWritePort_23_bits_mask = vrfWritePort_23_bits_mask_0;
  assign vrfWritePort_23_bits_data = vrfWritePort_23_bits_data_0;
  assign vrfWritePort_23_bits_last = vrfWritePort_23_bits_last_0;
  assign vrfWritePort_23_bits_instructionIndex = vrfWritePort_23_bits_instructionIndex_0;
  assign vrfWritePort_24_valid = vrfWritePort_24_valid_0;
  assign vrfWritePort_24_bits_vd = vrfWritePort_24_bits_vd_0;
  assign vrfWritePort_24_bits_mask = vrfWritePort_24_bits_mask_0;
  assign vrfWritePort_24_bits_data = vrfWritePort_24_bits_data_0;
  assign vrfWritePort_24_bits_last = vrfWritePort_24_bits_last_0;
  assign vrfWritePort_24_bits_instructionIndex = vrfWritePort_24_bits_instructionIndex_0;
  assign vrfWritePort_25_valid = vrfWritePort_25_valid_0;
  assign vrfWritePort_25_bits_vd = vrfWritePort_25_bits_vd_0;
  assign vrfWritePort_25_bits_mask = vrfWritePort_25_bits_mask_0;
  assign vrfWritePort_25_bits_data = vrfWritePort_25_bits_data_0;
  assign vrfWritePort_25_bits_last = vrfWritePort_25_bits_last_0;
  assign vrfWritePort_25_bits_instructionIndex = vrfWritePort_25_bits_instructionIndex_0;
  assign vrfWritePort_26_valid = vrfWritePort_26_valid_0;
  assign vrfWritePort_26_bits_vd = vrfWritePort_26_bits_vd_0;
  assign vrfWritePort_26_bits_mask = vrfWritePort_26_bits_mask_0;
  assign vrfWritePort_26_bits_data = vrfWritePort_26_bits_data_0;
  assign vrfWritePort_26_bits_last = vrfWritePort_26_bits_last_0;
  assign vrfWritePort_26_bits_instructionIndex = vrfWritePort_26_bits_instructionIndex_0;
  assign vrfWritePort_27_valid = vrfWritePort_27_valid_0;
  assign vrfWritePort_27_bits_vd = vrfWritePort_27_bits_vd_0;
  assign vrfWritePort_27_bits_mask = vrfWritePort_27_bits_mask_0;
  assign vrfWritePort_27_bits_data = vrfWritePort_27_bits_data_0;
  assign vrfWritePort_27_bits_last = vrfWritePort_27_bits_last_0;
  assign vrfWritePort_27_bits_instructionIndex = vrfWritePort_27_bits_instructionIndex_0;
  assign vrfWritePort_28_valid = vrfWritePort_28_valid_0;
  assign vrfWritePort_28_bits_vd = vrfWritePort_28_bits_vd_0;
  assign vrfWritePort_28_bits_mask = vrfWritePort_28_bits_mask_0;
  assign vrfWritePort_28_bits_data = vrfWritePort_28_bits_data_0;
  assign vrfWritePort_28_bits_last = vrfWritePort_28_bits_last_0;
  assign vrfWritePort_28_bits_instructionIndex = vrfWritePort_28_bits_instructionIndex_0;
  assign vrfWritePort_29_valid = vrfWritePort_29_valid_0;
  assign vrfWritePort_29_bits_vd = vrfWritePort_29_bits_vd_0;
  assign vrfWritePort_29_bits_mask = vrfWritePort_29_bits_mask_0;
  assign vrfWritePort_29_bits_data = vrfWritePort_29_bits_data_0;
  assign vrfWritePort_29_bits_last = vrfWritePort_29_bits_last_0;
  assign vrfWritePort_29_bits_instructionIndex = vrfWritePort_29_bits_instructionIndex_0;
  assign vrfWritePort_30_valid = vrfWritePort_30_valid_0;
  assign vrfWritePort_30_bits_vd = vrfWritePort_30_bits_vd_0;
  assign vrfWritePort_30_bits_mask = vrfWritePort_30_bits_mask_0;
  assign vrfWritePort_30_bits_data = vrfWritePort_30_bits_data_0;
  assign vrfWritePort_30_bits_last = vrfWritePort_30_bits_last_0;
  assign vrfWritePort_30_bits_instructionIndex = vrfWritePort_30_bits_instructionIndex_0;
  assign vrfWritePort_31_valid = vrfWritePort_31_valid_0;
  assign vrfWritePort_31_bits_vd = vrfWritePort_31_bits_vd_0;
  assign vrfWritePort_31_bits_mask = vrfWritePort_31_bits_mask_0;
  assign vrfWritePort_31_bits_data = vrfWritePort_31_bits_data_0;
  assign vrfWritePort_31_bits_last = vrfWritePort_31_bits_last_0;
  assign vrfWritePort_31_bits_instructionIndex = vrfWritePort_31_bits_instructionIndex_0;
  assign dataInWriteQueue_0 = {dataInWriteQueue_0_hi, dataInWriteQueue_0_lo} | dataInMSHR;
  assign dataInWriteQueue_1 = {dataInWriteQueue_1_hi, dataInWriteQueue_1_lo} | dataInMSHR;
  assign dataInWriteQueue_2 = {dataInWriteQueue_2_hi, dataInWriteQueue_2_lo} | dataInMSHR;
  assign dataInWriteQueue_3 = {dataInWriteQueue_3_hi, dataInWriteQueue_3_lo} | dataInMSHR;
  assign dataInWriteQueue_4 = {dataInWriteQueue_4_hi, dataInWriteQueue_4_lo} | dataInMSHR;
  assign dataInWriteQueue_5 = {dataInWriteQueue_5_hi, dataInWriteQueue_5_lo} | dataInMSHR;
  assign dataInWriteQueue_6 = {dataInWriteQueue_6_hi, dataInWriteQueue_6_lo} | dataInMSHR;
  assign dataInWriteQueue_7 = {dataInWriteQueue_7_hi, dataInWriteQueue_7_lo} | dataInMSHR;
  assign dataInWriteQueue_8 = {dataInWriteQueue_8_hi, dataInWriteQueue_8_lo} | dataInMSHR;
  assign dataInWriteQueue_9 = {dataInWriteQueue_9_hi, dataInWriteQueue_9_lo} | dataInMSHR;
  assign dataInWriteQueue_10 = {dataInWriteQueue_10_hi, dataInWriteQueue_10_lo} | dataInMSHR;
  assign dataInWriteQueue_11 = {dataInWriteQueue_11_hi, dataInWriteQueue_11_lo} | dataInMSHR;
  assign dataInWriteQueue_12 = {dataInWriteQueue_12_hi, dataInWriteQueue_12_lo} | dataInMSHR;
  assign dataInWriteQueue_13 = {dataInWriteQueue_13_hi, dataInWriteQueue_13_lo} | dataInMSHR;
  assign dataInWriteQueue_14 = {dataInWriteQueue_14_hi, dataInWriteQueue_14_lo} | dataInMSHR;
  assign dataInWriteQueue_15 = {dataInWriteQueue_15_hi, dataInWriteQueue_15_lo} | dataInMSHR;
  assign dataInWriteQueue_16 = {dataInWriteQueue_16_hi, dataInWriteQueue_16_lo} | dataInMSHR;
  assign dataInWriteQueue_17 = {dataInWriteQueue_17_hi, dataInWriteQueue_17_lo} | dataInMSHR;
  assign dataInWriteQueue_18 = {dataInWriteQueue_18_hi, dataInWriteQueue_18_lo} | dataInMSHR;
  assign dataInWriteQueue_19 = {dataInWriteQueue_19_hi, dataInWriteQueue_19_lo} | dataInMSHR;
  assign dataInWriteQueue_20 = {dataInWriteQueue_20_hi, dataInWriteQueue_20_lo} | dataInMSHR;
  assign dataInWriteQueue_21 = {dataInWriteQueue_21_hi, dataInWriteQueue_21_lo} | dataInMSHR;
  assign dataInWriteQueue_22 = {dataInWriteQueue_22_hi, dataInWriteQueue_22_lo} | dataInMSHR;
  assign dataInWriteQueue_23 = {dataInWriteQueue_23_hi, dataInWriteQueue_23_lo} | dataInMSHR;
  assign dataInWriteQueue_24 = {dataInWriteQueue_24_hi, dataInWriteQueue_24_lo} | dataInMSHR;
  assign dataInWriteQueue_25 = {dataInWriteQueue_25_hi, dataInWriteQueue_25_lo} | dataInMSHR;
  assign dataInWriteQueue_26 = {dataInWriteQueue_26_hi, dataInWriteQueue_26_lo} | dataInMSHR;
  assign dataInWriteQueue_27 = {dataInWriteQueue_27_hi, dataInWriteQueue_27_lo} | dataInMSHR;
  assign dataInWriteQueue_28 = {dataInWriteQueue_28_hi, dataInWriteQueue_28_lo} | dataInMSHR;
  assign dataInWriteQueue_29 = {dataInWriteQueue_29_hi, dataInWriteQueue_29_lo} | dataInMSHR;
  assign dataInWriteQueue_30 = {dataInWriteQueue_30_hi, dataInWriteQueue_30_lo} | dataInMSHR;
  assign dataInWriteQueue_31 = {dataInWriteQueue_31_hi, dataInWriteQueue_31_lo} | dataInMSHR;
  assign lastReport = (_loadUnit_status_last ? 8'h1 << _GEN_18 : 8'h0) | (_storeUnit_status_last ? 8'h1 << _storeUnit_status_instructionIndex : 8'h0) | (_otherUnit_status_last ? 8'h1 << _GEN_19 : 8'h0);
  assign tokenIO_offsetGroupRelease = {tokenIO_offsetGroupRelease_hi, tokenIO_offsetGroupRelease_lo};
endmodule

