
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module T1TokenManager(
  input        clock,
               reset,
               instructionIssue_valid,
  input  [2:0] instructionIssue_bits_instructionIndex,
  input        instructionIssue_bits_writeV0,
               instructionIssue_bits_useV0AsMask,
               instructionIssue_bits_toLane,
               instructionIssue_bits_toMask,
               lsuWriteV0_0_valid,
  input  [2:0] lsuWriteV0_0_bits,
  input        lsuWriteV0_1_valid,
  input  [2:0] lsuWriteV0_1_bits,
  input        lsuWriteV0_2_valid,
  input  [2:0] lsuWriteV0_2_bits,
  input        lsuWriteV0_3_valid,
  input  [2:0] lsuWriteV0_3_bits,
  input        lsuWriteV0_4_valid,
  input  [2:0] lsuWriteV0_4_bits,
  input        lsuWriteV0_5_valid,
  input  [2:0] lsuWriteV0_5_bits,
  input        lsuWriteV0_6_valid,
  input  [2:0] lsuWriteV0_6_bits,
  input        lsuWriteV0_7_valid,
  input  [2:0] lsuWriteV0_7_bits,
  input        lsuWriteV0_8_valid,
  input  [2:0] lsuWriteV0_8_bits,
  input        lsuWriteV0_9_valid,
  input  [2:0] lsuWriteV0_9_bits,
  input        lsuWriteV0_10_valid,
  input  [2:0] lsuWriteV0_10_bits,
  input        lsuWriteV0_11_valid,
  input  [2:0] lsuWriteV0_11_bits,
  input        lsuWriteV0_12_valid,
  input  [2:0] lsuWriteV0_12_bits,
  input        lsuWriteV0_13_valid,
  input  [2:0] lsuWriteV0_13_bits,
  input        lsuWriteV0_14_valid,
  input  [2:0] lsuWriteV0_14_bits,
  input        lsuWriteV0_15_valid,
  input  [2:0] lsuWriteV0_15_bits,
  input        lsuWriteV0_16_valid,
  input  [2:0] lsuWriteV0_16_bits,
  input        lsuWriteV0_17_valid,
  input  [2:0] lsuWriteV0_17_bits,
  input        lsuWriteV0_18_valid,
  input  [2:0] lsuWriteV0_18_bits,
  input        lsuWriteV0_19_valid,
  input  [2:0] lsuWriteV0_19_bits,
  input        lsuWriteV0_20_valid,
  input  [2:0] lsuWriteV0_20_bits,
  input        lsuWriteV0_21_valid,
  input  [2:0] lsuWriteV0_21_bits,
  input        lsuWriteV0_22_valid,
  input  [2:0] lsuWriteV0_22_bits,
  input        lsuWriteV0_23_valid,
  input  [2:0] lsuWriteV0_23_bits,
  input        lsuWriteV0_24_valid,
  input  [2:0] lsuWriteV0_24_bits,
  input        lsuWriteV0_25_valid,
  input  [2:0] lsuWriteV0_25_bits,
  input        lsuWriteV0_26_valid,
  input  [2:0] lsuWriteV0_26_bits,
  input        lsuWriteV0_27_valid,
  input  [2:0] lsuWriteV0_27_bits,
  input        lsuWriteV0_28_valid,
  input  [2:0] lsuWriteV0_28_bits,
  input        lsuWriteV0_29_valid,
  input  [2:0] lsuWriteV0_29_bits,
  input        lsuWriteV0_30_valid,
  input  [2:0] lsuWriteV0_30_bits,
  input        lsuWriteV0_31_valid,
  input  [2:0] lsuWriteV0_31_bits,
  output       issueAllow,
  input  [7:0] instructionFinish_0,
               instructionFinish_1,
               instructionFinish_2,
               instructionFinish_3,
               instructionFinish_4,
               instructionFinish_5,
               instructionFinish_6,
               instructionFinish_7,
               instructionFinish_8,
               instructionFinish_9,
               instructionFinish_10,
               instructionFinish_11,
               instructionFinish_12,
               instructionFinish_13,
               instructionFinish_14,
               instructionFinish_15,
               instructionFinish_16,
               instructionFinish_17,
               instructionFinish_18,
               instructionFinish_19,
               instructionFinish_20,
               instructionFinish_21,
               instructionFinish_22,
               instructionFinish_23,
               instructionFinish_24,
               instructionFinish_25,
               instructionFinish_26,
               instructionFinish_27,
               instructionFinish_28,
               instructionFinish_29,
               instructionFinish_30,
               instructionFinish_31,
  output [7:0] v0WriteValid,
  input        maskUnitFree
);

  wire [7:0] issueIndex1H = 8'h1 << instructionIssue_bits_instructionIndex;
  wire [7:0] v0WriteValidVec_lsuWriteSet = lsuWriteV0_0_valid ? 8'h1 << lsuWriteV0_0_bits : 8'h0;
  wire       _maskUnitWriteV0_set_T = instructionIssue_valid & instructionIssue_bits_writeV0;
  wire       _GEN = _maskUnitWriteV0_set_T & instructionIssue_bits_toLane;
  wire       v0WriteValidVec_v0WriteIssue;
  assign v0WriteValidVec_v0WriteIssue = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_1;
  assign v0WriteValidVec_v0WriteIssue_1 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_2;
  assign v0WriteValidVec_v0WriteIssue_2 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_3;
  assign v0WriteValidVec_v0WriteIssue_3 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_4;
  assign v0WriteValidVec_v0WriteIssue_4 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_5;
  assign v0WriteValidVec_v0WriteIssue_5 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_6;
  assign v0WriteValidVec_v0WriteIssue_6 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_7;
  assign v0WriteValidVec_v0WriteIssue_7 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_8;
  assign v0WriteValidVec_v0WriteIssue_8 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_9;
  assign v0WriteValidVec_v0WriteIssue_9 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_10;
  assign v0WriteValidVec_v0WriteIssue_10 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_11;
  assign v0WriteValidVec_v0WriteIssue_11 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_12;
  assign v0WriteValidVec_v0WriteIssue_12 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_13;
  assign v0WriteValidVec_v0WriteIssue_13 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_14;
  assign v0WriteValidVec_v0WriteIssue_14 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_15;
  assign v0WriteValidVec_v0WriteIssue_15 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_16;
  assign v0WriteValidVec_v0WriteIssue_16 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_17;
  assign v0WriteValidVec_v0WriteIssue_17 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_18;
  assign v0WriteValidVec_v0WriteIssue_18 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_19;
  assign v0WriteValidVec_v0WriteIssue_19 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_20;
  assign v0WriteValidVec_v0WriteIssue_20 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_21;
  assign v0WriteValidVec_v0WriteIssue_21 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_22;
  assign v0WriteValidVec_v0WriteIssue_22 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_23;
  assign v0WriteValidVec_v0WriteIssue_23 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_24;
  assign v0WriteValidVec_v0WriteIssue_24 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_25;
  assign v0WriteValidVec_v0WriteIssue_25 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_26;
  assign v0WriteValidVec_v0WriteIssue_26 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_27;
  assign v0WriteValidVec_v0WriteIssue_27 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_28;
  assign v0WriteValidVec_v0WriteIssue_28 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_29;
  assign v0WriteValidVec_v0WriteIssue_29 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_30;
  assign v0WriteValidVec_v0WriteIssue_30 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_31;
  assign v0WriteValidVec_v0WriteIssue_31 = _GEN;
  wire [7:0] v0WriteValidVec_updateOH = v0WriteValidVec_v0WriteIssue ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res;
  reg        v0WriteValidVec_res_1;
  reg        v0WriteValidVec_res_2;
  reg        v0WriteValidVec_res_3;
  reg        v0WriteValidVec_res_4;
  reg        v0WriteValidVec_res_5;
  reg        v0WriteValidVec_res_6;
  reg        v0WriteValidVec_res_7;
  wire [1:0] v0WriteValidVec_lo_lo = {v0WriteValidVec_res_1, v0WriteValidVec_res};
  wire [1:0] v0WriteValidVec_lo_hi = {v0WriteValidVec_res_3, v0WriteValidVec_res_2};
  wire [3:0] v0WriteValidVec_lo = {v0WriteValidVec_lo_hi, v0WriteValidVec_lo_lo};
  wire [1:0] v0WriteValidVec_hi_lo = {v0WriteValidVec_res_5, v0WriteValidVec_res_4};
  wire [1:0] v0WriteValidVec_hi_hi = {v0WriteValidVec_res_7, v0WriteValidVec_res_6};
  wire [3:0] v0WriteValidVec_hi = {v0WriteValidVec_hi_hi, v0WriteValidVec_hi_lo};
  wire [7:0] v0WriteValidVec_0 = {v0WriteValidVec_hi, v0WriteValidVec_lo};
  wire [7:0] v0WriteValidVec_lsuWriteSet_1 = lsuWriteV0_1_valid ? 8'h1 << lsuWriteV0_1_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_1 = v0WriteValidVec_v0WriteIssue_1 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_8;
  reg        v0WriteValidVec_res_9;
  reg        v0WriteValidVec_res_10;
  reg        v0WriteValidVec_res_11;
  reg        v0WriteValidVec_res_12;
  reg        v0WriteValidVec_res_13;
  reg        v0WriteValidVec_res_14;
  reg        v0WriteValidVec_res_15;
  wire [1:0] v0WriteValidVec_lo_lo_1 = {v0WriteValidVec_res_9, v0WriteValidVec_res_8};
  wire [1:0] v0WriteValidVec_lo_hi_1 = {v0WriteValidVec_res_11, v0WriteValidVec_res_10};
  wire [3:0] v0WriteValidVec_lo_1 = {v0WriteValidVec_lo_hi_1, v0WriteValidVec_lo_lo_1};
  wire [1:0] v0WriteValidVec_hi_lo_1 = {v0WriteValidVec_res_13, v0WriteValidVec_res_12};
  wire [1:0] v0WriteValidVec_hi_hi_1 = {v0WriteValidVec_res_15, v0WriteValidVec_res_14};
  wire [3:0] v0WriteValidVec_hi_1 = {v0WriteValidVec_hi_hi_1, v0WriteValidVec_hi_lo_1};
  wire [7:0] v0WriteValidVec_1 = {v0WriteValidVec_hi_1, v0WriteValidVec_lo_1};
  wire [7:0] v0WriteValidVec_lsuWriteSet_2 = lsuWriteV0_2_valid ? 8'h1 << lsuWriteV0_2_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_2 = v0WriteValidVec_v0WriteIssue_2 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_16;
  reg        v0WriteValidVec_res_17;
  reg        v0WriteValidVec_res_18;
  reg        v0WriteValidVec_res_19;
  reg        v0WriteValidVec_res_20;
  reg        v0WriteValidVec_res_21;
  reg        v0WriteValidVec_res_22;
  reg        v0WriteValidVec_res_23;
  wire [1:0] v0WriteValidVec_lo_lo_2 = {v0WriteValidVec_res_17, v0WriteValidVec_res_16};
  wire [1:0] v0WriteValidVec_lo_hi_2 = {v0WriteValidVec_res_19, v0WriteValidVec_res_18};
  wire [3:0] v0WriteValidVec_lo_2 = {v0WriteValidVec_lo_hi_2, v0WriteValidVec_lo_lo_2};
  wire [1:0] v0WriteValidVec_hi_lo_2 = {v0WriteValidVec_res_21, v0WriteValidVec_res_20};
  wire [1:0] v0WriteValidVec_hi_hi_2 = {v0WriteValidVec_res_23, v0WriteValidVec_res_22};
  wire [3:0] v0WriteValidVec_hi_2 = {v0WriteValidVec_hi_hi_2, v0WriteValidVec_hi_lo_2};
  wire [7:0] v0WriteValidVec_2 = {v0WriteValidVec_hi_2, v0WriteValidVec_lo_2};
  wire [7:0] v0WriteValidVec_lsuWriteSet_3 = lsuWriteV0_3_valid ? 8'h1 << lsuWriteV0_3_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_3 = v0WriteValidVec_v0WriteIssue_3 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_24;
  reg        v0WriteValidVec_res_25;
  reg        v0WriteValidVec_res_26;
  reg        v0WriteValidVec_res_27;
  reg        v0WriteValidVec_res_28;
  reg        v0WriteValidVec_res_29;
  reg        v0WriteValidVec_res_30;
  reg        v0WriteValidVec_res_31;
  wire [1:0] v0WriteValidVec_lo_lo_3 = {v0WriteValidVec_res_25, v0WriteValidVec_res_24};
  wire [1:0] v0WriteValidVec_lo_hi_3 = {v0WriteValidVec_res_27, v0WriteValidVec_res_26};
  wire [3:0] v0WriteValidVec_lo_3 = {v0WriteValidVec_lo_hi_3, v0WriteValidVec_lo_lo_3};
  wire [1:0] v0WriteValidVec_hi_lo_3 = {v0WriteValidVec_res_29, v0WriteValidVec_res_28};
  wire [1:0] v0WriteValidVec_hi_hi_3 = {v0WriteValidVec_res_31, v0WriteValidVec_res_30};
  wire [3:0] v0WriteValidVec_hi_3 = {v0WriteValidVec_hi_hi_3, v0WriteValidVec_hi_lo_3};
  wire [7:0] v0WriteValidVec_3 = {v0WriteValidVec_hi_3, v0WriteValidVec_lo_3};
  wire [7:0] v0WriteValidVec_lsuWriteSet_4 = lsuWriteV0_4_valid ? 8'h1 << lsuWriteV0_4_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_4 = v0WriteValidVec_v0WriteIssue_4 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_32;
  reg        v0WriteValidVec_res_33;
  reg        v0WriteValidVec_res_34;
  reg        v0WriteValidVec_res_35;
  reg        v0WriteValidVec_res_36;
  reg        v0WriteValidVec_res_37;
  reg        v0WriteValidVec_res_38;
  reg        v0WriteValidVec_res_39;
  wire [1:0] v0WriteValidVec_lo_lo_4 = {v0WriteValidVec_res_33, v0WriteValidVec_res_32};
  wire [1:0] v0WriteValidVec_lo_hi_4 = {v0WriteValidVec_res_35, v0WriteValidVec_res_34};
  wire [3:0] v0WriteValidVec_lo_4 = {v0WriteValidVec_lo_hi_4, v0WriteValidVec_lo_lo_4};
  wire [1:0] v0WriteValidVec_hi_lo_4 = {v0WriteValidVec_res_37, v0WriteValidVec_res_36};
  wire [1:0] v0WriteValidVec_hi_hi_4 = {v0WriteValidVec_res_39, v0WriteValidVec_res_38};
  wire [3:0] v0WriteValidVec_hi_4 = {v0WriteValidVec_hi_hi_4, v0WriteValidVec_hi_lo_4};
  wire [7:0] v0WriteValidVec_4 = {v0WriteValidVec_hi_4, v0WriteValidVec_lo_4};
  wire [7:0] v0WriteValidVec_lsuWriteSet_5 = lsuWriteV0_5_valid ? 8'h1 << lsuWriteV0_5_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_5 = v0WriteValidVec_v0WriteIssue_5 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_40;
  reg        v0WriteValidVec_res_41;
  reg        v0WriteValidVec_res_42;
  reg        v0WriteValidVec_res_43;
  reg        v0WriteValidVec_res_44;
  reg        v0WriteValidVec_res_45;
  reg        v0WriteValidVec_res_46;
  reg        v0WriteValidVec_res_47;
  wire [1:0] v0WriteValidVec_lo_lo_5 = {v0WriteValidVec_res_41, v0WriteValidVec_res_40};
  wire [1:0] v0WriteValidVec_lo_hi_5 = {v0WriteValidVec_res_43, v0WriteValidVec_res_42};
  wire [3:0] v0WriteValidVec_lo_5 = {v0WriteValidVec_lo_hi_5, v0WriteValidVec_lo_lo_5};
  wire [1:0] v0WriteValidVec_hi_lo_5 = {v0WriteValidVec_res_45, v0WriteValidVec_res_44};
  wire [1:0] v0WriteValidVec_hi_hi_5 = {v0WriteValidVec_res_47, v0WriteValidVec_res_46};
  wire [3:0] v0WriteValidVec_hi_5 = {v0WriteValidVec_hi_hi_5, v0WriteValidVec_hi_lo_5};
  wire [7:0] v0WriteValidVec_5 = {v0WriteValidVec_hi_5, v0WriteValidVec_lo_5};
  wire [7:0] v0WriteValidVec_lsuWriteSet_6 = lsuWriteV0_6_valid ? 8'h1 << lsuWriteV0_6_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_6 = v0WriteValidVec_v0WriteIssue_6 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_48;
  reg        v0WriteValidVec_res_49;
  reg        v0WriteValidVec_res_50;
  reg        v0WriteValidVec_res_51;
  reg        v0WriteValidVec_res_52;
  reg        v0WriteValidVec_res_53;
  reg        v0WriteValidVec_res_54;
  reg        v0WriteValidVec_res_55;
  wire [1:0] v0WriteValidVec_lo_lo_6 = {v0WriteValidVec_res_49, v0WriteValidVec_res_48};
  wire [1:0] v0WriteValidVec_lo_hi_6 = {v0WriteValidVec_res_51, v0WriteValidVec_res_50};
  wire [3:0] v0WriteValidVec_lo_6 = {v0WriteValidVec_lo_hi_6, v0WriteValidVec_lo_lo_6};
  wire [1:0] v0WriteValidVec_hi_lo_6 = {v0WriteValidVec_res_53, v0WriteValidVec_res_52};
  wire [1:0] v0WriteValidVec_hi_hi_6 = {v0WriteValidVec_res_55, v0WriteValidVec_res_54};
  wire [3:0] v0WriteValidVec_hi_6 = {v0WriteValidVec_hi_hi_6, v0WriteValidVec_hi_lo_6};
  wire [7:0] v0WriteValidVec_6 = {v0WriteValidVec_hi_6, v0WriteValidVec_lo_6};
  wire [7:0] v0WriteValidVec_lsuWriteSet_7 = lsuWriteV0_7_valid ? 8'h1 << lsuWriteV0_7_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_7 = v0WriteValidVec_v0WriteIssue_7 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_56;
  reg        v0WriteValidVec_res_57;
  reg        v0WriteValidVec_res_58;
  reg        v0WriteValidVec_res_59;
  reg        v0WriteValidVec_res_60;
  reg        v0WriteValidVec_res_61;
  reg        v0WriteValidVec_res_62;
  reg        v0WriteValidVec_res_63;
  wire [1:0] v0WriteValidVec_lo_lo_7 = {v0WriteValidVec_res_57, v0WriteValidVec_res_56};
  wire [1:0] v0WriteValidVec_lo_hi_7 = {v0WriteValidVec_res_59, v0WriteValidVec_res_58};
  wire [3:0] v0WriteValidVec_lo_7 = {v0WriteValidVec_lo_hi_7, v0WriteValidVec_lo_lo_7};
  wire [1:0] v0WriteValidVec_hi_lo_7 = {v0WriteValidVec_res_61, v0WriteValidVec_res_60};
  wire [1:0] v0WriteValidVec_hi_hi_7 = {v0WriteValidVec_res_63, v0WriteValidVec_res_62};
  wire [3:0] v0WriteValidVec_hi_7 = {v0WriteValidVec_hi_hi_7, v0WriteValidVec_hi_lo_7};
  wire [7:0] v0WriteValidVec_7 = {v0WriteValidVec_hi_7, v0WriteValidVec_lo_7};
  wire [7:0] v0WriteValidVec_lsuWriteSet_8 = lsuWriteV0_8_valid ? 8'h1 << lsuWriteV0_8_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_8 = v0WriteValidVec_v0WriteIssue_8 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_64;
  reg        v0WriteValidVec_res_65;
  reg        v0WriteValidVec_res_66;
  reg        v0WriteValidVec_res_67;
  reg        v0WriteValidVec_res_68;
  reg        v0WriteValidVec_res_69;
  reg        v0WriteValidVec_res_70;
  reg        v0WriteValidVec_res_71;
  wire [1:0] v0WriteValidVec_lo_lo_8 = {v0WriteValidVec_res_65, v0WriteValidVec_res_64};
  wire [1:0] v0WriteValidVec_lo_hi_8 = {v0WriteValidVec_res_67, v0WriteValidVec_res_66};
  wire [3:0] v0WriteValidVec_lo_8 = {v0WriteValidVec_lo_hi_8, v0WriteValidVec_lo_lo_8};
  wire [1:0] v0WriteValidVec_hi_lo_8 = {v0WriteValidVec_res_69, v0WriteValidVec_res_68};
  wire [1:0] v0WriteValidVec_hi_hi_8 = {v0WriteValidVec_res_71, v0WriteValidVec_res_70};
  wire [3:0] v0WriteValidVec_hi_8 = {v0WriteValidVec_hi_hi_8, v0WriteValidVec_hi_lo_8};
  wire [7:0] v0WriteValidVec_8 = {v0WriteValidVec_hi_8, v0WriteValidVec_lo_8};
  wire [7:0] v0WriteValidVec_lsuWriteSet_9 = lsuWriteV0_9_valid ? 8'h1 << lsuWriteV0_9_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_9 = v0WriteValidVec_v0WriteIssue_9 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_72;
  reg        v0WriteValidVec_res_73;
  reg        v0WriteValidVec_res_74;
  reg        v0WriteValidVec_res_75;
  reg        v0WriteValidVec_res_76;
  reg        v0WriteValidVec_res_77;
  reg        v0WriteValidVec_res_78;
  reg        v0WriteValidVec_res_79;
  wire [1:0] v0WriteValidVec_lo_lo_9 = {v0WriteValidVec_res_73, v0WriteValidVec_res_72};
  wire [1:0] v0WriteValidVec_lo_hi_9 = {v0WriteValidVec_res_75, v0WriteValidVec_res_74};
  wire [3:0] v0WriteValidVec_lo_9 = {v0WriteValidVec_lo_hi_9, v0WriteValidVec_lo_lo_9};
  wire [1:0] v0WriteValidVec_hi_lo_9 = {v0WriteValidVec_res_77, v0WriteValidVec_res_76};
  wire [1:0] v0WriteValidVec_hi_hi_9 = {v0WriteValidVec_res_79, v0WriteValidVec_res_78};
  wire [3:0] v0WriteValidVec_hi_9 = {v0WriteValidVec_hi_hi_9, v0WriteValidVec_hi_lo_9};
  wire [7:0] v0WriteValidVec_9 = {v0WriteValidVec_hi_9, v0WriteValidVec_lo_9};
  wire [7:0] v0WriteValidVec_lsuWriteSet_10 = lsuWriteV0_10_valid ? 8'h1 << lsuWriteV0_10_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_10 = v0WriteValidVec_v0WriteIssue_10 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_80;
  reg        v0WriteValidVec_res_81;
  reg        v0WriteValidVec_res_82;
  reg        v0WriteValidVec_res_83;
  reg        v0WriteValidVec_res_84;
  reg        v0WriteValidVec_res_85;
  reg        v0WriteValidVec_res_86;
  reg        v0WriteValidVec_res_87;
  wire [1:0] v0WriteValidVec_lo_lo_10 = {v0WriteValidVec_res_81, v0WriteValidVec_res_80};
  wire [1:0] v0WriteValidVec_lo_hi_10 = {v0WriteValidVec_res_83, v0WriteValidVec_res_82};
  wire [3:0] v0WriteValidVec_lo_10 = {v0WriteValidVec_lo_hi_10, v0WriteValidVec_lo_lo_10};
  wire [1:0] v0WriteValidVec_hi_lo_10 = {v0WriteValidVec_res_85, v0WriteValidVec_res_84};
  wire [1:0] v0WriteValidVec_hi_hi_10 = {v0WriteValidVec_res_87, v0WriteValidVec_res_86};
  wire [3:0] v0WriteValidVec_hi_10 = {v0WriteValidVec_hi_hi_10, v0WriteValidVec_hi_lo_10};
  wire [7:0] v0WriteValidVec_10 = {v0WriteValidVec_hi_10, v0WriteValidVec_lo_10};
  wire [7:0] v0WriteValidVec_lsuWriteSet_11 = lsuWriteV0_11_valid ? 8'h1 << lsuWriteV0_11_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_11 = v0WriteValidVec_v0WriteIssue_11 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_88;
  reg        v0WriteValidVec_res_89;
  reg        v0WriteValidVec_res_90;
  reg        v0WriteValidVec_res_91;
  reg        v0WriteValidVec_res_92;
  reg        v0WriteValidVec_res_93;
  reg        v0WriteValidVec_res_94;
  reg        v0WriteValidVec_res_95;
  wire [1:0] v0WriteValidVec_lo_lo_11 = {v0WriteValidVec_res_89, v0WriteValidVec_res_88};
  wire [1:0] v0WriteValidVec_lo_hi_11 = {v0WriteValidVec_res_91, v0WriteValidVec_res_90};
  wire [3:0] v0WriteValidVec_lo_11 = {v0WriteValidVec_lo_hi_11, v0WriteValidVec_lo_lo_11};
  wire [1:0] v0WriteValidVec_hi_lo_11 = {v0WriteValidVec_res_93, v0WriteValidVec_res_92};
  wire [1:0] v0WriteValidVec_hi_hi_11 = {v0WriteValidVec_res_95, v0WriteValidVec_res_94};
  wire [3:0] v0WriteValidVec_hi_11 = {v0WriteValidVec_hi_hi_11, v0WriteValidVec_hi_lo_11};
  wire [7:0] v0WriteValidVec_11 = {v0WriteValidVec_hi_11, v0WriteValidVec_lo_11};
  wire [7:0] v0WriteValidVec_lsuWriteSet_12 = lsuWriteV0_12_valid ? 8'h1 << lsuWriteV0_12_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_12 = v0WriteValidVec_v0WriteIssue_12 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_96;
  reg        v0WriteValidVec_res_97;
  reg        v0WriteValidVec_res_98;
  reg        v0WriteValidVec_res_99;
  reg        v0WriteValidVec_res_100;
  reg        v0WriteValidVec_res_101;
  reg        v0WriteValidVec_res_102;
  reg        v0WriteValidVec_res_103;
  wire [1:0] v0WriteValidVec_lo_lo_12 = {v0WriteValidVec_res_97, v0WriteValidVec_res_96};
  wire [1:0] v0WriteValidVec_lo_hi_12 = {v0WriteValidVec_res_99, v0WriteValidVec_res_98};
  wire [3:0] v0WriteValidVec_lo_12 = {v0WriteValidVec_lo_hi_12, v0WriteValidVec_lo_lo_12};
  wire [1:0] v0WriteValidVec_hi_lo_12 = {v0WriteValidVec_res_101, v0WriteValidVec_res_100};
  wire [1:0] v0WriteValidVec_hi_hi_12 = {v0WriteValidVec_res_103, v0WriteValidVec_res_102};
  wire [3:0] v0WriteValidVec_hi_12 = {v0WriteValidVec_hi_hi_12, v0WriteValidVec_hi_lo_12};
  wire [7:0] v0WriteValidVec_12 = {v0WriteValidVec_hi_12, v0WriteValidVec_lo_12};
  wire [7:0] v0WriteValidVec_lsuWriteSet_13 = lsuWriteV0_13_valid ? 8'h1 << lsuWriteV0_13_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_13 = v0WriteValidVec_v0WriteIssue_13 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_104;
  reg        v0WriteValidVec_res_105;
  reg        v0WriteValidVec_res_106;
  reg        v0WriteValidVec_res_107;
  reg        v0WriteValidVec_res_108;
  reg        v0WriteValidVec_res_109;
  reg        v0WriteValidVec_res_110;
  reg        v0WriteValidVec_res_111;
  wire [1:0] v0WriteValidVec_lo_lo_13 = {v0WriteValidVec_res_105, v0WriteValidVec_res_104};
  wire [1:0] v0WriteValidVec_lo_hi_13 = {v0WriteValidVec_res_107, v0WriteValidVec_res_106};
  wire [3:0] v0WriteValidVec_lo_13 = {v0WriteValidVec_lo_hi_13, v0WriteValidVec_lo_lo_13};
  wire [1:0] v0WriteValidVec_hi_lo_13 = {v0WriteValidVec_res_109, v0WriteValidVec_res_108};
  wire [1:0] v0WriteValidVec_hi_hi_13 = {v0WriteValidVec_res_111, v0WriteValidVec_res_110};
  wire [3:0] v0WriteValidVec_hi_13 = {v0WriteValidVec_hi_hi_13, v0WriteValidVec_hi_lo_13};
  wire [7:0] v0WriteValidVec_13 = {v0WriteValidVec_hi_13, v0WriteValidVec_lo_13};
  wire [7:0] v0WriteValidVec_lsuWriteSet_14 = lsuWriteV0_14_valid ? 8'h1 << lsuWriteV0_14_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_14 = v0WriteValidVec_v0WriteIssue_14 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_112;
  reg        v0WriteValidVec_res_113;
  reg        v0WriteValidVec_res_114;
  reg        v0WriteValidVec_res_115;
  reg        v0WriteValidVec_res_116;
  reg        v0WriteValidVec_res_117;
  reg        v0WriteValidVec_res_118;
  reg        v0WriteValidVec_res_119;
  wire [1:0] v0WriteValidVec_lo_lo_14 = {v0WriteValidVec_res_113, v0WriteValidVec_res_112};
  wire [1:0] v0WriteValidVec_lo_hi_14 = {v0WriteValidVec_res_115, v0WriteValidVec_res_114};
  wire [3:0] v0WriteValidVec_lo_14 = {v0WriteValidVec_lo_hi_14, v0WriteValidVec_lo_lo_14};
  wire [1:0] v0WriteValidVec_hi_lo_14 = {v0WriteValidVec_res_117, v0WriteValidVec_res_116};
  wire [1:0] v0WriteValidVec_hi_hi_14 = {v0WriteValidVec_res_119, v0WriteValidVec_res_118};
  wire [3:0] v0WriteValidVec_hi_14 = {v0WriteValidVec_hi_hi_14, v0WriteValidVec_hi_lo_14};
  wire [7:0] v0WriteValidVec_14 = {v0WriteValidVec_hi_14, v0WriteValidVec_lo_14};
  wire [7:0] v0WriteValidVec_lsuWriteSet_15 = lsuWriteV0_15_valid ? 8'h1 << lsuWriteV0_15_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_15 = v0WriteValidVec_v0WriteIssue_15 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_120;
  reg        v0WriteValidVec_res_121;
  reg        v0WriteValidVec_res_122;
  reg        v0WriteValidVec_res_123;
  reg        v0WriteValidVec_res_124;
  reg        v0WriteValidVec_res_125;
  reg        v0WriteValidVec_res_126;
  reg        v0WriteValidVec_res_127;
  wire [1:0] v0WriteValidVec_lo_lo_15 = {v0WriteValidVec_res_121, v0WriteValidVec_res_120};
  wire [1:0] v0WriteValidVec_lo_hi_15 = {v0WriteValidVec_res_123, v0WriteValidVec_res_122};
  wire [3:0] v0WriteValidVec_lo_15 = {v0WriteValidVec_lo_hi_15, v0WriteValidVec_lo_lo_15};
  wire [1:0] v0WriteValidVec_hi_lo_15 = {v0WriteValidVec_res_125, v0WriteValidVec_res_124};
  wire [1:0] v0WriteValidVec_hi_hi_15 = {v0WriteValidVec_res_127, v0WriteValidVec_res_126};
  wire [3:0] v0WriteValidVec_hi_15 = {v0WriteValidVec_hi_hi_15, v0WriteValidVec_hi_lo_15};
  wire [7:0] v0WriteValidVec_15 = {v0WriteValidVec_hi_15, v0WriteValidVec_lo_15};
  wire [7:0] v0WriteValidVec_lsuWriteSet_16 = lsuWriteV0_16_valid ? 8'h1 << lsuWriteV0_16_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_16 = v0WriteValidVec_v0WriteIssue_16 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_128;
  reg        v0WriteValidVec_res_129;
  reg        v0WriteValidVec_res_130;
  reg        v0WriteValidVec_res_131;
  reg        v0WriteValidVec_res_132;
  reg        v0WriteValidVec_res_133;
  reg        v0WriteValidVec_res_134;
  reg        v0WriteValidVec_res_135;
  wire [1:0] v0WriteValidVec_lo_lo_16 = {v0WriteValidVec_res_129, v0WriteValidVec_res_128};
  wire [1:0] v0WriteValidVec_lo_hi_16 = {v0WriteValidVec_res_131, v0WriteValidVec_res_130};
  wire [3:0] v0WriteValidVec_lo_16 = {v0WriteValidVec_lo_hi_16, v0WriteValidVec_lo_lo_16};
  wire [1:0] v0WriteValidVec_hi_lo_16 = {v0WriteValidVec_res_133, v0WriteValidVec_res_132};
  wire [1:0] v0WriteValidVec_hi_hi_16 = {v0WriteValidVec_res_135, v0WriteValidVec_res_134};
  wire [3:0] v0WriteValidVec_hi_16 = {v0WriteValidVec_hi_hi_16, v0WriteValidVec_hi_lo_16};
  wire [7:0] v0WriteValidVec_16 = {v0WriteValidVec_hi_16, v0WriteValidVec_lo_16};
  wire [7:0] v0WriteValidVec_lsuWriteSet_17 = lsuWriteV0_17_valid ? 8'h1 << lsuWriteV0_17_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_17 = v0WriteValidVec_v0WriteIssue_17 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_136;
  reg        v0WriteValidVec_res_137;
  reg        v0WriteValidVec_res_138;
  reg        v0WriteValidVec_res_139;
  reg        v0WriteValidVec_res_140;
  reg        v0WriteValidVec_res_141;
  reg        v0WriteValidVec_res_142;
  reg        v0WriteValidVec_res_143;
  wire [1:0] v0WriteValidVec_lo_lo_17 = {v0WriteValidVec_res_137, v0WriteValidVec_res_136};
  wire [1:0] v0WriteValidVec_lo_hi_17 = {v0WriteValidVec_res_139, v0WriteValidVec_res_138};
  wire [3:0] v0WriteValidVec_lo_17 = {v0WriteValidVec_lo_hi_17, v0WriteValidVec_lo_lo_17};
  wire [1:0] v0WriteValidVec_hi_lo_17 = {v0WriteValidVec_res_141, v0WriteValidVec_res_140};
  wire [1:0] v0WriteValidVec_hi_hi_17 = {v0WriteValidVec_res_143, v0WriteValidVec_res_142};
  wire [3:0] v0WriteValidVec_hi_17 = {v0WriteValidVec_hi_hi_17, v0WriteValidVec_hi_lo_17};
  wire [7:0] v0WriteValidVec_17 = {v0WriteValidVec_hi_17, v0WriteValidVec_lo_17};
  wire [7:0] v0WriteValidVec_lsuWriteSet_18 = lsuWriteV0_18_valid ? 8'h1 << lsuWriteV0_18_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_18 = v0WriteValidVec_v0WriteIssue_18 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_144;
  reg        v0WriteValidVec_res_145;
  reg        v0WriteValidVec_res_146;
  reg        v0WriteValidVec_res_147;
  reg        v0WriteValidVec_res_148;
  reg        v0WriteValidVec_res_149;
  reg        v0WriteValidVec_res_150;
  reg        v0WriteValidVec_res_151;
  wire [1:0] v0WriteValidVec_lo_lo_18 = {v0WriteValidVec_res_145, v0WriteValidVec_res_144};
  wire [1:0] v0WriteValidVec_lo_hi_18 = {v0WriteValidVec_res_147, v0WriteValidVec_res_146};
  wire [3:0] v0WriteValidVec_lo_18 = {v0WriteValidVec_lo_hi_18, v0WriteValidVec_lo_lo_18};
  wire [1:0] v0WriteValidVec_hi_lo_18 = {v0WriteValidVec_res_149, v0WriteValidVec_res_148};
  wire [1:0] v0WriteValidVec_hi_hi_18 = {v0WriteValidVec_res_151, v0WriteValidVec_res_150};
  wire [3:0] v0WriteValidVec_hi_18 = {v0WriteValidVec_hi_hi_18, v0WriteValidVec_hi_lo_18};
  wire [7:0] v0WriteValidVec_18 = {v0WriteValidVec_hi_18, v0WriteValidVec_lo_18};
  wire [7:0] v0WriteValidVec_lsuWriteSet_19 = lsuWriteV0_19_valid ? 8'h1 << lsuWriteV0_19_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_19 = v0WriteValidVec_v0WriteIssue_19 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_152;
  reg        v0WriteValidVec_res_153;
  reg        v0WriteValidVec_res_154;
  reg        v0WriteValidVec_res_155;
  reg        v0WriteValidVec_res_156;
  reg        v0WriteValidVec_res_157;
  reg        v0WriteValidVec_res_158;
  reg        v0WriteValidVec_res_159;
  wire [1:0] v0WriteValidVec_lo_lo_19 = {v0WriteValidVec_res_153, v0WriteValidVec_res_152};
  wire [1:0] v0WriteValidVec_lo_hi_19 = {v0WriteValidVec_res_155, v0WriteValidVec_res_154};
  wire [3:0] v0WriteValidVec_lo_19 = {v0WriteValidVec_lo_hi_19, v0WriteValidVec_lo_lo_19};
  wire [1:0] v0WriteValidVec_hi_lo_19 = {v0WriteValidVec_res_157, v0WriteValidVec_res_156};
  wire [1:0] v0WriteValidVec_hi_hi_19 = {v0WriteValidVec_res_159, v0WriteValidVec_res_158};
  wire [3:0] v0WriteValidVec_hi_19 = {v0WriteValidVec_hi_hi_19, v0WriteValidVec_hi_lo_19};
  wire [7:0] v0WriteValidVec_19 = {v0WriteValidVec_hi_19, v0WriteValidVec_lo_19};
  wire [7:0] v0WriteValidVec_lsuWriteSet_20 = lsuWriteV0_20_valid ? 8'h1 << lsuWriteV0_20_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_20 = v0WriteValidVec_v0WriteIssue_20 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_160;
  reg        v0WriteValidVec_res_161;
  reg        v0WriteValidVec_res_162;
  reg        v0WriteValidVec_res_163;
  reg        v0WriteValidVec_res_164;
  reg        v0WriteValidVec_res_165;
  reg        v0WriteValidVec_res_166;
  reg        v0WriteValidVec_res_167;
  wire [1:0] v0WriteValidVec_lo_lo_20 = {v0WriteValidVec_res_161, v0WriteValidVec_res_160};
  wire [1:0] v0WriteValidVec_lo_hi_20 = {v0WriteValidVec_res_163, v0WriteValidVec_res_162};
  wire [3:0] v0WriteValidVec_lo_20 = {v0WriteValidVec_lo_hi_20, v0WriteValidVec_lo_lo_20};
  wire [1:0] v0WriteValidVec_hi_lo_20 = {v0WriteValidVec_res_165, v0WriteValidVec_res_164};
  wire [1:0] v0WriteValidVec_hi_hi_20 = {v0WriteValidVec_res_167, v0WriteValidVec_res_166};
  wire [3:0] v0WriteValidVec_hi_20 = {v0WriteValidVec_hi_hi_20, v0WriteValidVec_hi_lo_20};
  wire [7:0] v0WriteValidVec_20 = {v0WriteValidVec_hi_20, v0WriteValidVec_lo_20};
  wire [7:0] v0WriteValidVec_lsuWriteSet_21 = lsuWriteV0_21_valid ? 8'h1 << lsuWriteV0_21_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_21 = v0WriteValidVec_v0WriteIssue_21 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_168;
  reg        v0WriteValidVec_res_169;
  reg        v0WriteValidVec_res_170;
  reg        v0WriteValidVec_res_171;
  reg        v0WriteValidVec_res_172;
  reg        v0WriteValidVec_res_173;
  reg        v0WriteValidVec_res_174;
  reg        v0WriteValidVec_res_175;
  wire [1:0] v0WriteValidVec_lo_lo_21 = {v0WriteValidVec_res_169, v0WriteValidVec_res_168};
  wire [1:0] v0WriteValidVec_lo_hi_21 = {v0WriteValidVec_res_171, v0WriteValidVec_res_170};
  wire [3:0] v0WriteValidVec_lo_21 = {v0WriteValidVec_lo_hi_21, v0WriteValidVec_lo_lo_21};
  wire [1:0] v0WriteValidVec_hi_lo_21 = {v0WriteValidVec_res_173, v0WriteValidVec_res_172};
  wire [1:0] v0WriteValidVec_hi_hi_21 = {v0WriteValidVec_res_175, v0WriteValidVec_res_174};
  wire [3:0] v0WriteValidVec_hi_21 = {v0WriteValidVec_hi_hi_21, v0WriteValidVec_hi_lo_21};
  wire [7:0] v0WriteValidVec_21 = {v0WriteValidVec_hi_21, v0WriteValidVec_lo_21};
  wire [7:0] v0WriteValidVec_lsuWriteSet_22 = lsuWriteV0_22_valid ? 8'h1 << lsuWriteV0_22_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_22 = v0WriteValidVec_v0WriteIssue_22 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_176;
  reg        v0WriteValidVec_res_177;
  reg        v0WriteValidVec_res_178;
  reg        v0WriteValidVec_res_179;
  reg        v0WriteValidVec_res_180;
  reg        v0WriteValidVec_res_181;
  reg        v0WriteValidVec_res_182;
  reg        v0WriteValidVec_res_183;
  wire [1:0] v0WriteValidVec_lo_lo_22 = {v0WriteValidVec_res_177, v0WriteValidVec_res_176};
  wire [1:0] v0WriteValidVec_lo_hi_22 = {v0WriteValidVec_res_179, v0WriteValidVec_res_178};
  wire [3:0] v0WriteValidVec_lo_22 = {v0WriteValidVec_lo_hi_22, v0WriteValidVec_lo_lo_22};
  wire [1:0] v0WriteValidVec_hi_lo_22 = {v0WriteValidVec_res_181, v0WriteValidVec_res_180};
  wire [1:0] v0WriteValidVec_hi_hi_22 = {v0WriteValidVec_res_183, v0WriteValidVec_res_182};
  wire [3:0] v0WriteValidVec_hi_22 = {v0WriteValidVec_hi_hi_22, v0WriteValidVec_hi_lo_22};
  wire [7:0] v0WriteValidVec_22 = {v0WriteValidVec_hi_22, v0WriteValidVec_lo_22};
  wire [7:0] v0WriteValidVec_lsuWriteSet_23 = lsuWriteV0_23_valid ? 8'h1 << lsuWriteV0_23_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_23 = v0WriteValidVec_v0WriteIssue_23 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_184;
  reg        v0WriteValidVec_res_185;
  reg        v0WriteValidVec_res_186;
  reg        v0WriteValidVec_res_187;
  reg        v0WriteValidVec_res_188;
  reg        v0WriteValidVec_res_189;
  reg        v0WriteValidVec_res_190;
  reg        v0WriteValidVec_res_191;
  wire [1:0] v0WriteValidVec_lo_lo_23 = {v0WriteValidVec_res_185, v0WriteValidVec_res_184};
  wire [1:0] v0WriteValidVec_lo_hi_23 = {v0WriteValidVec_res_187, v0WriteValidVec_res_186};
  wire [3:0] v0WriteValidVec_lo_23 = {v0WriteValidVec_lo_hi_23, v0WriteValidVec_lo_lo_23};
  wire [1:0] v0WriteValidVec_hi_lo_23 = {v0WriteValidVec_res_189, v0WriteValidVec_res_188};
  wire [1:0] v0WriteValidVec_hi_hi_23 = {v0WriteValidVec_res_191, v0WriteValidVec_res_190};
  wire [3:0] v0WriteValidVec_hi_23 = {v0WriteValidVec_hi_hi_23, v0WriteValidVec_hi_lo_23};
  wire [7:0] v0WriteValidVec_23 = {v0WriteValidVec_hi_23, v0WriteValidVec_lo_23};
  wire [7:0] v0WriteValidVec_lsuWriteSet_24 = lsuWriteV0_24_valid ? 8'h1 << lsuWriteV0_24_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_24 = v0WriteValidVec_v0WriteIssue_24 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_192;
  reg        v0WriteValidVec_res_193;
  reg        v0WriteValidVec_res_194;
  reg        v0WriteValidVec_res_195;
  reg        v0WriteValidVec_res_196;
  reg        v0WriteValidVec_res_197;
  reg        v0WriteValidVec_res_198;
  reg        v0WriteValidVec_res_199;
  wire [1:0] v0WriteValidVec_lo_lo_24 = {v0WriteValidVec_res_193, v0WriteValidVec_res_192};
  wire [1:0] v0WriteValidVec_lo_hi_24 = {v0WriteValidVec_res_195, v0WriteValidVec_res_194};
  wire [3:0] v0WriteValidVec_lo_24 = {v0WriteValidVec_lo_hi_24, v0WriteValidVec_lo_lo_24};
  wire [1:0] v0WriteValidVec_hi_lo_24 = {v0WriteValidVec_res_197, v0WriteValidVec_res_196};
  wire [1:0] v0WriteValidVec_hi_hi_24 = {v0WriteValidVec_res_199, v0WriteValidVec_res_198};
  wire [3:0] v0WriteValidVec_hi_24 = {v0WriteValidVec_hi_hi_24, v0WriteValidVec_hi_lo_24};
  wire [7:0] v0WriteValidVec_24 = {v0WriteValidVec_hi_24, v0WriteValidVec_lo_24};
  wire [7:0] v0WriteValidVec_lsuWriteSet_25 = lsuWriteV0_25_valid ? 8'h1 << lsuWriteV0_25_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_25 = v0WriteValidVec_v0WriteIssue_25 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_200;
  reg        v0WriteValidVec_res_201;
  reg        v0WriteValidVec_res_202;
  reg        v0WriteValidVec_res_203;
  reg        v0WriteValidVec_res_204;
  reg        v0WriteValidVec_res_205;
  reg        v0WriteValidVec_res_206;
  reg        v0WriteValidVec_res_207;
  wire [1:0] v0WriteValidVec_lo_lo_25 = {v0WriteValidVec_res_201, v0WriteValidVec_res_200};
  wire [1:0] v0WriteValidVec_lo_hi_25 = {v0WriteValidVec_res_203, v0WriteValidVec_res_202};
  wire [3:0] v0WriteValidVec_lo_25 = {v0WriteValidVec_lo_hi_25, v0WriteValidVec_lo_lo_25};
  wire [1:0] v0WriteValidVec_hi_lo_25 = {v0WriteValidVec_res_205, v0WriteValidVec_res_204};
  wire [1:0] v0WriteValidVec_hi_hi_25 = {v0WriteValidVec_res_207, v0WriteValidVec_res_206};
  wire [3:0] v0WriteValidVec_hi_25 = {v0WriteValidVec_hi_hi_25, v0WriteValidVec_hi_lo_25};
  wire [7:0] v0WriteValidVec_25 = {v0WriteValidVec_hi_25, v0WriteValidVec_lo_25};
  wire [7:0] v0WriteValidVec_lsuWriteSet_26 = lsuWriteV0_26_valid ? 8'h1 << lsuWriteV0_26_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_26 = v0WriteValidVec_v0WriteIssue_26 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_208;
  reg        v0WriteValidVec_res_209;
  reg        v0WriteValidVec_res_210;
  reg        v0WriteValidVec_res_211;
  reg        v0WriteValidVec_res_212;
  reg        v0WriteValidVec_res_213;
  reg        v0WriteValidVec_res_214;
  reg        v0WriteValidVec_res_215;
  wire [1:0] v0WriteValidVec_lo_lo_26 = {v0WriteValidVec_res_209, v0WriteValidVec_res_208};
  wire [1:0] v0WriteValidVec_lo_hi_26 = {v0WriteValidVec_res_211, v0WriteValidVec_res_210};
  wire [3:0] v0WriteValidVec_lo_26 = {v0WriteValidVec_lo_hi_26, v0WriteValidVec_lo_lo_26};
  wire [1:0] v0WriteValidVec_hi_lo_26 = {v0WriteValidVec_res_213, v0WriteValidVec_res_212};
  wire [1:0] v0WriteValidVec_hi_hi_26 = {v0WriteValidVec_res_215, v0WriteValidVec_res_214};
  wire [3:0] v0WriteValidVec_hi_26 = {v0WriteValidVec_hi_hi_26, v0WriteValidVec_hi_lo_26};
  wire [7:0] v0WriteValidVec_26 = {v0WriteValidVec_hi_26, v0WriteValidVec_lo_26};
  wire [7:0] v0WriteValidVec_lsuWriteSet_27 = lsuWriteV0_27_valid ? 8'h1 << lsuWriteV0_27_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_27 = v0WriteValidVec_v0WriteIssue_27 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_216;
  reg        v0WriteValidVec_res_217;
  reg        v0WriteValidVec_res_218;
  reg        v0WriteValidVec_res_219;
  reg        v0WriteValidVec_res_220;
  reg        v0WriteValidVec_res_221;
  reg        v0WriteValidVec_res_222;
  reg        v0WriteValidVec_res_223;
  wire [1:0] v0WriteValidVec_lo_lo_27 = {v0WriteValidVec_res_217, v0WriteValidVec_res_216};
  wire [1:0] v0WriteValidVec_lo_hi_27 = {v0WriteValidVec_res_219, v0WriteValidVec_res_218};
  wire [3:0] v0WriteValidVec_lo_27 = {v0WriteValidVec_lo_hi_27, v0WriteValidVec_lo_lo_27};
  wire [1:0] v0WriteValidVec_hi_lo_27 = {v0WriteValidVec_res_221, v0WriteValidVec_res_220};
  wire [1:0] v0WriteValidVec_hi_hi_27 = {v0WriteValidVec_res_223, v0WriteValidVec_res_222};
  wire [3:0] v0WriteValidVec_hi_27 = {v0WriteValidVec_hi_hi_27, v0WriteValidVec_hi_lo_27};
  wire [7:0] v0WriteValidVec_27 = {v0WriteValidVec_hi_27, v0WriteValidVec_lo_27};
  wire [7:0] v0WriteValidVec_lsuWriteSet_28 = lsuWriteV0_28_valid ? 8'h1 << lsuWriteV0_28_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_28 = v0WriteValidVec_v0WriteIssue_28 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_224;
  reg        v0WriteValidVec_res_225;
  reg        v0WriteValidVec_res_226;
  reg        v0WriteValidVec_res_227;
  reg        v0WriteValidVec_res_228;
  reg        v0WriteValidVec_res_229;
  reg        v0WriteValidVec_res_230;
  reg        v0WriteValidVec_res_231;
  wire [1:0] v0WriteValidVec_lo_lo_28 = {v0WriteValidVec_res_225, v0WriteValidVec_res_224};
  wire [1:0] v0WriteValidVec_lo_hi_28 = {v0WriteValidVec_res_227, v0WriteValidVec_res_226};
  wire [3:0] v0WriteValidVec_lo_28 = {v0WriteValidVec_lo_hi_28, v0WriteValidVec_lo_lo_28};
  wire [1:0] v0WriteValidVec_hi_lo_28 = {v0WriteValidVec_res_229, v0WriteValidVec_res_228};
  wire [1:0] v0WriteValidVec_hi_hi_28 = {v0WriteValidVec_res_231, v0WriteValidVec_res_230};
  wire [3:0] v0WriteValidVec_hi_28 = {v0WriteValidVec_hi_hi_28, v0WriteValidVec_hi_lo_28};
  wire [7:0] v0WriteValidVec_28 = {v0WriteValidVec_hi_28, v0WriteValidVec_lo_28};
  wire [7:0] v0WriteValidVec_lsuWriteSet_29 = lsuWriteV0_29_valid ? 8'h1 << lsuWriteV0_29_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_29 = v0WriteValidVec_v0WriteIssue_29 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_232;
  reg        v0WriteValidVec_res_233;
  reg        v0WriteValidVec_res_234;
  reg        v0WriteValidVec_res_235;
  reg        v0WriteValidVec_res_236;
  reg        v0WriteValidVec_res_237;
  reg        v0WriteValidVec_res_238;
  reg        v0WriteValidVec_res_239;
  wire [1:0] v0WriteValidVec_lo_lo_29 = {v0WriteValidVec_res_233, v0WriteValidVec_res_232};
  wire [1:0] v0WriteValidVec_lo_hi_29 = {v0WriteValidVec_res_235, v0WriteValidVec_res_234};
  wire [3:0] v0WriteValidVec_lo_29 = {v0WriteValidVec_lo_hi_29, v0WriteValidVec_lo_lo_29};
  wire [1:0] v0WriteValidVec_hi_lo_29 = {v0WriteValidVec_res_237, v0WriteValidVec_res_236};
  wire [1:0] v0WriteValidVec_hi_hi_29 = {v0WriteValidVec_res_239, v0WriteValidVec_res_238};
  wire [3:0] v0WriteValidVec_hi_29 = {v0WriteValidVec_hi_hi_29, v0WriteValidVec_hi_lo_29};
  wire [7:0] v0WriteValidVec_29 = {v0WriteValidVec_hi_29, v0WriteValidVec_lo_29};
  wire [7:0] v0WriteValidVec_lsuWriteSet_30 = lsuWriteV0_30_valid ? 8'h1 << lsuWriteV0_30_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_30 = v0WriteValidVec_v0WriteIssue_30 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_240;
  reg        v0WriteValidVec_res_241;
  reg        v0WriteValidVec_res_242;
  reg        v0WriteValidVec_res_243;
  reg        v0WriteValidVec_res_244;
  reg        v0WriteValidVec_res_245;
  reg        v0WriteValidVec_res_246;
  reg        v0WriteValidVec_res_247;
  wire [1:0] v0WriteValidVec_lo_lo_30 = {v0WriteValidVec_res_241, v0WriteValidVec_res_240};
  wire [1:0] v0WriteValidVec_lo_hi_30 = {v0WriteValidVec_res_243, v0WriteValidVec_res_242};
  wire [3:0] v0WriteValidVec_lo_30 = {v0WriteValidVec_lo_hi_30, v0WriteValidVec_lo_lo_30};
  wire [1:0] v0WriteValidVec_hi_lo_30 = {v0WriteValidVec_res_245, v0WriteValidVec_res_244};
  wire [1:0] v0WriteValidVec_hi_hi_30 = {v0WriteValidVec_res_247, v0WriteValidVec_res_246};
  wire [3:0] v0WriteValidVec_hi_30 = {v0WriteValidVec_hi_hi_30, v0WriteValidVec_hi_lo_30};
  wire [7:0] v0WriteValidVec_30 = {v0WriteValidVec_hi_30, v0WriteValidVec_lo_30};
  wire [7:0] v0WriteValidVec_lsuWriteSet_31 = lsuWriteV0_31_valid ? 8'h1 << lsuWriteV0_31_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_31 = v0WriteValidVec_v0WriteIssue_31 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_248;
  reg        v0WriteValidVec_res_249;
  reg        v0WriteValidVec_res_250;
  reg        v0WriteValidVec_res_251;
  reg        v0WriteValidVec_res_252;
  reg        v0WriteValidVec_res_253;
  reg        v0WriteValidVec_res_254;
  reg        v0WriteValidVec_res_255;
  wire [1:0] v0WriteValidVec_lo_lo_31 = {v0WriteValidVec_res_249, v0WriteValidVec_res_248};
  wire [1:0] v0WriteValidVec_lo_hi_31 = {v0WriteValidVec_res_251, v0WriteValidVec_res_250};
  wire [3:0] v0WriteValidVec_lo_31 = {v0WriteValidVec_lo_hi_31, v0WriteValidVec_lo_lo_31};
  wire [1:0] v0WriteValidVec_hi_lo_31 = {v0WriteValidVec_res_253, v0WriteValidVec_res_252};
  wire [1:0] v0WriteValidVec_hi_hi_31 = {v0WriteValidVec_res_255, v0WriteValidVec_res_254};
  wire [3:0] v0WriteValidVec_hi_31 = {v0WriteValidVec_hi_hi_31, v0WriteValidVec_hi_lo_31};
  wire [7:0] v0WriteValidVec_31 = {v0WriteValidVec_hi_31, v0WriteValidVec_lo_31};
  wire       _GEN_0 = instructionIssue_valid & instructionIssue_bits_useV0AsMask & instructionIssue_bits_toLane;
  wire       useV0AsMaskToken_useV0Issue;
  assign useV0AsMaskToken_useV0Issue = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_1;
  assign useV0AsMaskToken_useV0Issue_1 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_2;
  assign useV0AsMaskToken_useV0Issue_2 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_3;
  assign useV0AsMaskToken_useV0Issue_3 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_4;
  assign useV0AsMaskToken_useV0Issue_4 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_5;
  assign useV0AsMaskToken_useV0Issue_5 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_6;
  assign useV0AsMaskToken_useV0Issue_6 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_7;
  assign useV0AsMaskToken_useV0Issue_7 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_8;
  assign useV0AsMaskToken_useV0Issue_8 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_9;
  assign useV0AsMaskToken_useV0Issue_9 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_10;
  assign useV0AsMaskToken_useV0Issue_10 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_11;
  assign useV0AsMaskToken_useV0Issue_11 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_12;
  assign useV0AsMaskToken_useV0Issue_12 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_13;
  assign useV0AsMaskToken_useV0Issue_13 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_14;
  assign useV0AsMaskToken_useV0Issue_14 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_15;
  assign useV0AsMaskToken_useV0Issue_15 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_16;
  assign useV0AsMaskToken_useV0Issue_16 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_17;
  assign useV0AsMaskToken_useV0Issue_17 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_18;
  assign useV0AsMaskToken_useV0Issue_18 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_19;
  assign useV0AsMaskToken_useV0Issue_19 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_20;
  assign useV0AsMaskToken_useV0Issue_20 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_21;
  assign useV0AsMaskToken_useV0Issue_21 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_22;
  assign useV0AsMaskToken_useV0Issue_22 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_23;
  assign useV0AsMaskToken_useV0Issue_23 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_24;
  assign useV0AsMaskToken_useV0Issue_24 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_25;
  assign useV0AsMaskToken_useV0Issue_25 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_26;
  assign useV0AsMaskToken_useV0Issue_26 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_27;
  assign useV0AsMaskToken_useV0Issue_27 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_28;
  assign useV0AsMaskToken_useV0Issue_28 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_29;
  assign useV0AsMaskToken_useV0Issue_29 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_30;
  assign useV0AsMaskToken_useV0Issue_30 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_31;
  assign useV0AsMaskToken_useV0Issue_31 = _GEN_0;
  wire [7:0] useV0AsMaskToken_updateOH = useV0AsMaskToken_useV0Issue ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res;
  reg        useV0AsMaskToken_res_1;
  reg        useV0AsMaskToken_res_2;
  reg        useV0AsMaskToken_res_3;
  reg        useV0AsMaskToken_res_4;
  reg        useV0AsMaskToken_res_5;
  reg        useV0AsMaskToken_res_6;
  reg        useV0AsMaskToken_res_7;
  wire [1:0] useV0AsMaskToken_lo_lo = {useV0AsMaskToken_res_1, useV0AsMaskToken_res};
  wire [1:0] useV0AsMaskToken_lo_hi = {useV0AsMaskToken_res_3, useV0AsMaskToken_res_2};
  wire [3:0] useV0AsMaskToken_lo = {useV0AsMaskToken_lo_hi, useV0AsMaskToken_lo_lo};
  wire [1:0] useV0AsMaskToken_hi_lo = {useV0AsMaskToken_res_5, useV0AsMaskToken_res_4};
  wire [1:0] useV0AsMaskToken_hi_hi = {useV0AsMaskToken_res_7, useV0AsMaskToken_res_6};
  wire [3:0] useV0AsMaskToken_hi = {useV0AsMaskToken_hi_hi, useV0AsMaskToken_hi_lo};
  wire [7:0] useV0AsMaskToken_updateOH_1 = useV0AsMaskToken_useV0Issue_1 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_8;
  reg        useV0AsMaskToken_res_9;
  reg        useV0AsMaskToken_res_10;
  reg        useV0AsMaskToken_res_11;
  reg        useV0AsMaskToken_res_12;
  reg        useV0AsMaskToken_res_13;
  reg        useV0AsMaskToken_res_14;
  reg        useV0AsMaskToken_res_15;
  wire [1:0] useV0AsMaskToken_lo_lo_1 = {useV0AsMaskToken_res_9, useV0AsMaskToken_res_8};
  wire [1:0] useV0AsMaskToken_lo_hi_1 = {useV0AsMaskToken_res_11, useV0AsMaskToken_res_10};
  wire [3:0] useV0AsMaskToken_lo_1 = {useV0AsMaskToken_lo_hi_1, useV0AsMaskToken_lo_lo_1};
  wire [1:0] useV0AsMaskToken_hi_lo_1 = {useV0AsMaskToken_res_13, useV0AsMaskToken_res_12};
  wire [1:0] useV0AsMaskToken_hi_hi_1 = {useV0AsMaskToken_res_15, useV0AsMaskToken_res_14};
  wire [3:0] useV0AsMaskToken_hi_1 = {useV0AsMaskToken_hi_hi_1, useV0AsMaskToken_hi_lo_1};
  wire [7:0] useV0AsMaskToken_updateOH_2 = useV0AsMaskToken_useV0Issue_2 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_16;
  reg        useV0AsMaskToken_res_17;
  reg        useV0AsMaskToken_res_18;
  reg        useV0AsMaskToken_res_19;
  reg        useV0AsMaskToken_res_20;
  reg        useV0AsMaskToken_res_21;
  reg        useV0AsMaskToken_res_22;
  reg        useV0AsMaskToken_res_23;
  wire [1:0] useV0AsMaskToken_lo_lo_2 = {useV0AsMaskToken_res_17, useV0AsMaskToken_res_16};
  wire [1:0] useV0AsMaskToken_lo_hi_2 = {useV0AsMaskToken_res_19, useV0AsMaskToken_res_18};
  wire [3:0] useV0AsMaskToken_lo_2 = {useV0AsMaskToken_lo_hi_2, useV0AsMaskToken_lo_lo_2};
  wire [1:0] useV0AsMaskToken_hi_lo_2 = {useV0AsMaskToken_res_21, useV0AsMaskToken_res_20};
  wire [1:0] useV0AsMaskToken_hi_hi_2 = {useV0AsMaskToken_res_23, useV0AsMaskToken_res_22};
  wire [3:0] useV0AsMaskToken_hi_2 = {useV0AsMaskToken_hi_hi_2, useV0AsMaskToken_hi_lo_2};
  wire [7:0] useV0AsMaskToken_updateOH_3 = useV0AsMaskToken_useV0Issue_3 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_24;
  reg        useV0AsMaskToken_res_25;
  reg        useV0AsMaskToken_res_26;
  reg        useV0AsMaskToken_res_27;
  reg        useV0AsMaskToken_res_28;
  reg        useV0AsMaskToken_res_29;
  reg        useV0AsMaskToken_res_30;
  reg        useV0AsMaskToken_res_31;
  wire [1:0] useV0AsMaskToken_lo_lo_3 = {useV0AsMaskToken_res_25, useV0AsMaskToken_res_24};
  wire [1:0] useV0AsMaskToken_lo_hi_3 = {useV0AsMaskToken_res_27, useV0AsMaskToken_res_26};
  wire [3:0] useV0AsMaskToken_lo_3 = {useV0AsMaskToken_lo_hi_3, useV0AsMaskToken_lo_lo_3};
  wire [1:0] useV0AsMaskToken_hi_lo_3 = {useV0AsMaskToken_res_29, useV0AsMaskToken_res_28};
  wire [1:0] useV0AsMaskToken_hi_hi_3 = {useV0AsMaskToken_res_31, useV0AsMaskToken_res_30};
  wire [3:0] useV0AsMaskToken_hi_3 = {useV0AsMaskToken_hi_hi_3, useV0AsMaskToken_hi_lo_3};
  wire [7:0] useV0AsMaskToken_updateOH_4 = useV0AsMaskToken_useV0Issue_4 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_32;
  reg        useV0AsMaskToken_res_33;
  reg        useV0AsMaskToken_res_34;
  reg        useV0AsMaskToken_res_35;
  reg        useV0AsMaskToken_res_36;
  reg        useV0AsMaskToken_res_37;
  reg        useV0AsMaskToken_res_38;
  reg        useV0AsMaskToken_res_39;
  wire [1:0] useV0AsMaskToken_lo_lo_4 = {useV0AsMaskToken_res_33, useV0AsMaskToken_res_32};
  wire [1:0] useV0AsMaskToken_lo_hi_4 = {useV0AsMaskToken_res_35, useV0AsMaskToken_res_34};
  wire [3:0] useV0AsMaskToken_lo_4 = {useV0AsMaskToken_lo_hi_4, useV0AsMaskToken_lo_lo_4};
  wire [1:0] useV0AsMaskToken_hi_lo_4 = {useV0AsMaskToken_res_37, useV0AsMaskToken_res_36};
  wire [1:0] useV0AsMaskToken_hi_hi_4 = {useV0AsMaskToken_res_39, useV0AsMaskToken_res_38};
  wire [3:0] useV0AsMaskToken_hi_4 = {useV0AsMaskToken_hi_hi_4, useV0AsMaskToken_hi_lo_4};
  wire [7:0] useV0AsMaskToken_updateOH_5 = useV0AsMaskToken_useV0Issue_5 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_40;
  reg        useV0AsMaskToken_res_41;
  reg        useV0AsMaskToken_res_42;
  reg        useV0AsMaskToken_res_43;
  reg        useV0AsMaskToken_res_44;
  reg        useV0AsMaskToken_res_45;
  reg        useV0AsMaskToken_res_46;
  reg        useV0AsMaskToken_res_47;
  wire [1:0] useV0AsMaskToken_lo_lo_5 = {useV0AsMaskToken_res_41, useV0AsMaskToken_res_40};
  wire [1:0] useV0AsMaskToken_lo_hi_5 = {useV0AsMaskToken_res_43, useV0AsMaskToken_res_42};
  wire [3:0] useV0AsMaskToken_lo_5 = {useV0AsMaskToken_lo_hi_5, useV0AsMaskToken_lo_lo_5};
  wire [1:0] useV0AsMaskToken_hi_lo_5 = {useV0AsMaskToken_res_45, useV0AsMaskToken_res_44};
  wire [1:0] useV0AsMaskToken_hi_hi_5 = {useV0AsMaskToken_res_47, useV0AsMaskToken_res_46};
  wire [3:0] useV0AsMaskToken_hi_5 = {useV0AsMaskToken_hi_hi_5, useV0AsMaskToken_hi_lo_5};
  wire [7:0] useV0AsMaskToken_updateOH_6 = useV0AsMaskToken_useV0Issue_6 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_48;
  reg        useV0AsMaskToken_res_49;
  reg        useV0AsMaskToken_res_50;
  reg        useV0AsMaskToken_res_51;
  reg        useV0AsMaskToken_res_52;
  reg        useV0AsMaskToken_res_53;
  reg        useV0AsMaskToken_res_54;
  reg        useV0AsMaskToken_res_55;
  wire [1:0] useV0AsMaskToken_lo_lo_6 = {useV0AsMaskToken_res_49, useV0AsMaskToken_res_48};
  wire [1:0] useV0AsMaskToken_lo_hi_6 = {useV0AsMaskToken_res_51, useV0AsMaskToken_res_50};
  wire [3:0] useV0AsMaskToken_lo_6 = {useV0AsMaskToken_lo_hi_6, useV0AsMaskToken_lo_lo_6};
  wire [1:0] useV0AsMaskToken_hi_lo_6 = {useV0AsMaskToken_res_53, useV0AsMaskToken_res_52};
  wire [1:0] useV0AsMaskToken_hi_hi_6 = {useV0AsMaskToken_res_55, useV0AsMaskToken_res_54};
  wire [3:0] useV0AsMaskToken_hi_6 = {useV0AsMaskToken_hi_hi_6, useV0AsMaskToken_hi_lo_6};
  wire [7:0] useV0AsMaskToken_updateOH_7 = useV0AsMaskToken_useV0Issue_7 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_56;
  reg        useV0AsMaskToken_res_57;
  reg        useV0AsMaskToken_res_58;
  reg        useV0AsMaskToken_res_59;
  reg        useV0AsMaskToken_res_60;
  reg        useV0AsMaskToken_res_61;
  reg        useV0AsMaskToken_res_62;
  reg        useV0AsMaskToken_res_63;
  wire [1:0] useV0AsMaskToken_lo_lo_7 = {useV0AsMaskToken_res_57, useV0AsMaskToken_res_56};
  wire [1:0] useV0AsMaskToken_lo_hi_7 = {useV0AsMaskToken_res_59, useV0AsMaskToken_res_58};
  wire [3:0] useV0AsMaskToken_lo_7 = {useV0AsMaskToken_lo_hi_7, useV0AsMaskToken_lo_lo_7};
  wire [1:0] useV0AsMaskToken_hi_lo_7 = {useV0AsMaskToken_res_61, useV0AsMaskToken_res_60};
  wire [1:0] useV0AsMaskToken_hi_hi_7 = {useV0AsMaskToken_res_63, useV0AsMaskToken_res_62};
  wire [3:0] useV0AsMaskToken_hi_7 = {useV0AsMaskToken_hi_hi_7, useV0AsMaskToken_hi_lo_7};
  wire [7:0] useV0AsMaskToken_updateOH_8 = useV0AsMaskToken_useV0Issue_8 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_64;
  reg        useV0AsMaskToken_res_65;
  reg        useV0AsMaskToken_res_66;
  reg        useV0AsMaskToken_res_67;
  reg        useV0AsMaskToken_res_68;
  reg        useV0AsMaskToken_res_69;
  reg        useV0AsMaskToken_res_70;
  reg        useV0AsMaskToken_res_71;
  wire [1:0] useV0AsMaskToken_lo_lo_8 = {useV0AsMaskToken_res_65, useV0AsMaskToken_res_64};
  wire [1:0] useV0AsMaskToken_lo_hi_8 = {useV0AsMaskToken_res_67, useV0AsMaskToken_res_66};
  wire [3:0] useV0AsMaskToken_lo_8 = {useV0AsMaskToken_lo_hi_8, useV0AsMaskToken_lo_lo_8};
  wire [1:0] useV0AsMaskToken_hi_lo_8 = {useV0AsMaskToken_res_69, useV0AsMaskToken_res_68};
  wire [1:0] useV0AsMaskToken_hi_hi_8 = {useV0AsMaskToken_res_71, useV0AsMaskToken_res_70};
  wire [3:0] useV0AsMaskToken_hi_8 = {useV0AsMaskToken_hi_hi_8, useV0AsMaskToken_hi_lo_8};
  wire [7:0] useV0AsMaskToken_updateOH_9 = useV0AsMaskToken_useV0Issue_9 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_72;
  reg        useV0AsMaskToken_res_73;
  reg        useV0AsMaskToken_res_74;
  reg        useV0AsMaskToken_res_75;
  reg        useV0AsMaskToken_res_76;
  reg        useV0AsMaskToken_res_77;
  reg        useV0AsMaskToken_res_78;
  reg        useV0AsMaskToken_res_79;
  wire [1:0] useV0AsMaskToken_lo_lo_9 = {useV0AsMaskToken_res_73, useV0AsMaskToken_res_72};
  wire [1:0] useV0AsMaskToken_lo_hi_9 = {useV0AsMaskToken_res_75, useV0AsMaskToken_res_74};
  wire [3:0] useV0AsMaskToken_lo_9 = {useV0AsMaskToken_lo_hi_9, useV0AsMaskToken_lo_lo_9};
  wire [1:0] useV0AsMaskToken_hi_lo_9 = {useV0AsMaskToken_res_77, useV0AsMaskToken_res_76};
  wire [1:0] useV0AsMaskToken_hi_hi_9 = {useV0AsMaskToken_res_79, useV0AsMaskToken_res_78};
  wire [3:0] useV0AsMaskToken_hi_9 = {useV0AsMaskToken_hi_hi_9, useV0AsMaskToken_hi_lo_9};
  wire [7:0] useV0AsMaskToken_updateOH_10 = useV0AsMaskToken_useV0Issue_10 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_80;
  reg        useV0AsMaskToken_res_81;
  reg        useV0AsMaskToken_res_82;
  reg        useV0AsMaskToken_res_83;
  reg        useV0AsMaskToken_res_84;
  reg        useV0AsMaskToken_res_85;
  reg        useV0AsMaskToken_res_86;
  reg        useV0AsMaskToken_res_87;
  wire [1:0] useV0AsMaskToken_lo_lo_10 = {useV0AsMaskToken_res_81, useV0AsMaskToken_res_80};
  wire [1:0] useV0AsMaskToken_lo_hi_10 = {useV0AsMaskToken_res_83, useV0AsMaskToken_res_82};
  wire [3:0] useV0AsMaskToken_lo_10 = {useV0AsMaskToken_lo_hi_10, useV0AsMaskToken_lo_lo_10};
  wire [1:0] useV0AsMaskToken_hi_lo_10 = {useV0AsMaskToken_res_85, useV0AsMaskToken_res_84};
  wire [1:0] useV0AsMaskToken_hi_hi_10 = {useV0AsMaskToken_res_87, useV0AsMaskToken_res_86};
  wire [3:0] useV0AsMaskToken_hi_10 = {useV0AsMaskToken_hi_hi_10, useV0AsMaskToken_hi_lo_10};
  wire [7:0] useV0AsMaskToken_updateOH_11 = useV0AsMaskToken_useV0Issue_11 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_88;
  reg        useV0AsMaskToken_res_89;
  reg        useV0AsMaskToken_res_90;
  reg        useV0AsMaskToken_res_91;
  reg        useV0AsMaskToken_res_92;
  reg        useV0AsMaskToken_res_93;
  reg        useV0AsMaskToken_res_94;
  reg        useV0AsMaskToken_res_95;
  wire [1:0] useV0AsMaskToken_lo_lo_11 = {useV0AsMaskToken_res_89, useV0AsMaskToken_res_88};
  wire [1:0] useV0AsMaskToken_lo_hi_11 = {useV0AsMaskToken_res_91, useV0AsMaskToken_res_90};
  wire [3:0] useV0AsMaskToken_lo_11 = {useV0AsMaskToken_lo_hi_11, useV0AsMaskToken_lo_lo_11};
  wire [1:0] useV0AsMaskToken_hi_lo_11 = {useV0AsMaskToken_res_93, useV0AsMaskToken_res_92};
  wire [1:0] useV0AsMaskToken_hi_hi_11 = {useV0AsMaskToken_res_95, useV0AsMaskToken_res_94};
  wire [3:0] useV0AsMaskToken_hi_11 = {useV0AsMaskToken_hi_hi_11, useV0AsMaskToken_hi_lo_11};
  wire [7:0] useV0AsMaskToken_updateOH_12 = useV0AsMaskToken_useV0Issue_12 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_96;
  reg        useV0AsMaskToken_res_97;
  reg        useV0AsMaskToken_res_98;
  reg        useV0AsMaskToken_res_99;
  reg        useV0AsMaskToken_res_100;
  reg        useV0AsMaskToken_res_101;
  reg        useV0AsMaskToken_res_102;
  reg        useV0AsMaskToken_res_103;
  wire [1:0] useV0AsMaskToken_lo_lo_12 = {useV0AsMaskToken_res_97, useV0AsMaskToken_res_96};
  wire [1:0] useV0AsMaskToken_lo_hi_12 = {useV0AsMaskToken_res_99, useV0AsMaskToken_res_98};
  wire [3:0] useV0AsMaskToken_lo_12 = {useV0AsMaskToken_lo_hi_12, useV0AsMaskToken_lo_lo_12};
  wire [1:0] useV0AsMaskToken_hi_lo_12 = {useV0AsMaskToken_res_101, useV0AsMaskToken_res_100};
  wire [1:0] useV0AsMaskToken_hi_hi_12 = {useV0AsMaskToken_res_103, useV0AsMaskToken_res_102};
  wire [3:0] useV0AsMaskToken_hi_12 = {useV0AsMaskToken_hi_hi_12, useV0AsMaskToken_hi_lo_12};
  wire [7:0] useV0AsMaskToken_updateOH_13 = useV0AsMaskToken_useV0Issue_13 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_104;
  reg        useV0AsMaskToken_res_105;
  reg        useV0AsMaskToken_res_106;
  reg        useV0AsMaskToken_res_107;
  reg        useV0AsMaskToken_res_108;
  reg        useV0AsMaskToken_res_109;
  reg        useV0AsMaskToken_res_110;
  reg        useV0AsMaskToken_res_111;
  wire [1:0] useV0AsMaskToken_lo_lo_13 = {useV0AsMaskToken_res_105, useV0AsMaskToken_res_104};
  wire [1:0] useV0AsMaskToken_lo_hi_13 = {useV0AsMaskToken_res_107, useV0AsMaskToken_res_106};
  wire [3:0] useV0AsMaskToken_lo_13 = {useV0AsMaskToken_lo_hi_13, useV0AsMaskToken_lo_lo_13};
  wire [1:0] useV0AsMaskToken_hi_lo_13 = {useV0AsMaskToken_res_109, useV0AsMaskToken_res_108};
  wire [1:0] useV0AsMaskToken_hi_hi_13 = {useV0AsMaskToken_res_111, useV0AsMaskToken_res_110};
  wire [3:0] useV0AsMaskToken_hi_13 = {useV0AsMaskToken_hi_hi_13, useV0AsMaskToken_hi_lo_13};
  wire [7:0] useV0AsMaskToken_updateOH_14 = useV0AsMaskToken_useV0Issue_14 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_112;
  reg        useV0AsMaskToken_res_113;
  reg        useV0AsMaskToken_res_114;
  reg        useV0AsMaskToken_res_115;
  reg        useV0AsMaskToken_res_116;
  reg        useV0AsMaskToken_res_117;
  reg        useV0AsMaskToken_res_118;
  reg        useV0AsMaskToken_res_119;
  wire [1:0] useV0AsMaskToken_lo_lo_14 = {useV0AsMaskToken_res_113, useV0AsMaskToken_res_112};
  wire [1:0] useV0AsMaskToken_lo_hi_14 = {useV0AsMaskToken_res_115, useV0AsMaskToken_res_114};
  wire [3:0] useV0AsMaskToken_lo_14 = {useV0AsMaskToken_lo_hi_14, useV0AsMaskToken_lo_lo_14};
  wire [1:0] useV0AsMaskToken_hi_lo_14 = {useV0AsMaskToken_res_117, useV0AsMaskToken_res_116};
  wire [1:0] useV0AsMaskToken_hi_hi_14 = {useV0AsMaskToken_res_119, useV0AsMaskToken_res_118};
  wire [3:0] useV0AsMaskToken_hi_14 = {useV0AsMaskToken_hi_hi_14, useV0AsMaskToken_hi_lo_14};
  wire [7:0] useV0AsMaskToken_updateOH_15 = useV0AsMaskToken_useV0Issue_15 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_120;
  reg        useV0AsMaskToken_res_121;
  reg        useV0AsMaskToken_res_122;
  reg        useV0AsMaskToken_res_123;
  reg        useV0AsMaskToken_res_124;
  reg        useV0AsMaskToken_res_125;
  reg        useV0AsMaskToken_res_126;
  reg        useV0AsMaskToken_res_127;
  wire [1:0] useV0AsMaskToken_lo_lo_15 = {useV0AsMaskToken_res_121, useV0AsMaskToken_res_120};
  wire [1:0] useV0AsMaskToken_lo_hi_15 = {useV0AsMaskToken_res_123, useV0AsMaskToken_res_122};
  wire [3:0] useV0AsMaskToken_lo_15 = {useV0AsMaskToken_lo_hi_15, useV0AsMaskToken_lo_lo_15};
  wire [1:0] useV0AsMaskToken_hi_lo_15 = {useV0AsMaskToken_res_125, useV0AsMaskToken_res_124};
  wire [1:0] useV0AsMaskToken_hi_hi_15 = {useV0AsMaskToken_res_127, useV0AsMaskToken_res_126};
  wire [3:0] useV0AsMaskToken_hi_15 = {useV0AsMaskToken_hi_hi_15, useV0AsMaskToken_hi_lo_15};
  wire [7:0] useV0AsMaskToken_updateOH_16 = useV0AsMaskToken_useV0Issue_16 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_128;
  reg        useV0AsMaskToken_res_129;
  reg        useV0AsMaskToken_res_130;
  reg        useV0AsMaskToken_res_131;
  reg        useV0AsMaskToken_res_132;
  reg        useV0AsMaskToken_res_133;
  reg        useV0AsMaskToken_res_134;
  reg        useV0AsMaskToken_res_135;
  wire [1:0] useV0AsMaskToken_lo_lo_16 = {useV0AsMaskToken_res_129, useV0AsMaskToken_res_128};
  wire [1:0] useV0AsMaskToken_lo_hi_16 = {useV0AsMaskToken_res_131, useV0AsMaskToken_res_130};
  wire [3:0] useV0AsMaskToken_lo_16 = {useV0AsMaskToken_lo_hi_16, useV0AsMaskToken_lo_lo_16};
  wire [1:0] useV0AsMaskToken_hi_lo_16 = {useV0AsMaskToken_res_133, useV0AsMaskToken_res_132};
  wire [1:0] useV0AsMaskToken_hi_hi_16 = {useV0AsMaskToken_res_135, useV0AsMaskToken_res_134};
  wire [3:0] useV0AsMaskToken_hi_16 = {useV0AsMaskToken_hi_hi_16, useV0AsMaskToken_hi_lo_16};
  wire [7:0] useV0AsMaskToken_updateOH_17 = useV0AsMaskToken_useV0Issue_17 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_136;
  reg        useV0AsMaskToken_res_137;
  reg        useV0AsMaskToken_res_138;
  reg        useV0AsMaskToken_res_139;
  reg        useV0AsMaskToken_res_140;
  reg        useV0AsMaskToken_res_141;
  reg        useV0AsMaskToken_res_142;
  reg        useV0AsMaskToken_res_143;
  wire [1:0] useV0AsMaskToken_lo_lo_17 = {useV0AsMaskToken_res_137, useV0AsMaskToken_res_136};
  wire [1:0] useV0AsMaskToken_lo_hi_17 = {useV0AsMaskToken_res_139, useV0AsMaskToken_res_138};
  wire [3:0] useV0AsMaskToken_lo_17 = {useV0AsMaskToken_lo_hi_17, useV0AsMaskToken_lo_lo_17};
  wire [1:0] useV0AsMaskToken_hi_lo_17 = {useV0AsMaskToken_res_141, useV0AsMaskToken_res_140};
  wire [1:0] useV0AsMaskToken_hi_hi_17 = {useV0AsMaskToken_res_143, useV0AsMaskToken_res_142};
  wire [3:0] useV0AsMaskToken_hi_17 = {useV0AsMaskToken_hi_hi_17, useV0AsMaskToken_hi_lo_17};
  wire [7:0] useV0AsMaskToken_updateOH_18 = useV0AsMaskToken_useV0Issue_18 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_144;
  reg        useV0AsMaskToken_res_145;
  reg        useV0AsMaskToken_res_146;
  reg        useV0AsMaskToken_res_147;
  reg        useV0AsMaskToken_res_148;
  reg        useV0AsMaskToken_res_149;
  reg        useV0AsMaskToken_res_150;
  reg        useV0AsMaskToken_res_151;
  wire [1:0] useV0AsMaskToken_lo_lo_18 = {useV0AsMaskToken_res_145, useV0AsMaskToken_res_144};
  wire [1:0] useV0AsMaskToken_lo_hi_18 = {useV0AsMaskToken_res_147, useV0AsMaskToken_res_146};
  wire [3:0] useV0AsMaskToken_lo_18 = {useV0AsMaskToken_lo_hi_18, useV0AsMaskToken_lo_lo_18};
  wire [1:0] useV0AsMaskToken_hi_lo_18 = {useV0AsMaskToken_res_149, useV0AsMaskToken_res_148};
  wire [1:0] useV0AsMaskToken_hi_hi_18 = {useV0AsMaskToken_res_151, useV0AsMaskToken_res_150};
  wire [3:0] useV0AsMaskToken_hi_18 = {useV0AsMaskToken_hi_hi_18, useV0AsMaskToken_hi_lo_18};
  wire [7:0] useV0AsMaskToken_updateOH_19 = useV0AsMaskToken_useV0Issue_19 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_152;
  reg        useV0AsMaskToken_res_153;
  reg        useV0AsMaskToken_res_154;
  reg        useV0AsMaskToken_res_155;
  reg        useV0AsMaskToken_res_156;
  reg        useV0AsMaskToken_res_157;
  reg        useV0AsMaskToken_res_158;
  reg        useV0AsMaskToken_res_159;
  wire [1:0] useV0AsMaskToken_lo_lo_19 = {useV0AsMaskToken_res_153, useV0AsMaskToken_res_152};
  wire [1:0] useV0AsMaskToken_lo_hi_19 = {useV0AsMaskToken_res_155, useV0AsMaskToken_res_154};
  wire [3:0] useV0AsMaskToken_lo_19 = {useV0AsMaskToken_lo_hi_19, useV0AsMaskToken_lo_lo_19};
  wire [1:0] useV0AsMaskToken_hi_lo_19 = {useV0AsMaskToken_res_157, useV0AsMaskToken_res_156};
  wire [1:0] useV0AsMaskToken_hi_hi_19 = {useV0AsMaskToken_res_159, useV0AsMaskToken_res_158};
  wire [3:0] useV0AsMaskToken_hi_19 = {useV0AsMaskToken_hi_hi_19, useV0AsMaskToken_hi_lo_19};
  wire [7:0] useV0AsMaskToken_updateOH_20 = useV0AsMaskToken_useV0Issue_20 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_160;
  reg        useV0AsMaskToken_res_161;
  reg        useV0AsMaskToken_res_162;
  reg        useV0AsMaskToken_res_163;
  reg        useV0AsMaskToken_res_164;
  reg        useV0AsMaskToken_res_165;
  reg        useV0AsMaskToken_res_166;
  reg        useV0AsMaskToken_res_167;
  wire [1:0] useV0AsMaskToken_lo_lo_20 = {useV0AsMaskToken_res_161, useV0AsMaskToken_res_160};
  wire [1:0] useV0AsMaskToken_lo_hi_20 = {useV0AsMaskToken_res_163, useV0AsMaskToken_res_162};
  wire [3:0] useV0AsMaskToken_lo_20 = {useV0AsMaskToken_lo_hi_20, useV0AsMaskToken_lo_lo_20};
  wire [1:0] useV0AsMaskToken_hi_lo_20 = {useV0AsMaskToken_res_165, useV0AsMaskToken_res_164};
  wire [1:0] useV0AsMaskToken_hi_hi_20 = {useV0AsMaskToken_res_167, useV0AsMaskToken_res_166};
  wire [3:0] useV0AsMaskToken_hi_20 = {useV0AsMaskToken_hi_hi_20, useV0AsMaskToken_hi_lo_20};
  wire [7:0] useV0AsMaskToken_updateOH_21 = useV0AsMaskToken_useV0Issue_21 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_168;
  reg        useV0AsMaskToken_res_169;
  reg        useV0AsMaskToken_res_170;
  reg        useV0AsMaskToken_res_171;
  reg        useV0AsMaskToken_res_172;
  reg        useV0AsMaskToken_res_173;
  reg        useV0AsMaskToken_res_174;
  reg        useV0AsMaskToken_res_175;
  wire [1:0] useV0AsMaskToken_lo_lo_21 = {useV0AsMaskToken_res_169, useV0AsMaskToken_res_168};
  wire [1:0] useV0AsMaskToken_lo_hi_21 = {useV0AsMaskToken_res_171, useV0AsMaskToken_res_170};
  wire [3:0] useV0AsMaskToken_lo_21 = {useV0AsMaskToken_lo_hi_21, useV0AsMaskToken_lo_lo_21};
  wire [1:0] useV0AsMaskToken_hi_lo_21 = {useV0AsMaskToken_res_173, useV0AsMaskToken_res_172};
  wire [1:0] useV0AsMaskToken_hi_hi_21 = {useV0AsMaskToken_res_175, useV0AsMaskToken_res_174};
  wire [3:0] useV0AsMaskToken_hi_21 = {useV0AsMaskToken_hi_hi_21, useV0AsMaskToken_hi_lo_21};
  wire [7:0] useV0AsMaskToken_updateOH_22 = useV0AsMaskToken_useV0Issue_22 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_176;
  reg        useV0AsMaskToken_res_177;
  reg        useV0AsMaskToken_res_178;
  reg        useV0AsMaskToken_res_179;
  reg        useV0AsMaskToken_res_180;
  reg        useV0AsMaskToken_res_181;
  reg        useV0AsMaskToken_res_182;
  reg        useV0AsMaskToken_res_183;
  wire [1:0] useV0AsMaskToken_lo_lo_22 = {useV0AsMaskToken_res_177, useV0AsMaskToken_res_176};
  wire [1:0] useV0AsMaskToken_lo_hi_22 = {useV0AsMaskToken_res_179, useV0AsMaskToken_res_178};
  wire [3:0] useV0AsMaskToken_lo_22 = {useV0AsMaskToken_lo_hi_22, useV0AsMaskToken_lo_lo_22};
  wire [1:0] useV0AsMaskToken_hi_lo_22 = {useV0AsMaskToken_res_181, useV0AsMaskToken_res_180};
  wire [1:0] useV0AsMaskToken_hi_hi_22 = {useV0AsMaskToken_res_183, useV0AsMaskToken_res_182};
  wire [3:0] useV0AsMaskToken_hi_22 = {useV0AsMaskToken_hi_hi_22, useV0AsMaskToken_hi_lo_22};
  wire [7:0] useV0AsMaskToken_updateOH_23 = useV0AsMaskToken_useV0Issue_23 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_184;
  reg        useV0AsMaskToken_res_185;
  reg        useV0AsMaskToken_res_186;
  reg        useV0AsMaskToken_res_187;
  reg        useV0AsMaskToken_res_188;
  reg        useV0AsMaskToken_res_189;
  reg        useV0AsMaskToken_res_190;
  reg        useV0AsMaskToken_res_191;
  wire [1:0] useV0AsMaskToken_lo_lo_23 = {useV0AsMaskToken_res_185, useV0AsMaskToken_res_184};
  wire [1:0] useV0AsMaskToken_lo_hi_23 = {useV0AsMaskToken_res_187, useV0AsMaskToken_res_186};
  wire [3:0] useV0AsMaskToken_lo_23 = {useV0AsMaskToken_lo_hi_23, useV0AsMaskToken_lo_lo_23};
  wire [1:0] useV0AsMaskToken_hi_lo_23 = {useV0AsMaskToken_res_189, useV0AsMaskToken_res_188};
  wire [1:0] useV0AsMaskToken_hi_hi_23 = {useV0AsMaskToken_res_191, useV0AsMaskToken_res_190};
  wire [3:0] useV0AsMaskToken_hi_23 = {useV0AsMaskToken_hi_hi_23, useV0AsMaskToken_hi_lo_23};
  wire [7:0] useV0AsMaskToken_updateOH_24 = useV0AsMaskToken_useV0Issue_24 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_192;
  reg        useV0AsMaskToken_res_193;
  reg        useV0AsMaskToken_res_194;
  reg        useV0AsMaskToken_res_195;
  reg        useV0AsMaskToken_res_196;
  reg        useV0AsMaskToken_res_197;
  reg        useV0AsMaskToken_res_198;
  reg        useV0AsMaskToken_res_199;
  wire [1:0] useV0AsMaskToken_lo_lo_24 = {useV0AsMaskToken_res_193, useV0AsMaskToken_res_192};
  wire [1:0] useV0AsMaskToken_lo_hi_24 = {useV0AsMaskToken_res_195, useV0AsMaskToken_res_194};
  wire [3:0] useV0AsMaskToken_lo_24 = {useV0AsMaskToken_lo_hi_24, useV0AsMaskToken_lo_lo_24};
  wire [1:0] useV0AsMaskToken_hi_lo_24 = {useV0AsMaskToken_res_197, useV0AsMaskToken_res_196};
  wire [1:0] useV0AsMaskToken_hi_hi_24 = {useV0AsMaskToken_res_199, useV0AsMaskToken_res_198};
  wire [3:0] useV0AsMaskToken_hi_24 = {useV0AsMaskToken_hi_hi_24, useV0AsMaskToken_hi_lo_24};
  wire [7:0] useV0AsMaskToken_updateOH_25 = useV0AsMaskToken_useV0Issue_25 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_200;
  reg        useV0AsMaskToken_res_201;
  reg        useV0AsMaskToken_res_202;
  reg        useV0AsMaskToken_res_203;
  reg        useV0AsMaskToken_res_204;
  reg        useV0AsMaskToken_res_205;
  reg        useV0AsMaskToken_res_206;
  reg        useV0AsMaskToken_res_207;
  wire [1:0] useV0AsMaskToken_lo_lo_25 = {useV0AsMaskToken_res_201, useV0AsMaskToken_res_200};
  wire [1:0] useV0AsMaskToken_lo_hi_25 = {useV0AsMaskToken_res_203, useV0AsMaskToken_res_202};
  wire [3:0] useV0AsMaskToken_lo_25 = {useV0AsMaskToken_lo_hi_25, useV0AsMaskToken_lo_lo_25};
  wire [1:0] useV0AsMaskToken_hi_lo_25 = {useV0AsMaskToken_res_205, useV0AsMaskToken_res_204};
  wire [1:0] useV0AsMaskToken_hi_hi_25 = {useV0AsMaskToken_res_207, useV0AsMaskToken_res_206};
  wire [3:0] useV0AsMaskToken_hi_25 = {useV0AsMaskToken_hi_hi_25, useV0AsMaskToken_hi_lo_25};
  wire [7:0] useV0AsMaskToken_updateOH_26 = useV0AsMaskToken_useV0Issue_26 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_208;
  reg        useV0AsMaskToken_res_209;
  reg        useV0AsMaskToken_res_210;
  reg        useV0AsMaskToken_res_211;
  reg        useV0AsMaskToken_res_212;
  reg        useV0AsMaskToken_res_213;
  reg        useV0AsMaskToken_res_214;
  reg        useV0AsMaskToken_res_215;
  wire [1:0] useV0AsMaskToken_lo_lo_26 = {useV0AsMaskToken_res_209, useV0AsMaskToken_res_208};
  wire [1:0] useV0AsMaskToken_lo_hi_26 = {useV0AsMaskToken_res_211, useV0AsMaskToken_res_210};
  wire [3:0] useV0AsMaskToken_lo_26 = {useV0AsMaskToken_lo_hi_26, useV0AsMaskToken_lo_lo_26};
  wire [1:0] useV0AsMaskToken_hi_lo_26 = {useV0AsMaskToken_res_213, useV0AsMaskToken_res_212};
  wire [1:0] useV0AsMaskToken_hi_hi_26 = {useV0AsMaskToken_res_215, useV0AsMaskToken_res_214};
  wire [3:0] useV0AsMaskToken_hi_26 = {useV0AsMaskToken_hi_hi_26, useV0AsMaskToken_hi_lo_26};
  wire [7:0] useV0AsMaskToken_updateOH_27 = useV0AsMaskToken_useV0Issue_27 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_216;
  reg        useV0AsMaskToken_res_217;
  reg        useV0AsMaskToken_res_218;
  reg        useV0AsMaskToken_res_219;
  reg        useV0AsMaskToken_res_220;
  reg        useV0AsMaskToken_res_221;
  reg        useV0AsMaskToken_res_222;
  reg        useV0AsMaskToken_res_223;
  wire [1:0] useV0AsMaskToken_lo_lo_27 = {useV0AsMaskToken_res_217, useV0AsMaskToken_res_216};
  wire [1:0] useV0AsMaskToken_lo_hi_27 = {useV0AsMaskToken_res_219, useV0AsMaskToken_res_218};
  wire [3:0] useV0AsMaskToken_lo_27 = {useV0AsMaskToken_lo_hi_27, useV0AsMaskToken_lo_lo_27};
  wire [1:0] useV0AsMaskToken_hi_lo_27 = {useV0AsMaskToken_res_221, useV0AsMaskToken_res_220};
  wire [1:0] useV0AsMaskToken_hi_hi_27 = {useV0AsMaskToken_res_223, useV0AsMaskToken_res_222};
  wire [3:0] useV0AsMaskToken_hi_27 = {useV0AsMaskToken_hi_hi_27, useV0AsMaskToken_hi_lo_27};
  wire [7:0] useV0AsMaskToken_updateOH_28 = useV0AsMaskToken_useV0Issue_28 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_224;
  reg        useV0AsMaskToken_res_225;
  reg        useV0AsMaskToken_res_226;
  reg        useV0AsMaskToken_res_227;
  reg        useV0AsMaskToken_res_228;
  reg        useV0AsMaskToken_res_229;
  reg        useV0AsMaskToken_res_230;
  reg        useV0AsMaskToken_res_231;
  wire [1:0] useV0AsMaskToken_lo_lo_28 = {useV0AsMaskToken_res_225, useV0AsMaskToken_res_224};
  wire [1:0] useV0AsMaskToken_lo_hi_28 = {useV0AsMaskToken_res_227, useV0AsMaskToken_res_226};
  wire [3:0] useV0AsMaskToken_lo_28 = {useV0AsMaskToken_lo_hi_28, useV0AsMaskToken_lo_lo_28};
  wire [1:0] useV0AsMaskToken_hi_lo_28 = {useV0AsMaskToken_res_229, useV0AsMaskToken_res_228};
  wire [1:0] useV0AsMaskToken_hi_hi_28 = {useV0AsMaskToken_res_231, useV0AsMaskToken_res_230};
  wire [3:0] useV0AsMaskToken_hi_28 = {useV0AsMaskToken_hi_hi_28, useV0AsMaskToken_hi_lo_28};
  wire [7:0] useV0AsMaskToken_updateOH_29 = useV0AsMaskToken_useV0Issue_29 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_232;
  reg        useV0AsMaskToken_res_233;
  reg        useV0AsMaskToken_res_234;
  reg        useV0AsMaskToken_res_235;
  reg        useV0AsMaskToken_res_236;
  reg        useV0AsMaskToken_res_237;
  reg        useV0AsMaskToken_res_238;
  reg        useV0AsMaskToken_res_239;
  wire [1:0] useV0AsMaskToken_lo_lo_29 = {useV0AsMaskToken_res_233, useV0AsMaskToken_res_232};
  wire [1:0] useV0AsMaskToken_lo_hi_29 = {useV0AsMaskToken_res_235, useV0AsMaskToken_res_234};
  wire [3:0] useV0AsMaskToken_lo_29 = {useV0AsMaskToken_lo_hi_29, useV0AsMaskToken_lo_lo_29};
  wire [1:0] useV0AsMaskToken_hi_lo_29 = {useV0AsMaskToken_res_237, useV0AsMaskToken_res_236};
  wire [1:0] useV0AsMaskToken_hi_hi_29 = {useV0AsMaskToken_res_239, useV0AsMaskToken_res_238};
  wire [3:0] useV0AsMaskToken_hi_29 = {useV0AsMaskToken_hi_hi_29, useV0AsMaskToken_hi_lo_29};
  wire [7:0] useV0AsMaskToken_updateOH_30 = useV0AsMaskToken_useV0Issue_30 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_240;
  reg        useV0AsMaskToken_res_241;
  reg        useV0AsMaskToken_res_242;
  reg        useV0AsMaskToken_res_243;
  reg        useV0AsMaskToken_res_244;
  reg        useV0AsMaskToken_res_245;
  reg        useV0AsMaskToken_res_246;
  reg        useV0AsMaskToken_res_247;
  wire [1:0] useV0AsMaskToken_lo_lo_30 = {useV0AsMaskToken_res_241, useV0AsMaskToken_res_240};
  wire [1:0] useV0AsMaskToken_lo_hi_30 = {useV0AsMaskToken_res_243, useV0AsMaskToken_res_242};
  wire [3:0] useV0AsMaskToken_lo_30 = {useV0AsMaskToken_lo_hi_30, useV0AsMaskToken_lo_lo_30};
  wire [1:0] useV0AsMaskToken_hi_lo_30 = {useV0AsMaskToken_res_245, useV0AsMaskToken_res_244};
  wire [1:0] useV0AsMaskToken_hi_hi_30 = {useV0AsMaskToken_res_247, useV0AsMaskToken_res_246};
  wire [3:0] useV0AsMaskToken_hi_30 = {useV0AsMaskToken_hi_hi_30, useV0AsMaskToken_hi_lo_30};
  wire [7:0] useV0AsMaskToken_updateOH_31 = useV0AsMaskToken_useV0Issue_31 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_248;
  reg        useV0AsMaskToken_res_249;
  reg        useV0AsMaskToken_res_250;
  reg        useV0AsMaskToken_res_251;
  reg        useV0AsMaskToken_res_252;
  reg        useV0AsMaskToken_res_253;
  reg        useV0AsMaskToken_res_254;
  reg        useV0AsMaskToken_res_255;
  wire [1:0] useV0AsMaskToken_lo_lo_31 = {useV0AsMaskToken_res_249, useV0AsMaskToken_res_248};
  wire [1:0] useV0AsMaskToken_lo_hi_31 = {useV0AsMaskToken_res_251, useV0AsMaskToken_res_250};
  wire [3:0] useV0AsMaskToken_lo_31 = {useV0AsMaskToken_lo_hi_31, useV0AsMaskToken_lo_lo_31};
  wire [1:0] useV0AsMaskToken_hi_lo_31 = {useV0AsMaskToken_res_253, useV0AsMaskToken_res_252};
  wire [1:0] useV0AsMaskToken_hi_hi_31 = {useV0AsMaskToken_res_255, useV0AsMaskToken_res_254};
  wire [3:0] useV0AsMaskToken_hi_31 = {useV0AsMaskToken_hi_hi_31, useV0AsMaskToken_hi_lo_31};
  wire [7:0] useV0AsMaskToken =
    {useV0AsMaskToken_hi, useV0AsMaskToken_lo} | {useV0AsMaskToken_hi_1, useV0AsMaskToken_lo_1} | {useV0AsMaskToken_hi_2, useV0AsMaskToken_lo_2} | {useV0AsMaskToken_hi_3, useV0AsMaskToken_lo_3}
    | {useV0AsMaskToken_hi_4, useV0AsMaskToken_lo_4} | {useV0AsMaskToken_hi_5, useV0AsMaskToken_lo_5} | {useV0AsMaskToken_hi_6, useV0AsMaskToken_lo_6} | {useV0AsMaskToken_hi_7, useV0AsMaskToken_lo_7}
    | {useV0AsMaskToken_hi_8, useV0AsMaskToken_lo_8} | {useV0AsMaskToken_hi_9, useV0AsMaskToken_lo_9} | {useV0AsMaskToken_hi_10, useV0AsMaskToken_lo_10} | {useV0AsMaskToken_hi_11, useV0AsMaskToken_lo_11}
    | {useV0AsMaskToken_hi_12, useV0AsMaskToken_lo_12} | {useV0AsMaskToken_hi_13, useV0AsMaskToken_lo_13} | {useV0AsMaskToken_hi_14, useV0AsMaskToken_lo_14} | {useV0AsMaskToken_hi_15, useV0AsMaskToken_lo_15}
    | {useV0AsMaskToken_hi_16, useV0AsMaskToken_lo_16} | {useV0AsMaskToken_hi_17, useV0AsMaskToken_lo_17} | {useV0AsMaskToken_hi_18, useV0AsMaskToken_lo_18} | {useV0AsMaskToken_hi_19, useV0AsMaskToken_lo_19}
    | {useV0AsMaskToken_hi_20, useV0AsMaskToken_lo_20} | {useV0AsMaskToken_hi_21, useV0AsMaskToken_lo_21} | {useV0AsMaskToken_hi_22, useV0AsMaskToken_lo_22} | {useV0AsMaskToken_hi_23, useV0AsMaskToken_lo_23}
    | {useV0AsMaskToken_hi_24, useV0AsMaskToken_lo_24} | {useV0AsMaskToken_hi_25, useV0AsMaskToken_lo_25} | {useV0AsMaskToken_hi_26, useV0AsMaskToken_lo_26} | {useV0AsMaskToken_hi_27, useV0AsMaskToken_lo_27}
    | {useV0AsMaskToken_hi_28, useV0AsMaskToken_lo_28} | {useV0AsMaskToken_hi_29, useV0AsMaskToken_lo_29} | {useV0AsMaskToken_hi_30, useV0AsMaskToken_lo_30} | {useV0AsMaskToken_hi_31, useV0AsMaskToken_lo_31};
  wire       maskUnitWriteV0_set = _maskUnitWriteV0_set_T & instructionIssue_bits_toMask;
  reg        maskUnitWriteV0;
  wire [7:0] _v0WriteValid_output =
    v0WriteValidVec_0 | v0WriteValidVec_1 | v0WriteValidVec_2 | v0WriteValidVec_3 | v0WriteValidVec_4 | v0WriteValidVec_5 | v0WriteValidVec_6 | v0WriteValidVec_7 | v0WriteValidVec_8 | v0WriteValidVec_9 | v0WriteValidVec_10
    | v0WriteValidVec_11 | v0WriteValidVec_12 | v0WriteValidVec_13 | v0WriteValidVec_14 | v0WriteValidVec_15 | v0WriteValidVec_16 | v0WriteValidVec_17 | v0WriteValidVec_18 | v0WriteValidVec_19 | v0WriteValidVec_20 | v0WriteValidVec_21
    | v0WriteValidVec_22 | v0WriteValidVec_23 | v0WriteValidVec_24 | v0WriteValidVec_25 | v0WriteValidVec_26 | v0WriteValidVec_27 | v0WriteValidVec_28 | v0WriteValidVec_29 | v0WriteValidVec_30 | v0WriteValidVec_31;
  wire       v0Conflict = instructionIssue_bits_writeV0 & (|useV0AsMaskToken) | instructionIssue_bits_useV0AsMask & ((|_v0WriteValid_output) | maskUnitWriteV0);
  always @(posedge clock) begin
    if (reset) begin
      v0WriteValidVec_res <= 1'h0;
      v0WriteValidVec_res_1 <= 1'h0;
      v0WriteValidVec_res_2 <= 1'h0;
      v0WriteValidVec_res_3 <= 1'h0;
      v0WriteValidVec_res_4 <= 1'h0;
      v0WriteValidVec_res_5 <= 1'h0;
      v0WriteValidVec_res_6 <= 1'h0;
      v0WriteValidVec_res_7 <= 1'h0;
      v0WriteValidVec_res_8 <= 1'h0;
      v0WriteValidVec_res_9 <= 1'h0;
      v0WriteValidVec_res_10 <= 1'h0;
      v0WriteValidVec_res_11 <= 1'h0;
      v0WriteValidVec_res_12 <= 1'h0;
      v0WriteValidVec_res_13 <= 1'h0;
      v0WriteValidVec_res_14 <= 1'h0;
      v0WriteValidVec_res_15 <= 1'h0;
      v0WriteValidVec_res_16 <= 1'h0;
      v0WriteValidVec_res_17 <= 1'h0;
      v0WriteValidVec_res_18 <= 1'h0;
      v0WriteValidVec_res_19 <= 1'h0;
      v0WriteValidVec_res_20 <= 1'h0;
      v0WriteValidVec_res_21 <= 1'h0;
      v0WriteValidVec_res_22 <= 1'h0;
      v0WriteValidVec_res_23 <= 1'h0;
      v0WriteValidVec_res_24 <= 1'h0;
      v0WriteValidVec_res_25 <= 1'h0;
      v0WriteValidVec_res_26 <= 1'h0;
      v0WriteValidVec_res_27 <= 1'h0;
      v0WriteValidVec_res_28 <= 1'h0;
      v0WriteValidVec_res_29 <= 1'h0;
      v0WriteValidVec_res_30 <= 1'h0;
      v0WriteValidVec_res_31 <= 1'h0;
      v0WriteValidVec_res_32 <= 1'h0;
      v0WriteValidVec_res_33 <= 1'h0;
      v0WriteValidVec_res_34 <= 1'h0;
      v0WriteValidVec_res_35 <= 1'h0;
      v0WriteValidVec_res_36 <= 1'h0;
      v0WriteValidVec_res_37 <= 1'h0;
      v0WriteValidVec_res_38 <= 1'h0;
      v0WriteValidVec_res_39 <= 1'h0;
      v0WriteValidVec_res_40 <= 1'h0;
      v0WriteValidVec_res_41 <= 1'h0;
      v0WriteValidVec_res_42 <= 1'h0;
      v0WriteValidVec_res_43 <= 1'h0;
      v0WriteValidVec_res_44 <= 1'h0;
      v0WriteValidVec_res_45 <= 1'h0;
      v0WriteValidVec_res_46 <= 1'h0;
      v0WriteValidVec_res_47 <= 1'h0;
      v0WriteValidVec_res_48 <= 1'h0;
      v0WriteValidVec_res_49 <= 1'h0;
      v0WriteValidVec_res_50 <= 1'h0;
      v0WriteValidVec_res_51 <= 1'h0;
      v0WriteValidVec_res_52 <= 1'h0;
      v0WriteValidVec_res_53 <= 1'h0;
      v0WriteValidVec_res_54 <= 1'h0;
      v0WriteValidVec_res_55 <= 1'h0;
      v0WriteValidVec_res_56 <= 1'h0;
      v0WriteValidVec_res_57 <= 1'h0;
      v0WriteValidVec_res_58 <= 1'h0;
      v0WriteValidVec_res_59 <= 1'h0;
      v0WriteValidVec_res_60 <= 1'h0;
      v0WriteValidVec_res_61 <= 1'h0;
      v0WriteValidVec_res_62 <= 1'h0;
      v0WriteValidVec_res_63 <= 1'h0;
      v0WriteValidVec_res_64 <= 1'h0;
      v0WriteValidVec_res_65 <= 1'h0;
      v0WriteValidVec_res_66 <= 1'h0;
      v0WriteValidVec_res_67 <= 1'h0;
      v0WriteValidVec_res_68 <= 1'h0;
      v0WriteValidVec_res_69 <= 1'h0;
      v0WriteValidVec_res_70 <= 1'h0;
      v0WriteValidVec_res_71 <= 1'h0;
      v0WriteValidVec_res_72 <= 1'h0;
      v0WriteValidVec_res_73 <= 1'h0;
      v0WriteValidVec_res_74 <= 1'h0;
      v0WriteValidVec_res_75 <= 1'h0;
      v0WriteValidVec_res_76 <= 1'h0;
      v0WriteValidVec_res_77 <= 1'h0;
      v0WriteValidVec_res_78 <= 1'h0;
      v0WriteValidVec_res_79 <= 1'h0;
      v0WriteValidVec_res_80 <= 1'h0;
      v0WriteValidVec_res_81 <= 1'h0;
      v0WriteValidVec_res_82 <= 1'h0;
      v0WriteValidVec_res_83 <= 1'h0;
      v0WriteValidVec_res_84 <= 1'h0;
      v0WriteValidVec_res_85 <= 1'h0;
      v0WriteValidVec_res_86 <= 1'h0;
      v0WriteValidVec_res_87 <= 1'h0;
      v0WriteValidVec_res_88 <= 1'h0;
      v0WriteValidVec_res_89 <= 1'h0;
      v0WriteValidVec_res_90 <= 1'h0;
      v0WriteValidVec_res_91 <= 1'h0;
      v0WriteValidVec_res_92 <= 1'h0;
      v0WriteValidVec_res_93 <= 1'h0;
      v0WriteValidVec_res_94 <= 1'h0;
      v0WriteValidVec_res_95 <= 1'h0;
      v0WriteValidVec_res_96 <= 1'h0;
      v0WriteValidVec_res_97 <= 1'h0;
      v0WriteValidVec_res_98 <= 1'h0;
      v0WriteValidVec_res_99 <= 1'h0;
      v0WriteValidVec_res_100 <= 1'h0;
      v0WriteValidVec_res_101 <= 1'h0;
      v0WriteValidVec_res_102 <= 1'h0;
      v0WriteValidVec_res_103 <= 1'h0;
      v0WriteValidVec_res_104 <= 1'h0;
      v0WriteValidVec_res_105 <= 1'h0;
      v0WriteValidVec_res_106 <= 1'h0;
      v0WriteValidVec_res_107 <= 1'h0;
      v0WriteValidVec_res_108 <= 1'h0;
      v0WriteValidVec_res_109 <= 1'h0;
      v0WriteValidVec_res_110 <= 1'h0;
      v0WriteValidVec_res_111 <= 1'h0;
      v0WriteValidVec_res_112 <= 1'h0;
      v0WriteValidVec_res_113 <= 1'h0;
      v0WriteValidVec_res_114 <= 1'h0;
      v0WriteValidVec_res_115 <= 1'h0;
      v0WriteValidVec_res_116 <= 1'h0;
      v0WriteValidVec_res_117 <= 1'h0;
      v0WriteValidVec_res_118 <= 1'h0;
      v0WriteValidVec_res_119 <= 1'h0;
      v0WriteValidVec_res_120 <= 1'h0;
      v0WriteValidVec_res_121 <= 1'h0;
      v0WriteValidVec_res_122 <= 1'h0;
      v0WriteValidVec_res_123 <= 1'h0;
      v0WriteValidVec_res_124 <= 1'h0;
      v0WriteValidVec_res_125 <= 1'h0;
      v0WriteValidVec_res_126 <= 1'h0;
      v0WriteValidVec_res_127 <= 1'h0;
      v0WriteValidVec_res_128 <= 1'h0;
      v0WriteValidVec_res_129 <= 1'h0;
      v0WriteValidVec_res_130 <= 1'h0;
      v0WriteValidVec_res_131 <= 1'h0;
      v0WriteValidVec_res_132 <= 1'h0;
      v0WriteValidVec_res_133 <= 1'h0;
      v0WriteValidVec_res_134 <= 1'h0;
      v0WriteValidVec_res_135 <= 1'h0;
      v0WriteValidVec_res_136 <= 1'h0;
      v0WriteValidVec_res_137 <= 1'h0;
      v0WriteValidVec_res_138 <= 1'h0;
      v0WriteValidVec_res_139 <= 1'h0;
      v0WriteValidVec_res_140 <= 1'h0;
      v0WriteValidVec_res_141 <= 1'h0;
      v0WriteValidVec_res_142 <= 1'h0;
      v0WriteValidVec_res_143 <= 1'h0;
      v0WriteValidVec_res_144 <= 1'h0;
      v0WriteValidVec_res_145 <= 1'h0;
      v0WriteValidVec_res_146 <= 1'h0;
      v0WriteValidVec_res_147 <= 1'h0;
      v0WriteValidVec_res_148 <= 1'h0;
      v0WriteValidVec_res_149 <= 1'h0;
      v0WriteValidVec_res_150 <= 1'h0;
      v0WriteValidVec_res_151 <= 1'h0;
      v0WriteValidVec_res_152 <= 1'h0;
      v0WriteValidVec_res_153 <= 1'h0;
      v0WriteValidVec_res_154 <= 1'h0;
      v0WriteValidVec_res_155 <= 1'h0;
      v0WriteValidVec_res_156 <= 1'h0;
      v0WriteValidVec_res_157 <= 1'h0;
      v0WriteValidVec_res_158 <= 1'h0;
      v0WriteValidVec_res_159 <= 1'h0;
      v0WriteValidVec_res_160 <= 1'h0;
      v0WriteValidVec_res_161 <= 1'h0;
      v0WriteValidVec_res_162 <= 1'h0;
      v0WriteValidVec_res_163 <= 1'h0;
      v0WriteValidVec_res_164 <= 1'h0;
      v0WriteValidVec_res_165 <= 1'h0;
      v0WriteValidVec_res_166 <= 1'h0;
      v0WriteValidVec_res_167 <= 1'h0;
      v0WriteValidVec_res_168 <= 1'h0;
      v0WriteValidVec_res_169 <= 1'h0;
      v0WriteValidVec_res_170 <= 1'h0;
      v0WriteValidVec_res_171 <= 1'h0;
      v0WriteValidVec_res_172 <= 1'h0;
      v0WriteValidVec_res_173 <= 1'h0;
      v0WriteValidVec_res_174 <= 1'h0;
      v0WriteValidVec_res_175 <= 1'h0;
      v0WriteValidVec_res_176 <= 1'h0;
      v0WriteValidVec_res_177 <= 1'h0;
      v0WriteValidVec_res_178 <= 1'h0;
      v0WriteValidVec_res_179 <= 1'h0;
      v0WriteValidVec_res_180 <= 1'h0;
      v0WriteValidVec_res_181 <= 1'h0;
      v0WriteValidVec_res_182 <= 1'h0;
      v0WriteValidVec_res_183 <= 1'h0;
      v0WriteValidVec_res_184 <= 1'h0;
      v0WriteValidVec_res_185 <= 1'h0;
      v0WriteValidVec_res_186 <= 1'h0;
      v0WriteValidVec_res_187 <= 1'h0;
      v0WriteValidVec_res_188 <= 1'h0;
      v0WriteValidVec_res_189 <= 1'h0;
      v0WriteValidVec_res_190 <= 1'h0;
      v0WriteValidVec_res_191 <= 1'h0;
      v0WriteValidVec_res_192 <= 1'h0;
      v0WriteValidVec_res_193 <= 1'h0;
      v0WriteValidVec_res_194 <= 1'h0;
      v0WriteValidVec_res_195 <= 1'h0;
      v0WriteValidVec_res_196 <= 1'h0;
      v0WriteValidVec_res_197 <= 1'h0;
      v0WriteValidVec_res_198 <= 1'h0;
      v0WriteValidVec_res_199 <= 1'h0;
      v0WriteValidVec_res_200 <= 1'h0;
      v0WriteValidVec_res_201 <= 1'h0;
      v0WriteValidVec_res_202 <= 1'h0;
      v0WriteValidVec_res_203 <= 1'h0;
      v0WriteValidVec_res_204 <= 1'h0;
      v0WriteValidVec_res_205 <= 1'h0;
      v0WriteValidVec_res_206 <= 1'h0;
      v0WriteValidVec_res_207 <= 1'h0;
      v0WriteValidVec_res_208 <= 1'h0;
      v0WriteValidVec_res_209 <= 1'h0;
      v0WriteValidVec_res_210 <= 1'h0;
      v0WriteValidVec_res_211 <= 1'h0;
      v0WriteValidVec_res_212 <= 1'h0;
      v0WriteValidVec_res_213 <= 1'h0;
      v0WriteValidVec_res_214 <= 1'h0;
      v0WriteValidVec_res_215 <= 1'h0;
      v0WriteValidVec_res_216 <= 1'h0;
      v0WriteValidVec_res_217 <= 1'h0;
      v0WriteValidVec_res_218 <= 1'h0;
      v0WriteValidVec_res_219 <= 1'h0;
      v0WriteValidVec_res_220 <= 1'h0;
      v0WriteValidVec_res_221 <= 1'h0;
      v0WriteValidVec_res_222 <= 1'h0;
      v0WriteValidVec_res_223 <= 1'h0;
      v0WriteValidVec_res_224 <= 1'h0;
      v0WriteValidVec_res_225 <= 1'h0;
      v0WriteValidVec_res_226 <= 1'h0;
      v0WriteValidVec_res_227 <= 1'h0;
      v0WriteValidVec_res_228 <= 1'h0;
      v0WriteValidVec_res_229 <= 1'h0;
      v0WriteValidVec_res_230 <= 1'h0;
      v0WriteValidVec_res_231 <= 1'h0;
      v0WriteValidVec_res_232 <= 1'h0;
      v0WriteValidVec_res_233 <= 1'h0;
      v0WriteValidVec_res_234 <= 1'h0;
      v0WriteValidVec_res_235 <= 1'h0;
      v0WriteValidVec_res_236 <= 1'h0;
      v0WriteValidVec_res_237 <= 1'h0;
      v0WriteValidVec_res_238 <= 1'h0;
      v0WriteValidVec_res_239 <= 1'h0;
      v0WriteValidVec_res_240 <= 1'h0;
      v0WriteValidVec_res_241 <= 1'h0;
      v0WriteValidVec_res_242 <= 1'h0;
      v0WriteValidVec_res_243 <= 1'h0;
      v0WriteValidVec_res_244 <= 1'h0;
      v0WriteValidVec_res_245 <= 1'h0;
      v0WriteValidVec_res_246 <= 1'h0;
      v0WriteValidVec_res_247 <= 1'h0;
      v0WriteValidVec_res_248 <= 1'h0;
      v0WriteValidVec_res_249 <= 1'h0;
      v0WriteValidVec_res_250 <= 1'h0;
      v0WriteValidVec_res_251 <= 1'h0;
      v0WriteValidVec_res_252 <= 1'h0;
      v0WriteValidVec_res_253 <= 1'h0;
      v0WriteValidVec_res_254 <= 1'h0;
      v0WriteValidVec_res_255 <= 1'h0;
      useV0AsMaskToken_res <= 1'h0;
      useV0AsMaskToken_res_1 <= 1'h0;
      useV0AsMaskToken_res_2 <= 1'h0;
      useV0AsMaskToken_res_3 <= 1'h0;
      useV0AsMaskToken_res_4 <= 1'h0;
      useV0AsMaskToken_res_5 <= 1'h0;
      useV0AsMaskToken_res_6 <= 1'h0;
      useV0AsMaskToken_res_7 <= 1'h0;
      useV0AsMaskToken_res_8 <= 1'h0;
      useV0AsMaskToken_res_9 <= 1'h0;
      useV0AsMaskToken_res_10 <= 1'h0;
      useV0AsMaskToken_res_11 <= 1'h0;
      useV0AsMaskToken_res_12 <= 1'h0;
      useV0AsMaskToken_res_13 <= 1'h0;
      useV0AsMaskToken_res_14 <= 1'h0;
      useV0AsMaskToken_res_15 <= 1'h0;
      useV0AsMaskToken_res_16 <= 1'h0;
      useV0AsMaskToken_res_17 <= 1'h0;
      useV0AsMaskToken_res_18 <= 1'h0;
      useV0AsMaskToken_res_19 <= 1'h0;
      useV0AsMaskToken_res_20 <= 1'h0;
      useV0AsMaskToken_res_21 <= 1'h0;
      useV0AsMaskToken_res_22 <= 1'h0;
      useV0AsMaskToken_res_23 <= 1'h0;
      useV0AsMaskToken_res_24 <= 1'h0;
      useV0AsMaskToken_res_25 <= 1'h0;
      useV0AsMaskToken_res_26 <= 1'h0;
      useV0AsMaskToken_res_27 <= 1'h0;
      useV0AsMaskToken_res_28 <= 1'h0;
      useV0AsMaskToken_res_29 <= 1'h0;
      useV0AsMaskToken_res_30 <= 1'h0;
      useV0AsMaskToken_res_31 <= 1'h0;
      useV0AsMaskToken_res_32 <= 1'h0;
      useV0AsMaskToken_res_33 <= 1'h0;
      useV0AsMaskToken_res_34 <= 1'h0;
      useV0AsMaskToken_res_35 <= 1'h0;
      useV0AsMaskToken_res_36 <= 1'h0;
      useV0AsMaskToken_res_37 <= 1'h0;
      useV0AsMaskToken_res_38 <= 1'h0;
      useV0AsMaskToken_res_39 <= 1'h0;
      useV0AsMaskToken_res_40 <= 1'h0;
      useV0AsMaskToken_res_41 <= 1'h0;
      useV0AsMaskToken_res_42 <= 1'h0;
      useV0AsMaskToken_res_43 <= 1'h0;
      useV0AsMaskToken_res_44 <= 1'h0;
      useV0AsMaskToken_res_45 <= 1'h0;
      useV0AsMaskToken_res_46 <= 1'h0;
      useV0AsMaskToken_res_47 <= 1'h0;
      useV0AsMaskToken_res_48 <= 1'h0;
      useV0AsMaskToken_res_49 <= 1'h0;
      useV0AsMaskToken_res_50 <= 1'h0;
      useV0AsMaskToken_res_51 <= 1'h0;
      useV0AsMaskToken_res_52 <= 1'h0;
      useV0AsMaskToken_res_53 <= 1'h0;
      useV0AsMaskToken_res_54 <= 1'h0;
      useV0AsMaskToken_res_55 <= 1'h0;
      useV0AsMaskToken_res_56 <= 1'h0;
      useV0AsMaskToken_res_57 <= 1'h0;
      useV0AsMaskToken_res_58 <= 1'h0;
      useV0AsMaskToken_res_59 <= 1'h0;
      useV0AsMaskToken_res_60 <= 1'h0;
      useV0AsMaskToken_res_61 <= 1'h0;
      useV0AsMaskToken_res_62 <= 1'h0;
      useV0AsMaskToken_res_63 <= 1'h0;
      useV0AsMaskToken_res_64 <= 1'h0;
      useV0AsMaskToken_res_65 <= 1'h0;
      useV0AsMaskToken_res_66 <= 1'h0;
      useV0AsMaskToken_res_67 <= 1'h0;
      useV0AsMaskToken_res_68 <= 1'h0;
      useV0AsMaskToken_res_69 <= 1'h0;
      useV0AsMaskToken_res_70 <= 1'h0;
      useV0AsMaskToken_res_71 <= 1'h0;
      useV0AsMaskToken_res_72 <= 1'h0;
      useV0AsMaskToken_res_73 <= 1'h0;
      useV0AsMaskToken_res_74 <= 1'h0;
      useV0AsMaskToken_res_75 <= 1'h0;
      useV0AsMaskToken_res_76 <= 1'h0;
      useV0AsMaskToken_res_77 <= 1'h0;
      useV0AsMaskToken_res_78 <= 1'h0;
      useV0AsMaskToken_res_79 <= 1'h0;
      useV0AsMaskToken_res_80 <= 1'h0;
      useV0AsMaskToken_res_81 <= 1'h0;
      useV0AsMaskToken_res_82 <= 1'h0;
      useV0AsMaskToken_res_83 <= 1'h0;
      useV0AsMaskToken_res_84 <= 1'h0;
      useV0AsMaskToken_res_85 <= 1'h0;
      useV0AsMaskToken_res_86 <= 1'h0;
      useV0AsMaskToken_res_87 <= 1'h0;
      useV0AsMaskToken_res_88 <= 1'h0;
      useV0AsMaskToken_res_89 <= 1'h0;
      useV0AsMaskToken_res_90 <= 1'h0;
      useV0AsMaskToken_res_91 <= 1'h0;
      useV0AsMaskToken_res_92 <= 1'h0;
      useV0AsMaskToken_res_93 <= 1'h0;
      useV0AsMaskToken_res_94 <= 1'h0;
      useV0AsMaskToken_res_95 <= 1'h0;
      useV0AsMaskToken_res_96 <= 1'h0;
      useV0AsMaskToken_res_97 <= 1'h0;
      useV0AsMaskToken_res_98 <= 1'h0;
      useV0AsMaskToken_res_99 <= 1'h0;
      useV0AsMaskToken_res_100 <= 1'h0;
      useV0AsMaskToken_res_101 <= 1'h0;
      useV0AsMaskToken_res_102 <= 1'h0;
      useV0AsMaskToken_res_103 <= 1'h0;
      useV0AsMaskToken_res_104 <= 1'h0;
      useV0AsMaskToken_res_105 <= 1'h0;
      useV0AsMaskToken_res_106 <= 1'h0;
      useV0AsMaskToken_res_107 <= 1'h0;
      useV0AsMaskToken_res_108 <= 1'h0;
      useV0AsMaskToken_res_109 <= 1'h0;
      useV0AsMaskToken_res_110 <= 1'h0;
      useV0AsMaskToken_res_111 <= 1'h0;
      useV0AsMaskToken_res_112 <= 1'h0;
      useV0AsMaskToken_res_113 <= 1'h0;
      useV0AsMaskToken_res_114 <= 1'h0;
      useV0AsMaskToken_res_115 <= 1'h0;
      useV0AsMaskToken_res_116 <= 1'h0;
      useV0AsMaskToken_res_117 <= 1'h0;
      useV0AsMaskToken_res_118 <= 1'h0;
      useV0AsMaskToken_res_119 <= 1'h0;
      useV0AsMaskToken_res_120 <= 1'h0;
      useV0AsMaskToken_res_121 <= 1'h0;
      useV0AsMaskToken_res_122 <= 1'h0;
      useV0AsMaskToken_res_123 <= 1'h0;
      useV0AsMaskToken_res_124 <= 1'h0;
      useV0AsMaskToken_res_125 <= 1'h0;
      useV0AsMaskToken_res_126 <= 1'h0;
      useV0AsMaskToken_res_127 <= 1'h0;
      useV0AsMaskToken_res_128 <= 1'h0;
      useV0AsMaskToken_res_129 <= 1'h0;
      useV0AsMaskToken_res_130 <= 1'h0;
      useV0AsMaskToken_res_131 <= 1'h0;
      useV0AsMaskToken_res_132 <= 1'h0;
      useV0AsMaskToken_res_133 <= 1'h0;
      useV0AsMaskToken_res_134 <= 1'h0;
      useV0AsMaskToken_res_135 <= 1'h0;
      useV0AsMaskToken_res_136 <= 1'h0;
      useV0AsMaskToken_res_137 <= 1'h0;
      useV0AsMaskToken_res_138 <= 1'h0;
      useV0AsMaskToken_res_139 <= 1'h0;
      useV0AsMaskToken_res_140 <= 1'h0;
      useV0AsMaskToken_res_141 <= 1'h0;
      useV0AsMaskToken_res_142 <= 1'h0;
      useV0AsMaskToken_res_143 <= 1'h0;
      useV0AsMaskToken_res_144 <= 1'h0;
      useV0AsMaskToken_res_145 <= 1'h0;
      useV0AsMaskToken_res_146 <= 1'h0;
      useV0AsMaskToken_res_147 <= 1'h0;
      useV0AsMaskToken_res_148 <= 1'h0;
      useV0AsMaskToken_res_149 <= 1'h0;
      useV0AsMaskToken_res_150 <= 1'h0;
      useV0AsMaskToken_res_151 <= 1'h0;
      useV0AsMaskToken_res_152 <= 1'h0;
      useV0AsMaskToken_res_153 <= 1'h0;
      useV0AsMaskToken_res_154 <= 1'h0;
      useV0AsMaskToken_res_155 <= 1'h0;
      useV0AsMaskToken_res_156 <= 1'h0;
      useV0AsMaskToken_res_157 <= 1'h0;
      useV0AsMaskToken_res_158 <= 1'h0;
      useV0AsMaskToken_res_159 <= 1'h0;
      useV0AsMaskToken_res_160 <= 1'h0;
      useV0AsMaskToken_res_161 <= 1'h0;
      useV0AsMaskToken_res_162 <= 1'h0;
      useV0AsMaskToken_res_163 <= 1'h0;
      useV0AsMaskToken_res_164 <= 1'h0;
      useV0AsMaskToken_res_165 <= 1'h0;
      useV0AsMaskToken_res_166 <= 1'h0;
      useV0AsMaskToken_res_167 <= 1'h0;
      useV0AsMaskToken_res_168 <= 1'h0;
      useV0AsMaskToken_res_169 <= 1'h0;
      useV0AsMaskToken_res_170 <= 1'h0;
      useV0AsMaskToken_res_171 <= 1'h0;
      useV0AsMaskToken_res_172 <= 1'h0;
      useV0AsMaskToken_res_173 <= 1'h0;
      useV0AsMaskToken_res_174 <= 1'h0;
      useV0AsMaskToken_res_175 <= 1'h0;
      useV0AsMaskToken_res_176 <= 1'h0;
      useV0AsMaskToken_res_177 <= 1'h0;
      useV0AsMaskToken_res_178 <= 1'h0;
      useV0AsMaskToken_res_179 <= 1'h0;
      useV0AsMaskToken_res_180 <= 1'h0;
      useV0AsMaskToken_res_181 <= 1'h0;
      useV0AsMaskToken_res_182 <= 1'h0;
      useV0AsMaskToken_res_183 <= 1'h0;
      useV0AsMaskToken_res_184 <= 1'h0;
      useV0AsMaskToken_res_185 <= 1'h0;
      useV0AsMaskToken_res_186 <= 1'h0;
      useV0AsMaskToken_res_187 <= 1'h0;
      useV0AsMaskToken_res_188 <= 1'h0;
      useV0AsMaskToken_res_189 <= 1'h0;
      useV0AsMaskToken_res_190 <= 1'h0;
      useV0AsMaskToken_res_191 <= 1'h0;
      useV0AsMaskToken_res_192 <= 1'h0;
      useV0AsMaskToken_res_193 <= 1'h0;
      useV0AsMaskToken_res_194 <= 1'h0;
      useV0AsMaskToken_res_195 <= 1'h0;
      useV0AsMaskToken_res_196 <= 1'h0;
      useV0AsMaskToken_res_197 <= 1'h0;
      useV0AsMaskToken_res_198 <= 1'h0;
      useV0AsMaskToken_res_199 <= 1'h0;
      useV0AsMaskToken_res_200 <= 1'h0;
      useV0AsMaskToken_res_201 <= 1'h0;
      useV0AsMaskToken_res_202 <= 1'h0;
      useV0AsMaskToken_res_203 <= 1'h0;
      useV0AsMaskToken_res_204 <= 1'h0;
      useV0AsMaskToken_res_205 <= 1'h0;
      useV0AsMaskToken_res_206 <= 1'h0;
      useV0AsMaskToken_res_207 <= 1'h0;
      useV0AsMaskToken_res_208 <= 1'h0;
      useV0AsMaskToken_res_209 <= 1'h0;
      useV0AsMaskToken_res_210 <= 1'h0;
      useV0AsMaskToken_res_211 <= 1'h0;
      useV0AsMaskToken_res_212 <= 1'h0;
      useV0AsMaskToken_res_213 <= 1'h0;
      useV0AsMaskToken_res_214 <= 1'h0;
      useV0AsMaskToken_res_215 <= 1'h0;
      useV0AsMaskToken_res_216 <= 1'h0;
      useV0AsMaskToken_res_217 <= 1'h0;
      useV0AsMaskToken_res_218 <= 1'h0;
      useV0AsMaskToken_res_219 <= 1'h0;
      useV0AsMaskToken_res_220 <= 1'h0;
      useV0AsMaskToken_res_221 <= 1'h0;
      useV0AsMaskToken_res_222 <= 1'h0;
      useV0AsMaskToken_res_223 <= 1'h0;
      useV0AsMaskToken_res_224 <= 1'h0;
      useV0AsMaskToken_res_225 <= 1'h0;
      useV0AsMaskToken_res_226 <= 1'h0;
      useV0AsMaskToken_res_227 <= 1'h0;
      useV0AsMaskToken_res_228 <= 1'h0;
      useV0AsMaskToken_res_229 <= 1'h0;
      useV0AsMaskToken_res_230 <= 1'h0;
      useV0AsMaskToken_res_231 <= 1'h0;
      useV0AsMaskToken_res_232 <= 1'h0;
      useV0AsMaskToken_res_233 <= 1'h0;
      useV0AsMaskToken_res_234 <= 1'h0;
      useV0AsMaskToken_res_235 <= 1'h0;
      useV0AsMaskToken_res_236 <= 1'h0;
      useV0AsMaskToken_res_237 <= 1'h0;
      useV0AsMaskToken_res_238 <= 1'h0;
      useV0AsMaskToken_res_239 <= 1'h0;
      useV0AsMaskToken_res_240 <= 1'h0;
      useV0AsMaskToken_res_241 <= 1'h0;
      useV0AsMaskToken_res_242 <= 1'h0;
      useV0AsMaskToken_res_243 <= 1'h0;
      useV0AsMaskToken_res_244 <= 1'h0;
      useV0AsMaskToken_res_245 <= 1'h0;
      useV0AsMaskToken_res_246 <= 1'h0;
      useV0AsMaskToken_res_247 <= 1'h0;
      useV0AsMaskToken_res_248 <= 1'h0;
      useV0AsMaskToken_res_249 <= 1'h0;
      useV0AsMaskToken_res_250 <= 1'h0;
      useV0AsMaskToken_res_251 <= 1'h0;
      useV0AsMaskToken_res_252 <= 1'h0;
      useV0AsMaskToken_res_253 <= 1'h0;
      useV0AsMaskToken_res_254 <= 1'h0;
      useV0AsMaskToken_res_255 <= 1'h0;
      maskUnitWriteV0 <= 1'h0;
    end
    else begin
      automatic logic [7:0] _v0WriteValidVec_T = v0WriteValidVec_updateOH | v0WriteValidVec_lsuWriteSet;
      automatic logic [7:0] _v0WriteValidVec_T_25 = v0WriteValidVec_updateOH_1 | v0WriteValidVec_lsuWriteSet_1;
      automatic logic [7:0] _v0WriteValidVec_T_50 = v0WriteValidVec_updateOH_2 | v0WriteValidVec_lsuWriteSet_2;
      automatic logic [7:0] _v0WriteValidVec_T_75 = v0WriteValidVec_updateOH_3 | v0WriteValidVec_lsuWriteSet_3;
      automatic logic [7:0] _v0WriteValidVec_T_100 = v0WriteValidVec_updateOH_4 | v0WriteValidVec_lsuWriteSet_4;
      automatic logic [7:0] _v0WriteValidVec_T_125 = v0WriteValidVec_updateOH_5 | v0WriteValidVec_lsuWriteSet_5;
      automatic logic [7:0] _v0WriteValidVec_T_150 = v0WriteValidVec_updateOH_6 | v0WriteValidVec_lsuWriteSet_6;
      automatic logic [7:0] _v0WriteValidVec_T_175 = v0WriteValidVec_updateOH_7 | v0WriteValidVec_lsuWriteSet_7;
      automatic logic [7:0] _v0WriteValidVec_T_200 = v0WriteValidVec_updateOH_8 | v0WriteValidVec_lsuWriteSet_8;
      automatic logic [7:0] _v0WriteValidVec_T_225 = v0WriteValidVec_updateOH_9 | v0WriteValidVec_lsuWriteSet_9;
      automatic logic [7:0] _v0WriteValidVec_T_250 = v0WriteValidVec_updateOH_10 | v0WriteValidVec_lsuWriteSet_10;
      automatic logic [7:0] _v0WriteValidVec_T_275 = v0WriteValidVec_updateOH_11 | v0WriteValidVec_lsuWriteSet_11;
      automatic logic [7:0] _v0WriteValidVec_T_300 = v0WriteValidVec_updateOH_12 | v0WriteValidVec_lsuWriteSet_12;
      automatic logic [7:0] _v0WriteValidVec_T_325 = v0WriteValidVec_updateOH_13 | v0WriteValidVec_lsuWriteSet_13;
      automatic logic [7:0] _v0WriteValidVec_T_350 = v0WriteValidVec_updateOH_14 | v0WriteValidVec_lsuWriteSet_14;
      automatic logic [7:0] _v0WriteValidVec_T_375 = v0WriteValidVec_updateOH_15 | v0WriteValidVec_lsuWriteSet_15;
      automatic logic [7:0] _v0WriteValidVec_T_400 = v0WriteValidVec_updateOH_16 | v0WriteValidVec_lsuWriteSet_16;
      automatic logic [7:0] _v0WriteValidVec_T_425 = v0WriteValidVec_updateOH_17 | v0WriteValidVec_lsuWriteSet_17;
      automatic logic [7:0] _v0WriteValidVec_T_450 = v0WriteValidVec_updateOH_18 | v0WriteValidVec_lsuWriteSet_18;
      automatic logic [7:0] _v0WriteValidVec_T_475 = v0WriteValidVec_updateOH_19 | v0WriteValidVec_lsuWriteSet_19;
      automatic logic [7:0] _v0WriteValidVec_T_500 = v0WriteValidVec_updateOH_20 | v0WriteValidVec_lsuWriteSet_20;
      automatic logic [7:0] _v0WriteValidVec_T_525 = v0WriteValidVec_updateOH_21 | v0WriteValidVec_lsuWriteSet_21;
      automatic logic [7:0] _v0WriteValidVec_T_550 = v0WriteValidVec_updateOH_22 | v0WriteValidVec_lsuWriteSet_22;
      automatic logic [7:0] _v0WriteValidVec_T_575 = v0WriteValidVec_updateOH_23 | v0WriteValidVec_lsuWriteSet_23;
      automatic logic [7:0] _v0WriteValidVec_T_600 = v0WriteValidVec_updateOH_24 | v0WriteValidVec_lsuWriteSet_24;
      automatic logic [7:0] _v0WriteValidVec_T_625 = v0WriteValidVec_updateOH_25 | v0WriteValidVec_lsuWriteSet_25;
      automatic logic [7:0] _v0WriteValidVec_T_650 = v0WriteValidVec_updateOH_26 | v0WriteValidVec_lsuWriteSet_26;
      automatic logic [7:0] _v0WriteValidVec_T_675 = v0WriteValidVec_updateOH_27 | v0WriteValidVec_lsuWriteSet_27;
      automatic logic [7:0] _v0WriteValidVec_T_700 = v0WriteValidVec_updateOH_28 | v0WriteValidVec_lsuWriteSet_28;
      automatic logic [7:0] _v0WriteValidVec_T_725 = v0WriteValidVec_updateOH_29 | v0WriteValidVec_lsuWriteSet_29;
      automatic logic [7:0] _v0WriteValidVec_T_750 = v0WriteValidVec_updateOH_30 | v0WriteValidVec_lsuWriteSet_30;
      automatic logic [7:0] _v0WriteValidVec_T_775 = v0WriteValidVec_updateOH_31 | v0WriteValidVec_lsuWriteSet_31;
      if (_v0WriteValidVec_T[0] | instructionFinish_0[0])
        v0WriteValidVec_res <= _v0WriteValidVec_T[0];
      if (_v0WriteValidVec_T[1] | instructionFinish_0[1])
        v0WriteValidVec_res_1 <= _v0WriteValidVec_T[1];
      if (_v0WriteValidVec_T[2] | instructionFinish_0[2])
        v0WriteValidVec_res_2 <= _v0WriteValidVec_T[2];
      if (_v0WriteValidVec_T[3] | instructionFinish_0[3])
        v0WriteValidVec_res_3 <= _v0WriteValidVec_T[3];
      if (_v0WriteValidVec_T[4] | instructionFinish_0[4])
        v0WriteValidVec_res_4 <= _v0WriteValidVec_T[4];
      if (_v0WriteValidVec_T[5] | instructionFinish_0[5])
        v0WriteValidVec_res_5 <= _v0WriteValidVec_T[5];
      if (_v0WriteValidVec_T[6] | instructionFinish_0[6])
        v0WriteValidVec_res_6 <= _v0WriteValidVec_T[6];
      if (_v0WriteValidVec_T[7] | instructionFinish_0[7])
        v0WriteValidVec_res_7 <= _v0WriteValidVec_T[7];
      if (_v0WriteValidVec_T_25[0] | instructionFinish_1[0])
        v0WriteValidVec_res_8 <= _v0WriteValidVec_T_25[0];
      if (_v0WriteValidVec_T_25[1] | instructionFinish_1[1])
        v0WriteValidVec_res_9 <= _v0WriteValidVec_T_25[1];
      if (_v0WriteValidVec_T_25[2] | instructionFinish_1[2])
        v0WriteValidVec_res_10 <= _v0WriteValidVec_T_25[2];
      if (_v0WriteValidVec_T_25[3] | instructionFinish_1[3])
        v0WriteValidVec_res_11 <= _v0WriteValidVec_T_25[3];
      if (_v0WriteValidVec_T_25[4] | instructionFinish_1[4])
        v0WriteValidVec_res_12 <= _v0WriteValidVec_T_25[4];
      if (_v0WriteValidVec_T_25[5] | instructionFinish_1[5])
        v0WriteValidVec_res_13 <= _v0WriteValidVec_T_25[5];
      if (_v0WriteValidVec_T_25[6] | instructionFinish_1[6])
        v0WriteValidVec_res_14 <= _v0WriteValidVec_T_25[6];
      if (_v0WriteValidVec_T_25[7] | instructionFinish_1[7])
        v0WriteValidVec_res_15 <= _v0WriteValidVec_T_25[7];
      if (_v0WriteValidVec_T_50[0] | instructionFinish_2[0])
        v0WriteValidVec_res_16 <= _v0WriteValidVec_T_50[0];
      if (_v0WriteValidVec_T_50[1] | instructionFinish_2[1])
        v0WriteValidVec_res_17 <= _v0WriteValidVec_T_50[1];
      if (_v0WriteValidVec_T_50[2] | instructionFinish_2[2])
        v0WriteValidVec_res_18 <= _v0WriteValidVec_T_50[2];
      if (_v0WriteValidVec_T_50[3] | instructionFinish_2[3])
        v0WriteValidVec_res_19 <= _v0WriteValidVec_T_50[3];
      if (_v0WriteValidVec_T_50[4] | instructionFinish_2[4])
        v0WriteValidVec_res_20 <= _v0WriteValidVec_T_50[4];
      if (_v0WriteValidVec_T_50[5] | instructionFinish_2[5])
        v0WriteValidVec_res_21 <= _v0WriteValidVec_T_50[5];
      if (_v0WriteValidVec_T_50[6] | instructionFinish_2[6])
        v0WriteValidVec_res_22 <= _v0WriteValidVec_T_50[6];
      if (_v0WriteValidVec_T_50[7] | instructionFinish_2[7])
        v0WriteValidVec_res_23 <= _v0WriteValidVec_T_50[7];
      if (_v0WriteValidVec_T_75[0] | instructionFinish_3[0])
        v0WriteValidVec_res_24 <= _v0WriteValidVec_T_75[0];
      if (_v0WriteValidVec_T_75[1] | instructionFinish_3[1])
        v0WriteValidVec_res_25 <= _v0WriteValidVec_T_75[1];
      if (_v0WriteValidVec_T_75[2] | instructionFinish_3[2])
        v0WriteValidVec_res_26 <= _v0WriteValidVec_T_75[2];
      if (_v0WriteValidVec_T_75[3] | instructionFinish_3[3])
        v0WriteValidVec_res_27 <= _v0WriteValidVec_T_75[3];
      if (_v0WriteValidVec_T_75[4] | instructionFinish_3[4])
        v0WriteValidVec_res_28 <= _v0WriteValidVec_T_75[4];
      if (_v0WriteValidVec_T_75[5] | instructionFinish_3[5])
        v0WriteValidVec_res_29 <= _v0WriteValidVec_T_75[5];
      if (_v0WriteValidVec_T_75[6] | instructionFinish_3[6])
        v0WriteValidVec_res_30 <= _v0WriteValidVec_T_75[6];
      if (_v0WriteValidVec_T_75[7] | instructionFinish_3[7])
        v0WriteValidVec_res_31 <= _v0WriteValidVec_T_75[7];
      if (_v0WriteValidVec_T_100[0] | instructionFinish_4[0])
        v0WriteValidVec_res_32 <= _v0WriteValidVec_T_100[0];
      if (_v0WriteValidVec_T_100[1] | instructionFinish_4[1])
        v0WriteValidVec_res_33 <= _v0WriteValidVec_T_100[1];
      if (_v0WriteValidVec_T_100[2] | instructionFinish_4[2])
        v0WriteValidVec_res_34 <= _v0WriteValidVec_T_100[2];
      if (_v0WriteValidVec_T_100[3] | instructionFinish_4[3])
        v0WriteValidVec_res_35 <= _v0WriteValidVec_T_100[3];
      if (_v0WriteValidVec_T_100[4] | instructionFinish_4[4])
        v0WriteValidVec_res_36 <= _v0WriteValidVec_T_100[4];
      if (_v0WriteValidVec_T_100[5] | instructionFinish_4[5])
        v0WriteValidVec_res_37 <= _v0WriteValidVec_T_100[5];
      if (_v0WriteValidVec_T_100[6] | instructionFinish_4[6])
        v0WriteValidVec_res_38 <= _v0WriteValidVec_T_100[6];
      if (_v0WriteValidVec_T_100[7] | instructionFinish_4[7])
        v0WriteValidVec_res_39 <= _v0WriteValidVec_T_100[7];
      if (_v0WriteValidVec_T_125[0] | instructionFinish_5[0])
        v0WriteValidVec_res_40 <= _v0WriteValidVec_T_125[0];
      if (_v0WriteValidVec_T_125[1] | instructionFinish_5[1])
        v0WriteValidVec_res_41 <= _v0WriteValidVec_T_125[1];
      if (_v0WriteValidVec_T_125[2] | instructionFinish_5[2])
        v0WriteValidVec_res_42 <= _v0WriteValidVec_T_125[2];
      if (_v0WriteValidVec_T_125[3] | instructionFinish_5[3])
        v0WriteValidVec_res_43 <= _v0WriteValidVec_T_125[3];
      if (_v0WriteValidVec_T_125[4] | instructionFinish_5[4])
        v0WriteValidVec_res_44 <= _v0WriteValidVec_T_125[4];
      if (_v0WriteValidVec_T_125[5] | instructionFinish_5[5])
        v0WriteValidVec_res_45 <= _v0WriteValidVec_T_125[5];
      if (_v0WriteValidVec_T_125[6] | instructionFinish_5[6])
        v0WriteValidVec_res_46 <= _v0WriteValidVec_T_125[6];
      if (_v0WriteValidVec_T_125[7] | instructionFinish_5[7])
        v0WriteValidVec_res_47 <= _v0WriteValidVec_T_125[7];
      if (_v0WriteValidVec_T_150[0] | instructionFinish_6[0])
        v0WriteValidVec_res_48 <= _v0WriteValidVec_T_150[0];
      if (_v0WriteValidVec_T_150[1] | instructionFinish_6[1])
        v0WriteValidVec_res_49 <= _v0WriteValidVec_T_150[1];
      if (_v0WriteValidVec_T_150[2] | instructionFinish_6[2])
        v0WriteValidVec_res_50 <= _v0WriteValidVec_T_150[2];
      if (_v0WriteValidVec_T_150[3] | instructionFinish_6[3])
        v0WriteValidVec_res_51 <= _v0WriteValidVec_T_150[3];
      if (_v0WriteValidVec_T_150[4] | instructionFinish_6[4])
        v0WriteValidVec_res_52 <= _v0WriteValidVec_T_150[4];
      if (_v0WriteValidVec_T_150[5] | instructionFinish_6[5])
        v0WriteValidVec_res_53 <= _v0WriteValidVec_T_150[5];
      if (_v0WriteValidVec_T_150[6] | instructionFinish_6[6])
        v0WriteValidVec_res_54 <= _v0WriteValidVec_T_150[6];
      if (_v0WriteValidVec_T_150[7] | instructionFinish_6[7])
        v0WriteValidVec_res_55 <= _v0WriteValidVec_T_150[7];
      if (_v0WriteValidVec_T_175[0] | instructionFinish_7[0])
        v0WriteValidVec_res_56 <= _v0WriteValidVec_T_175[0];
      if (_v0WriteValidVec_T_175[1] | instructionFinish_7[1])
        v0WriteValidVec_res_57 <= _v0WriteValidVec_T_175[1];
      if (_v0WriteValidVec_T_175[2] | instructionFinish_7[2])
        v0WriteValidVec_res_58 <= _v0WriteValidVec_T_175[2];
      if (_v0WriteValidVec_T_175[3] | instructionFinish_7[3])
        v0WriteValidVec_res_59 <= _v0WriteValidVec_T_175[3];
      if (_v0WriteValidVec_T_175[4] | instructionFinish_7[4])
        v0WriteValidVec_res_60 <= _v0WriteValidVec_T_175[4];
      if (_v0WriteValidVec_T_175[5] | instructionFinish_7[5])
        v0WriteValidVec_res_61 <= _v0WriteValidVec_T_175[5];
      if (_v0WriteValidVec_T_175[6] | instructionFinish_7[6])
        v0WriteValidVec_res_62 <= _v0WriteValidVec_T_175[6];
      if (_v0WriteValidVec_T_175[7] | instructionFinish_7[7])
        v0WriteValidVec_res_63 <= _v0WriteValidVec_T_175[7];
      if (_v0WriteValidVec_T_200[0] | instructionFinish_8[0])
        v0WriteValidVec_res_64 <= _v0WriteValidVec_T_200[0];
      if (_v0WriteValidVec_T_200[1] | instructionFinish_8[1])
        v0WriteValidVec_res_65 <= _v0WriteValidVec_T_200[1];
      if (_v0WriteValidVec_T_200[2] | instructionFinish_8[2])
        v0WriteValidVec_res_66 <= _v0WriteValidVec_T_200[2];
      if (_v0WriteValidVec_T_200[3] | instructionFinish_8[3])
        v0WriteValidVec_res_67 <= _v0WriteValidVec_T_200[3];
      if (_v0WriteValidVec_T_200[4] | instructionFinish_8[4])
        v0WriteValidVec_res_68 <= _v0WriteValidVec_T_200[4];
      if (_v0WriteValidVec_T_200[5] | instructionFinish_8[5])
        v0WriteValidVec_res_69 <= _v0WriteValidVec_T_200[5];
      if (_v0WriteValidVec_T_200[6] | instructionFinish_8[6])
        v0WriteValidVec_res_70 <= _v0WriteValidVec_T_200[6];
      if (_v0WriteValidVec_T_200[7] | instructionFinish_8[7])
        v0WriteValidVec_res_71 <= _v0WriteValidVec_T_200[7];
      if (_v0WriteValidVec_T_225[0] | instructionFinish_9[0])
        v0WriteValidVec_res_72 <= _v0WriteValidVec_T_225[0];
      if (_v0WriteValidVec_T_225[1] | instructionFinish_9[1])
        v0WriteValidVec_res_73 <= _v0WriteValidVec_T_225[1];
      if (_v0WriteValidVec_T_225[2] | instructionFinish_9[2])
        v0WriteValidVec_res_74 <= _v0WriteValidVec_T_225[2];
      if (_v0WriteValidVec_T_225[3] | instructionFinish_9[3])
        v0WriteValidVec_res_75 <= _v0WriteValidVec_T_225[3];
      if (_v0WriteValidVec_T_225[4] | instructionFinish_9[4])
        v0WriteValidVec_res_76 <= _v0WriteValidVec_T_225[4];
      if (_v0WriteValidVec_T_225[5] | instructionFinish_9[5])
        v0WriteValidVec_res_77 <= _v0WriteValidVec_T_225[5];
      if (_v0WriteValidVec_T_225[6] | instructionFinish_9[6])
        v0WriteValidVec_res_78 <= _v0WriteValidVec_T_225[6];
      if (_v0WriteValidVec_T_225[7] | instructionFinish_9[7])
        v0WriteValidVec_res_79 <= _v0WriteValidVec_T_225[7];
      if (_v0WriteValidVec_T_250[0] | instructionFinish_10[0])
        v0WriteValidVec_res_80 <= _v0WriteValidVec_T_250[0];
      if (_v0WriteValidVec_T_250[1] | instructionFinish_10[1])
        v0WriteValidVec_res_81 <= _v0WriteValidVec_T_250[1];
      if (_v0WriteValidVec_T_250[2] | instructionFinish_10[2])
        v0WriteValidVec_res_82 <= _v0WriteValidVec_T_250[2];
      if (_v0WriteValidVec_T_250[3] | instructionFinish_10[3])
        v0WriteValidVec_res_83 <= _v0WriteValidVec_T_250[3];
      if (_v0WriteValidVec_T_250[4] | instructionFinish_10[4])
        v0WriteValidVec_res_84 <= _v0WriteValidVec_T_250[4];
      if (_v0WriteValidVec_T_250[5] | instructionFinish_10[5])
        v0WriteValidVec_res_85 <= _v0WriteValidVec_T_250[5];
      if (_v0WriteValidVec_T_250[6] | instructionFinish_10[6])
        v0WriteValidVec_res_86 <= _v0WriteValidVec_T_250[6];
      if (_v0WriteValidVec_T_250[7] | instructionFinish_10[7])
        v0WriteValidVec_res_87 <= _v0WriteValidVec_T_250[7];
      if (_v0WriteValidVec_T_275[0] | instructionFinish_11[0])
        v0WriteValidVec_res_88 <= _v0WriteValidVec_T_275[0];
      if (_v0WriteValidVec_T_275[1] | instructionFinish_11[1])
        v0WriteValidVec_res_89 <= _v0WriteValidVec_T_275[1];
      if (_v0WriteValidVec_T_275[2] | instructionFinish_11[2])
        v0WriteValidVec_res_90 <= _v0WriteValidVec_T_275[2];
      if (_v0WriteValidVec_T_275[3] | instructionFinish_11[3])
        v0WriteValidVec_res_91 <= _v0WriteValidVec_T_275[3];
      if (_v0WriteValidVec_T_275[4] | instructionFinish_11[4])
        v0WriteValidVec_res_92 <= _v0WriteValidVec_T_275[4];
      if (_v0WriteValidVec_T_275[5] | instructionFinish_11[5])
        v0WriteValidVec_res_93 <= _v0WriteValidVec_T_275[5];
      if (_v0WriteValidVec_T_275[6] | instructionFinish_11[6])
        v0WriteValidVec_res_94 <= _v0WriteValidVec_T_275[6];
      if (_v0WriteValidVec_T_275[7] | instructionFinish_11[7])
        v0WriteValidVec_res_95 <= _v0WriteValidVec_T_275[7];
      if (_v0WriteValidVec_T_300[0] | instructionFinish_12[0])
        v0WriteValidVec_res_96 <= _v0WriteValidVec_T_300[0];
      if (_v0WriteValidVec_T_300[1] | instructionFinish_12[1])
        v0WriteValidVec_res_97 <= _v0WriteValidVec_T_300[1];
      if (_v0WriteValidVec_T_300[2] | instructionFinish_12[2])
        v0WriteValidVec_res_98 <= _v0WriteValidVec_T_300[2];
      if (_v0WriteValidVec_T_300[3] | instructionFinish_12[3])
        v0WriteValidVec_res_99 <= _v0WriteValidVec_T_300[3];
      if (_v0WriteValidVec_T_300[4] | instructionFinish_12[4])
        v0WriteValidVec_res_100 <= _v0WriteValidVec_T_300[4];
      if (_v0WriteValidVec_T_300[5] | instructionFinish_12[5])
        v0WriteValidVec_res_101 <= _v0WriteValidVec_T_300[5];
      if (_v0WriteValidVec_T_300[6] | instructionFinish_12[6])
        v0WriteValidVec_res_102 <= _v0WriteValidVec_T_300[6];
      if (_v0WriteValidVec_T_300[7] | instructionFinish_12[7])
        v0WriteValidVec_res_103 <= _v0WriteValidVec_T_300[7];
      if (_v0WriteValidVec_T_325[0] | instructionFinish_13[0])
        v0WriteValidVec_res_104 <= _v0WriteValidVec_T_325[0];
      if (_v0WriteValidVec_T_325[1] | instructionFinish_13[1])
        v0WriteValidVec_res_105 <= _v0WriteValidVec_T_325[1];
      if (_v0WriteValidVec_T_325[2] | instructionFinish_13[2])
        v0WriteValidVec_res_106 <= _v0WriteValidVec_T_325[2];
      if (_v0WriteValidVec_T_325[3] | instructionFinish_13[3])
        v0WriteValidVec_res_107 <= _v0WriteValidVec_T_325[3];
      if (_v0WriteValidVec_T_325[4] | instructionFinish_13[4])
        v0WriteValidVec_res_108 <= _v0WriteValidVec_T_325[4];
      if (_v0WriteValidVec_T_325[5] | instructionFinish_13[5])
        v0WriteValidVec_res_109 <= _v0WriteValidVec_T_325[5];
      if (_v0WriteValidVec_T_325[6] | instructionFinish_13[6])
        v0WriteValidVec_res_110 <= _v0WriteValidVec_T_325[6];
      if (_v0WriteValidVec_T_325[7] | instructionFinish_13[7])
        v0WriteValidVec_res_111 <= _v0WriteValidVec_T_325[7];
      if (_v0WriteValidVec_T_350[0] | instructionFinish_14[0])
        v0WriteValidVec_res_112 <= _v0WriteValidVec_T_350[0];
      if (_v0WriteValidVec_T_350[1] | instructionFinish_14[1])
        v0WriteValidVec_res_113 <= _v0WriteValidVec_T_350[1];
      if (_v0WriteValidVec_T_350[2] | instructionFinish_14[2])
        v0WriteValidVec_res_114 <= _v0WriteValidVec_T_350[2];
      if (_v0WriteValidVec_T_350[3] | instructionFinish_14[3])
        v0WriteValidVec_res_115 <= _v0WriteValidVec_T_350[3];
      if (_v0WriteValidVec_T_350[4] | instructionFinish_14[4])
        v0WriteValidVec_res_116 <= _v0WriteValidVec_T_350[4];
      if (_v0WriteValidVec_T_350[5] | instructionFinish_14[5])
        v0WriteValidVec_res_117 <= _v0WriteValidVec_T_350[5];
      if (_v0WriteValidVec_T_350[6] | instructionFinish_14[6])
        v0WriteValidVec_res_118 <= _v0WriteValidVec_T_350[6];
      if (_v0WriteValidVec_T_350[7] | instructionFinish_14[7])
        v0WriteValidVec_res_119 <= _v0WriteValidVec_T_350[7];
      if (_v0WriteValidVec_T_375[0] | instructionFinish_15[0])
        v0WriteValidVec_res_120 <= _v0WriteValidVec_T_375[0];
      if (_v0WriteValidVec_T_375[1] | instructionFinish_15[1])
        v0WriteValidVec_res_121 <= _v0WriteValidVec_T_375[1];
      if (_v0WriteValidVec_T_375[2] | instructionFinish_15[2])
        v0WriteValidVec_res_122 <= _v0WriteValidVec_T_375[2];
      if (_v0WriteValidVec_T_375[3] | instructionFinish_15[3])
        v0WriteValidVec_res_123 <= _v0WriteValidVec_T_375[3];
      if (_v0WriteValidVec_T_375[4] | instructionFinish_15[4])
        v0WriteValidVec_res_124 <= _v0WriteValidVec_T_375[4];
      if (_v0WriteValidVec_T_375[5] | instructionFinish_15[5])
        v0WriteValidVec_res_125 <= _v0WriteValidVec_T_375[5];
      if (_v0WriteValidVec_T_375[6] | instructionFinish_15[6])
        v0WriteValidVec_res_126 <= _v0WriteValidVec_T_375[6];
      if (_v0WriteValidVec_T_375[7] | instructionFinish_15[7])
        v0WriteValidVec_res_127 <= _v0WriteValidVec_T_375[7];
      if (_v0WriteValidVec_T_400[0] | instructionFinish_16[0])
        v0WriteValidVec_res_128 <= _v0WriteValidVec_T_400[0];
      if (_v0WriteValidVec_T_400[1] | instructionFinish_16[1])
        v0WriteValidVec_res_129 <= _v0WriteValidVec_T_400[1];
      if (_v0WriteValidVec_T_400[2] | instructionFinish_16[2])
        v0WriteValidVec_res_130 <= _v0WriteValidVec_T_400[2];
      if (_v0WriteValidVec_T_400[3] | instructionFinish_16[3])
        v0WriteValidVec_res_131 <= _v0WriteValidVec_T_400[3];
      if (_v0WriteValidVec_T_400[4] | instructionFinish_16[4])
        v0WriteValidVec_res_132 <= _v0WriteValidVec_T_400[4];
      if (_v0WriteValidVec_T_400[5] | instructionFinish_16[5])
        v0WriteValidVec_res_133 <= _v0WriteValidVec_T_400[5];
      if (_v0WriteValidVec_T_400[6] | instructionFinish_16[6])
        v0WriteValidVec_res_134 <= _v0WriteValidVec_T_400[6];
      if (_v0WriteValidVec_T_400[7] | instructionFinish_16[7])
        v0WriteValidVec_res_135 <= _v0WriteValidVec_T_400[7];
      if (_v0WriteValidVec_T_425[0] | instructionFinish_17[0])
        v0WriteValidVec_res_136 <= _v0WriteValidVec_T_425[0];
      if (_v0WriteValidVec_T_425[1] | instructionFinish_17[1])
        v0WriteValidVec_res_137 <= _v0WriteValidVec_T_425[1];
      if (_v0WriteValidVec_T_425[2] | instructionFinish_17[2])
        v0WriteValidVec_res_138 <= _v0WriteValidVec_T_425[2];
      if (_v0WriteValidVec_T_425[3] | instructionFinish_17[3])
        v0WriteValidVec_res_139 <= _v0WriteValidVec_T_425[3];
      if (_v0WriteValidVec_T_425[4] | instructionFinish_17[4])
        v0WriteValidVec_res_140 <= _v0WriteValidVec_T_425[4];
      if (_v0WriteValidVec_T_425[5] | instructionFinish_17[5])
        v0WriteValidVec_res_141 <= _v0WriteValidVec_T_425[5];
      if (_v0WriteValidVec_T_425[6] | instructionFinish_17[6])
        v0WriteValidVec_res_142 <= _v0WriteValidVec_T_425[6];
      if (_v0WriteValidVec_T_425[7] | instructionFinish_17[7])
        v0WriteValidVec_res_143 <= _v0WriteValidVec_T_425[7];
      if (_v0WriteValidVec_T_450[0] | instructionFinish_18[0])
        v0WriteValidVec_res_144 <= _v0WriteValidVec_T_450[0];
      if (_v0WriteValidVec_T_450[1] | instructionFinish_18[1])
        v0WriteValidVec_res_145 <= _v0WriteValidVec_T_450[1];
      if (_v0WriteValidVec_T_450[2] | instructionFinish_18[2])
        v0WriteValidVec_res_146 <= _v0WriteValidVec_T_450[2];
      if (_v0WriteValidVec_T_450[3] | instructionFinish_18[3])
        v0WriteValidVec_res_147 <= _v0WriteValidVec_T_450[3];
      if (_v0WriteValidVec_T_450[4] | instructionFinish_18[4])
        v0WriteValidVec_res_148 <= _v0WriteValidVec_T_450[4];
      if (_v0WriteValidVec_T_450[5] | instructionFinish_18[5])
        v0WriteValidVec_res_149 <= _v0WriteValidVec_T_450[5];
      if (_v0WriteValidVec_T_450[6] | instructionFinish_18[6])
        v0WriteValidVec_res_150 <= _v0WriteValidVec_T_450[6];
      if (_v0WriteValidVec_T_450[7] | instructionFinish_18[7])
        v0WriteValidVec_res_151 <= _v0WriteValidVec_T_450[7];
      if (_v0WriteValidVec_T_475[0] | instructionFinish_19[0])
        v0WriteValidVec_res_152 <= _v0WriteValidVec_T_475[0];
      if (_v0WriteValidVec_T_475[1] | instructionFinish_19[1])
        v0WriteValidVec_res_153 <= _v0WriteValidVec_T_475[1];
      if (_v0WriteValidVec_T_475[2] | instructionFinish_19[2])
        v0WriteValidVec_res_154 <= _v0WriteValidVec_T_475[2];
      if (_v0WriteValidVec_T_475[3] | instructionFinish_19[3])
        v0WriteValidVec_res_155 <= _v0WriteValidVec_T_475[3];
      if (_v0WriteValidVec_T_475[4] | instructionFinish_19[4])
        v0WriteValidVec_res_156 <= _v0WriteValidVec_T_475[4];
      if (_v0WriteValidVec_T_475[5] | instructionFinish_19[5])
        v0WriteValidVec_res_157 <= _v0WriteValidVec_T_475[5];
      if (_v0WriteValidVec_T_475[6] | instructionFinish_19[6])
        v0WriteValidVec_res_158 <= _v0WriteValidVec_T_475[6];
      if (_v0WriteValidVec_T_475[7] | instructionFinish_19[7])
        v0WriteValidVec_res_159 <= _v0WriteValidVec_T_475[7];
      if (_v0WriteValidVec_T_500[0] | instructionFinish_20[0])
        v0WriteValidVec_res_160 <= _v0WriteValidVec_T_500[0];
      if (_v0WriteValidVec_T_500[1] | instructionFinish_20[1])
        v0WriteValidVec_res_161 <= _v0WriteValidVec_T_500[1];
      if (_v0WriteValidVec_T_500[2] | instructionFinish_20[2])
        v0WriteValidVec_res_162 <= _v0WriteValidVec_T_500[2];
      if (_v0WriteValidVec_T_500[3] | instructionFinish_20[3])
        v0WriteValidVec_res_163 <= _v0WriteValidVec_T_500[3];
      if (_v0WriteValidVec_T_500[4] | instructionFinish_20[4])
        v0WriteValidVec_res_164 <= _v0WriteValidVec_T_500[4];
      if (_v0WriteValidVec_T_500[5] | instructionFinish_20[5])
        v0WriteValidVec_res_165 <= _v0WriteValidVec_T_500[5];
      if (_v0WriteValidVec_T_500[6] | instructionFinish_20[6])
        v0WriteValidVec_res_166 <= _v0WriteValidVec_T_500[6];
      if (_v0WriteValidVec_T_500[7] | instructionFinish_20[7])
        v0WriteValidVec_res_167 <= _v0WriteValidVec_T_500[7];
      if (_v0WriteValidVec_T_525[0] | instructionFinish_21[0])
        v0WriteValidVec_res_168 <= _v0WriteValidVec_T_525[0];
      if (_v0WriteValidVec_T_525[1] | instructionFinish_21[1])
        v0WriteValidVec_res_169 <= _v0WriteValidVec_T_525[1];
      if (_v0WriteValidVec_T_525[2] | instructionFinish_21[2])
        v0WriteValidVec_res_170 <= _v0WriteValidVec_T_525[2];
      if (_v0WriteValidVec_T_525[3] | instructionFinish_21[3])
        v0WriteValidVec_res_171 <= _v0WriteValidVec_T_525[3];
      if (_v0WriteValidVec_T_525[4] | instructionFinish_21[4])
        v0WriteValidVec_res_172 <= _v0WriteValidVec_T_525[4];
      if (_v0WriteValidVec_T_525[5] | instructionFinish_21[5])
        v0WriteValidVec_res_173 <= _v0WriteValidVec_T_525[5];
      if (_v0WriteValidVec_T_525[6] | instructionFinish_21[6])
        v0WriteValidVec_res_174 <= _v0WriteValidVec_T_525[6];
      if (_v0WriteValidVec_T_525[7] | instructionFinish_21[7])
        v0WriteValidVec_res_175 <= _v0WriteValidVec_T_525[7];
      if (_v0WriteValidVec_T_550[0] | instructionFinish_22[0])
        v0WriteValidVec_res_176 <= _v0WriteValidVec_T_550[0];
      if (_v0WriteValidVec_T_550[1] | instructionFinish_22[1])
        v0WriteValidVec_res_177 <= _v0WriteValidVec_T_550[1];
      if (_v0WriteValidVec_T_550[2] | instructionFinish_22[2])
        v0WriteValidVec_res_178 <= _v0WriteValidVec_T_550[2];
      if (_v0WriteValidVec_T_550[3] | instructionFinish_22[3])
        v0WriteValidVec_res_179 <= _v0WriteValidVec_T_550[3];
      if (_v0WriteValidVec_T_550[4] | instructionFinish_22[4])
        v0WriteValidVec_res_180 <= _v0WriteValidVec_T_550[4];
      if (_v0WriteValidVec_T_550[5] | instructionFinish_22[5])
        v0WriteValidVec_res_181 <= _v0WriteValidVec_T_550[5];
      if (_v0WriteValidVec_T_550[6] | instructionFinish_22[6])
        v0WriteValidVec_res_182 <= _v0WriteValidVec_T_550[6];
      if (_v0WriteValidVec_T_550[7] | instructionFinish_22[7])
        v0WriteValidVec_res_183 <= _v0WriteValidVec_T_550[7];
      if (_v0WriteValidVec_T_575[0] | instructionFinish_23[0])
        v0WriteValidVec_res_184 <= _v0WriteValidVec_T_575[0];
      if (_v0WriteValidVec_T_575[1] | instructionFinish_23[1])
        v0WriteValidVec_res_185 <= _v0WriteValidVec_T_575[1];
      if (_v0WriteValidVec_T_575[2] | instructionFinish_23[2])
        v0WriteValidVec_res_186 <= _v0WriteValidVec_T_575[2];
      if (_v0WriteValidVec_T_575[3] | instructionFinish_23[3])
        v0WriteValidVec_res_187 <= _v0WriteValidVec_T_575[3];
      if (_v0WriteValidVec_T_575[4] | instructionFinish_23[4])
        v0WriteValidVec_res_188 <= _v0WriteValidVec_T_575[4];
      if (_v0WriteValidVec_T_575[5] | instructionFinish_23[5])
        v0WriteValidVec_res_189 <= _v0WriteValidVec_T_575[5];
      if (_v0WriteValidVec_T_575[6] | instructionFinish_23[6])
        v0WriteValidVec_res_190 <= _v0WriteValidVec_T_575[6];
      if (_v0WriteValidVec_T_575[7] | instructionFinish_23[7])
        v0WriteValidVec_res_191 <= _v0WriteValidVec_T_575[7];
      if (_v0WriteValidVec_T_600[0] | instructionFinish_24[0])
        v0WriteValidVec_res_192 <= _v0WriteValidVec_T_600[0];
      if (_v0WriteValidVec_T_600[1] | instructionFinish_24[1])
        v0WriteValidVec_res_193 <= _v0WriteValidVec_T_600[1];
      if (_v0WriteValidVec_T_600[2] | instructionFinish_24[2])
        v0WriteValidVec_res_194 <= _v0WriteValidVec_T_600[2];
      if (_v0WriteValidVec_T_600[3] | instructionFinish_24[3])
        v0WriteValidVec_res_195 <= _v0WriteValidVec_T_600[3];
      if (_v0WriteValidVec_T_600[4] | instructionFinish_24[4])
        v0WriteValidVec_res_196 <= _v0WriteValidVec_T_600[4];
      if (_v0WriteValidVec_T_600[5] | instructionFinish_24[5])
        v0WriteValidVec_res_197 <= _v0WriteValidVec_T_600[5];
      if (_v0WriteValidVec_T_600[6] | instructionFinish_24[6])
        v0WriteValidVec_res_198 <= _v0WriteValidVec_T_600[6];
      if (_v0WriteValidVec_T_600[7] | instructionFinish_24[7])
        v0WriteValidVec_res_199 <= _v0WriteValidVec_T_600[7];
      if (_v0WriteValidVec_T_625[0] | instructionFinish_25[0])
        v0WriteValidVec_res_200 <= _v0WriteValidVec_T_625[0];
      if (_v0WriteValidVec_T_625[1] | instructionFinish_25[1])
        v0WriteValidVec_res_201 <= _v0WriteValidVec_T_625[1];
      if (_v0WriteValidVec_T_625[2] | instructionFinish_25[2])
        v0WriteValidVec_res_202 <= _v0WriteValidVec_T_625[2];
      if (_v0WriteValidVec_T_625[3] | instructionFinish_25[3])
        v0WriteValidVec_res_203 <= _v0WriteValidVec_T_625[3];
      if (_v0WriteValidVec_T_625[4] | instructionFinish_25[4])
        v0WriteValidVec_res_204 <= _v0WriteValidVec_T_625[4];
      if (_v0WriteValidVec_T_625[5] | instructionFinish_25[5])
        v0WriteValidVec_res_205 <= _v0WriteValidVec_T_625[5];
      if (_v0WriteValidVec_T_625[6] | instructionFinish_25[6])
        v0WriteValidVec_res_206 <= _v0WriteValidVec_T_625[6];
      if (_v0WriteValidVec_T_625[7] | instructionFinish_25[7])
        v0WriteValidVec_res_207 <= _v0WriteValidVec_T_625[7];
      if (_v0WriteValidVec_T_650[0] | instructionFinish_26[0])
        v0WriteValidVec_res_208 <= _v0WriteValidVec_T_650[0];
      if (_v0WriteValidVec_T_650[1] | instructionFinish_26[1])
        v0WriteValidVec_res_209 <= _v0WriteValidVec_T_650[1];
      if (_v0WriteValidVec_T_650[2] | instructionFinish_26[2])
        v0WriteValidVec_res_210 <= _v0WriteValidVec_T_650[2];
      if (_v0WriteValidVec_T_650[3] | instructionFinish_26[3])
        v0WriteValidVec_res_211 <= _v0WriteValidVec_T_650[3];
      if (_v0WriteValidVec_T_650[4] | instructionFinish_26[4])
        v0WriteValidVec_res_212 <= _v0WriteValidVec_T_650[4];
      if (_v0WriteValidVec_T_650[5] | instructionFinish_26[5])
        v0WriteValidVec_res_213 <= _v0WriteValidVec_T_650[5];
      if (_v0WriteValidVec_T_650[6] | instructionFinish_26[6])
        v0WriteValidVec_res_214 <= _v0WriteValidVec_T_650[6];
      if (_v0WriteValidVec_T_650[7] | instructionFinish_26[7])
        v0WriteValidVec_res_215 <= _v0WriteValidVec_T_650[7];
      if (_v0WriteValidVec_T_675[0] | instructionFinish_27[0])
        v0WriteValidVec_res_216 <= _v0WriteValidVec_T_675[0];
      if (_v0WriteValidVec_T_675[1] | instructionFinish_27[1])
        v0WriteValidVec_res_217 <= _v0WriteValidVec_T_675[1];
      if (_v0WriteValidVec_T_675[2] | instructionFinish_27[2])
        v0WriteValidVec_res_218 <= _v0WriteValidVec_T_675[2];
      if (_v0WriteValidVec_T_675[3] | instructionFinish_27[3])
        v0WriteValidVec_res_219 <= _v0WriteValidVec_T_675[3];
      if (_v0WriteValidVec_T_675[4] | instructionFinish_27[4])
        v0WriteValidVec_res_220 <= _v0WriteValidVec_T_675[4];
      if (_v0WriteValidVec_T_675[5] | instructionFinish_27[5])
        v0WriteValidVec_res_221 <= _v0WriteValidVec_T_675[5];
      if (_v0WriteValidVec_T_675[6] | instructionFinish_27[6])
        v0WriteValidVec_res_222 <= _v0WriteValidVec_T_675[6];
      if (_v0WriteValidVec_T_675[7] | instructionFinish_27[7])
        v0WriteValidVec_res_223 <= _v0WriteValidVec_T_675[7];
      if (_v0WriteValidVec_T_700[0] | instructionFinish_28[0])
        v0WriteValidVec_res_224 <= _v0WriteValidVec_T_700[0];
      if (_v0WriteValidVec_T_700[1] | instructionFinish_28[1])
        v0WriteValidVec_res_225 <= _v0WriteValidVec_T_700[1];
      if (_v0WriteValidVec_T_700[2] | instructionFinish_28[2])
        v0WriteValidVec_res_226 <= _v0WriteValidVec_T_700[2];
      if (_v0WriteValidVec_T_700[3] | instructionFinish_28[3])
        v0WriteValidVec_res_227 <= _v0WriteValidVec_T_700[3];
      if (_v0WriteValidVec_T_700[4] | instructionFinish_28[4])
        v0WriteValidVec_res_228 <= _v0WriteValidVec_T_700[4];
      if (_v0WriteValidVec_T_700[5] | instructionFinish_28[5])
        v0WriteValidVec_res_229 <= _v0WriteValidVec_T_700[5];
      if (_v0WriteValidVec_T_700[6] | instructionFinish_28[6])
        v0WriteValidVec_res_230 <= _v0WriteValidVec_T_700[6];
      if (_v0WriteValidVec_T_700[7] | instructionFinish_28[7])
        v0WriteValidVec_res_231 <= _v0WriteValidVec_T_700[7];
      if (_v0WriteValidVec_T_725[0] | instructionFinish_29[0])
        v0WriteValidVec_res_232 <= _v0WriteValidVec_T_725[0];
      if (_v0WriteValidVec_T_725[1] | instructionFinish_29[1])
        v0WriteValidVec_res_233 <= _v0WriteValidVec_T_725[1];
      if (_v0WriteValidVec_T_725[2] | instructionFinish_29[2])
        v0WriteValidVec_res_234 <= _v0WriteValidVec_T_725[2];
      if (_v0WriteValidVec_T_725[3] | instructionFinish_29[3])
        v0WriteValidVec_res_235 <= _v0WriteValidVec_T_725[3];
      if (_v0WriteValidVec_T_725[4] | instructionFinish_29[4])
        v0WriteValidVec_res_236 <= _v0WriteValidVec_T_725[4];
      if (_v0WriteValidVec_T_725[5] | instructionFinish_29[5])
        v0WriteValidVec_res_237 <= _v0WriteValidVec_T_725[5];
      if (_v0WriteValidVec_T_725[6] | instructionFinish_29[6])
        v0WriteValidVec_res_238 <= _v0WriteValidVec_T_725[6];
      if (_v0WriteValidVec_T_725[7] | instructionFinish_29[7])
        v0WriteValidVec_res_239 <= _v0WriteValidVec_T_725[7];
      if (_v0WriteValidVec_T_750[0] | instructionFinish_30[0])
        v0WriteValidVec_res_240 <= _v0WriteValidVec_T_750[0];
      if (_v0WriteValidVec_T_750[1] | instructionFinish_30[1])
        v0WriteValidVec_res_241 <= _v0WriteValidVec_T_750[1];
      if (_v0WriteValidVec_T_750[2] | instructionFinish_30[2])
        v0WriteValidVec_res_242 <= _v0WriteValidVec_T_750[2];
      if (_v0WriteValidVec_T_750[3] | instructionFinish_30[3])
        v0WriteValidVec_res_243 <= _v0WriteValidVec_T_750[3];
      if (_v0WriteValidVec_T_750[4] | instructionFinish_30[4])
        v0WriteValidVec_res_244 <= _v0WriteValidVec_T_750[4];
      if (_v0WriteValidVec_T_750[5] | instructionFinish_30[5])
        v0WriteValidVec_res_245 <= _v0WriteValidVec_T_750[5];
      if (_v0WriteValidVec_T_750[6] | instructionFinish_30[6])
        v0WriteValidVec_res_246 <= _v0WriteValidVec_T_750[6];
      if (_v0WriteValidVec_T_750[7] | instructionFinish_30[7])
        v0WriteValidVec_res_247 <= _v0WriteValidVec_T_750[7];
      if (_v0WriteValidVec_T_775[0] | instructionFinish_31[0])
        v0WriteValidVec_res_248 <= _v0WriteValidVec_T_775[0];
      if (_v0WriteValidVec_T_775[1] | instructionFinish_31[1])
        v0WriteValidVec_res_249 <= _v0WriteValidVec_T_775[1];
      if (_v0WriteValidVec_T_775[2] | instructionFinish_31[2])
        v0WriteValidVec_res_250 <= _v0WriteValidVec_T_775[2];
      if (_v0WriteValidVec_T_775[3] | instructionFinish_31[3])
        v0WriteValidVec_res_251 <= _v0WriteValidVec_T_775[3];
      if (_v0WriteValidVec_T_775[4] | instructionFinish_31[4])
        v0WriteValidVec_res_252 <= _v0WriteValidVec_T_775[4];
      if (_v0WriteValidVec_T_775[5] | instructionFinish_31[5])
        v0WriteValidVec_res_253 <= _v0WriteValidVec_T_775[5];
      if (_v0WriteValidVec_T_775[6] | instructionFinish_31[6])
        v0WriteValidVec_res_254 <= _v0WriteValidVec_T_775[6];
      if (_v0WriteValidVec_T_775[7] | instructionFinish_31[7])
        v0WriteValidVec_res_255 <= _v0WriteValidVec_T_775[7];
      if (useV0AsMaskToken_updateOH[0] | instructionFinish_0[0])
        useV0AsMaskToken_res <= useV0AsMaskToken_updateOH[0];
      if (useV0AsMaskToken_updateOH[1] | instructionFinish_0[1])
        useV0AsMaskToken_res_1 <= useV0AsMaskToken_updateOH[1];
      if (useV0AsMaskToken_updateOH[2] | instructionFinish_0[2])
        useV0AsMaskToken_res_2 <= useV0AsMaskToken_updateOH[2];
      if (useV0AsMaskToken_updateOH[3] | instructionFinish_0[3])
        useV0AsMaskToken_res_3 <= useV0AsMaskToken_updateOH[3];
      if (useV0AsMaskToken_updateOH[4] | instructionFinish_0[4])
        useV0AsMaskToken_res_4 <= useV0AsMaskToken_updateOH[4];
      if (useV0AsMaskToken_updateOH[5] | instructionFinish_0[5])
        useV0AsMaskToken_res_5 <= useV0AsMaskToken_updateOH[5];
      if (useV0AsMaskToken_updateOH[6] | instructionFinish_0[6])
        useV0AsMaskToken_res_6 <= useV0AsMaskToken_updateOH[6];
      if (useV0AsMaskToken_updateOH[7] | instructionFinish_0[7])
        useV0AsMaskToken_res_7 <= useV0AsMaskToken_updateOH[7];
      if (useV0AsMaskToken_updateOH_1[0] | instructionFinish_1[0])
        useV0AsMaskToken_res_8 <= useV0AsMaskToken_updateOH_1[0];
      if (useV0AsMaskToken_updateOH_1[1] | instructionFinish_1[1])
        useV0AsMaskToken_res_9 <= useV0AsMaskToken_updateOH_1[1];
      if (useV0AsMaskToken_updateOH_1[2] | instructionFinish_1[2])
        useV0AsMaskToken_res_10 <= useV0AsMaskToken_updateOH_1[2];
      if (useV0AsMaskToken_updateOH_1[3] | instructionFinish_1[3])
        useV0AsMaskToken_res_11 <= useV0AsMaskToken_updateOH_1[3];
      if (useV0AsMaskToken_updateOH_1[4] | instructionFinish_1[4])
        useV0AsMaskToken_res_12 <= useV0AsMaskToken_updateOH_1[4];
      if (useV0AsMaskToken_updateOH_1[5] | instructionFinish_1[5])
        useV0AsMaskToken_res_13 <= useV0AsMaskToken_updateOH_1[5];
      if (useV0AsMaskToken_updateOH_1[6] | instructionFinish_1[6])
        useV0AsMaskToken_res_14 <= useV0AsMaskToken_updateOH_1[6];
      if (useV0AsMaskToken_updateOH_1[7] | instructionFinish_1[7])
        useV0AsMaskToken_res_15 <= useV0AsMaskToken_updateOH_1[7];
      if (useV0AsMaskToken_updateOH_2[0] | instructionFinish_2[0])
        useV0AsMaskToken_res_16 <= useV0AsMaskToken_updateOH_2[0];
      if (useV0AsMaskToken_updateOH_2[1] | instructionFinish_2[1])
        useV0AsMaskToken_res_17 <= useV0AsMaskToken_updateOH_2[1];
      if (useV0AsMaskToken_updateOH_2[2] | instructionFinish_2[2])
        useV0AsMaskToken_res_18 <= useV0AsMaskToken_updateOH_2[2];
      if (useV0AsMaskToken_updateOH_2[3] | instructionFinish_2[3])
        useV0AsMaskToken_res_19 <= useV0AsMaskToken_updateOH_2[3];
      if (useV0AsMaskToken_updateOH_2[4] | instructionFinish_2[4])
        useV0AsMaskToken_res_20 <= useV0AsMaskToken_updateOH_2[4];
      if (useV0AsMaskToken_updateOH_2[5] | instructionFinish_2[5])
        useV0AsMaskToken_res_21 <= useV0AsMaskToken_updateOH_2[5];
      if (useV0AsMaskToken_updateOH_2[6] | instructionFinish_2[6])
        useV0AsMaskToken_res_22 <= useV0AsMaskToken_updateOH_2[6];
      if (useV0AsMaskToken_updateOH_2[7] | instructionFinish_2[7])
        useV0AsMaskToken_res_23 <= useV0AsMaskToken_updateOH_2[7];
      if (useV0AsMaskToken_updateOH_3[0] | instructionFinish_3[0])
        useV0AsMaskToken_res_24 <= useV0AsMaskToken_updateOH_3[0];
      if (useV0AsMaskToken_updateOH_3[1] | instructionFinish_3[1])
        useV0AsMaskToken_res_25 <= useV0AsMaskToken_updateOH_3[1];
      if (useV0AsMaskToken_updateOH_3[2] | instructionFinish_3[2])
        useV0AsMaskToken_res_26 <= useV0AsMaskToken_updateOH_3[2];
      if (useV0AsMaskToken_updateOH_3[3] | instructionFinish_3[3])
        useV0AsMaskToken_res_27 <= useV0AsMaskToken_updateOH_3[3];
      if (useV0AsMaskToken_updateOH_3[4] | instructionFinish_3[4])
        useV0AsMaskToken_res_28 <= useV0AsMaskToken_updateOH_3[4];
      if (useV0AsMaskToken_updateOH_3[5] | instructionFinish_3[5])
        useV0AsMaskToken_res_29 <= useV0AsMaskToken_updateOH_3[5];
      if (useV0AsMaskToken_updateOH_3[6] | instructionFinish_3[6])
        useV0AsMaskToken_res_30 <= useV0AsMaskToken_updateOH_3[6];
      if (useV0AsMaskToken_updateOH_3[7] | instructionFinish_3[7])
        useV0AsMaskToken_res_31 <= useV0AsMaskToken_updateOH_3[7];
      if (useV0AsMaskToken_updateOH_4[0] | instructionFinish_4[0])
        useV0AsMaskToken_res_32 <= useV0AsMaskToken_updateOH_4[0];
      if (useV0AsMaskToken_updateOH_4[1] | instructionFinish_4[1])
        useV0AsMaskToken_res_33 <= useV0AsMaskToken_updateOH_4[1];
      if (useV0AsMaskToken_updateOH_4[2] | instructionFinish_4[2])
        useV0AsMaskToken_res_34 <= useV0AsMaskToken_updateOH_4[2];
      if (useV0AsMaskToken_updateOH_4[3] | instructionFinish_4[3])
        useV0AsMaskToken_res_35 <= useV0AsMaskToken_updateOH_4[3];
      if (useV0AsMaskToken_updateOH_4[4] | instructionFinish_4[4])
        useV0AsMaskToken_res_36 <= useV0AsMaskToken_updateOH_4[4];
      if (useV0AsMaskToken_updateOH_4[5] | instructionFinish_4[5])
        useV0AsMaskToken_res_37 <= useV0AsMaskToken_updateOH_4[5];
      if (useV0AsMaskToken_updateOH_4[6] | instructionFinish_4[6])
        useV0AsMaskToken_res_38 <= useV0AsMaskToken_updateOH_4[6];
      if (useV0AsMaskToken_updateOH_4[7] | instructionFinish_4[7])
        useV0AsMaskToken_res_39 <= useV0AsMaskToken_updateOH_4[7];
      if (useV0AsMaskToken_updateOH_5[0] | instructionFinish_5[0])
        useV0AsMaskToken_res_40 <= useV0AsMaskToken_updateOH_5[0];
      if (useV0AsMaskToken_updateOH_5[1] | instructionFinish_5[1])
        useV0AsMaskToken_res_41 <= useV0AsMaskToken_updateOH_5[1];
      if (useV0AsMaskToken_updateOH_5[2] | instructionFinish_5[2])
        useV0AsMaskToken_res_42 <= useV0AsMaskToken_updateOH_5[2];
      if (useV0AsMaskToken_updateOH_5[3] | instructionFinish_5[3])
        useV0AsMaskToken_res_43 <= useV0AsMaskToken_updateOH_5[3];
      if (useV0AsMaskToken_updateOH_5[4] | instructionFinish_5[4])
        useV0AsMaskToken_res_44 <= useV0AsMaskToken_updateOH_5[4];
      if (useV0AsMaskToken_updateOH_5[5] | instructionFinish_5[5])
        useV0AsMaskToken_res_45 <= useV0AsMaskToken_updateOH_5[5];
      if (useV0AsMaskToken_updateOH_5[6] | instructionFinish_5[6])
        useV0AsMaskToken_res_46 <= useV0AsMaskToken_updateOH_5[6];
      if (useV0AsMaskToken_updateOH_5[7] | instructionFinish_5[7])
        useV0AsMaskToken_res_47 <= useV0AsMaskToken_updateOH_5[7];
      if (useV0AsMaskToken_updateOH_6[0] | instructionFinish_6[0])
        useV0AsMaskToken_res_48 <= useV0AsMaskToken_updateOH_6[0];
      if (useV0AsMaskToken_updateOH_6[1] | instructionFinish_6[1])
        useV0AsMaskToken_res_49 <= useV0AsMaskToken_updateOH_6[1];
      if (useV0AsMaskToken_updateOH_6[2] | instructionFinish_6[2])
        useV0AsMaskToken_res_50 <= useV0AsMaskToken_updateOH_6[2];
      if (useV0AsMaskToken_updateOH_6[3] | instructionFinish_6[3])
        useV0AsMaskToken_res_51 <= useV0AsMaskToken_updateOH_6[3];
      if (useV0AsMaskToken_updateOH_6[4] | instructionFinish_6[4])
        useV0AsMaskToken_res_52 <= useV0AsMaskToken_updateOH_6[4];
      if (useV0AsMaskToken_updateOH_6[5] | instructionFinish_6[5])
        useV0AsMaskToken_res_53 <= useV0AsMaskToken_updateOH_6[5];
      if (useV0AsMaskToken_updateOH_6[6] | instructionFinish_6[6])
        useV0AsMaskToken_res_54 <= useV0AsMaskToken_updateOH_6[6];
      if (useV0AsMaskToken_updateOH_6[7] | instructionFinish_6[7])
        useV0AsMaskToken_res_55 <= useV0AsMaskToken_updateOH_6[7];
      if (useV0AsMaskToken_updateOH_7[0] | instructionFinish_7[0])
        useV0AsMaskToken_res_56 <= useV0AsMaskToken_updateOH_7[0];
      if (useV0AsMaskToken_updateOH_7[1] | instructionFinish_7[1])
        useV0AsMaskToken_res_57 <= useV0AsMaskToken_updateOH_7[1];
      if (useV0AsMaskToken_updateOH_7[2] | instructionFinish_7[2])
        useV0AsMaskToken_res_58 <= useV0AsMaskToken_updateOH_7[2];
      if (useV0AsMaskToken_updateOH_7[3] | instructionFinish_7[3])
        useV0AsMaskToken_res_59 <= useV0AsMaskToken_updateOH_7[3];
      if (useV0AsMaskToken_updateOH_7[4] | instructionFinish_7[4])
        useV0AsMaskToken_res_60 <= useV0AsMaskToken_updateOH_7[4];
      if (useV0AsMaskToken_updateOH_7[5] | instructionFinish_7[5])
        useV0AsMaskToken_res_61 <= useV0AsMaskToken_updateOH_7[5];
      if (useV0AsMaskToken_updateOH_7[6] | instructionFinish_7[6])
        useV0AsMaskToken_res_62 <= useV0AsMaskToken_updateOH_7[6];
      if (useV0AsMaskToken_updateOH_7[7] | instructionFinish_7[7])
        useV0AsMaskToken_res_63 <= useV0AsMaskToken_updateOH_7[7];
      if (useV0AsMaskToken_updateOH_8[0] | instructionFinish_8[0])
        useV0AsMaskToken_res_64 <= useV0AsMaskToken_updateOH_8[0];
      if (useV0AsMaskToken_updateOH_8[1] | instructionFinish_8[1])
        useV0AsMaskToken_res_65 <= useV0AsMaskToken_updateOH_8[1];
      if (useV0AsMaskToken_updateOH_8[2] | instructionFinish_8[2])
        useV0AsMaskToken_res_66 <= useV0AsMaskToken_updateOH_8[2];
      if (useV0AsMaskToken_updateOH_8[3] | instructionFinish_8[3])
        useV0AsMaskToken_res_67 <= useV0AsMaskToken_updateOH_8[3];
      if (useV0AsMaskToken_updateOH_8[4] | instructionFinish_8[4])
        useV0AsMaskToken_res_68 <= useV0AsMaskToken_updateOH_8[4];
      if (useV0AsMaskToken_updateOH_8[5] | instructionFinish_8[5])
        useV0AsMaskToken_res_69 <= useV0AsMaskToken_updateOH_8[5];
      if (useV0AsMaskToken_updateOH_8[6] | instructionFinish_8[6])
        useV0AsMaskToken_res_70 <= useV0AsMaskToken_updateOH_8[6];
      if (useV0AsMaskToken_updateOH_8[7] | instructionFinish_8[7])
        useV0AsMaskToken_res_71 <= useV0AsMaskToken_updateOH_8[7];
      if (useV0AsMaskToken_updateOH_9[0] | instructionFinish_9[0])
        useV0AsMaskToken_res_72 <= useV0AsMaskToken_updateOH_9[0];
      if (useV0AsMaskToken_updateOH_9[1] | instructionFinish_9[1])
        useV0AsMaskToken_res_73 <= useV0AsMaskToken_updateOH_9[1];
      if (useV0AsMaskToken_updateOH_9[2] | instructionFinish_9[2])
        useV0AsMaskToken_res_74 <= useV0AsMaskToken_updateOH_9[2];
      if (useV0AsMaskToken_updateOH_9[3] | instructionFinish_9[3])
        useV0AsMaskToken_res_75 <= useV0AsMaskToken_updateOH_9[3];
      if (useV0AsMaskToken_updateOH_9[4] | instructionFinish_9[4])
        useV0AsMaskToken_res_76 <= useV0AsMaskToken_updateOH_9[4];
      if (useV0AsMaskToken_updateOH_9[5] | instructionFinish_9[5])
        useV0AsMaskToken_res_77 <= useV0AsMaskToken_updateOH_9[5];
      if (useV0AsMaskToken_updateOH_9[6] | instructionFinish_9[6])
        useV0AsMaskToken_res_78 <= useV0AsMaskToken_updateOH_9[6];
      if (useV0AsMaskToken_updateOH_9[7] | instructionFinish_9[7])
        useV0AsMaskToken_res_79 <= useV0AsMaskToken_updateOH_9[7];
      if (useV0AsMaskToken_updateOH_10[0] | instructionFinish_10[0])
        useV0AsMaskToken_res_80 <= useV0AsMaskToken_updateOH_10[0];
      if (useV0AsMaskToken_updateOH_10[1] | instructionFinish_10[1])
        useV0AsMaskToken_res_81 <= useV0AsMaskToken_updateOH_10[1];
      if (useV0AsMaskToken_updateOH_10[2] | instructionFinish_10[2])
        useV0AsMaskToken_res_82 <= useV0AsMaskToken_updateOH_10[2];
      if (useV0AsMaskToken_updateOH_10[3] | instructionFinish_10[3])
        useV0AsMaskToken_res_83 <= useV0AsMaskToken_updateOH_10[3];
      if (useV0AsMaskToken_updateOH_10[4] | instructionFinish_10[4])
        useV0AsMaskToken_res_84 <= useV0AsMaskToken_updateOH_10[4];
      if (useV0AsMaskToken_updateOH_10[5] | instructionFinish_10[5])
        useV0AsMaskToken_res_85 <= useV0AsMaskToken_updateOH_10[5];
      if (useV0AsMaskToken_updateOH_10[6] | instructionFinish_10[6])
        useV0AsMaskToken_res_86 <= useV0AsMaskToken_updateOH_10[6];
      if (useV0AsMaskToken_updateOH_10[7] | instructionFinish_10[7])
        useV0AsMaskToken_res_87 <= useV0AsMaskToken_updateOH_10[7];
      if (useV0AsMaskToken_updateOH_11[0] | instructionFinish_11[0])
        useV0AsMaskToken_res_88 <= useV0AsMaskToken_updateOH_11[0];
      if (useV0AsMaskToken_updateOH_11[1] | instructionFinish_11[1])
        useV0AsMaskToken_res_89 <= useV0AsMaskToken_updateOH_11[1];
      if (useV0AsMaskToken_updateOH_11[2] | instructionFinish_11[2])
        useV0AsMaskToken_res_90 <= useV0AsMaskToken_updateOH_11[2];
      if (useV0AsMaskToken_updateOH_11[3] | instructionFinish_11[3])
        useV0AsMaskToken_res_91 <= useV0AsMaskToken_updateOH_11[3];
      if (useV0AsMaskToken_updateOH_11[4] | instructionFinish_11[4])
        useV0AsMaskToken_res_92 <= useV0AsMaskToken_updateOH_11[4];
      if (useV0AsMaskToken_updateOH_11[5] | instructionFinish_11[5])
        useV0AsMaskToken_res_93 <= useV0AsMaskToken_updateOH_11[5];
      if (useV0AsMaskToken_updateOH_11[6] | instructionFinish_11[6])
        useV0AsMaskToken_res_94 <= useV0AsMaskToken_updateOH_11[6];
      if (useV0AsMaskToken_updateOH_11[7] | instructionFinish_11[7])
        useV0AsMaskToken_res_95 <= useV0AsMaskToken_updateOH_11[7];
      if (useV0AsMaskToken_updateOH_12[0] | instructionFinish_12[0])
        useV0AsMaskToken_res_96 <= useV0AsMaskToken_updateOH_12[0];
      if (useV0AsMaskToken_updateOH_12[1] | instructionFinish_12[1])
        useV0AsMaskToken_res_97 <= useV0AsMaskToken_updateOH_12[1];
      if (useV0AsMaskToken_updateOH_12[2] | instructionFinish_12[2])
        useV0AsMaskToken_res_98 <= useV0AsMaskToken_updateOH_12[2];
      if (useV0AsMaskToken_updateOH_12[3] | instructionFinish_12[3])
        useV0AsMaskToken_res_99 <= useV0AsMaskToken_updateOH_12[3];
      if (useV0AsMaskToken_updateOH_12[4] | instructionFinish_12[4])
        useV0AsMaskToken_res_100 <= useV0AsMaskToken_updateOH_12[4];
      if (useV0AsMaskToken_updateOH_12[5] | instructionFinish_12[5])
        useV0AsMaskToken_res_101 <= useV0AsMaskToken_updateOH_12[5];
      if (useV0AsMaskToken_updateOH_12[6] | instructionFinish_12[6])
        useV0AsMaskToken_res_102 <= useV0AsMaskToken_updateOH_12[6];
      if (useV0AsMaskToken_updateOH_12[7] | instructionFinish_12[7])
        useV0AsMaskToken_res_103 <= useV0AsMaskToken_updateOH_12[7];
      if (useV0AsMaskToken_updateOH_13[0] | instructionFinish_13[0])
        useV0AsMaskToken_res_104 <= useV0AsMaskToken_updateOH_13[0];
      if (useV0AsMaskToken_updateOH_13[1] | instructionFinish_13[1])
        useV0AsMaskToken_res_105 <= useV0AsMaskToken_updateOH_13[1];
      if (useV0AsMaskToken_updateOH_13[2] | instructionFinish_13[2])
        useV0AsMaskToken_res_106 <= useV0AsMaskToken_updateOH_13[2];
      if (useV0AsMaskToken_updateOH_13[3] | instructionFinish_13[3])
        useV0AsMaskToken_res_107 <= useV0AsMaskToken_updateOH_13[3];
      if (useV0AsMaskToken_updateOH_13[4] | instructionFinish_13[4])
        useV0AsMaskToken_res_108 <= useV0AsMaskToken_updateOH_13[4];
      if (useV0AsMaskToken_updateOH_13[5] | instructionFinish_13[5])
        useV0AsMaskToken_res_109 <= useV0AsMaskToken_updateOH_13[5];
      if (useV0AsMaskToken_updateOH_13[6] | instructionFinish_13[6])
        useV0AsMaskToken_res_110 <= useV0AsMaskToken_updateOH_13[6];
      if (useV0AsMaskToken_updateOH_13[7] | instructionFinish_13[7])
        useV0AsMaskToken_res_111 <= useV0AsMaskToken_updateOH_13[7];
      if (useV0AsMaskToken_updateOH_14[0] | instructionFinish_14[0])
        useV0AsMaskToken_res_112 <= useV0AsMaskToken_updateOH_14[0];
      if (useV0AsMaskToken_updateOH_14[1] | instructionFinish_14[1])
        useV0AsMaskToken_res_113 <= useV0AsMaskToken_updateOH_14[1];
      if (useV0AsMaskToken_updateOH_14[2] | instructionFinish_14[2])
        useV0AsMaskToken_res_114 <= useV0AsMaskToken_updateOH_14[2];
      if (useV0AsMaskToken_updateOH_14[3] | instructionFinish_14[3])
        useV0AsMaskToken_res_115 <= useV0AsMaskToken_updateOH_14[3];
      if (useV0AsMaskToken_updateOH_14[4] | instructionFinish_14[4])
        useV0AsMaskToken_res_116 <= useV0AsMaskToken_updateOH_14[4];
      if (useV0AsMaskToken_updateOH_14[5] | instructionFinish_14[5])
        useV0AsMaskToken_res_117 <= useV0AsMaskToken_updateOH_14[5];
      if (useV0AsMaskToken_updateOH_14[6] | instructionFinish_14[6])
        useV0AsMaskToken_res_118 <= useV0AsMaskToken_updateOH_14[6];
      if (useV0AsMaskToken_updateOH_14[7] | instructionFinish_14[7])
        useV0AsMaskToken_res_119 <= useV0AsMaskToken_updateOH_14[7];
      if (useV0AsMaskToken_updateOH_15[0] | instructionFinish_15[0])
        useV0AsMaskToken_res_120 <= useV0AsMaskToken_updateOH_15[0];
      if (useV0AsMaskToken_updateOH_15[1] | instructionFinish_15[1])
        useV0AsMaskToken_res_121 <= useV0AsMaskToken_updateOH_15[1];
      if (useV0AsMaskToken_updateOH_15[2] | instructionFinish_15[2])
        useV0AsMaskToken_res_122 <= useV0AsMaskToken_updateOH_15[2];
      if (useV0AsMaskToken_updateOH_15[3] | instructionFinish_15[3])
        useV0AsMaskToken_res_123 <= useV0AsMaskToken_updateOH_15[3];
      if (useV0AsMaskToken_updateOH_15[4] | instructionFinish_15[4])
        useV0AsMaskToken_res_124 <= useV0AsMaskToken_updateOH_15[4];
      if (useV0AsMaskToken_updateOH_15[5] | instructionFinish_15[5])
        useV0AsMaskToken_res_125 <= useV0AsMaskToken_updateOH_15[5];
      if (useV0AsMaskToken_updateOH_15[6] | instructionFinish_15[6])
        useV0AsMaskToken_res_126 <= useV0AsMaskToken_updateOH_15[6];
      if (useV0AsMaskToken_updateOH_15[7] | instructionFinish_15[7])
        useV0AsMaskToken_res_127 <= useV0AsMaskToken_updateOH_15[7];
      if (useV0AsMaskToken_updateOH_16[0] | instructionFinish_16[0])
        useV0AsMaskToken_res_128 <= useV0AsMaskToken_updateOH_16[0];
      if (useV0AsMaskToken_updateOH_16[1] | instructionFinish_16[1])
        useV0AsMaskToken_res_129 <= useV0AsMaskToken_updateOH_16[1];
      if (useV0AsMaskToken_updateOH_16[2] | instructionFinish_16[2])
        useV0AsMaskToken_res_130 <= useV0AsMaskToken_updateOH_16[2];
      if (useV0AsMaskToken_updateOH_16[3] | instructionFinish_16[3])
        useV0AsMaskToken_res_131 <= useV0AsMaskToken_updateOH_16[3];
      if (useV0AsMaskToken_updateOH_16[4] | instructionFinish_16[4])
        useV0AsMaskToken_res_132 <= useV0AsMaskToken_updateOH_16[4];
      if (useV0AsMaskToken_updateOH_16[5] | instructionFinish_16[5])
        useV0AsMaskToken_res_133 <= useV0AsMaskToken_updateOH_16[5];
      if (useV0AsMaskToken_updateOH_16[6] | instructionFinish_16[6])
        useV0AsMaskToken_res_134 <= useV0AsMaskToken_updateOH_16[6];
      if (useV0AsMaskToken_updateOH_16[7] | instructionFinish_16[7])
        useV0AsMaskToken_res_135 <= useV0AsMaskToken_updateOH_16[7];
      if (useV0AsMaskToken_updateOH_17[0] | instructionFinish_17[0])
        useV0AsMaskToken_res_136 <= useV0AsMaskToken_updateOH_17[0];
      if (useV0AsMaskToken_updateOH_17[1] | instructionFinish_17[1])
        useV0AsMaskToken_res_137 <= useV0AsMaskToken_updateOH_17[1];
      if (useV0AsMaskToken_updateOH_17[2] | instructionFinish_17[2])
        useV0AsMaskToken_res_138 <= useV0AsMaskToken_updateOH_17[2];
      if (useV0AsMaskToken_updateOH_17[3] | instructionFinish_17[3])
        useV0AsMaskToken_res_139 <= useV0AsMaskToken_updateOH_17[3];
      if (useV0AsMaskToken_updateOH_17[4] | instructionFinish_17[4])
        useV0AsMaskToken_res_140 <= useV0AsMaskToken_updateOH_17[4];
      if (useV0AsMaskToken_updateOH_17[5] | instructionFinish_17[5])
        useV0AsMaskToken_res_141 <= useV0AsMaskToken_updateOH_17[5];
      if (useV0AsMaskToken_updateOH_17[6] | instructionFinish_17[6])
        useV0AsMaskToken_res_142 <= useV0AsMaskToken_updateOH_17[6];
      if (useV0AsMaskToken_updateOH_17[7] | instructionFinish_17[7])
        useV0AsMaskToken_res_143 <= useV0AsMaskToken_updateOH_17[7];
      if (useV0AsMaskToken_updateOH_18[0] | instructionFinish_18[0])
        useV0AsMaskToken_res_144 <= useV0AsMaskToken_updateOH_18[0];
      if (useV0AsMaskToken_updateOH_18[1] | instructionFinish_18[1])
        useV0AsMaskToken_res_145 <= useV0AsMaskToken_updateOH_18[1];
      if (useV0AsMaskToken_updateOH_18[2] | instructionFinish_18[2])
        useV0AsMaskToken_res_146 <= useV0AsMaskToken_updateOH_18[2];
      if (useV0AsMaskToken_updateOH_18[3] | instructionFinish_18[3])
        useV0AsMaskToken_res_147 <= useV0AsMaskToken_updateOH_18[3];
      if (useV0AsMaskToken_updateOH_18[4] | instructionFinish_18[4])
        useV0AsMaskToken_res_148 <= useV0AsMaskToken_updateOH_18[4];
      if (useV0AsMaskToken_updateOH_18[5] | instructionFinish_18[5])
        useV0AsMaskToken_res_149 <= useV0AsMaskToken_updateOH_18[5];
      if (useV0AsMaskToken_updateOH_18[6] | instructionFinish_18[6])
        useV0AsMaskToken_res_150 <= useV0AsMaskToken_updateOH_18[6];
      if (useV0AsMaskToken_updateOH_18[7] | instructionFinish_18[7])
        useV0AsMaskToken_res_151 <= useV0AsMaskToken_updateOH_18[7];
      if (useV0AsMaskToken_updateOH_19[0] | instructionFinish_19[0])
        useV0AsMaskToken_res_152 <= useV0AsMaskToken_updateOH_19[0];
      if (useV0AsMaskToken_updateOH_19[1] | instructionFinish_19[1])
        useV0AsMaskToken_res_153 <= useV0AsMaskToken_updateOH_19[1];
      if (useV0AsMaskToken_updateOH_19[2] | instructionFinish_19[2])
        useV0AsMaskToken_res_154 <= useV0AsMaskToken_updateOH_19[2];
      if (useV0AsMaskToken_updateOH_19[3] | instructionFinish_19[3])
        useV0AsMaskToken_res_155 <= useV0AsMaskToken_updateOH_19[3];
      if (useV0AsMaskToken_updateOH_19[4] | instructionFinish_19[4])
        useV0AsMaskToken_res_156 <= useV0AsMaskToken_updateOH_19[4];
      if (useV0AsMaskToken_updateOH_19[5] | instructionFinish_19[5])
        useV0AsMaskToken_res_157 <= useV0AsMaskToken_updateOH_19[5];
      if (useV0AsMaskToken_updateOH_19[6] | instructionFinish_19[6])
        useV0AsMaskToken_res_158 <= useV0AsMaskToken_updateOH_19[6];
      if (useV0AsMaskToken_updateOH_19[7] | instructionFinish_19[7])
        useV0AsMaskToken_res_159 <= useV0AsMaskToken_updateOH_19[7];
      if (useV0AsMaskToken_updateOH_20[0] | instructionFinish_20[0])
        useV0AsMaskToken_res_160 <= useV0AsMaskToken_updateOH_20[0];
      if (useV0AsMaskToken_updateOH_20[1] | instructionFinish_20[1])
        useV0AsMaskToken_res_161 <= useV0AsMaskToken_updateOH_20[1];
      if (useV0AsMaskToken_updateOH_20[2] | instructionFinish_20[2])
        useV0AsMaskToken_res_162 <= useV0AsMaskToken_updateOH_20[2];
      if (useV0AsMaskToken_updateOH_20[3] | instructionFinish_20[3])
        useV0AsMaskToken_res_163 <= useV0AsMaskToken_updateOH_20[3];
      if (useV0AsMaskToken_updateOH_20[4] | instructionFinish_20[4])
        useV0AsMaskToken_res_164 <= useV0AsMaskToken_updateOH_20[4];
      if (useV0AsMaskToken_updateOH_20[5] | instructionFinish_20[5])
        useV0AsMaskToken_res_165 <= useV0AsMaskToken_updateOH_20[5];
      if (useV0AsMaskToken_updateOH_20[6] | instructionFinish_20[6])
        useV0AsMaskToken_res_166 <= useV0AsMaskToken_updateOH_20[6];
      if (useV0AsMaskToken_updateOH_20[7] | instructionFinish_20[7])
        useV0AsMaskToken_res_167 <= useV0AsMaskToken_updateOH_20[7];
      if (useV0AsMaskToken_updateOH_21[0] | instructionFinish_21[0])
        useV0AsMaskToken_res_168 <= useV0AsMaskToken_updateOH_21[0];
      if (useV0AsMaskToken_updateOH_21[1] | instructionFinish_21[1])
        useV0AsMaskToken_res_169 <= useV0AsMaskToken_updateOH_21[1];
      if (useV0AsMaskToken_updateOH_21[2] | instructionFinish_21[2])
        useV0AsMaskToken_res_170 <= useV0AsMaskToken_updateOH_21[2];
      if (useV0AsMaskToken_updateOH_21[3] | instructionFinish_21[3])
        useV0AsMaskToken_res_171 <= useV0AsMaskToken_updateOH_21[3];
      if (useV0AsMaskToken_updateOH_21[4] | instructionFinish_21[4])
        useV0AsMaskToken_res_172 <= useV0AsMaskToken_updateOH_21[4];
      if (useV0AsMaskToken_updateOH_21[5] | instructionFinish_21[5])
        useV0AsMaskToken_res_173 <= useV0AsMaskToken_updateOH_21[5];
      if (useV0AsMaskToken_updateOH_21[6] | instructionFinish_21[6])
        useV0AsMaskToken_res_174 <= useV0AsMaskToken_updateOH_21[6];
      if (useV0AsMaskToken_updateOH_21[7] | instructionFinish_21[7])
        useV0AsMaskToken_res_175 <= useV0AsMaskToken_updateOH_21[7];
      if (useV0AsMaskToken_updateOH_22[0] | instructionFinish_22[0])
        useV0AsMaskToken_res_176 <= useV0AsMaskToken_updateOH_22[0];
      if (useV0AsMaskToken_updateOH_22[1] | instructionFinish_22[1])
        useV0AsMaskToken_res_177 <= useV0AsMaskToken_updateOH_22[1];
      if (useV0AsMaskToken_updateOH_22[2] | instructionFinish_22[2])
        useV0AsMaskToken_res_178 <= useV0AsMaskToken_updateOH_22[2];
      if (useV0AsMaskToken_updateOH_22[3] | instructionFinish_22[3])
        useV0AsMaskToken_res_179 <= useV0AsMaskToken_updateOH_22[3];
      if (useV0AsMaskToken_updateOH_22[4] | instructionFinish_22[4])
        useV0AsMaskToken_res_180 <= useV0AsMaskToken_updateOH_22[4];
      if (useV0AsMaskToken_updateOH_22[5] | instructionFinish_22[5])
        useV0AsMaskToken_res_181 <= useV0AsMaskToken_updateOH_22[5];
      if (useV0AsMaskToken_updateOH_22[6] | instructionFinish_22[6])
        useV0AsMaskToken_res_182 <= useV0AsMaskToken_updateOH_22[6];
      if (useV0AsMaskToken_updateOH_22[7] | instructionFinish_22[7])
        useV0AsMaskToken_res_183 <= useV0AsMaskToken_updateOH_22[7];
      if (useV0AsMaskToken_updateOH_23[0] | instructionFinish_23[0])
        useV0AsMaskToken_res_184 <= useV0AsMaskToken_updateOH_23[0];
      if (useV0AsMaskToken_updateOH_23[1] | instructionFinish_23[1])
        useV0AsMaskToken_res_185 <= useV0AsMaskToken_updateOH_23[1];
      if (useV0AsMaskToken_updateOH_23[2] | instructionFinish_23[2])
        useV0AsMaskToken_res_186 <= useV0AsMaskToken_updateOH_23[2];
      if (useV0AsMaskToken_updateOH_23[3] | instructionFinish_23[3])
        useV0AsMaskToken_res_187 <= useV0AsMaskToken_updateOH_23[3];
      if (useV0AsMaskToken_updateOH_23[4] | instructionFinish_23[4])
        useV0AsMaskToken_res_188 <= useV0AsMaskToken_updateOH_23[4];
      if (useV0AsMaskToken_updateOH_23[5] | instructionFinish_23[5])
        useV0AsMaskToken_res_189 <= useV0AsMaskToken_updateOH_23[5];
      if (useV0AsMaskToken_updateOH_23[6] | instructionFinish_23[6])
        useV0AsMaskToken_res_190 <= useV0AsMaskToken_updateOH_23[6];
      if (useV0AsMaskToken_updateOH_23[7] | instructionFinish_23[7])
        useV0AsMaskToken_res_191 <= useV0AsMaskToken_updateOH_23[7];
      if (useV0AsMaskToken_updateOH_24[0] | instructionFinish_24[0])
        useV0AsMaskToken_res_192 <= useV0AsMaskToken_updateOH_24[0];
      if (useV0AsMaskToken_updateOH_24[1] | instructionFinish_24[1])
        useV0AsMaskToken_res_193 <= useV0AsMaskToken_updateOH_24[1];
      if (useV0AsMaskToken_updateOH_24[2] | instructionFinish_24[2])
        useV0AsMaskToken_res_194 <= useV0AsMaskToken_updateOH_24[2];
      if (useV0AsMaskToken_updateOH_24[3] | instructionFinish_24[3])
        useV0AsMaskToken_res_195 <= useV0AsMaskToken_updateOH_24[3];
      if (useV0AsMaskToken_updateOH_24[4] | instructionFinish_24[4])
        useV0AsMaskToken_res_196 <= useV0AsMaskToken_updateOH_24[4];
      if (useV0AsMaskToken_updateOH_24[5] | instructionFinish_24[5])
        useV0AsMaskToken_res_197 <= useV0AsMaskToken_updateOH_24[5];
      if (useV0AsMaskToken_updateOH_24[6] | instructionFinish_24[6])
        useV0AsMaskToken_res_198 <= useV0AsMaskToken_updateOH_24[6];
      if (useV0AsMaskToken_updateOH_24[7] | instructionFinish_24[7])
        useV0AsMaskToken_res_199 <= useV0AsMaskToken_updateOH_24[7];
      if (useV0AsMaskToken_updateOH_25[0] | instructionFinish_25[0])
        useV0AsMaskToken_res_200 <= useV0AsMaskToken_updateOH_25[0];
      if (useV0AsMaskToken_updateOH_25[1] | instructionFinish_25[1])
        useV0AsMaskToken_res_201 <= useV0AsMaskToken_updateOH_25[1];
      if (useV0AsMaskToken_updateOH_25[2] | instructionFinish_25[2])
        useV0AsMaskToken_res_202 <= useV0AsMaskToken_updateOH_25[2];
      if (useV0AsMaskToken_updateOH_25[3] | instructionFinish_25[3])
        useV0AsMaskToken_res_203 <= useV0AsMaskToken_updateOH_25[3];
      if (useV0AsMaskToken_updateOH_25[4] | instructionFinish_25[4])
        useV0AsMaskToken_res_204 <= useV0AsMaskToken_updateOH_25[4];
      if (useV0AsMaskToken_updateOH_25[5] | instructionFinish_25[5])
        useV0AsMaskToken_res_205 <= useV0AsMaskToken_updateOH_25[5];
      if (useV0AsMaskToken_updateOH_25[6] | instructionFinish_25[6])
        useV0AsMaskToken_res_206 <= useV0AsMaskToken_updateOH_25[6];
      if (useV0AsMaskToken_updateOH_25[7] | instructionFinish_25[7])
        useV0AsMaskToken_res_207 <= useV0AsMaskToken_updateOH_25[7];
      if (useV0AsMaskToken_updateOH_26[0] | instructionFinish_26[0])
        useV0AsMaskToken_res_208 <= useV0AsMaskToken_updateOH_26[0];
      if (useV0AsMaskToken_updateOH_26[1] | instructionFinish_26[1])
        useV0AsMaskToken_res_209 <= useV0AsMaskToken_updateOH_26[1];
      if (useV0AsMaskToken_updateOH_26[2] | instructionFinish_26[2])
        useV0AsMaskToken_res_210 <= useV0AsMaskToken_updateOH_26[2];
      if (useV0AsMaskToken_updateOH_26[3] | instructionFinish_26[3])
        useV0AsMaskToken_res_211 <= useV0AsMaskToken_updateOH_26[3];
      if (useV0AsMaskToken_updateOH_26[4] | instructionFinish_26[4])
        useV0AsMaskToken_res_212 <= useV0AsMaskToken_updateOH_26[4];
      if (useV0AsMaskToken_updateOH_26[5] | instructionFinish_26[5])
        useV0AsMaskToken_res_213 <= useV0AsMaskToken_updateOH_26[5];
      if (useV0AsMaskToken_updateOH_26[6] | instructionFinish_26[6])
        useV0AsMaskToken_res_214 <= useV0AsMaskToken_updateOH_26[6];
      if (useV0AsMaskToken_updateOH_26[7] | instructionFinish_26[7])
        useV0AsMaskToken_res_215 <= useV0AsMaskToken_updateOH_26[7];
      if (useV0AsMaskToken_updateOH_27[0] | instructionFinish_27[0])
        useV0AsMaskToken_res_216 <= useV0AsMaskToken_updateOH_27[0];
      if (useV0AsMaskToken_updateOH_27[1] | instructionFinish_27[1])
        useV0AsMaskToken_res_217 <= useV0AsMaskToken_updateOH_27[1];
      if (useV0AsMaskToken_updateOH_27[2] | instructionFinish_27[2])
        useV0AsMaskToken_res_218 <= useV0AsMaskToken_updateOH_27[2];
      if (useV0AsMaskToken_updateOH_27[3] | instructionFinish_27[3])
        useV0AsMaskToken_res_219 <= useV0AsMaskToken_updateOH_27[3];
      if (useV0AsMaskToken_updateOH_27[4] | instructionFinish_27[4])
        useV0AsMaskToken_res_220 <= useV0AsMaskToken_updateOH_27[4];
      if (useV0AsMaskToken_updateOH_27[5] | instructionFinish_27[5])
        useV0AsMaskToken_res_221 <= useV0AsMaskToken_updateOH_27[5];
      if (useV0AsMaskToken_updateOH_27[6] | instructionFinish_27[6])
        useV0AsMaskToken_res_222 <= useV0AsMaskToken_updateOH_27[6];
      if (useV0AsMaskToken_updateOH_27[7] | instructionFinish_27[7])
        useV0AsMaskToken_res_223 <= useV0AsMaskToken_updateOH_27[7];
      if (useV0AsMaskToken_updateOH_28[0] | instructionFinish_28[0])
        useV0AsMaskToken_res_224 <= useV0AsMaskToken_updateOH_28[0];
      if (useV0AsMaskToken_updateOH_28[1] | instructionFinish_28[1])
        useV0AsMaskToken_res_225 <= useV0AsMaskToken_updateOH_28[1];
      if (useV0AsMaskToken_updateOH_28[2] | instructionFinish_28[2])
        useV0AsMaskToken_res_226 <= useV0AsMaskToken_updateOH_28[2];
      if (useV0AsMaskToken_updateOH_28[3] | instructionFinish_28[3])
        useV0AsMaskToken_res_227 <= useV0AsMaskToken_updateOH_28[3];
      if (useV0AsMaskToken_updateOH_28[4] | instructionFinish_28[4])
        useV0AsMaskToken_res_228 <= useV0AsMaskToken_updateOH_28[4];
      if (useV0AsMaskToken_updateOH_28[5] | instructionFinish_28[5])
        useV0AsMaskToken_res_229 <= useV0AsMaskToken_updateOH_28[5];
      if (useV0AsMaskToken_updateOH_28[6] | instructionFinish_28[6])
        useV0AsMaskToken_res_230 <= useV0AsMaskToken_updateOH_28[6];
      if (useV0AsMaskToken_updateOH_28[7] | instructionFinish_28[7])
        useV0AsMaskToken_res_231 <= useV0AsMaskToken_updateOH_28[7];
      if (useV0AsMaskToken_updateOH_29[0] | instructionFinish_29[0])
        useV0AsMaskToken_res_232 <= useV0AsMaskToken_updateOH_29[0];
      if (useV0AsMaskToken_updateOH_29[1] | instructionFinish_29[1])
        useV0AsMaskToken_res_233 <= useV0AsMaskToken_updateOH_29[1];
      if (useV0AsMaskToken_updateOH_29[2] | instructionFinish_29[2])
        useV0AsMaskToken_res_234 <= useV0AsMaskToken_updateOH_29[2];
      if (useV0AsMaskToken_updateOH_29[3] | instructionFinish_29[3])
        useV0AsMaskToken_res_235 <= useV0AsMaskToken_updateOH_29[3];
      if (useV0AsMaskToken_updateOH_29[4] | instructionFinish_29[4])
        useV0AsMaskToken_res_236 <= useV0AsMaskToken_updateOH_29[4];
      if (useV0AsMaskToken_updateOH_29[5] | instructionFinish_29[5])
        useV0AsMaskToken_res_237 <= useV0AsMaskToken_updateOH_29[5];
      if (useV0AsMaskToken_updateOH_29[6] | instructionFinish_29[6])
        useV0AsMaskToken_res_238 <= useV0AsMaskToken_updateOH_29[6];
      if (useV0AsMaskToken_updateOH_29[7] | instructionFinish_29[7])
        useV0AsMaskToken_res_239 <= useV0AsMaskToken_updateOH_29[7];
      if (useV0AsMaskToken_updateOH_30[0] | instructionFinish_30[0])
        useV0AsMaskToken_res_240 <= useV0AsMaskToken_updateOH_30[0];
      if (useV0AsMaskToken_updateOH_30[1] | instructionFinish_30[1])
        useV0AsMaskToken_res_241 <= useV0AsMaskToken_updateOH_30[1];
      if (useV0AsMaskToken_updateOH_30[2] | instructionFinish_30[2])
        useV0AsMaskToken_res_242 <= useV0AsMaskToken_updateOH_30[2];
      if (useV0AsMaskToken_updateOH_30[3] | instructionFinish_30[3])
        useV0AsMaskToken_res_243 <= useV0AsMaskToken_updateOH_30[3];
      if (useV0AsMaskToken_updateOH_30[4] | instructionFinish_30[4])
        useV0AsMaskToken_res_244 <= useV0AsMaskToken_updateOH_30[4];
      if (useV0AsMaskToken_updateOH_30[5] | instructionFinish_30[5])
        useV0AsMaskToken_res_245 <= useV0AsMaskToken_updateOH_30[5];
      if (useV0AsMaskToken_updateOH_30[6] | instructionFinish_30[6])
        useV0AsMaskToken_res_246 <= useV0AsMaskToken_updateOH_30[6];
      if (useV0AsMaskToken_updateOH_30[7] | instructionFinish_30[7])
        useV0AsMaskToken_res_247 <= useV0AsMaskToken_updateOH_30[7];
      if (useV0AsMaskToken_updateOH_31[0] | instructionFinish_31[0])
        useV0AsMaskToken_res_248 <= useV0AsMaskToken_updateOH_31[0];
      if (useV0AsMaskToken_updateOH_31[1] | instructionFinish_31[1])
        useV0AsMaskToken_res_249 <= useV0AsMaskToken_updateOH_31[1];
      if (useV0AsMaskToken_updateOH_31[2] | instructionFinish_31[2])
        useV0AsMaskToken_res_250 <= useV0AsMaskToken_updateOH_31[2];
      if (useV0AsMaskToken_updateOH_31[3] | instructionFinish_31[3])
        useV0AsMaskToken_res_251 <= useV0AsMaskToken_updateOH_31[3];
      if (useV0AsMaskToken_updateOH_31[4] | instructionFinish_31[4])
        useV0AsMaskToken_res_252 <= useV0AsMaskToken_updateOH_31[4];
      if (useV0AsMaskToken_updateOH_31[5] | instructionFinish_31[5])
        useV0AsMaskToken_res_253 <= useV0AsMaskToken_updateOH_31[5];
      if (useV0AsMaskToken_updateOH_31[6] | instructionFinish_31[6])
        useV0AsMaskToken_res_254 <= useV0AsMaskToken_updateOH_31[6];
      if (useV0AsMaskToken_updateOH_31[7] | instructionFinish_31[7])
        useV0AsMaskToken_res_255 <= useV0AsMaskToken_updateOH_31[7];
      if (maskUnitWriteV0_set | maskUnitFree)
        maskUnitWriteV0 <= maskUnitWriteV0_set;
    end
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:16];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [4:0] i = 5'h0; i < 5'h11; i += 5'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        v0WriteValidVec_res = _RANDOM[5'h0][0];
        v0WriteValidVec_res_1 = _RANDOM[5'h0][1];
        v0WriteValidVec_res_2 = _RANDOM[5'h0][2];
        v0WriteValidVec_res_3 = _RANDOM[5'h0][3];
        v0WriteValidVec_res_4 = _RANDOM[5'h0][4];
        v0WriteValidVec_res_5 = _RANDOM[5'h0][5];
        v0WriteValidVec_res_6 = _RANDOM[5'h0][6];
        v0WriteValidVec_res_7 = _RANDOM[5'h0][7];
        v0WriteValidVec_res_8 = _RANDOM[5'h0][8];
        v0WriteValidVec_res_9 = _RANDOM[5'h0][9];
        v0WriteValidVec_res_10 = _RANDOM[5'h0][10];
        v0WriteValidVec_res_11 = _RANDOM[5'h0][11];
        v0WriteValidVec_res_12 = _RANDOM[5'h0][12];
        v0WriteValidVec_res_13 = _RANDOM[5'h0][13];
        v0WriteValidVec_res_14 = _RANDOM[5'h0][14];
        v0WriteValidVec_res_15 = _RANDOM[5'h0][15];
        v0WriteValidVec_res_16 = _RANDOM[5'h0][16];
        v0WriteValidVec_res_17 = _RANDOM[5'h0][17];
        v0WriteValidVec_res_18 = _RANDOM[5'h0][18];
        v0WriteValidVec_res_19 = _RANDOM[5'h0][19];
        v0WriteValidVec_res_20 = _RANDOM[5'h0][20];
        v0WriteValidVec_res_21 = _RANDOM[5'h0][21];
        v0WriteValidVec_res_22 = _RANDOM[5'h0][22];
        v0WriteValidVec_res_23 = _RANDOM[5'h0][23];
        v0WriteValidVec_res_24 = _RANDOM[5'h0][24];
        v0WriteValidVec_res_25 = _RANDOM[5'h0][25];
        v0WriteValidVec_res_26 = _RANDOM[5'h0][26];
        v0WriteValidVec_res_27 = _RANDOM[5'h0][27];
        v0WriteValidVec_res_28 = _RANDOM[5'h0][28];
        v0WriteValidVec_res_29 = _RANDOM[5'h0][29];
        v0WriteValidVec_res_30 = _RANDOM[5'h0][30];
        v0WriteValidVec_res_31 = _RANDOM[5'h0][31];
        v0WriteValidVec_res_32 = _RANDOM[5'h1][0];
        v0WriteValidVec_res_33 = _RANDOM[5'h1][1];
        v0WriteValidVec_res_34 = _RANDOM[5'h1][2];
        v0WriteValidVec_res_35 = _RANDOM[5'h1][3];
        v0WriteValidVec_res_36 = _RANDOM[5'h1][4];
        v0WriteValidVec_res_37 = _RANDOM[5'h1][5];
        v0WriteValidVec_res_38 = _RANDOM[5'h1][6];
        v0WriteValidVec_res_39 = _RANDOM[5'h1][7];
        v0WriteValidVec_res_40 = _RANDOM[5'h1][8];
        v0WriteValidVec_res_41 = _RANDOM[5'h1][9];
        v0WriteValidVec_res_42 = _RANDOM[5'h1][10];
        v0WriteValidVec_res_43 = _RANDOM[5'h1][11];
        v0WriteValidVec_res_44 = _RANDOM[5'h1][12];
        v0WriteValidVec_res_45 = _RANDOM[5'h1][13];
        v0WriteValidVec_res_46 = _RANDOM[5'h1][14];
        v0WriteValidVec_res_47 = _RANDOM[5'h1][15];
        v0WriteValidVec_res_48 = _RANDOM[5'h1][16];
        v0WriteValidVec_res_49 = _RANDOM[5'h1][17];
        v0WriteValidVec_res_50 = _RANDOM[5'h1][18];
        v0WriteValidVec_res_51 = _RANDOM[5'h1][19];
        v0WriteValidVec_res_52 = _RANDOM[5'h1][20];
        v0WriteValidVec_res_53 = _RANDOM[5'h1][21];
        v0WriteValidVec_res_54 = _RANDOM[5'h1][22];
        v0WriteValidVec_res_55 = _RANDOM[5'h1][23];
        v0WriteValidVec_res_56 = _RANDOM[5'h1][24];
        v0WriteValidVec_res_57 = _RANDOM[5'h1][25];
        v0WriteValidVec_res_58 = _RANDOM[5'h1][26];
        v0WriteValidVec_res_59 = _RANDOM[5'h1][27];
        v0WriteValidVec_res_60 = _RANDOM[5'h1][28];
        v0WriteValidVec_res_61 = _RANDOM[5'h1][29];
        v0WriteValidVec_res_62 = _RANDOM[5'h1][30];
        v0WriteValidVec_res_63 = _RANDOM[5'h1][31];
        v0WriteValidVec_res_64 = _RANDOM[5'h2][0];
        v0WriteValidVec_res_65 = _RANDOM[5'h2][1];
        v0WriteValidVec_res_66 = _RANDOM[5'h2][2];
        v0WriteValidVec_res_67 = _RANDOM[5'h2][3];
        v0WriteValidVec_res_68 = _RANDOM[5'h2][4];
        v0WriteValidVec_res_69 = _RANDOM[5'h2][5];
        v0WriteValidVec_res_70 = _RANDOM[5'h2][6];
        v0WriteValidVec_res_71 = _RANDOM[5'h2][7];
        v0WriteValidVec_res_72 = _RANDOM[5'h2][8];
        v0WriteValidVec_res_73 = _RANDOM[5'h2][9];
        v0WriteValidVec_res_74 = _RANDOM[5'h2][10];
        v0WriteValidVec_res_75 = _RANDOM[5'h2][11];
        v0WriteValidVec_res_76 = _RANDOM[5'h2][12];
        v0WriteValidVec_res_77 = _RANDOM[5'h2][13];
        v0WriteValidVec_res_78 = _RANDOM[5'h2][14];
        v0WriteValidVec_res_79 = _RANDOM[5'h2][15];
        v0WriteValidVec_res_80 = _RANDOM[5'h2][16];
        v0WriteValidVec_res_81 = _RANDOM[5'h2][17];
        v0WriteValidVec_res_82 = _RANDOM[5'h2][18];
        v0WriteValidVec_res_83 = _RANDOM[5'h2][19];
        v0WriteValidVec_res_84 = _RANDOM[5'h2][20];
        v0WriteValidVec_res_85 = _RANDOM[5'h2][21];
        v0WriteValidVec_res_86 = _RANDOM[5'h2][22];
        v0WriteValidVec_res_87 = _RANDOM[5'h2][23];
        v0WriteValidVec_res_88 = _RANDOM[5'h2][24];
        v0WriteValidVec_res_89 = _RANDOM[5'h2][25];
        v0WriteValidVec_res_90 = _RANDOM[5'h2][26];
        v0WriteValidVec_res_91 = _RANDOM[5'h2][27];
        v0WriteValidVec_res_92 = _RANDOM[5'h2][28];
        v0WriteValidVec_res_93 = _RANDOM[5'h2][29];
        v0WriteValidVec_res_94 = _RANDOM[5'h2][30];
        v0WriteValidVec_res_95 = _RANDOM[5'h2][31];
        v0WriteValidVec_res_96 = _RANDOM[5'h3][0];
        v0WriteValidVec_res_97 = _RANDOM[5'h3][1];
        v0WriteValidVec_res_98 = _RANDOM[5'h3][2];
        v0WriteValidVec_res_99 = _RANDOM[5'h3][3];
        v0WriteValidVec_res_100 = _RANDOM[5'h3][4];
        v0WriteValidVec_res_101 = _RANDOM[5'h3][5];
        v0WriteValidVec_res_102 = _RANDOM[5'h3][6];
        v0WriteValidVec_res_103 = _RANDOM[5'h3][7];
        v0WriteValidVec_res_104 = _RANDOM[5'h3][8];
        v0WriteValidVec_res_105 = _RANDOM[5'h3][9];
        v0WriteValidVec_res_106 = _RANDOM[5'h3][10];
        v0WriteValidVec_res_107 = _RANDOM[5'h3][11];
        v0WriteValidVec_res_108 = _RANDOM[5'h3][12];
        v0WriteValidVec_res_109 = _RANDOM[5'h3][13];
        v0WriteValidVec_res_110 = _RANDOM[5'h3][14];
        v0WriteValidVec_res_111 = _RANDOM[5'h3][15];
        v0WriteValidVec_res_112 = _RANDOM[5'h3][16];
        v0WriteValidVec_res_113 = _RANDOM[5'h3][17];
        v0WriteValidVec_res_114 = _RANDOM[5'h3][18];
        v0WriteValidVec_res_115 = _RANDOM[5'h3][19];
        v0WriteValidVec_res_116 = _RANDOM[5'h3][20];
        v0WriteValidVec_res_117 = _RANDOM[5'h3][21];
        v0WriteValidVec_res_118 = _RANDOM[5'h3][22];
        v0WriteValidVec_res_119 = _RANDOM[5'h3][23];
        v0WriteValidVec_res_120 = _RANDOM[5'h3][24];
        v0WriteValidVec_res_121 = _RANDOM[5'h3][25];
        v0WriteValidVec_res_122 = _RANDOM[5'h3][26];
        v0WriteValidVec_res_123 = _RANDOM[5'h3][27];
        v0WriteValidVec_res_124 = _RANDOM[5'h3][28];
        v0WriteValidVec_res_125 = _RANDOM[5'h3][29];
        v0WriteValidVec_res_126 = _RANDOM[5'h3][30];
        v0WriteValidVec_res_127 = _RANDOM[5'h3][31];
        v0WriteValidVec_res_128 = _RANDOM[5'h4][0];
        v0WriteValidVec_res_129 = _RANDOM[5'h4][1];
        v0WriteValidVec_res_130 = _RANDOM[5'h4][2];
        v0WriteValidVec_res_131 = _RANDOM[5'h4][3];
        v0WriteValidVec_res_132 = _RANDOM[5'h4][4];
        v0WriteValidVec_res_133 = _RANDOM[5'h4][5];
        v0WriteValidVec_res_134 = _RANDOM[5'h4][6];
        v0WriteValidVec_res_135 = _RANDOM[5'h4][7];
        v0WriteValidVec_res_136 = _RANDOM[5'h4][8];
        v0WriteValidVec_res_137 = _RANDOM[5'h4][9];
        v0WriteValidVec_res_138 = _RANDOM[5'h4][10];
        v0WriteValidVec_res_139 = _RANDOM[5'h4][11];
        v0WriteValidVec_res_140 = _RANDOM[5'h4][12];
        v0WriteValidVec_res_141 = _RANDOM[5'h4][13];
        v0WriteValidVec_res_142 = _RANDOM[5'h4][14];
        v0WriteValidVec_res_143 = _RANDOM[5'h4][15];
        v0WriteValidVec_res_144 = _RANDOM[5'h4][16];
        v0WriteValidVec_res_145 = _RANDOM[5'h4][17];
        v0WriteValidVec_res_146 = _RANDOM[5'h4][18];
        v0WriteValidVec_res_147 = _RANDOM[5'h4][19];
        v0WriteValidVec_res_148 = _RANDOM[5'h4][20];
        v0WriteValidVec_res_149 = _RANDOM[5'h4][21];
        v0WriteValidVec_res_150 = _RANDOM[5'h4][22];
        v0WriteValidVec_res_151 = _RANDOM[5'h4][23];
        v0WriteValidVec_res_152 = _RANDOM[5'h4][24];
        v0WriteValidVec_res_153 = _RANDOM[5'h4][25];
        v0WriteValidVec_res_154 = _RANDOM[5'h4][26];
        v0WriteValidVec_res_155 = _RANDOM[5'h4][27];
        v0WriteValidVec_res_156 = _RANDOM[5'h4][28];
        v0WriteValidVec_res_157 = _RANDOM[5'h4][29];
        v0WriteValidVec_res_158 = _RANDOM[5'h4][30];
        v0WriteValidVec_res_159 = _RANDOM[5'h4][31];
        v0WriteValidVec_res_160 = _RANDOM[5'h5][0];
        v0WriteValidVec_res_161 = _RANDOM[5'h5][1];
        v0WriteValidVec_res_162 = _RANDOM[5'h5][2];
        v0WriteValidVec_res_163 = _RANDOM[5'h5][3];
        v0WriteValidVec_res_164 = _RANDOM[5'h5][4];
        v0WriteValidVec_res_165 = _RANDOM[5'h5][5];
        v0WriteValidVec_res_166 = _RANDOM[5'h5][6];
        v0WriteValidVec_res_167 = _RANDOM[5'h5][7];
        v0WriteValidVec_res_168 = _RANDOM[5'h5][8];
        v0WriteValidVec_res_169 = _RANDOM[5'h5][9];
        v0WriteValidVec_res_170 = _RANDOM[5'h5][10];
        v0WriteValidVec_res_171 = _RANDOM[5'h5][11];
        v0WriteValidVec_res_172 = _RANDOM[5'h5][12];
        v0WriteValidVec_res_173 = _RANDOM[5'h5][13];
        v0WriteValidVec_res_174 = _RANDOM[5'h5][14];
        v0WriteValidVec_res_175 = _RANDOM[5'h5][15];
        v0WriteValidVec_res_176 = _RANDOM[5'h5][16];
        v0WriteValidVec_res_177 = _RANDOM[5'h5][17];
        v0WriteValidVec_res_178 = _RANDOM[5'h5][18];
        v0WriteValidVec_res_179 = _RANDOM[5'h5][19];
        v0WriteValidVec_res_180 = _RANDOM[5'h5][20];
        v0WriteValidVec_res_181 = _RANDOM[5'h5][21];
        v0WriteValidVec_res_182 = _RANDOM[5'h5][22];
        v0WriteValidVec_res_183 = _RANDOM[5'h5][23];
        v0WriteValidVec_res_184 = _RANDOM[5'h5][24];
        v0WriteValidVec_res_185 = _RANDOM[5'h5][25];
        v0WriteValidVec_res_186 = _RANDOM[5'h5][26];
        v0WriteValidVec_res_187 = _RANDOM[5'h5][27];
        v0WriteValidVec_res_188 = _RANDOM[5'h5][28];
        v0WriteValidVec_res_189 = _RANDOM[5'h5][29];
        v0WriteValidVec_res_190 = _RANDOM[5'h5][30];
        v0WriteValidVec_res_191 = _RANDOM[5'h5][31];
        v0WriteValidVec_res_192 = _RANDOM[5'h6][0];
        v0WriteValidVec_res_193 = _RANDOM[5'h6][1];
        v0WriteValidVec_res_194 = _RANDOM[5'h6][2];
        v0WriteValidVec_res_195 = _RANDOM[5'h6][3];
        v0WriteValidVec_res_196 = _RANDOM[5'h6][4];
        v0WriteValidVec_res_197 = _RANDOM[5'h6][5];
        v0WriteValidVec_res_198 = _RANDOM[5'h6][6];
        v0WriteValidVec_res_199 = _RANDOM[5'h6][7];
        v0WriteValidVec_res_200 = _RANDOM[5'h6][8];
        v0WriteValidVec_res_201 = _RANDOM[5'h6][9];
        v0WriteValidVec_res_202 = _RANDOM[5'h6][10];
        v0WriteValidVec_res_203 = _RANDOM[5'h6][11];
        v0WriteValidVec_res_204 = _RANDOM[5'h6][12];
        v0WriteValidVec_res_205 = _RANDOM[5'h6][13];
        v0WriteValidVec_res_206 = _RANDOM[5'h6][14];
        v0WriteValidVec_res_207 = _RANDOM[5'h6][15];
        v0WriteValidVec_res_208 = _RANDOM[5'h6][16];
        v0WriteValidVec_res_209 = _RANDOM[5'h6][17];
        v0WriteValidVec_res_210 = _RANDOM[5'h6][18];
        v0WriteValidVec_res_211 = _RANDOM[5'h6][19];
        v0WriteValidVec_res_212 = _RANDOM[5'h6][20];
        v0WriteValidVec_res_213 = _RANDOM[5'h6][21];
        v0WriteValidVec_res_214 = _RANDOM[5'h6][22];
        v0WriteValidVec_res_215 = _RANDOM[5'h6][23];
        v0WriteValidVec_res_216 = _RANDOM[5'h6][24];
        v0WriteValidVec_res_217 = _RANDOM[5'h6][25];
        v0WriteValidVec_res_218 = _RANDOM[5'h6][26];
        v0WriteValidVec_res_219 = _RANDOM[5'h6][27];
        v0WriteValidVec_res_220 = _RANDOM[5'h6][28];
        v0WriteValidVec_res_221 = _RANDOM[5'h6][29];
        v0WriteValidVec_res_222 = _RANDOM[5'h6][30];
        v0WriteValidVec_res_223 = _RANDOM[5'h6][31];
        v0WriteValidVec_res_224 = _RANDOM[5'h7][0];
        v0WriteValidVec_res_225 = _RANDOM[5'h7][1];
        v0WriteValidVec_res_226 = _RANDOM[5'h7][2];
        v0WriteValidVec_res_227 = _RANDOM[5'h7][3];
        v0WriteValidVec_res_228 = _RANDOM[5'h7][4];
        v0WriteValidVec_res_229 = _RANDOM[5'h7][5];
        v0WriteValidVec_res_230 = _RANDOM[5'h7][6];
        v0WriteValidVec_res_231 = _RANDOM[5'h7][7];
        v0WriteValidVec_res_232 = _RANDOM[5'h7][8];
        v0WriteValidVec_res_233 = _RANDOM[5'h7][9];
        v0WriteValidVec_res_234 = _RANDOM[5'h7][10];
        v0WriteValidVec_res_235 = _RANDOM[5'h7][11];
        v0WriteValidVec_res_236 = _RANDOM[5'h7][12];
        v0WriteValidVec_res_237 = _RANDOM[5'h7][13];
        v0WriteValidVec_res_238 = _RANDOM[5'h7][14];
        v0WriteValidVec_res_239 = _RANDOM[5'h7][15];
        v0WriteValidVec_res_240 = _RANDOM[5'h7][16];
        v0WriteValidVec_res_241 = _RANDOM[5'h7][17];
        v0WriteValidVec_res_242 = _RANDOM[5'h7][18];
        v0WriteValidVec_res_243 = _RANDOM[5'h7][19];
        v0WriteValidVec_res_244 = _RANDOM[5'h7][20];
        v0WriteValidVec_res_245 = _RANDOM[5'h7][21];
        v0WriteValidVec_res_246 = _RANDOM[5'h7][22];
        v0WriteValidVec_res_247 = _RANDOM[5'h7][23];
        v0WriteValidVec_res_248 = _RANDOM[5'h7][24];
        v0WriteValidVec_res_249 = _RANDOM[5'h7][25];
        v0WriteValidVec_res_250 = _RANDOM[5'h7][26];
        v0WriteValidVec_res_251 = _RANDOM[5'h7][27];
        v0WriteValidVec_res_252 = _RANDOM[5'h7][28];
        v0WriteValidVec_res_253 = _RANDOM[5'h7][29];
        v0WriteValidVec_res_254 = _RANDOM[5'h7][30];
        v0WriteValidVec_res_255 = _RANDOM[5'h7][31];
        useV0AsMaskToken_res = _RANDOM[5'h8][0];
        useV0AsMaskToken_res_1 = _RANDOM[5'h8][1];
        useV0AsMaskToken_res_2 = _RANDOM[5'h8][2];
        useV0AsMaskToken_res_3 = _RANDOM[5'h8][3];
        useV0AsMaskToken_res_4 = _RANDOM[5'h8][4];
        useV0AsMaskToken_res_5 = _RANDOM[5'h8][5];
        useV0AsMaskToken_res_6 = _RANDOM[5'h8][6];
        useV0AsMaskToken_res_7 = _RANDOM[5'h8][7];
        useV0AsMaskToken_res_8 = _RANDOM[5'h8][8];
        useV0AsMaskToken_res_9 = _RANDOM[5'h8][9];
        useV0AsMaskToken_res_10 = _RANDOM[5'h8][10];
        useV0AsMaskToken_res_11 = _RANDOM[5'h8][11];
        useV0AsMaskToken_res_12 = _RANDOM[5'h8][12];
        useV0AsMaskToken_res_13 = _RANDOM[5'h8][13];
        useV0AsMaskToken_res_14 = _RANDOM[5'h8][14];
        useV0AsMaskToken_res_15 = _RANDOM[5'h8][15];
        useV0AsMaskToken_res_16 = _RANDOM[5'h8][16];
        useV0AsMaskToken_res_17 = _RANDOM[5'h8][17];
        useV0AsMaskToken_res_18 = _RANDOM[5'h8][18];
        useV0AsMaskToken_res_19 = _RANDOM[5'h8][19];
        useV0AsMaskToken_res_20 = _RANDOM[5'h8][20];
        useV0AsMaskToken_res_21 = _RANDOM[5'h8][21];
        useV0AsMaskToken_res_22 = _RANDOM[5'h8][22];
        useV0AsMaskToken_res_23 = _RANDOM[5'h8][23];
        useV0AsMaskToken_res_24 = _RANDOM[5'h8][24];
        useV0AsMaskToken_res_25 = _RANDOM[5'h8][25];
        useV0AsMaskToken_res_26 = _RANDOM[5'h8][26];
        useV0AsMaskToken_res_27 = _RANDOM[5'h8][27];
        useV0AsMaskToken_res_28 = _RANDOM[5'h8][28];
        useV0AsMaskToken_res_29 = _RANDOM[5'h8][29];
        useV0AsMaskToken_res_30 = _RANDOM[5'h8][30];
        useV0AsMaskToken_res_31 = _RANDOM[5'h8][31];
        useV0AsMaskToken_res_32 = _RANDOM[5'h9][0];
        useV0AsMaskToken_res_33 = _RANDOM[5'h9][1];
        useV0AsMaskToken_res_34 = _RANDOM[5'h9][2];
        useV0AsMaskToken_res_35 = _RANDOM[5'h9][3];
        useV0AsMaskToken_res_36 = _RANDOM[5'h9][4];
        useV0AsMaskToken_res_37 = _RANDOM[5'h9][5];
        useV0AsMaskToken_res_38 = _RANDOM[5'h9][6];
        useV0AsMaskToken_res_39 = _RANDOM[5'h9][7];
        useV0AsMaskToken_res_40 = _RANDOM[5'h9][8];
        useV0AsMaskToken_res_41 = _RANDOM[5'h9][9];
        useV0AsMaskToken_res_42 = _RANDOM[5'h9][10];
        useV0AsMaskToken_res_43 = _RANDOM[5'h9][11];
        useV0AsMaskToken_res_44 = _RANDOM[5'h9][12];
        useV0AsMaskToken_res_45 = _RANDOM[5'h9][13];
        useV0AsMaskToken_res_46 = _RANDOM[5'h9][14];
        useV0AsMaskToken_res_47 = _RANDOM[5'h9][15];
        useV0AsMaskToken_res_48 = _RANDOM[5'h9][16];
        useV0AsMaskToken_res_49 = _RANDOM[5'h9][17];
        useV0AsMaskToken_res_50 = _RANDOM[5'h9][18];
        useV0AsMaskToken_res_51 = _RANDOM[5'h9][19];
        useV0AsMaskToken_res_52 = _RANDOM[5'h9][20];
        useV0AsMaskToken_res_53 = _RANDOM[5'h9][21];
        useV0AsMaskToken_res_54 = _RANDOM[5'h9][22];
        useV0AsMaskToken_res_55 = _RANDOM[5'h9][23];
        useV0AsMaskToken_res_56 = _RANDOM[5'h9][24];
        useV0AsMaskToken_res_57 = _RANDOM[5'h9][25];
        useV0AsMaskToken_res_58 = _RANDOM[5'h9][26];
        useV0AsMaskToken_res_59 = _RANDOM[5'h9][27];
        useV0AsMaskToken_res_60 = _RANDOM[5'h9][28];
        useV0AsMaskToken_res_61 = _RANDOM[5'h9][29];
        useV0AsMaskToken_res_62 = _RANDOM[5'h9][30];
        useV0AsMaskToken_res_63 = _RANDOM[5'h9][31];
        useV0AsMaskToken_res_64 = _RANDOM[5'hA][0];
        useV0AsMaskToken_res_65 = _RANDOM[5'hA][1];
        useV0AsMaskToken_res_66 = _RANDOM[5'hA][2];
        useV0AsMaskToken_res_67 = _RANDOM[5'hA][3];
        useV0AsMaskToken_res_68 = _RANDOM[5'hA][4];
        useV0AsMaskToken_res_69 = _RANDOM[5'hA][5];
        useV0AsMaskToken_res_70 = _RANDOM[5'hA][6];
        useV0AsMaskToken_res_71 = _RANDOM[5'hA][7];
        useV0AsMaskToken_res_72 = _RANDOM[5'hA][8];
        useV0AsMaskToken_res_73 = _RANDOM[5'hA][9];
        useV0AsMaskToken_res_74 = _RANDOM[5'hA][10];
        useV0AsMaskToken_res_75 = _RANDOM[5'hA][11];
        useV0AsMaskToken_res_76 = _RANDOM[5'hA][12];
        useV0AsMaskToken_res_77 = _RANDOM[5'hA][13];
        useV0AsMaskToken_res_78 = _RANDOM[5'hA][14];
        useV0AsMaskToken_res_79 = _RANDOM[5'hA][15];
        useV0AsMaskToken_res_80 = _RANDOM[5'hA][16];
        useV0AsMaskToken_res_81 = _RANDOM[5'hA][17];
        useV0AsMaskToken_res_82 = _RANDOM[5'hA][18];
        useV0AsMaskToken_res_83 = _RANDOM[5'hA][19];
        useV0AsMaskToken_res_84 = _RANDOM[5'hA][20];
        useV0AsMaskToken_res_85 = _RANDOM[5'hA][21];
        useV0AsMaskToken_res_86 = _RANDOM[5'hA][22];
        useV0AsMaskToken_res_87 = _RANDOM[5'hA][23];
        useV0AsMaskToken_res_88 = _RANDOM[5'hA][24];
        useV0AsMaskToken_res_89 = _RANDOM[5'hA][25];
        useV0AsMaskToken_res_90 = _RANDOM[5'hA][26];
        useV0AsMaskToken_res_91 = _RANDOM[5'hA][27];
        useV0AsMaskToken_res_92 = _RANDOM[5'hA][28];
        useV0AsMaskToken_res_93 = _RANDOM[5'hA][29];
        useV0AsMaskToken_res_94 = _RANDOM[5'hA][30];
        useV0AsMaskToken_res_95 = _RANDOM[5'hA][31];
        useV0AsMaskToken_res_96 = _RANDOM[5'hB][0];
        useV0AsMaskToken_res_97 = _RANDOM[5'hB][1];
        useV0AsMaskToken_res_98 = _RANDOM[5'hB][2];
        useV0AsMaskToken_res_99 = _RANDOM[5'hB][3];
        useV0AsMaskToken_res_100 = _RANDOM[5'hB][4];
        useV0AsMaskToken_res_101 = _RANDOM[5'hB][5];
        useV0AsMaskToken_res_102 = _RANDOM[5'hB][6];
        useV0AsMaskToken_res_103 = _RANDOM[5'hB][7];
        useV0AsMaskToken_res_104 = _RANDOM[5'hB][8];
        useV0AsMaskToken_res_105 = _RANDOM[5'hB][9];
        useV0AsMaskToken_res_106 = _RANDOM[5'hB][10];
        useV0AsMaskToken_res_107 = _RANDOM[5'hB][11];
        useV0AsMaskToken_res_108 = _RANDOM[5'hB][12];
        useV0AsMaskToken_res_109 = _RANDOM[5'hB][13];
        useV0AsMaskToken_res_110 = _RANDOM[5'hB][14];
        useV0AsMaskToken_res_111 = _RANDOM[5'hB][15];
        useV0AsMaskToken_res_112 = _RANDOM[5'hB][16];
        useV0AsMaskToken_res_113 = _RANDOM[5'hB][17];
        useV0AsMaskToken_res_114 = _RANDOM[5'hB][18];
        useV0AsMaskToken_res_115 = _RANDOM[5'hB][19];
        useV0AsMaskToken_res_116 = _RANDOM[5'hB][20];
        useV0AsMaskToken_res_117 = _RANDOM[5'hB][21];
        useV0AsMaskToken_res_118 = _RANDOM[5'hB][22];
        useV0AsMaskToken_res_119 = _RANDOM[5'hB][23];
        useV0AsMaskToken_res_120 = _RANDOM[5'hB][24];
        useV0AsMaskToken_res_121 = _RANDOM[5'hB][25];
        useV0AsMaskToken_res_122 = _RANDOM[5'hB][26];
        useV0AsMaskToken_res_123 = _RANDOM[5'hB][27];
        useV0AsMaskToken_res_124 = _RANDOM[5'hB][28];
        useV0AsMaskToken_res_125 = _RANDOM[5'hB][29];
        useV0AsMaskToken_res_126 = _RANDOM[5'hB][30];
        useV0AsMaskToken_res_127 = _RANDOM[5'hB][31];
        useV0AsMaskToken_res_128 = _RANDOM[5'hC][0];
        useV0AsMaskToken_res_129 = _RANDOM[5'hC][1];
        useV0AsMaskToken_res_130 = _RANDOM[5'hC][2];
        useV0AsMaskToken_res_131 = _RANDOM[5'hC][3];
        useV0AsMaskToken_res_132 = _RANDOM[5'hC][4];
        useV0AsMaskToken_res_133 = _RANDOM[5'hC][5];
        useV0AsMaskToken_res_134 = _RANDOM[5'hC][6];
        useV0AsMaskToken_res_135 = _RANDOM[5'hC][7];
        useV0AsMaskToken_res_136 = _RANDOM[5'hC][8];
        useV0AsMaskToken_res_137 = _RANDOM[5'hC][9];
        useV0AsMaskToken_res_138 = _RANDOM[5'hC][10];
        useV0AsMaskToken_res_139 = _RANDOM[5'hC][11];
        useV0AsMaskToken_res_140 = _RANDOM[5'hC][12];
        useV0AsMaskToken_res_141 = _RANDOM[5'hC][13];
        useV0AsMaskToken_res_142 = _RANDOM[5'hC][14];
        useV0AsMaskToken_res_143 = _RANDOM[5'hC][15];
        useV0AsMaskToken_res_144 = _RANDOM[5'hC][16];
        useV0AsMaskToken_res_145 = _RANDOM[5'hC][17];
        useV0AsMaskToken_res_146 = _RANDOM[5'hC][18];
        useV0AsMaskToken_res_147 = _RANDOM[5'hC][19];
        useV0AsMaskToken_res_148 = _RANDOM[5'hC][20];
        useV0AsMaskToken_res_149 = _RANDOM[5'hC][21];
        useV0AsMaskToken_res_150 = _RANDOM[5'hC][22];
        useV0AsMaskToken_res_151 = _RANDOM[5'hC][23];
        useV0AsMaskToken_res_152 = _RANDOM[5'hC][24];
        useV0AsMaskToken_res_153 = _RANDOM[5'hC][25];
        useV0AsMaskToken_res_154 = _RANDOM[5'hC][26];
        useV0AsMaskToken_res_155 = _RANDOM[5'hC][27];
        useV0AsMaskToken_res_156 = _RANDOM[5'hC][28];
        useV0AsMaskToken_res_157 = _RANDOM[5'hC][29];
        useV0AsMaskToken_res_158 = _RANDOM[5'hC][30];
        useV0AsMaskToken_res_159 = _RANDOM[5'hC][31];
        useV0AsMaskToken_res_160 = _RANDOM[5'hD][0];
        useV0AsMaskToken_res_161 = _RANDOM[5'hD][1];
        useV0AsMaskToken_res_162 = _RANDOM[5'hD][2];
        useV0AsMaskToken_res_163 = _RANDOM[5'hD][3];
        useV0AsMaskToken_res_164 = _RANDOM[5'hD][4];
        useV0AsMaskToken_res_165 = _RANDOM[5'hD][5];
        useV0AsMaskToken_res_166 = _RANDOM[5'hD][6];
        useV0AsMaskToken_res_167 = _RANDOM[5'hD][7];
        useV0AsMaskToken_res_168 = _RANDOM[5'hD][8];
        useV0AsMaskToken_res_169 = _RANDOM[5'hD][9];
        useV0AsMaskToken_res_170 = _RANDOM[5'hD][10];
        useV0AsMaskToken_res_171 = _RANDOM[5'hD][11];
        useV0AsMaskToken_res_172 = _RANDOM[5'hD][12];
        useV0AsMaskToken_res_173 = _RANDOM[5'hD][13];
        useV0AsMaskToken_res_174 = _RANDOM[5'hD][14];
        useV0AsMaskToken_res_175 = _RANDOM[5'hD][15];
        useV0AsMaskToken_res_176 = _RANDOM[5'hD][16];
        useV0AsMaskToken_res_177 = _RANDOM[5'hD][17];
        useV0AsMaskToken_res_178 = _RANDOM[5'hD][18];
        useV0AsMaskToken_res_179 = _RANDOM[5'hD][19];
        useV0AsMaskToken_res_180 = _RANDOM[5'hD][20];
        useV0AsMaskToken_res_181 = _RANDOM[5'hD][21];
        useV0AsMaskToken_res_182 = _RANDOM[5'hD][22];
        useV0AsMaskToken_res_183 = _RANDOM[5'hD][23];
        useV0AsMaskToken_res_184 = _RANDOM[5'hD][24];
        useV0AsMaskToken_res_185 = _RANDOM[5'hD][25];
        useV0AsMaskToken_res_186 = _RANDOM[5'hD][26];
        useV0AsMaskToken_res_187 = _RANDOM[5'hD][27];
        useV0AsMaskToken_res_188 = _RANDOM[5'hD][28];
        useV0AsMaskToken_res_189 = _RANDOM[5'hD][29];
        useV0AsMaskToken_res_190 = _RANDOM[5'hD][30];
        useV0AsMaskToken_res_191 = _RANDOM[5'hD][31];
        useV0AsMaskToken_res_192 = _RANDOM[5'hE][0];
        useV0AsMaskToken_res_193 = _RANDOM[5'hE][1];
        useV0AsMaskToken_res_194 = _RANDOM[5'hE][2];
        useV0AsMaskToken_res_195 = _RANDOM[5'hE][3];
        useV0AsMaskToken_res_196 = _RANDOM[5'hE][4];
        useV0AsMaskToken_res_197 = _RANDOM[5'hE][5];
        useV0AsMaskToken_res_198 = _RANDOM[5'hE][6];
        useV0AsMaskToken_res_199 = _RANDOM[5'hE][7];
        useV0AsMaskToken_res_200 = _RANDOM[5'hE][8];
        useV0AsMaskToken_res_201 = _RANDOM[5'hE][9];
        useV0AsMaskToken_res_202 = _RANDOM[5'hE][10];
        useV0AsMaskToken_res_203 = _RANDOM[5'hE][11];
        useV0AsMaskToken_res_204 = _RANDOM[5'hE][12];
        useV0AsMaskToken_res_205 = _RANDOM[5'hE][13];
        useV0AsMaskToken_res_206 = _RANDOM[5'hE][14];
        useV0AsMaskToken_res_207 = _RANDOM[5'hE][15];
        useV0AsMaskToken_res_208 = _RANDOM[5'hE][16];
        useV0AsMaskToken_res_209 = _RANDOM[5'hE][17];
        useV0AsMaskToken_res_210 = _RANDOM[5'hE][18];
        useV0AsMaskToken_res_211 = _RANDOM[5'hE][19];
        useV0AsMaskToken_res_212 = _RANDOM[5'hE][20];
        useV0AsMaskToken_res_213 = _RANDOM[5'hE][21];
        useV0AsMaskToken_res_214 = _RANDOM[5'hE][22];
        useV0AsMaskToken_res_215 = _RANDOM[5'hE][23];
        useV0AsMaskToken_res_216 = _RANDOM[5'hE][24];
        useV0AsMaskToken_res_217 = _RANDOM[5'hE][25];
        useV0AsMaskToken_res_218 = _RANDOM[5'hE][26];
        useV0AsMaskToken_res_219 = _RANDOM[5'hE][27];
        useV0AsMaskToken_res_220 = _RANDOM[5'hE][28];
        useV0AsMaskToken_res_221 = _RANDOM[5'hE][29];
        useV0AsMaskToken_res_222 = _RANDOM[5'hE][30];
        useV0AsMaskToken_res_223 = _RANDOM[5'hE][31];
        useV0AsMaskToken_res_224 = _RANDOM[5'hF][0];
        useV0AsMaskToken_res_225 = _RANDOM[5'hF][1];
        useV0AsMaskToken_res_226 = _RANDOM[5'hF][2];
        useV0AsMaskToken_res_227 = _RANDOM[5'hF][3];
        useV0AsMaskToken_res_228 = _RANDOM[5'hF][4];
        useV0AsMaskToken_res_229 = _RANDOM[5'hF][5];
        useV0AsMaskToken_res_230 = _RANDOM[5'hF][6];
        useV0AsMaskToken_res_231 = _RANDOM[5'hF][7];
        useV0AsMaskToken_res_232 = _RANDOM[5'hF][8];
        useV0AsMaskToken_res_233 = _RANDOM[5'hF][9];
        useV0AsMaskToken_res_234 = _RANDOM[5'hF][10];
        useV0AsMaskToken_res_235 = _RANDOM[5'hF][11];
        useV0AsMaskToken_res_236 = _RANDOM[5'hF][12];
        useV0AsMaskToken_res_237 = _RANDOM[5'hF][13];
        useV0AsMaskToken_res_238 = _RANDOM[5'hF][14];
        useV0AsMaskToken_res_239 = _RANDOM[5'hF][15];
        useV0AsMaskToken_res_240 = _RANDOM[5'hF][16];
        useV0AsMaskToken_res_241 = _RANDOM[5'hF][17];
        useV0AsMaskToken_res_242 = _RANDOM[5'hF][18];
        useV0AsMaskToken_res_243 = _RANDOM[5'hF][19];
        useV0AsMaskToken_res_244 = _RANDOM[5'hF][20];
        useV0AsMaskToken_res_245 = _RANDOM[5'hF][21];
        useV0AsMaskToken_res_246 = _RANDOM[5'hF][22];
        useV0AsMaskToken_res_247 = _RANDOM[5'hF][23];
        useV0AsMaskToken_res_248 = _RANDOM[5'hF][24];
        useV0AsMaskToken_res_249 = _RANDOM[5'hF][25];
        useV0AsMaskToken_res_250 = _RANDOM[5'hF][26];
        useV0AsMaskToken_res_251 = _RANDOM[5'hF][27];
        useV0AsMaskToken_res_252 = _RANDOM[5'hF][28];
        useV0AsMaskToken_res_253 = _RANDOM[5'hF][29];
        useV0AsMaskToken_res_254 = _RANDOM[5'hF][30];
        useV0AsMaskToken_res_255 = _RANDOM[5'hF][31];
        maskUnitWriteV0 = _RANDOM[5'h10][0];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  assign issueAllow = ~v0Conflict;
  assign v0WriteValid = _v0WriteValid_output;
endmodule

