
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module LSU(
  input          clock,
                 reset,
  output         request_ready,
  input          request_valid,
  input  [2:0]   request_bits_instructionInformation_nf,
  input          request_bits_instructionInformation_mew,
  input  [1:0]   request_bits_instructionInformation_mop,
  input  [4:0]   request_bits_instructionInformation_lumop,
  input  [1:0]   request_bits_instructionInformation_eew,
  input  [4:0]   request_bits_instructionInformation_vs3,
  input          request_bits_instructionInformation_isStore,
                 request_bits_instructionInformation_maskedLoadStore,
  input  [31:0]  request_bits_rs1Data,
                 request_bits_rs2Data,
  input  [2:0]   request_bits_instructionIndex,
  input          v0UpdateVec_0_valid,
  input  [31:0]  v0UpdateVec_0_bits_data,
  input  [1:0]   v0UpdateVec_0_bits_offset,
  input  [3:0]   v0UpdateVec_0_bits_mask,
  input          v0UpdateVec_1_valid,
  input  [31:0]  v0UpdateVec_1_bits_data,
  input  [1:0]   v0UpdateVec_1_bits_offset,
  input  [3:0]   v0UpdateVec_1_bits_mask,
  input          v0UpdateVec_2_valid,
  input  [31:0]  v0UpdateVec_2_bits_data,
  input  [1:0]   v0UpdateVec_2_bits_offset,
  input  [3:0]   v0UpdateVec_2_bits_mask,
  input          v0UpdateVec_3_valid,
  input  [31:0]  v0UpdateVec_3_bits_data,
  input  [1:0]   v0UpdateVec_3_bits_offset,
  input  [3:0]   v0UpdateVec_3_bits_mask,
  input          v0UpdateVec_4_valid,
  input  [31:0]  v0UpdateVec_4_bits_data,
  input  [1:0]   v0UpdateVec_4_bits_offset,
  input  [3:0]   v0UpdateVec_4_bits_mask,
  input          v0UpdateVec_5_valid,
  input  [31:0]  v0UpdateVec_5_bits_data,
  input  [1:0]   v0UpdateVec_5_bits_offset,
  input  [3:0]   v0UpdateVec_5_bits_mask,
  input          v0UpdateVec_6_valid,
  input  [31:0]  v0UpdateVec_6_bits_data,
  input  [1:0]   v0UpdateVec_6_bits_offset,
  input  [3:0]   v0UpdateVec_6_bits_mask,
  input          v0UpdateVec_7_valid,
  input  [31:0]  v0UpdateVec_7_bits_data,
  input  [1:0]   v0UpdateVec_7_bits_offset,
  input  [3:0]   v0UpdateVec_7_bits_mask,
  input          v0UpdateVec_8_valid,
  input  [31:0]  v0UpdateVec_8_bits_data,
  input  [1:0]   v0UpdateVec_8_bits_offset,
  input  [3:0]   v0UpdateVec_8_bits_mask,
  input          v0UpdateVec_9_valid,
  input  [31:0]  v0UpdateVec_9_bits_data,
  input  [1:0]   v0UpdateVec_9_bits_offset,
  input  [3:0]   v0UpdateVec_9_bits_mask,
  input          v0UpdateVec_10_valid,
  input  [31:0]  v0UpdateVec_10_bits_data,
  input  [1:0]   v0UpdateVec_10_bits_offset,
  input  [3:0]   v0UpdateVec_10_bits_mask,
  input          v0UpdateVec_11_valid,
  input  [31:0]  v0UpdateVec_11_bits_data,
  input  [1:0]   v0UpdateVec_11_bits_offset,
  input  [3:0]   v0UpdateVec_11_bits_mask,
  input          v0UpdateVec_12_valid,
  input  [31:0]  v0UpdateVec_12_bits_data,
  input  [1:0]   v0UpdateVec_12_bits_offset,
  input  [3:0]   v0UpdateVec_12_bits_mask,
  input          v0UpdateVec_13_valid,
  input  [31:0]  v0UpdateVec_13_bits_data,
  input  [1:0]   v0UpdateVec_13_bits_offset,
  input  [3:0]   v0UpdateVec_13_bits_mask,
  input          v0UpdateVec_14_valid,
  input  [31:0]  v0UpdateVec_14_bits_data,
  input  [1:0]   v0UpdateVec_14_bits_offset,
  input  [3:0]   v0UpdateVec_14_bits_mask,
  input          v0UpdateVec_15_valid,
  input  [31:0]  v0UpdateVec_15_bits_data,
  input  [1:0]   v0UpdateVec_15_bits_offset,
  input  [3:0]   v0UpdateVec_15_bits_mask,
  input          axi4Port_aw_ready,
  output         axi4Port_aw_valid,
  output [1:0]   axi4Port_aw_bits_id,
  output [31:0]  axi4Port_aw_bits_addr,
  input          axi4Port_w_ready,
  output         axi4Port_w_valid,
  output [511:0] axi4Port_w_bits_data,
  output [63:0]  axi4Port_w_bits_strb,
  input          axi4Port_b_valid,
  input  [1:0]   axi4Port_b_bits_id,
                 axi4Port_b_bits_resp,
  input          axi4Port_ar_ready,
  output         axi4Port_ar_valid,
  output [31:0]  axi4Port_ar_bits_addr,
  output         axi4Port_r_ready,
  input          axi4Port_r_valid,
  input  [1:0]   axi4Port_r_bits_id,
  input  [511:0] axi4Port_r_bits_data,
  input  [1:0]   axi4Port_r_bits_resp,
  input          axi4Port_r_bits_last,
                 simpleAccessPorts_aw_ready,
  output         simpleAccessPorts_aw_valid,
  output [1:0]   simpleAccessPorts_aw_bits_id,
  output [31:0]  simpleAccessPorts_aw_bits_addr,
  output [2:0]   simpleAccessPorts_aw_bits_size,
  input          simpleAccessPorts_w_ready,
  output         simpleAccessPorts_w_valid,
  output [31:0]  simpleAccessPorts_w_bits_data,
  output [3:0]   simpleAccessPorts_w_bits_strb,
  input          simpleAccessPorts_b_valid,
  input  [1:0]   simpleAccessPorts_b_bits_id,
                 simpleAccessPorts_b_bits_resp,
  input          simpleAccessPorts_ar_ready,
  output         simpleAccessPorts_ar_valid,
  output [31:0]  simpleAccessPorts_ar_bits_addr,
  output         simpleAccessPorts_r_ready,
  input          simpleAccessPorts_r_valid,
  input  [1:0]   simpleAccessPorts_r_bits_id,
  input  [31:0]  simpleAccessPorts_r_bits_data,
  input  [1:0]   simpleAccessPorts_r_bits_resp,
  input          simpleAccessPorts_r_bits_last,
                 vrfReadDataPorts_0_ready,
  output         vrfReadDataPorts_0_valid,
  output [4:0]   vrfReadDataPorts_0_bits_vs,
  output [1:0]   vrfReadDataPorts_0_bits_offset,
  output [2:0]   vrfReadDataPorts_0_bits_instructionIndex,
  input          vrfReadDataPorts_1_ready,
  output         vrfReadDataPorts_1_valid,
  output [4:0]   vrfReadDataPorts_1_bits_vs,
  output [1:0]   vrfReadDataPorts_1_bits_offset,
  output [2:0]   vrfReadDataPorts_1_bits_instructionIndex,
  input          vrfReadDataPorts_2_ready,
  output         vrfReadDataPorts_2_valid,
  output [4:0]   vrfReadDataPorts_2_bits_vs,
  output [1:0]   vrfReadDataPorts_2_bits_offset,
  output [2:0]   vrfReadDataPorts_2_bits_instructionIndex,
  input          vrfReadDataPorts_3_ready,
  output         vrfReadDataPorts_3_valid,
  output [4:0]   vrfReadDataPorts_3_bits_vs,
  output [1:0]   vrfReadDataPorts_3_bits_offset,
  output [2:0]   vrfReadDataPorts_3_bits_instructionIndex,
  input          vrfReadDataPorts_4_ready,
  output         vrfReadDataPorts_4_valid,
  output [4:0]   vrfReadDataPorts_4_bits_vs,
  output [1:0]   vrfReadDataPorts_4_bits_offset,
  output [2:0]   vrfReadDataPorts_4_bits_instructionIndex,
  input          vrfReadDataPorts_5_ready,
  output         vrfReadDataPorts_5_valid,
  output [4:0]   vrfReadDataPorts_5_bits_vs,
  output [1:0]   vrfReadDataPorts_5_bits_offset,
  output [2:0]   vrfReadDataPorts_5_bits_instructionIndex,
  input          vrfReadDataPorts_6_ready,
  output         vrfReadDataPorts_6_valid,
  output [4:0]   vrfReadDataPorts_6_bits_vs,
  output [1:0]   vrfReadDataPorts_6_bits_offset,
  output [2:0]   vrfReadDataPorts_6_bits_instructionIndex,
  input          vrfReadDataPorts_7_ready,
  output         vrfReadDataPorts_7_valid,
  output [4:0]   vrfReadDataPorts_7_bits_vs,
  output [1:0]   vrfReadDataPorts_7_bits_offset,
  output [2:0]   vrfReadDataPorts_7_bits_instructionIndex,
  input          vrfReadDataPorts_8_ready,
  output         vrfReadDataPorts_8_valid,
  output [4:0]   vrfReadDataPorts_8_bits_vs,
  output [1:0]   vrfReadDataPorts_8_bits_offset,
  output [2:0]   vrfReadDataPorts_8_bits_instructionIndex,
  input          vrfReadDataPorts_9_ready,
  output         vrfReadDataPorts_9_valid,
  output [4:0]   vrfReadDataPorts_9_bits_vs,
  output [1:0]   vrfReadDataPorts_9_bits_offset,
  output [2:0]   vrfReadDataPorts_9_bits_instructionIndex,
  input          vrfReadDataPorts_10_ready,
  output         vrfReadDataPorts_10_valid,
  output [4:0]   vrfReadDataPorts_10_bits_vs,
  output [1:0]   vrfReadDataPorts_10_bits_offset,
  output [2:0]   vrfReadDataPorts_10_bits_instructionIndex,
  input          vrfReadDataPorts_11_ready,
  output         vrfReadDataPorts_11_valid,
  output [4:0]   vrfReadDataPorts_11_bits_vs,
  output [1:0]   vrfReadDataPorts_11_bits_offset,
  output [2:0]   vrfReadDataPorts_11_bits_instructionIndex,
  input          vrfReadDataPorts_12_ready,
  output         vrfReadDataPorts_12_valid,
  output [4:0]   vrfReadDataPorts_12_bits_vs,
  output [1:0]   vrfReadDataPorts_12_bits_offset,
  output [2:0]   vrfReadDataPorts_12_bits_instructionIndex,
  input          vrfReadDataPorts_13_ready,
  output         vrfReadDataPorts_13_valid,
  output [4:0]   vrfReadDataPorts_13_bits_vs,
  output [1:0]   vrfReadDataPorts_13_bits_offset,
  output [2:0]   vrfReadDataPorts_13_bits_instructionIndex,
  input          vrfReadDataPorts_14_ready,
  output         vrfReadDataPorts_14_valid,
  output [4:0]   vrfReadDataPorts_14_bits_vs,
  output [1:0]   vrfReadDataPorts_14_bits_offset,
  output [2:0]   vrfReadDataPorts_14_bits_instructionIndex,
  input          vrfReadDataPorts_15_ready,
  output         vrfReadDataPorts_15_valid,
  output [4:0]   vrfReadDataPorts_15_bits_vs,
  output [1:0]   vrfReadDataPorts_15_bits_offset,
  output [2:0]   vrfReadDataPorts_15_bits_instructionIndex,
  input          vrfReadResults_0_valid,
  input  [31:0]  vrfReadResults_0_bits,
  input          vrfReadResults_1_valid,
  input  [31:0]  vrfReadResults_1_bits,
  input          vrfReadResults_2_valid,
  input  [31:0]  vrfReadResults_2_bits,
  input          vrfReadResults_3_valid,
  input  [31:0]  vrfReadResults_3_bits,
  input          vrfReadResults_4_valid,
  input  [31:0]  vrfReadResults_4_bits,
  input          vrfReadResults_5_valid,
  input  [31:0]  vrfReadResults_5_bits,
  input          vrfReadResults_6_valid,
  input  [31:0]  vrfReadResults_6_bits,
  input          vrfReadResults_7_valid,
  input  [31:0]  vrfReadResults_7_bits,
  input          vrfReadResults_8_valid,
  input  [31:0]  vrfReadResults_8_bits,
  input          vrfReadResults_9_valid,
  input  [31:0]  vrfReadResults_9_bits,
  input          vrfReadResults_10_valid,
  input  [31:0]  vrfReadResults_10_bits,
  input          vrfReadResults_11_valid,
  input  [31:0]  vrfReadResults_11_bits,
  input          vrfReadResults_12_valid,
  input  [31:0]  vrfReadResults_12_bits,
  input          vrfReadResults_13_valid,
  input  [31:0]  vrfReadResults_13_bits,
  input          vrfReadResults_14_valid,
  input  [31:0]  vrfReadResults_14_bits,
  input          vrfReadResults_15_valid,
  input  [31:0]  vrfReadResults_15_bits,
  input          vrfWritePort_0_ready,
  output         vrfWritePort_0_valid,
  output [4:0]   vrfWritePort_0_bits_vd,
  output [1:0]   vrfWritePort_0_bits_offset,
  output [3:0]   vrfWritePort_0_bits_mask,
  output [31:0]  vrfWritePort_0_bits_data,
  output         vrfWritePort_0_bits_last,
  output [2:0]   vrfWritePort_0_bits_instructionIndex,
  input          vrfWritePort_1_ready,
  output         vrfWritePort_1_valid,
  output [4:0]   vrfWritePort_1_bits_vd,
  output [1:0]   vrfWritePort_1_bits_offset,
  output [3:0]   vrfWritePort_1_bits_mask,
  output [31:0]  vrfWritePort_1_bits_data,
  output         vrfWritePort_1_bits_last,
  output [2:0]   vrfWritePort_1_bits_instructionIndex,
  input          vrfWritePort_2_ready,
  output         vrfWritePort_2_valid,
  output [4:0]   vrfWritePort_2_bits_vd,
  output [1:0]   vrfWritePort_2_bits_offset,
  output [3:0]   vrfWritePort_2_bits_mask,
  output [31:0]  vrfWritePort_2_bits_data,
  output         vrfWritePort_2_bits_last,
  output [2:0]   vrfWritePort_2_bits_instructionIndex,
  input          vrfWritePort_3_ready,
  output         vrfWritePort_3_valid,
  output [4:0]   vrfWritePort_3_bits_vd,
  output [1:0]   vrfWritePort_3_bits_offset,
  output [3:0]   vrfWritePort_3_bits_mask,
  output [31:0]  vrfWritePort_3_bits_data,
  output         vrfWritePort_3_bits_last,
  output [2:0]   vrfWritePort_3_bits_instructionIndex,
  input          vrfWritePort_4_ready,
  output         vrfWritePort_4_valid,
  output [4:0]   vrfWritePort_4_bits_vd,
  output [1:0]   vrfWritePort_4_bits_offset,
  output [3:0]   vrfWritePort_4_bits_mask,
  output [31:0]  vrfWritePort_4_bits_data,
  output         vrfWritePort_4_bits_last,
  output [2:0]   vrfWritePort_4_bits_instructionIndex,
  input          vrfWritePort_5_ready,
  output         vrfWritePort_5_valid,
  output [4:0]   vrfWritePort_5_bits_vd,
  output [1:0]   vrfWritePort_5_bits_offset,
  output [3:0]   vrfWritePort_5_bits_mask,
  output [31:0]  vrfWritePort_5_bits_data,
  output         vrfWritePort_5_bits_last,
  output [2:0]   vrfWritePort_5_bits_instructionIndex,
  input          vrfWritePort_6_ready,
  output         vrfWritePort_6_valid,
  output [4:0]   vrfWritePort_6_bits_vd,
  output [1:0]   vrfWritePort_6_bits_offset,
  output [3:0]   vrfWritePort_6_bits_mask,
  output [31:0]  vrfWritePort_6_bits_data,
  output         vrfWritePort_6_bits_last,
  output [2:0]   vrfWritePort_6_bits_instructionIndex,
  input          vrfWritePort_7_ready,
  output         vrfWritePort_7_valid,
  output [4:0]   vrfWritePort_7_bits_vd,
  output [1:0]   vrfWritePort_7_bits_offset,
  output [3:0]   vrfWritePort_7_bits_mask,
  output [31:0]  vrfWritePort_7_bits_data,
  output         vrfWritePort_7_bits_last,
  output [2:0]   vrfWritePort_7_bits_instructionIndex,
  input          vrfWritePort_8_ready,
  output         vrfWritePort_8_valid,
  output [4:0]   vrfWritePort_8_bits_vd,
  output [1:0]   vrfWritePort_8_bits_offset,
  output [3:0]   vrfWritePort_8_bits_mask,
  output [31:0]  vrfWritePort_8_bits_data,
  output         vrfWritePort_8_bits_last,
  output [2:0]   vrfWritePort_8_bits_instructionIndex,
  input          vrfWritePort_9_ready,
  output         vrfWritePort_9_valid,
  output [4:0]   vrfWritePort_9_bits_vd,
  output [1:0]   vrfWritePort_9_bits_offset,
  output [3:0]   vrfWritePort_9_bits_mask,
  output [31:0]  vrfWritePort_9_bits_data,
  output         vrfWritePort_9_bits_last,
  output [2:0]   vrfWritePort_9_bits_instructionIndex,
  input          vrfWritePort_10_ready,
  output         vrfWritePort_10_valid,
  output [4:0]   vrfWritePort_10_bits_vd,
  output [1:0]   vrfWritePort_10_bits_offset,
  output [3:0]   vrfWritePort_10_bits_mask,
  output [31:0]  vrfWritePort_10_bits_data,
  output         vrfWritePort_10_bits_last,
  output [2:0]   vrfWritePort_10_bits_instructionIndex,
  input          vrfWritePort_11_ready,
  output         vrfWritePort_11_valid,
  output [4:0]   vrfWritePort_11_bits_vd,
  output [1:0]   vrfWritePort_11_bits_offset,
  output [3:0]   vrfWritePort_11_bits_mask,
  output [31:0]  vrfWritePort_11_bits_data,
  output         vrfWritePort_11_bits_last,
  output [2:0]   vrfWritePort_11_bits_instructionIndex,
  input          vrfWritePort_12_ready,
  output         vrfWritePort_12_valid,
  output [4:0]   vrfWritePort_12_bits_vd,
  output [1:0]   vrfWritePort_12_bits_offset,
  output [3:0]   vrfWritePort_12_bits_mask,
  output [31:0]  vrfWritePort_12_bits_data,
  output         vrfWritePort_12_bits_last,
  output [2:0]   vrfWritePort_12_bits_instructionIndex,
  input          vrfWritePort_13_ready,
  output         vrfWritePort_13_valid,
  output [4:0]   vrfWritePort_13_bits_vd,
  output [1:0]   vrfWritePort_13_bits_offset,
  output [3:0]   vrfWritePort_13_bits_mask,
  output [31:0]  vrfWritePort_13_bits_data,
  output         vrfWritePort_13_bits_last,
  output [2:0]   vrfWritePort_13_bits_instructionIndex,
  input          vrfWritePort_14_ready,
  output         vrfWritePort_14_valid,
  output [4:0]   vrfWritePort_14_bits_vd,
  output [1:0]   vrfWritePort_14_bits_offset,
  output [3:0]   vrfWritePort_14_bits_mask,
  output [31:0]  vrfWritePort_14_bits_data,
  output         vrfWritePort_14_bits_last,
  output [2:0]   vrfWritePort_14_bits_instructionIndex,
  input          vrfWritePort_15_ready,
  output         vrfWritePort_15_valid,
  output [4:0]   vrfWritePort_15_bits_vd,
  output [1:0]   vrfWritePort_15_bits_offset,
  output [3:0]   vrfWritePort_15_bits_mask,
  output [31:0]  vrfWritePort_15_bits_data,
  output         vrfWritePort_15_bits_last,
  output [2:0]   vrfWritePort_15_bits_instructionIndex,
  input          writeRelease_0,
                 writeRelease_1,
                 writeRelease_2,
                 writeRelease_3,
                 writeRelease_4,
                 writeRelease_5,
                 writeRelease_6,
                 writeRelease_7,
                 writeRelease_8,
                 writeRelease_9,
                 writeRelease_10,
                 writeRelease_11,
                 writeRelease_12,
                 writeRelease_13,
                 writeRelease_14,
                 writeRelease_15,
  output [7:0]   dataInWriteQueue_0,
                 dataInWriteQueue_1,
                 dataInWriteQueue_2,
                 dataInWriteQueue_3,
                 dataInWriteQueue_4,
                 dataInWriteQueue_5,
                 dataInWriteQueue_6,
                 dataInWriteQueue_7,
                 dataInWriteQueue_8,
                 dataInWriteQueue_9,
                 dataInWriteQueue_10,
                 dataInWriteQueue_11,
                 dataInWriteQueue_12,
                 dataInWriteQueue_13,
                 dataInWriteQueue_14,
                 dataInWriteQueue_15,
  input  [11:0]  csrInterface_vl,
                 csrInterface_vStart,
  input  [2:0]   csrInterface_vlmul,
  input  [1:0]   csrInterface_vSew,
                 csrInterface_vxrm,
  input          csrInterface_vta,
                 csrInterface_vma,
                 offsetReadResult_0_valid,
  input  [31:0]  offsetReadResult_0_bits,
  input          offsetReadResult_1_valid,
  input  [31:0]  offsetReadResult_1_bits,
  input          offsetReadResult_2_valid,
  input  [31:0]  offsetReadResult_2_bits,
  input          offsetReadResult_3_valid,
  input  [31:0]  offsetReadResult_3_bits,
  input          offsetReadResult_4_valid,
  input  [31:0]  offsetReadResult_4_bits,
  input          offsetReadResult_5_valid,
  input  [31:0]  offsetReadResult_5_bits,
  input          offsetReadResult_6_valid,
  input  [31:0]  offsetReadResult_6_bits,
  input          offsetReadResult_7_valid,
  input  [31:0]  offsetReadResult_7_bits,
  input          offsetReadResult_8_valid,
  input  [31:0]  offsetReadResult_8_bits,
  input          offsetReadResult_9_valid,
  input  [31:0]  offsetReadResult_9_bits,
  input          offsetReadResult_10_valid,
  input  [31:0]  offsetReadResult_10_bits,
  input          offsetReadResult_11_valid,
  input  [31:0]  offsetReadResult_11_bits,
  input          offsetReadResult_12_valid,
  input  [31:0]  offsetReadResult_12_bits,
  input          offsetReadResult_13_valid,
  input  [31:0]  offsetReadResult_13_bits,
  input          offsetReadResult_14_valid,
  input  [31:0]  offsetReadResult_14_bits,
  input          offsetReadResult_15_valid,
  input  [31:0]  offsetReadResult_15_bits,
  output [7:0]   lastReport,
  output [15:0]  tokenIO_offsetGroupRelease
);

  wire              _simpleDataQueue_fifo_empty;
  wire              _simpleDataQueue_fifo_full;
  wire              _simpleDataQueue_fifo_error;
  wire [77:0]       _simpleDataQueue_fifo_data_out;
  wire              _simpleSourceQueue_fifo_empty;
  wire              _simpleSourceQueue_fifo_full;
  wire              _simpleSourceQueue_fifo_error;
  wire              _dataQueue_fifo_empty;
  wire              _dataQueue_fifo_full;
  wire              _dataQueue_fifo_error;
  wire [613:0]      _dataQueue_fifo_data_out;
  wire              _sourceQueue_fifo_empty;
  wire              _sourceQueue_fifo_full;
  wire              _sourceQueue_fifo_error;
  wire              _writeIndexQueue_fifo_15_empty;
  wire              _writeIndexQueue_fifo_15_full;
  wire              _writeIndexQueue_fifo_15_error;
  wire              _writeIndexQueue_fifo_14_empty;
  wire              _writeIndexQueue_fifo_14_full;
  wire              _writeIndexQueue_fifo_14_error;
  wire              _writeIndexQueue_fifo_13_empty;
  wire              _writeIndexQueue_fifo_13_full;
  wire              _writeIndexQueue_fifo_13_error;
  wire              _writeIndexQueue_fifo_12_empty;
  wire              _writeIndexQueue_fifo_12_full;
  wire              _writeIndexQueue_fifo_12_error;
  wire              _writeIndexQueue_fifo_11_empty;
  wire              _writeIndexQueue_fifo_11_full;
  wire              _writeIndexQueue_fifo_11_error;
  wire              _writeIndexQueue_fifo_10_empty;
  wire              _writeIndexQueue_fifo_10_full;
  wire              _writeIndexQueue_fifo_10_error;
  wire              _writeIndexQueue_fifo_9_empty;
  wire              _writeIndexQueue_fifo_9_full;
  wire              _writeIndexQueue_fifo_9_error;
  wire              _writeIndexQueue_fifo_8_empty;
  wire              _writeIndexQueue_fifo_8_full;
  wire              _writeIndexQueue_fifo_8_error;
  wire              _writeIndexQueue_fifo_7_empty;
  wire              _writeIndexQueue_fifo_7_full;
  wire              _writeIndexQueue_fifo_7_error;
  wire              _writeIndexQueue_fifo_6_empty;
  wire              _writeIndexQueue_fifo_6_full;
  wire              _writeIndexQueue_fifo_6_error;
  wire              _writeIndexQueue_fifo_5_empty;
  wire              _writeIndexQueue_fifo_5_full;
  wire              _writeIndexQueue_fifo_5_error;
  wire              _writeIndexQueue_fifo_4_empty;
  wire              _writeIndexQueue_fifo_4_full;
  wire              _writeIndexQueue_fifo_4_error;
  wire              _writeIndexQueue_fifo_3_empty;
  wire              _writeIndexQueue_fifo_3_full;
  wire              _writeIndexQueue_fifo_3_error;
  wire              _writeIndexQueue_fifo_2_empty;
  wire              _writeIndexQueue_fifo_2_full;
  wire              _writeIndexQueue_fifo_2_error;
  wire              _writeIndexQueue_fifo_1_empty;
  wire              _writeIndexQueue_fifo_1_full;
  wire              _writeIndexQueue_fifo_1_error;
  wire              _writeIndexQueue_fifo_empty;
  wire              _writeIndexQueue_fifo_full;
  wire              _writeIndexQueue_fifo_error;
  wire              _otherUnitDataQueueVec_fifo_15_empty;
  wire              _otherUnitDataQueueVec_fifo_15_full;
  wire              _otherUnitDataQueueVec_fifo_15_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_15_data_out;
  wire              _otherUnitDataQueueVec_fifo_14_empty;
  wire              _otherUnitDataQueueVec_fifo_14_full;
  wire              _otherUnitDataQueueVec_fifo_14_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_14_data_out;
  wire              _otherUnitDataQueueVec_fifo_13_empty;
  wire              _otherUnitDataQueueVec_fifo_13_full;
  wire              _otherUnitDataQueueVec_fifo_13_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_13_data_out;
  wire              _otherUnitDataQueueVec_fifo_12_empty;
  wire              _otherUnitDataQueueVec_fifo_12_full;
  wire              _otherUnitDataQueueVec_fifo_12_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_12_data_out;
  wire              _otherUnitDataQueueVec_fifo_11_empty;
  wire              _otherUnitDataQueueVec_fifo_11_full;
  wire              _otherUnitDataQueueVec_fifo_11_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_11_data_out;
  wire              _otherUnitDataQueueVec_fifo_10_empty;
  wire              _otherUnitDataQueueVec_fifo_10_full;
  wire              _otherUnitDataQueueVec_fifo_10_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_10_data_out;
  wire              _otherUnitDataQueueVec_fifo_9_empty;
  wire              _otherUnitDataQueueVec_fifo_9_full;
  wire              _otherUnitDataQueueVec_fifo_9_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_9_data_out;
  wire              _otherUnitDataQueueVec_fifo_8_empty;
  wire              _otherUnitDataQueueVec_fifo_8_full;
  wire              _otherUnitDataQueueVec_fifo_8_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_8_data_out;
  wire              _otherUnitDataQueueVec_fifo_7_empty;
  wire              _otherUnitDataQueueVec_fifo_7_full;
  wire              _otherUnitDataQueueVec_fifo_7_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_7_data_out;
  wire              _otherUnitDataQueueVec_fifo_6_empty;
  wire              _otherUnitDataQueueVec_fifo_6_full;
  wire              _otherUnitDataQueueVec_fifo_6_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_6_data_out;
  wire              _otherUnitDataQueueVec_fifo_5_empty;
  wire              _otherUnitDataQueueVec_fifo_5_full;
  wire              _otherUnitDataQueueVec_fifo_5_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_5_data_out;
  wire              _otherUnitDataQueueVec_fifo_4_empty;
  wire              _otherUnitDataQueueVec_fifo_4_full;
  wire              _otherUnitDataQueueVec_fifo_4_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_4_data_out;
  wire              _otherUnitDataQueueVec_fifo_3_empty;
  wire              _otherUnitDataQueueVec_fifo_3_full;
  wire              _otherUnitDataQueueVec_fifo_3_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_3_data_out;
  wire              _otherUnitDataQueueVec_fifo_2_empty;
  wire              _otherUnitDataQueueVec_fifo_2_full;
  wire              _otherUnitDataQueueVec_fifo_2_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_2_data_out;
  wire              _otherUnitDataQueueVec_fifo_1_empty;
  wire              _otherUnitDataQueueVec_fifo_1_full;
  wire              _otherUnitDataQueueVec_fifo_1_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_1_data_out;
  wire              _otherUnitDataQueueVec_fifo_empty;
  wire              _otherUnitDataQueueVec_fifo_full;
  wire              _otherUnitDataQueueVec_fifo_error;
  wire [31:0]       _otherUnitDataQueueVec_fifo_data_out;
  wire              _otherUnitTargetQueue_fifo_empty;
  wire              _otherUnitTargetQueue_fifo_full;
  wire              _otherUnitTargetQueue_fifo_error;
  wire              _writeQueueVec_fifo_15_empty;
  wire              _writeQueueVec_fifo_15_full;
  wire              _writeQueueVec_fifo_15_error;
  wire [62:0]       _writeQueueVec_fifo_15_data_out;
  wire              _writeQueueVec_fifo_14_empty;
  wire              _writeQueueVec_fifo_14_full;
  wire              _writeQueueVec_fifo_14_error;
  wire [62:0]       _writeQueueVec_fifo_14_data_out;
  wire              _writeQueueVec_fifo_13_empty;
  wire              _writeQueueVec_fifo_13_full;
  wire              _writeQueueVec_fifo_13_error;
  wire [62:0]       _writeQueueVec_fifo_13_data_out;
  wire              _writeQueueVec_fifo_12_empty;
  wire              _writeQueueVec_fifo_12_full;
  wire              _writeQueueVec_fifo_12_error;
  wire [62:0]       _writeQueueVec_fifo_12_data_out;
  wire              _writeQueueVec_fifo_11_empty;
  wire              _writeQueueVec_fifo_11_full;
  wire              _writeQueueVec_fifo_11_error;
  wire [62:0]       _writeQueueVec_fifo_11_data_out;
  wire              _writeQueueVec_fifo_10_empty;
  wire              _writeQueueVec_fifo_10_full;
  wire              _writeQueueVec_fifo_10_error;
  wire [62:0]       _writeQueueVec_fifo_10_data_out;
  wire              _writeQueueVec_fifo_9_empty;
  wire              _writeQueueVec_fifo_9_full;
  wire              _writeQueueVec_fifo_9_error;
  wire [62:0]       _writeQueueVec_fifo_9_data_out;
  wire              _writeQueueVec_fifo_8_empty;
  wire              _writeQueueVec_fifo_8_full;
  wire              _writeQueueVec_fifo_8_error;
  wire [62:0]       _writeQueueVec_fifo_8_data_out;
  wire              _writeQueueVec_fifo_7_empty;
  wire              _writeQueueVec_fifo_7_full;
  wire              _writeQueueVec_fifo_7_error;
  wire [62:0]       _writeQueueVec_fifo_7_data_out;
  wire              _writeQueueVec_fifo_6_empty;
  wire              _writeQueueVec_fifo_6_full;
  wire              _writeQueueVec_fifo_6_error;
  wire [62:0]       _writeQueueVec_fifo_6_data_out;
  wire              _writeQueueVec_fifo_5_empty;
  wire              _writeQueueVec_fifo_5_full;
  wire              _writeQueueVec_fifo_5_error;
  wire [62:0]       _writeQueueVec_fifo_5_data_out;
  wire              _writeQueueVec_fifo_4_empty;
  wire              _writeQueueVec_fifo_4_full;
  wire              _writeQueueVec_fifo_4_error;
  wire [62:0]       _writeQueueVec_fifo_4_data_out;
  wire              _writeQueueVec_fifo_3_empty;
  wire              _writeQueueVec_fifo_3_full;
  wire              _writeQueueVec_fifo_3_error;
  wire [62:0]       _writeQueueVec_fifo_3_data_out;
  wire              _writeQueueVec_fifo_2_empty;
  wire              _writeQueueVec_fifo_2_full;
  wire              _writeQueueVec_fifo_2_error;
  wire [62:0]       _writeQueueVec_fifo_2_data_out;
  wire              _writeQueueVec_fifo_1_empty;
  wire              _writeQueueVec_fifo_1_full;
  wire              _writeQueueVec_fifo_1_error;
  wire [62:0]       _writeQueueVec_fifo_1_data_out;
  wire              _writeQueueVec_fifo_empty;
  wire              _writeQueueVec_fifo_full;
  wire              _writeQueueVec_fifo_error;
  wire [62:0]       _writeQueueVec_fifo_data_out;
  wire              _otherUnit_vrfReadDataPorts_valid;
  wire [4:0]        _otherUnit_vrfReadDataPorts_bits_vs;
  wire [1:0]        _otherUnit_vrfReadDataPorts_bits_offset;
  wire [2:0]        _otherUnit_vrfReadDataPorts_bits_instructionIndex;
  wire              _otherUnit_maskSelect_valid;
  wire [4:0]        _otherUnit_maskSelect_bits;
  wire              _otherUnit_memReadRequest_valid;
  wire              _otherUnit_memWriteRequest_valid;
  wire [7:0]        _otherUnit_memWriteRequest_bits_source;
  wire [31:0]       _otherUnit_memWriteRequest_bits_address;
  wire [1:0]        _otherUnit_memWriteRequest_bits_size;
  wire              _otherUnit_vrfWritePort_valid;
  wire [4:0]        _otherUnit_vrfWritePort_bits_vd;
  wire [1:0]        _otherUnit_vrfWritePort_bits_offset;
  wire [3:0]        _otherUnit_vrfWritePort_bits_mask;
  wire [31:0]       _otherUnit_vrfWritePort_bits_data;
  wire              _otherUnit_vrfWritePort_bits_last;
  wire [2:0]        _otherUnit_vrfWritePort_bits_instructionIndex;
  wire              _otherUnit_status_idle;
  wire              _otherUnit_status_last;
  wire [2:0]        _otherUnit_status_instructionIndex;
  wire [15:0]       _otherUnit_status_targetLane;
  wire              _otherUnit_status_isStore;
  wire              _otherUnit_offsetRelease_0;
  wire              _otherUnit_offsetRelease_1;
  wire              _otherUnit_offsetRelease_2;
  wire              _otherUnit_offsetRelease_3;
  wire              _otherUnit_offsetRelease_4;
  wire              _otherUnit_offsetRelease_5;
  wire              _otherUnit_offsetRelease_6;
  wire              _otherUnit_offsetRelease_7;
  wire              _otherUnit_offsetRelease_8;
  wire              _otherUnit_offsetRelease_9;
  wire              _otherUnit_offsetRelease_10;
  wire              _otherUnit_offsetRelease_11;
  wire              _otherUnit_offsetRelease_12;
  wire              _otherUnit_offsetRelease_13;
  wire              _otherUnit_offsetRelease_14;
  wire              _otherUnit_offsetRelease_15;
  wire              _storeUnit_maskSelect_valid;
  wire [4:0]        _storeUnit_maskSelect_bits;
  wire              _storeUnit_memRequest_valid;
  wire [5:0]        _storeUnit_memRequest_bits_index;
  wire [31:0]       _storeUnit_memRequest_bits_address;
  wire              _storeUnit_status_idle;
  wire              _storeUnit_status_last;
  wire [2:0]        _storeUnit_status_instructionIndex;
  wire [31:0]       _storeUnit_status_startAddress;
  wire [31:0]       _storeUnit_status_endAddress;
  wire              _storeUnit_vrfReadDataPorts_0_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_0_bits_vs;
  wire [1:0]        _storeUnit_vrfReadDataPorts_0_bits_offset;
  wire [2:0]        _storeUnit_vrfReadDataPorts_0_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_1_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_1_bits_vs;
  wire [1:0]        _storeUnit_vrfReadDataPorts_1_bits_offset;
  wire [2:0]        _storeUnit_vrfReadDataPorts_1_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_2_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_2_bits_vs;
  wire [1:0]        _storeUnit_vrfReadDataPorts_2_bits_offset;
  wire [2:0]        _storeUnit_vrfReadDataPorts_2_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_3_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_3_bits_vs;
  wire [1:0]        _storeUnit_vrfReadDataPorts_3_bits_offset;
  wire [2:0]        _storeUnit_vrfReadDataPorts_3_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_4_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_4_bits_vs;
  wire [1:0]        _storeUnit_vrfReadDataPorts_4_bits_offset;
  wire [2:0]        _storeUnit_vrfReadDataPorts_4_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_5_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_5_bits_vs;
  wire [1:0]        _storeUnit_vrfReadDataPorts_5_bits_offset;
  wire [2:0]        _storeUnit_vrfReadDataPorts_5_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_6_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_6_bits_vs;
  wire [1:0]        _storeUnit_vrfReadDataPorts_6_bits_offset;
  wire [2:0]        _storeUnit_vrfReadDataPorts_6_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_7_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_7_bits_vs;
  wire [1:0]        _storeUnit_vrfReadDataPorts_7_bits_offset;
  wire [2:0]        _storeUnit_vrfReadDataPorts_7_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_8_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_8_bits_vs;
  wire [1:0]        _storeUnit_vrfReadDataPorts_8_bits_offset;
  wire [2:0]        _storeUnit_vrfReadDataPorts_8_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_9_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_9_bits_vs;
  wire [1:0]        _storeUnit_vrfReadDataPorts_9_bits_offset;
  wire [2:0]        _storeUnit_vrfReadDataPorts_9_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_10_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_10_bits_vs;
  wire [1:0]        _storeUnit_vrfReadDataPorts_10_bits_offset;
  wire [2:0]        _storeUnit_vrfReadDataPorts_10_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_11_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_11_bits_vs;
  wire [1:0]        _storeUnit_vrfReadDataPorts_11_bits_offset;
  wire [2:0]        _storeUnit_vrfReadDataPorts_11_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_12_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_12_bits_vs;
  wire [1:0]        _storeUnit_vrfReadDataPorts_12_bits_offset;
  wire [2:0]        _storeUnit_vrfReadDataPorts_12_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_13_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_13_bits_vs;
  wire [1:0]        _storeUnit_vrfReadDataPorts_13_bits_offset;
  wire [2:0]        _storeUnit_vrfReadDataPorts_13_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_14_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_14_bits_vs;
  wire [1:0]        _storeUnit_vrfReadDataPorts_14_bits_offset;
  wire [2:0]        _storeUnit_vrfReadDataPorts_14_bits_instructionIndex;
  wire              _storeUnit_vrfReadDataPorts_15_valid;
  wire [4:0]        _storeUnit_vrfReadDataPorts_15_bits_vs;
  wire [1:0]        _storeUnit_vrfReadDataPorts_15_bits_offset;
  wire [2:0]        _storeUnit_vrfReadDataPorts_15_bits_instructionIndex;
  wire              _loadUnit_maskSelect_valid;
  wire [4:0]        _loadUnit_maskSelect_bits;
  wire              _loadUnit_memRequest_valid;
  wire              _loadUnit_status_idle;
  wire              _loadUnit_status_last;
  wire [2:0]        _loadUnit_status_instructionIndex;
  wire [31:0]       _loadUnit_status_startAddress;
  wire [31:0]       _loadUnit_status_endAddress;
  wire              _loadUnit_vrfWritePort_0_valid;
  wire [4:0]        _loadUnit_vrfWritePort_0_bits_vd;
  wire [1:0]        _loadUnit_vrfWritePort_0_bits_offset;
  wire [3:0]        _loadUnit_vrfWritePort_0_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_0_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_0_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_1_valid;
  wire [4:0]        _loadUnit_vrfWritePort_1_bits_vd;
  wire [1:0]        _loadUnit_vrfWritePort_1_bits_offset;
  wire [3:0]        _loadUnit_vrfWritePort_1_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_1_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_1_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_2_valid;
  wire [4:0]        _loadUnit_vrfWritePort_2_bits_vd;
  wire [1:0]        _loadUnit_vrfWritePort_2_bits_offset;
  wire [3:0]        _loadUnit_vrfWritePort_2_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_2_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_2_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_3_valid;
  wire [4:0]        _loadUnit_vrfWritePort_3_bits_vd;
  wire [1:0]        _loadUnit_vrfWritePort_3_bits_offset;
  wire [3:0]        _loadUnit_vrfWritePort_3_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_3_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_3_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_4_valid;
  wire [4:0]        _loadUnit_vrfWritePort_4_bits_vd;
  wire [1:0]        _loadUnit_vrfWritePort_4_bits_offset;
  wire [3:0]        _loadUnit_vrfWritePort_4_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_4_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_4_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_5_valid;
  wire [4:0]        _loadUnit_vrfWritePort_5_bits_vd;
  wire [1:0]        _loadUnit_vrfWritePort_5_bits_offset;
  wire [3:0]        _loadUnit_vrfWritePort_5_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_5_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_5_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_6_valid;
  wire [4:0]        _loadUnit_vrfWritePort_6_bits_vd;
  wire [1:0]        _loadUnit_vrfWritePort_6_bits_offset;
  wire [3:0]        _loadUnit_vrfWritePort_6_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_6_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_6_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_7_valid;
  wire [4:0]        _loadUnit_vrfWritePort_7_bits_vd;
  wire [1:0]        _loadUnit_vrfWritePort_7_bits_offset;
  wire [3:0]        _loadUnit_vrfWritePort_7_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_7_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_7_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_8_valid;
  wire [4:0]        _loadUnit_vrfWritePort_8_bits_vd;
  wire [1:0]        _loadUnit_vrfWritePort_8_bits_offset;
  wire [3:0]        _loadUnit_vrfWritePort_8_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_8_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_8_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_9_valid;
  wire [4:0]        _loadUnit_vrfWritePort_9_bits_vd;
  wire [1:0]        _loadUnit_vrfWritePort_9_bits_offset;
  wire [3:0]        _loadUnit_vrfWritePort_9_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_9_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_9_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_10_valid;
  wire [4:0]        _loadUnit_vrfWritePort_10_bits_vd;
  wire [1:0]        _loadUnit_vrfWritePort_10_bits_offset;
  wire [3:0]        _loadUnit_vrfWritePort_10_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_10_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_10_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_11_valid;
  wire [4:0]        _loadUnit_vrfWritePort_11_bits_vd;
  wire [1:0]        _loadUnit_vrfWritePort_11_bits_offset;
  wire [3:0]        _loadUnit_vrfWritePort_11_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_11_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_11_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_12_valid;
  wire [4:0]        _loadUnit_vrfWritePort_12_bits_vd;
  wire [1:0]        _loadUnit_vrfWritePort_12_bits_offset;
  wire [3:0]        _loadUnit_vrfWritePort_12_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_12_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_12_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_13_valid;
  wire [4:0]        _loadUnit_vrfWritePort_13_bits_vd;
  wire [1:0]        _loadUnit_vrfWritePort_13_bits_offset;
  wire [3:0]        _loadUnit_vrfWritePort_13_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_13_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_13_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_14_valid;
  wire [4:0]        _loadUnit_vrfWritePort_14_bits_vd;
  wire [1:0]        _loadUnit_vrfWritePort_14_bits_offset;
  wire [3:0]        _loadUnit_vrfWritePort_14_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_14_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_14_bits_instructionIndex;
  wire              _loadUnit_vrfWritePort_15_valid;
  wire [4:0]        _loadUnit_vrfWritePort_15_bits_vd;
  wire [1:0]        _loadUnit_vrfWritePort_15_bits_offset;
  wire [3:0]        _loadUnit_vrfWritePort_15_bits_mask;
  wire [31:0]       _loadUnit_vrfWritePort_15_bits_data;
  wire [2:0]        _loadUnit_vrfWritePort_15_bits_instructionIndex;
  wire              simpleDataQueue_almostFull;
  wire              simpleDataQueue_almostEmpty;
  wire              simpleSourceQueue_almostFull;
  wire              simpleSourceQueue_almostEmpty;
  wire              dataQueue_almostFull;
  wire              dataQueue_almostEmpty;
  wire              sourceQueue_almostFull;
  wire              sourceQueue_almostEmpty;
  wire              writeIndexQueue_15_almostFull;
  wire              writeIndexQueue_15_almostEmpty;
  wire              writeIndexQueue_14_almostFull;
  wire              writeIndexQueue_14_almostEmpty;
  wire              writeIndexQueue_13_almostFull;
  wire              writeIndexQueue_13_almostEmpty;
  wire              writeIndexQueue_12_almostFull;
  wire              writeIndexQueue_12_almostEmpty;
  wire              writeIndexQueue_11_almostFull;
  wire              writeIndexQueue_11_almostEmpty;
  wire              writeIndexQueue_10_almostFull;
  wire              writeIndexQueue_10_almostEmpty;
  wire              writeIndexQueue_9_almostFull;
  wire              writeIndexQueue_9_almostEmpty;
  wire              writeIndexQueue_8_almostFull;
  wire              writeIndexQueue_8_almostEmpty;
  wire              writeIndexQueue_7_almostFull;
  wire              writeIndexQueue_7_almostEmpty;
  wire              writeIndexQueue_6_almostFull;
  wire              writeIndexQueue_6_almostEmpty;
  wire              writeIndexQueue_5_almostFull;
  wire              writeIndexQueue_5_almostEmpty;
  wire              writeIndexQueue_4_almostFull;
  wire              writeIndexQueue_4_almostEmpty;
  wire              writeIndexQueue_3_almostFull;
  wire              writeIndexQueue_3_almostEmpty;
  wire              writeIndexQueue_2_almostFull;
  wire              writeIndexQueue_2_almostEmpty;
  wire              writeIndexQueue_1_almostFull;
  wire              writeIndexQueue_1_almostEmpty;
  wire              writeIndexQueue_almostFull;
  wire              writeIndexQueue_almostEmpty;
  wire              otherUnitDataQueueVec_15_almostFull;
  wire              otherUnitDataQueueVec_15_almostEmpty;
  wire              otherUnitDataQueueVec_14_almostFull;
  wire              otherUnitDataQueueVec_14_almostEmpty;
  wire              otherUnitDataQueueVec_13_almostFull;
  wire              otherUnitDataQueueVec_13_almostEmpty;
  wire              otherUnitDataQueueVec_12_almostFull;
  wire              otherUnitDataQueueVec_12_almostEmpty;
  wire              otherUnitDataQueueVec_11_almostFull;
  wire              otherUnitDataQueueVec_11_almostEmpty;
  wire              otherUnitDataQueueVec_10_almostFull;
  wire              otherUnitDataQueueVec_10_almostEmpty;
  wire              otherUnitDataQueueVec_9_almostFull;
  wire              otherUnitDataQueueVec_9_almostEmpty;
  wire              otherUnitDataQueueVec_8_almostFull;
  wire              otherUnitDataQueueVec_8_almostEmpty;
  wire              otherUnitDataQueueVec_7_almostFull;
  wire              otherUnitDataQueueVec_7_almostEmpty;
  wire              otherUnitDataQueueVec_6_almostFull;
  wire              otherUnitDataQueueVec_6_almostEmpty;
  wire              otherUnitDataQueueVec_5_almostFull;
  wire              otherUnitDataQueueVec_5_almostEmpty;
  wire              otherUnitDataQueueVec_4_almostFull;
  wire              otherUnitDataQueueVec_4_almostEmpty;
  wire              otherUnitDataQueueVec_3_almostFull;
  wire              otherUnitDataQueueVec_3_almostEmpty;
  wire              otherUnitDataQueueVec_2_almostFull;
  wire              otherUnitDataQueueVec_2_almostEmpty;
  wire              otherUnitDataQueueVec_1_almostFull;
  wire              otherUnitDataQueueVec_1_almostEmpty;
  wire              otherUnitDataQueueVec_0_almostFull;
  wire              otherUnitDataQueueVec_0_almostEmpty;
  wire              otherUnitTargetQueue_almostFull;
  wire              otherUnitTargetQueue_almostEmpty;
  wire              writeQueueVec_15_almostFull;
  wire              writeQueueVec_15_almostEmpty;
  wire              writeQueueVec_14_almostFull;
  wire              writeQueueVec_14_almostEmpty;
  wire              writeQueueVec_13_almostFull;
  wire              writeQueueVec_13_almostEmpty;
  wire              writeQueueVec_12_almostFull;
  wire              writeQueueVec_12_almostEmpty;
  wire              writeQueueVec_11_almostFull;
  wire              writeQueueVec_11_almostEmpty;
  wire              writeQueueVec_10_almostFull;
  wire              writeQueueVec_10_almostEmpty;
  wire              writeQueueVec_9_almostFull;
  wire              writeQueueVec_9_almostEmpty;
  wire              writeQueueVec_8_almostFull;
  wire              writeQueueVec_8_almostEmpty;
  wire              writeQueueVec_7_almostFull;
  wire              writeQueueVec_7_almostEmpty;
  wire              writeQueueVec_6_almostFull;
  wire              writeQueueVec_6_almostEmpty;
  wire              writeQueueVec_5_almostFull;
  wire              writeQueueVec_5_almostEmpty;
  wire              writeQueueVec_4_almostFull;
  wire              writeQueueVec_4_almostEmpty;
  wire              writeQueueVec_3_almostFull;
  wire              writeQueueVec_3_almostEmpty;
  wire              writeQueueVec_2_almostFull;
  wire              writeQueueVec_2_almostEmpty;
  wire              writeQueueVec_1_almostFull;
  wire              writeQueueVec_1_almostEmpty;
  wire              writeQueueVec_0_almostFull;
  wire              writeQueueVec_0_almostEmpty;
  wire [8:0]        simpleSourceQueue_enq_bits;
  wire [31:0]       simpleAccessPorts_ar_bits_addr_0;
  wire [5:0]        sourceQueue_enq_bits;
  wire [31:0]       axi4Port_ar_bits_addr_0;
  wire              request_valid_0 = request_valid;
  wire [2:0]        request_bits_instructionInformation_nf_0 = request_bits_instructionInformation_nf;
  wire              request_bits_instructionInformation_mew_0 = request_bits_instructionInformation_mew;
  wire [1:0]        request_bits_instructionInformation_mop_0 = request_bits_instructionInformation_mop;
  wire [4:0]        request_bits_instructionInformation_lumop_0 = request_bits_instructionInformation_lumop;
  wire [1:0]        request_bits_instructionInformation_eew_0 = request_bits_instructionInformation_eew;
  wire [4:0]        request_bits_instructionInformation_vs3_0 = request_bits_instructionInformation_vs3;
  wire              request_bits_instructionInformation_isStore_0 = request_bits_instructionInformation_isStore;
  wire              request_bits_instructionInformation_maskedLoadStore_0 = request_bits_instructionInformation_maskedLoadStore;
  wire [31:0]       request_bits_rs1Data_0 = request_bits_rs1Data;
  wire [31:0]       request_bits_rs2Data_0 = request_bits_rs2Data;
  wire [2:0]        request_bits_instructionIndex_0 = request_bits_instructionIndex;
  wire              axi4Port_aw_ready_0 = axi4Port_aw_ready;
  wire              axi4Port_w_ready_0 = axi4Port_w_ready;
  wire              axi4Port_b_valid_0 = axi4Port_b_valid;
  wire [1:0]        axi4Port_b_bits_id_0 = axi4Port_b_bits_id;
  wire [1:0]        axi4Port_b_bits_resp_0 = axi4Port_b_bits_resp;
  wire              axi4Port_ar_ready_0 = axi4Port_ar_ready;
  wire              axi4Port_r_valid_0 = axi4Port_r_valid;
  wire [1:0]        axi4Port_r_bits_id_0 = axi4Port_r_bits_id;
  wire [511:0]      axi4Port_r_bits_data_0 = axi4Port_r_bits_data;
  wire [1:0]        axi4Port_r_bits_resp_0 = axi4Port_r_bits_resp;
  wire              axi4Port_r_bits_last_0 = axi4Port_r_bits_last;
  wire              simpleAccessPorts_aw_ready_0 = simpleAccessPorts_aw_ready;
  wire              simpleAccessPorts_w_ready_0 = simpleAccessPorts_w_ready;
  wire              simpleAccessPorts_b_valid_0 = simpleAccessPorts_b_valid;
  wire [1:0]        simpleAccessPorts_b_bits_id_0 = simpleAccessPorts_b_bits_id;
  wire [1:0]        simpleAccessPorts_b_bits_resp_0 = simpleAccessPorts_b_bits_resp;
  wire              simpleAccessPorts_ar_ready_0 = simpleAccessPorts_ar_ready;
  wire              simpleAccessPorts_r_valid_0 = simpleAccessPorts_r_valid;
  wire [1:0]        simpleAccessPorts_r_bits_id_0 = simpleAccessPorts_r_bits_id;
  wire [31:0]       simpleAccessPorts_r_bits_data_0 = simpleAccessPorts_r_bits_data;
  wire [1:0]        simpleAccessPorts_r_bits_resp_0 = simpleAccessPorts_r_bits_resp;
  wire              simpleAccessPorts_r_bits_last_0 = simpleAccessPorts_r_bits_last;
  wire              vrfReadDataPorts_0_ready_0 = vrfReadDataPorts_0_ready;
  wire              vrfReadDataPorts_1_ready_0 = vrfReadDataPorts_1_ready;
  wire              vrfReadDataPorts_2_ready_0 = vrfReadDataPorts_2_ready;
  wire              vrfReadDataPorts_3_ready_0 = vrfReadDataPorts_3_ready;
  wire              vrfReadDataPorts_4_ready_0 = vrfReadDataPorts_4_ready;
  wire              vrfReadDataPorts_5_ready_0 = vrfReadDataPorts_5_ready;
  wire              vrfReadDataPorts_6_ready_0 = vrfReadDataPorts_6_ready;
  wire              vrfReadDataPorts_7_ready_0 = vrfReadDataPorts_7_ready;
  wire              vrfReadDataPorts_8_ready_0 = vrfReadDataPorts_8_ready;
  wire              vrfReadDataPorts_9_ready_0 = vrfReadDataPorts_9_ready;
  wire              vrfReadDataPorts_10_ready_0 = vrfReadDataPorts_10_ready;
  wire              vrfReadDataPorts_11_ready_0 = vrfReadDataPorts_11_ready;
  wire              vrfReadDataPorts_12_ready_0 = vrfReadDataPorts_12_ready;
  wire              vrfReadDataPorts_13_ready_0 = vrfReadDataPorts_13_ready;
  wire              vrfReadDataPorts_14_ready_0 = vrfReadDataPorts_14_ready;
  wire              vrfReadDataPorts_15_ready_0 = vrfReadDataPorts_15_ready;
  wire              vrfWritePort_0_ready_0 = vrfWritePort_0_ready;
  wire              vrfWritePort_1_ready_0 = vrfWritePort_1_ready;
  wire              vrfWritePort_2_ready_0 = vrfWritePort_2_ready;
  wire              vrfWritePort_3_ready_0 = vrfWritePort_3_ready;
  wire              vrfWritePort_4_ready_0 = vrfWritePort_4_ready;
  wire              vrfWritePort_5_ready_0 = vrfWritePort_5_ready;
  wire              vrfWritePort_6_ready_0 = vrfWritePort_6_ready;
  wire              vrfWritePort_7_ready_0 = vrfWritePort_7_ready;
  wire              vrfWritePort_8_ready_0 = vrfWritePort_8_ready;
  wire              vrfWritePort_9_ready_0 = vrfWritePort_9_ready;
  wire              vrfWritePort_10_ready_0 = vrfWritePort_10_ready;
  wire              vrfWritePort_11_ready_0 = vrfWritePort_11_ready;
  wire              vrfWritePort_12_ready_0 = vrfWritePort_12_ready;
  wire              vrfWritePort_13_ready_0 = vrfWritePort_13_ready;
  wire              vrfWritePort_14_ready_0 = vrfWritePort_14_ready;
  wire              vrfWritePort_15_ready_0 = vrfWritePort_15_ready;
  wire [31:0]       otherUnitDataQueueVec_0_enq_bits = vrfReadResults_0_bits;
  wire [31:0]       otherUnitDataQueueVec_1_enq_bits = vrfReadResults_1_bits;
  wire [31:0]       otherUnitDataQueueVec_2_enq_bits = vrfReadResults_2_bits;
  wire [31:0]       otherUnitDataQueueVec_3_enq_bits = vrfReadResults_3_bits;
  wire [31:0]       otherUnitDataQueueVec_4_enq_bits = vrfReadResults_4_bits;
  wire [31:0]       otherUnitDataQueueVec_5_enq_bits = vrfReadResults_5_bits;
  wire [31:0]       otherUnitDataQueueVec_6_enq_bits = vrfReadResults_6_bits;
  wire [31:0]       otherUnitDataQueueVec_7_enq_bits = vrfReadResults_7_bits;
  wire [31:0]       otherUnitDataQueueVec_8_enq_bits = vrfReadResults_8_bits;
  wire [31:0]       otherUnitDataQueueVec_9_enq_bits = vrfReadResults_9_bits;
  wire [31:0]       otherUnitDataQueueVec_10_enq_bits = vrfReadResults_10_bits;
  wire [31:0]       otherUnitDataQueueVec_11_enq_bits = vrfReadResults_11_bits;
  wire [31:0]       otherUnitDataQueueVec_12_enq_bits = vrfReadResults_12_bits;
  wire [31:0]       otherUnitDataQueueVec_13_enq_bits = vrfReadResults_13_bits;
  wire [31:0]       otherUnitDataQueueVec_14_enq_bits = vrfReadResults_14_bits;
  wire [31:0]       otherUnitDataQueueVec_15_enq_bits = vrfReadResults_15_bits;
  wire              writeIndexQueue_deq_ready = writeRelease_0;
  wire              writeIndexQueue_1_deq_ready = writeRelease_1;
  wire              writeIndexQueue_2_deq_ready = writeRelease_2;
  wire              writeIndexQueue_3_deq_ready = writeRelease_3;
  wire              writeIndexQueue_4_deq_ready = writeRelease_4;
  wire              writeIndexQueue_5_deq_ready = writeRelease_5;
  wire              writeIndexQueue_6_deq_ready = writeRelease_6;
  wire              writeIndexQueue_7_deq_ready = writeRelease_7;
  wire              writeIndexQueue_8_deq_ready = writeRelease_8;
  wire              writeIndexQueue_9_deq_ready = writeRelease_9;
  wire              writeIndexQueue_10_deq_ready = writeRelease_10;
  wire              writeIndexQueue_11_deq_ready = writeRelease_11;
  wire              writeIndexQueue_12_deq_ready = writeRelease_12;
  wire              writeIndexQueue_13_deq_ready = writeRelease_13;
  wire              writeIndexQueue_14_deq_ready = writeRelease_14;
  wire              writeIndexQueue_15_deq_ready = writeRelease_15;
  wire [3:0]        axi4Port_aw_bits_cache = 4'h0;
  wire [3:0]        axi4Port_aw_bits_qos = 4'h0;
  wire [3:0]        axi4Port_aw_bits_region = 4'h0;
  wire [3:0]        axi4Port_ar_bits_cache = 4'h0;
  wire [3:0]        axi4Port_ar_bits_qos = 4'h0;
  wire [3:0]        axi4Port_ar_bits_region = 4'h0;
  wire [3:0]        simpleAccessPorts_aw_bits_cache = 4'h0;
  wire [3:0]        simpleAccessPorts_aw_bits_qos = 4'h0;
  wire [3:0]        simpleAccessPorts_aw_bits_region = 4'h0;
  wire [3:0]        simpleAccessPorts_ar_bits_cache = 4'h0;
  wire [3:0]        simpleAccessPorts_ar_bits_qos = 4'h0;
  wire [3:0]        simpleAccessPorts_ar_bits_region = 4'h0;
  wire [15:0]       writeQueueVec_0_enq_bits_targetLane = 16'h1;
  wire [15:0]       writeQueueVec_1_enq_bits_targetLane = 16'h2;
  wire [15:0]       writeQueueVec_2_enq_bits_targetLane = 16'h4;
  wire [15:0]       writeQueueVec_3_enq_bits_targetLane = 16'h8;
  wire [15:0]       writeQueueVec_4_enq_bits_targetLane = 16'h10;
  wire [15:0]       writeQueueVec_5_enq_bits_targetLane = 16'h20;
  wire [15:0]       writeQueueVec_6_enq_bits_targetLane = 16'h40;
  wire [15:0]       writeQueueVec_7_enq_bits_targetLane = 16'h80;
  wire [15:0]       writeQueueVec_8_enq_bits_targetLane = 16'h100;
  wire [15:0]       writeQueueVec_9_enq_bits_targetLane = 16'h200;
  wire [15:0]       writeQueueVec_10_enq_bits_targetLane = 16'h400;
  wire [15:0]       writeQueueVec_11_enq_bits_targetLane = 16'h800;
  wire [15:0]       writeQueueVec_12_enq_bits_targetLane = 16'h1000;
  wire [15:0]       writeQueueVec_13_enq_bits_targetLane = 16'h2000;
  wire [15:0]       writeQueueVec_14_enq_bits_targetLane = 16'h4000;
  wire [15:0]       writeQueueVec_15_enq_bits_targetLane = 16'h8000;
  wire [7:0]        axi4Port_aw_bits_len = 8'h0;
  wire [7:0]        axi4Port_ar_bits_len = 8'h0;
  wire [7:0]        simpleAccessPorts_aw_bits_len = 8'h0;
  wire [7:0]        simpleAccessPorts_ar_bits_len = 8'h0;
  wire [2:0]        axi4Port_aw_bits_size = 3'h6;
  wire [2:0]        axi4Port_ar_bits_size = 3'h6;
  wire [1:0]        axi4Port_aw_bits_burst = 2'h1;
  wire [1:0]        axi4Port_ar_bits_burst = 2'h1;
  wire [1:0]        simpleAccessPorts_aw_bits_burst = 2'h1;
  wire [1:0]        simpleAccessPorts_ar_bits_burst = 2'h1;
  wire              axi4Port_aw_bits_lock = 1'h0;
  wire              axi4Port_ar_bits_lock = 1'h0;
  wire              simpleAccessPorts_aw_bits_lock = 1'h0;
  wire              simpleAccessPorts_ar_bits_lock = 1'h0;
  wire [2:0]        axi4Port_aw_bits_prot = 3'h0;
  wire [2:0]        axi4Port_ar_bits_prot = 3'h0;
  wire [2:0]        simpleAccessPorts_aw_bits_prot = 3'h0;
  wire [2:0]        simpleAccessPorts_ar_bits_prot = 3'h0;
  wire              axi4Port_w_bits_last = 1'h1;
  wire              axi4Port_b_ready = 1'h1;
  wire              simpleAccessPorts_w_bits_last = 1'h1;
  wire              simpleAccessPorts_b_ready = 1'h1;
  wire [1:0]        axi4Port_ar_bits_id = 2'h0;
  wire [1:0]        simpleAccessPorts_ar_bits_id = 2'h0;
  wire [2:0]        simpleAccessPorts_ar_bits_size = 3'h2;
  wire [1:0]        vrfReadDataPorts_0_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_1_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_2_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_3_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_4_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_5_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_6_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_7_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_8_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_9_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_10_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_11_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_12_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_13_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_14_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_15_bits_readSource = 2'h2;
  wire              dataQueue_deq_ready = axi4Port_w_ready_0;
  wire              dataQueue_deq_valid;
  wire [511:0]      dataQueue_deq_bits_data;
  wire [63:0]       dataQueue_deq_bits_mask;
  wire              simpleDataQueue_deq_ready = simpleAccessPorts_w_ready_0;
  wire              simpleDataQueue_deq_valid;
  wire [31:0]       simpleDataQueue_deq_bits_data;
  wire [3:0]        simpleDataQueue_deq_bits_mask;
  wire              writeQueueVec_0_deq_ready = vrfWritePort_0_ready_0;
  wire              writeQueueVec_0_deq_valid;
  wire [4:0]        writeQueueVec_0_deq_bits_data_vd;
  wire [1:0]        writeQueueVec_0_deq_bits_data_offset;
  wire [3:0]        writeQueueVec_0_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_0_deq_bits_data_data;
  wire              writeQueueVec_0_deq_bits_data_last;
  wire [2:0]        writeQueueVec_0_deq_bits_data_instructionIndex;
  wire              writeQueueVec_1_deq_ready = vrfWritePort_1_ready_0;
  wire              writeQueueVec_1_deq_valid;
  wire [4:0]        writeQueueVec_1_deq_bits_data_vd;
  wire [1:0]        writeQueueVec_1_deq_bits_data_offset;
  wire [3:0]        writeQueueVec_1_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_1_deq_bits_data_data;
  wire              writeQueueVec_1_deq_bits_data_last;
  wire [2:0]        writeQueueVec_1_deq_bits_data_instructionIndex;
  wire              writeQueueVec_2_deq_ready = vrfWritePort_2_ready_0;
  wire              writeQueueVec_2_deq_valid;
  wire [4:0]        writeQueueVec_2_deq_bits_data_vd;
  wire [1:0]        writeQueueVec_2_deq_bits_data_offset;
  wire [3:0]        writeQueueVec_2_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_2_deq_bits_data_data;
  wire              writeQueueVec_2_deq_bits_data_last;
  wire [2:0]        writeQueueVec_2_deq_bits_data_instructionIndex;
  wire              writeQueueVec_3_deq_ready = vrfWritePort_3_ready_0;
  wire              writeQueueVec_3_deq_valid;
  wire [4:0]        writeQueueVec_3_deq_bits_data_vd;
  wire [1:0]        writeQueueVec_3_deq_bits_data_offset;
  wire [3:0]        writeQueueVec_3_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_3_deq_bits_data_data;
  wire              writeQueueVec_3_deq_bits_data_last;
  wire [2:0]        writeQueueVec_3_deq_bits_data_instructionIndex;
  wire              writeQueueVec_4_deq_ready = vrfWritePort_4_ready_0;
  wire              writeQueueVec_4_deq_valid;
  wire [4:0]        writeQueueVec_4_deq_bits_data_vd;
  wire [1:0]        writeQueueVec_4_deq_bits_data_offset;
  wire [3:0]        writeQueueVec_4_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_4_deq_bits_data_data;
  wire              writeQueueVec_4_deq_bits_data_last;
  wire [2:0]        writeQueueVec_4_deq_bits_data_instructionIndex;
  wire              writeQueueVec_5_deq_ready = vrfWritePort_5_ready_0;
  wire              writeQueueVec_5_deq_valid;
  wire [4:0]        writeQueueVec_5_deq_bits_data_vd;
  wire [1:0]        writeQueueVec_5_deq_bits_data_offset;
  wire [3:0]        writeQueueVec_5_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_5_deq_bits_data_data;
  wire              writeQueueVec_5_deq_bits_data_last;
  wire [2:0]        writeQueueVec_5_deq_bits_data_instructionIndex;
  wire              writeQueueVec_6_deq_ready = vrfWritePort_6_ready_0;
  wire              writeQueueVec_6_deq_valid;
  wire [4:0]        writeQueueVec_6_deq_bits_data_vd;
  wire [1:0]        writeQueueVec_6_deq_bits_data_offset;
  wire [3:0]        writeQueueVec_6_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_6_deq_bits_data_data;
  wire              writeQueueVec_6_deq_bits_data_last;
  wire [2:0]        writeQueueVec_6_deq_bits_data_instructionIndex;
  wire              writeQueueVec_7_deq_ready = vrfWritePort_7_ready_0;
  wire              writeQueueVec_7_deq_valid;
  wire [4:0]        writeQueueVec_7_deq_bits_data_vd;
  wire [1:0]        writeQueueVec_7_deq_bits_data_offset;
  wire [3:0]        writeQueueVec_7_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_7_deq_bits_data_data;
  wire              writeQueueVec_7_deq_bits_data_last;
  wire [2:0]        writeQueueVec_7_deq_bits_data_instructionIndex;
  wire              writeQueueVec_8_deq_ready = vrfWritePort_8_ready_0;
  wire              writeQueueVec_8_deq_valid;
  wire [4:0]        writeQueueVec_8_deq_bits_data_vd;
  wire [1:0]        writeQueueVec_8_deq_bits_data_offset;
  wire [3:0]        writeQueueVec_8_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_8_deq_bits_data_data;
  wire              writeQueueVec_8_deq_bits_data_last;
  wire [2:0]        writeQueueVec_8_deq_bits_data_instructionIndex;
  wire              writeQueueVec_9_deq_ready = vrfWritePort_9_ready_0;
  wire              writeQueueVec_9_deq_valid;
  wire [4:0]        writeQueueVec_9_deq_bits_data_vd;
  wire [1:0]        writeQueueVec_9_deq_bits_data_offset;
  wire [3:0]        writeQueueVec_9_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_9_deq_bits_data_data;
  wire              writeQueueVec_9_deq_bits_data_last;
  wire [2:0]        writeQueueVec_9_deq_bits_data_instructionIndex;
  wire              writeQueueVec_10_deq_ready = vrfWritePort_10_ready_0;
  wire              writeQueueVec_10_deq_valid;
  wire [4:0]        writeQueueVec_10_deq_bits_data_vd;
  wire [1:0]        writeQueueVec_10_deq_bits_data_offset;
  wire [3:0]        writeQueueVec_10_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_10_deq_bits_data_data;
  wire              writeQueueVec_10_deq_bits_data_last;
  wire [2:0]        writeQueueVec_10_deq_bits_data_instructionIndex;
  wire              writeQueueVec_11_deq_ready = vrfWritePort_11_ready_0;
  wire              writeQueueVec_11_deq_valid;
  wire [4:0]        writeQueueVec_11_deq_bits_data_vd;
  wire [1:0]        writeQueueVec_11_deq_bits_data_offset;
  wire [3:0]        writeQueueVec_11_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_11_deq_bits_data_data;
  wire              writeQueueVec_11_deq_bits_data_last;
  wire [2:0]        writeQueueVec_11_deq_bits_data_instructionIndex;
  wire              writeQueueVec_12_deq_ready = vrfWritePort_12_ready_0;
  wire              writeQueueVec_12_deq_valid;
  wire [4:0]        writeQueueVec_12_deq_bits_data_vd;
  wire [1:0]        writeQueueVec_12_deq_bits_data_offset;
  wire [3:0]        writeQueueVec_12_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_12_deq_bits_data_data;
  wire              writeQueueVec_12_deq_bits_data_last;
  wire [2:0]        writeQueueVec_12_deq_bits_data_instructionIndex;
  wire              writeQueueVec_13_deq_ready = vrfWritePort_13_ready_0;
  wire              writeQueueVec_13_deq_valid;
  wire [4:0]        writeQueueVec_13_deq_bits_data_vd;
  wire [1:0]        writeQueueVec_13_deq_bits_data_offset;
  wire [3:0]        writeQueueVec_13_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_13_deq_bits_data_data;
  wire              writeQueueVec_13_deq_bits_data_last;
  wire [2:0]        writeQueueVec_13_deq_bits_data_instructionIndex;
  wire              writeQueueVec_14_deq_ready = vrfWritePort_14_ready_0;
  wire              writeQueueVec_14_deq_valid;
  wire [4:0]        writeQueueVec_14_deq_bits_data_vd;
  wire [1:0]        writeQueueVec_14_deq_bits_data_offset;
  wire [3:0]        writeQueueVec_14_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_14_deq_bits_data_data;
  wire              writeQueueVec_14_deq_bits_data_last;
  wire [2:0]        writeQueueVec_14_deq_bits_data_instructionIndex;
  wire              writeQueueVec_15_deq_ready = vrfWritePort_15_ready_0;
  wire              writeQueueVec_15_deq_valid;
  wire [4:0]        writeQueueVec_15_deq_bits_data_vd;
  wire [1:0]        writeQueueVec_15_deq_bits_data_offset;
  wire [3:0]        writeQueueVec_15_deq_bits_data_mask;
  wire [31:0]       writeQueueVec_15_deq_bits_data_data;
  wire              writeQueueVec_15_deq_bits_data_last;
  wire [2:0]        writeQueueVec_15_deq_bits_data_instructionIndex;
  reg  [31:0]       v0_0;
  reg  [31:0]       v0_1;
  reg  [31:0]       v0_2;
  reg  [31:0]       v0_3;
  reg  [31:0]       v0_4;
  reg  [31:0]       v0_5;
  reg  [31:0]       v0_6;
  reg  [31:0]       v0_7;
  reg  [31:0]       v0_8;
  reg  [31:0]       v0_9;
  reg  [31:0]       v0_10;
  reg  [31:0]       v0_11;
  reg  [31:0]       v0_12;
  reg  [31:0]       v0_13;
  reg  [31:0]       v0_14;
  reg  [31:0]       v0_15;
  reg  [31:0]       v0_16;
  reg  [31:0]       v0_17;
  reg  [31:0]       v0_18;
  reg  [31:0]       v0_19;
  reg  [31:0]       v0_20;
  reg  [31:0]       v0_21;
  reg  [31:0]       v0_22;
  reg  [31:0]       v0_23;
  reg  [31:0]       v0_24;
  reg  [31:0]       v0_25;
  reg  [31:0]       v0_26;
  reg  [31:0]       v0_27;
  reg  [31:0]       v0_28;
  reg  [31:0]       v0_29;
  reg  [31:0]       v0_30;
  reg  [31:0]       v0_31;
  reg  [31:0]       v0_32;
  reg  [31:0]       v0_33;
  reg  [31:0]       v0_34;
  reg  [31:0]       v0_35;
  reg  [31:0]       v0_36;
  reg  [31:0]       v0_37;
  reg  [31:0]       v0_38;
  reg  [31:0]       v0_39;
  reg  [31:0]       v0_40;
  reg  [31:0]       v0_41;
  reg  [31:0]       v0_42;
  reg  [31:0]       v0_43;
  reg  [31:0]       v0_44;
  reg  [31:0]       v0_45;
  reg  [31:0]       v0_46;
  reg  [31:0]       v0_47;
  reg  [31:0]       v0_48;
  reg  [31:0]       v0_49;
  reg  [31:0]       v0_50;
  reg  [31:0]       v0_51;
  reg  [31:0]       v0_52;
  reg  [31:0]       v0_53;
  reg  [31:0]       v0_54;
  reg  [31:0]       v0_55;
  reg  [31:0]       v0_56;
  reg  [31:0]       v0_57;
  reg  [31:0]       v0_58;
  reg  [31:0]       v0_59;
  reg  [31:0]       v0_60;
  reg  [31:0]       v0_61;
  reg  [31:0]       v0_62;
  reg  [31:0]       v0_63;
  wire [15:0]       maskExt_lo = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]       maskExt_hi = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]       maskExt = {maskExt_hi, maskExt_lo};
  wire [15:0]       maskExt_lo_1 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_1 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]       maskExt_1 = {maskExt_hi_1, maskExt_lo_1};
  wire [15:0]       maskExt_lo_2 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_2 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]       maskExt_2 = {maskExt_hi_2, maskExt_lo_2};
  wire [15:0]       maskExt_lo_3 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_3 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]       maskExt_3 = {maskExt_hi_3, maskExt_lo_3};
  wire [15:0]       maskExt_lo_4 = {{8{v0UpdateVec_4_bits_mask[1]}}, {8{v0UpdateVec_4_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_4 = {{8{v0UpdateVec_4_bits_mask[3]}}, {8{v0UpdateVec_4_bits_mask[2]}}};
  wire [31:0]       maskExt_4 = {maskExt_hi_4, maskExt_lo_4};
  wire [15:0]       maskExt_lo_5 = {{8{v0UpdateVec_5_bits_mask[1]}}, {8{v0UpdateVec_5_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_5 = {{8{v0UpdateVec_5_bits_mask[3]}}, {8{v0UpdateVec_5_bits_mask[2]}}};
  wire [31:0]       maskExt_5 = {maskExt_hi_5, maskExt_lo_5};
  wire [15:0]       maskExt_lo_6 = {{8{v0UpdateVec_6_bits_mask[1]}}, {8{v0UpdateVec_6_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_6 = {{8{v0UpdateVec_6_bits_mask[3]}}, {8{v0UpdateVec_6_bits_mask[2]}}};
  wire [31:0]       maskExt_6 = {maskExt_hi_6, maskExt_lo_6};
  wire [15:0]       maskExt_lo_7 = {{8{v0UpdateVec_7_bits_mask[1]}}, {8{v0UpdateVec_7_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_7 = {{8{v0UpdateVec_7_bits_mask[3]}}, {8{v0UpdateVec_7_bits_mask[2]}}};
  wire [31:0]       maskExt_7 = {maskExt_hi_7, maskExt_lo_7};
  wire [15:0]       maskExt_lo_8 = {{8{v0UpdateVec_8_bits_mask[1]}}, {8{v0UpdateVec_8_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_8 = {{8{v0UpdateVec_8_bits_mask[3]}}, {8{v0UpdateVec_8_bits_mask[2]}}};
  wire [31:0]       maskExt_8 = {maskExt_hi_8, maskExt_lo_8};
  wire [15:0]       maskExt_lo_9 = {{8{v0UpdateVec_9_bits_mask[1]}}, {8{v0UpdateVec_9_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_9 = {{8{v0UpdateVec_9_bits_mask[3]}}, {8{v0UpdateVec_9_bits_mask[2]}}};
  wire [31:0]       maskExt_9 = {maskExt_hi_9, maskExt_lo_9};
  wire [15:0]       maskExt_lo_10 = {{8{v0UpdateVec_10_bits_mask[1]}}, {8{v0UpdateVec_10_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_10 = {{8{v0UpdateVec_10_bits_mask[3]}}, {8{v0UpdateVec_10_bits_mask[2]}}};
  wire [31:0]       maskExt_10 = {maskExt_hi_10, maskExt_lo_10};
  wire [15:0]       maskExt_lo_11 = {{8{v0UpdateVec_11_bits_mask[1]}}, {8{v0UpdateVec_11_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_11 = {{8{v0UpdateVec_11_bits_mask[3]}}, {8{v0UpdateVec_11_bits_mask[2]}}};
  wire [31:0]       maskExt_11 = {maskExt_hi_11, maskExt_lo_11};
  wire [15:0]       maskExt_lo_12 = {{8{v0UpdateVec_12_bits_mask[1]}}, {8{v0UpdateVec_12_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_12 = {{8{v0UpdateVec_12_bits_mask[3]}}, {8{v0UpdateVec_12_bits_mask[2]}}};
  wire [31:0]       maskExt_12 = {maskExt_hi_12, maskExt_lo_12};
  wire [15:0]       maskExt_lo_13 = {{8{v0UpdateVec_13_bits_mask[1]}}, {8{v0UpdateVec_13_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_13 = {{8{v0UpdateVec_13_bits_mask[3]}}, {8{v0UpdateVec_13_bits_mask[2]}}};
  wire [31:0]       maskExt_13 = {maskExt_hi_13, maskExt_lo_13};
  wire [15:0]       maskExt_lo_14 = {{8{v0UpdateVec_14_bits_mask[1]}}, {8{v0UpdateVec_14_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_14 = {{8{v0UpdateVec_14_bits_mask[3]}}, {8{v0UpdateVec_14_bits_mask[2]}}};
  wire [31:0]       maskExt_14 = {maskExt_hi_14, maskExt_lo_14};
  wire [15:0]       maskExt_lo_15 = {{8{v0UpdateVec_15_bits_mask[1]}}, {8{v0UpdateVec_15_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_15 = {{8{v0UpdateVec_15_bits_mask[3]}}, {8{v0UpdateVec_15_bits_mask[2]}}};
  wire [31:0]       maskExt_15 = {maskExt_hi_15, maskExt_lo_15};
  wire [15:0]       maskExt_lo_16 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_16 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]       maskExt_16 = {maskExt_hi_16, maskExt_lo_16};
  wire [15:0]       maskExt_lo_17 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_17 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]       maskExt_17 = {maskExt_hi_17, maskExt_lo_17};
  wire [15:0]       maskExt_lo_18 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_18 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]       maskExt_18 = {maskExt_hi_18, maskExt_lo_18};
  wire [15:0]       maskExt_lo_19 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_19 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]       maskExt_19 = {maskExt_hi_19, maskExt_lo_19};
  wire [15:0]       maskExt_lo_20 = {{8{v0UpdateVec_4_bits_mask[1]}}, {8{v0UpdateVec_4_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_20 = {{8{v0UpdateVec_4_bits_mask[3]}}, {8{v0UpdateVec_4_bits_mask[2]}}};
  wire [31:0]       maskExt_20 = {maskExt_hi_20, maskExt_lo_20};
  wire [15:0]       maskExt_lo_21 = {{8{v0UpdateVec_5_bits_mask[1]}}, {8{v0UpdateVec_5_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_21 = {{8{v0UpdateVec_5_bits_mask[3]}}, {8{v0UpdateVec_5_bits_mask[2]}}};
  wire [31:0]       maskExt_21 = {maskExt_hi_21, maskExt_lo_21};
  wire [15:0]       maskExt_lo_22 = {{8{v0UpdateVec_6_bits_mask[1]}}, {8{v0UpdateVec_6_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_22 = {{8{v0UpdateVec_6_bits_mask[3]}}, {8{v0UpdateVec_6_bits_mask[2]}}};
  wire [31:0]       maskExt_22 = {maskExt_hi_22, maskExt_lo_22};
  wire [15:0]       maskExt_lo_23 = {{8{v0UpdateVec_7_bits_mask[1]}}, {8{v0UpdateVec_7_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_23 = {{8{v0UpdateVec_7_bits_mask[3]}}, {8{v0UpdateVec_7_bits_mask[2]}}};
  wire [31:0]       maskExt_23 = {maskExt_hi_23, maskExt_lo_23};
  wire [15:0]       maskExt_lo_24 = {{8{v0UpdateVec_8_bits_mask[1]}}, {8{v0UpdateVec_8_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_24 = {{8{v0UpdateVec_8_bits_mask[3]}}, {8{v0UpdateVec_8_bits_mask[2]}}};
  wire [31:0]       maskExt_24 = {maskExt_hi_24, maskExt_lo_24};
  wire [15:0]       maskExt_lo_25 = {{8{v0UpdateVec_9_bits_mask[1]}}, {8{v0UpdateVec_9_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_25 = {{8{v0UpdateVec_9_bits_mask[3]}}, {8{v0UpdateVec_9_bits_mask[2]}}};
  wire [31:0]       maskExt_25 = {maskExt_hi_25, maskExt_lo_25};
  wire [15:0]       maskExt_lo_26 = {{8{v0UpdateVec_10_bits_mask[1]}}, {8{v0UpdateVec_10_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_26 = {{8{v0UpdateVec_10_bits_mask[3]}}, {8{v0UpdateVec_10_bits_mask[2]}}};
  wire [31:0]       maskExt_26 = {maskExt_hi_26, maskExt_lo_26};
  wire [15:0]       maskExt_lo_27 = {{8{v0UpdateVec_11_bits_mask[1]}}, {8{v0UpdateVec_11_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_27 = {{8{v0UpdateVec_11_bits_mask[3]}}, {8{v0UpdateVec_11_bits_mask[2]}}};
  wire [31:0]       maskExt_27 = {maskExt_hi_27, maskExt_lo_27};
  wire [15:0]       maskExt_lo_28 = {{8{v0UpdateVec_12_bits_mask[1]}}, {8{v0UpdateVec_12_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_28 = {{8{v0UpdateVec_12_bits_mask[3]}}, {8{v0UpdateVec_12_bits_mask[2]}}};
  wire [31:0]       maskExt_28 = {maskExt_hi_28, maskExt_lo_28};
  wire [15:0]       maskExt_lo_29 = {{8{v0UpdateVec_13_bits_mask[1]}}, {8{v0UpdateVec_13_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_29 = {{8{v0UpdateVec_13_bits_mask[3]}}, {8{v0UpdateVec_13_bits_mask[2]}}};
  wire [31:0]       maskExt_29 = {maskExt_hi_29, maskExt_lo_29};
  wire [15:0]       maskExt_lo_30 = {{8{v0UpdateVec_14_bits_mask[1]}}, {8{v0UpdateVec_14_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_30 = {{8{v0UpdateVec_14_bits_mask[3]}}, {8{v0UpdateVec_14_bits_mask[2]}}};
  wire [31:0]       maskExt_30 = {maskExt_hi_30, maskExt_lo_30};
  wire [15:0]       maskExt_lo_31 = {{8{v0UpdateVec_15_bits_mask[1]}}, {8{v0UpdateVec_15_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_31 = {{8{v0UpdateVec_15_bits_mask[3]}}, {8{v0UpdateVec_15_bits_mask[2]}}};
  wire [31:0]       maskExt_31 = {maskExt_hi_31, maskExt_lo_31};
  wire [15:0]       maskExt_lo_32 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_32 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]       maskExt_32 = {maskExt_hi_32, maskExt_lo_32};
  wire [15:0]       maskExt_lo_33 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_33 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]       maskExt_33 = {maskExt_hi_33, maskExt_lo_33};
  wire [15:0]       maskExt_lo_34 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_34 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]       maskExt_34 = {maskExt_hi_34, maskExt_lo_34};
  wire [15:0]       maskExt_lo_35 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_35 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]       maskExt_35 = {maskExt_hi_35, maskExt_lo_35};
  wire [15:0]       maskExt_lo_36 = {{8{v0UpdateVec_4_bits_mask[1]}}, {8{v0UpdateVec_4_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_36 = {{8{v0UpdateVec_4_bits_mask[3]}}, {8{v0UpdateVec_4_bits_mask[2]}}};
  wire [31:0]       maskExt_36 = {maskExt_hi_36, maskExt_lo_36};
  wire [15:0]       maskExt_lo_37 = {{8{v0UpdateVec_5_bits_mask[1]}}, {8{v0UpdateVec_5_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_37 = {{8{v0UpdateVec_5_bits_mask[3]}}, {8{v0UpdateVec_5_bits_mask[2]}}};
  wire [31:0]       maskExt_37 = {maskExt_hi_37, maskExt_lo_37};
  wire [15:0]       maskExt_lo_38 = {{8{v0UpdateVec_6_bits_mask[1]}}, {8{v0UpdateVec_6_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_38 = {{8{v0UpdateVec_6_bits_mask[3]}}, {8{v0UpdateVec_6_bits_mask[2]}}};
  wire [31:0]       maskExt_38 = {maskExt_hi_38, maskExt_lo_38};
  wire [15:0]       maskExt_lo_39 = {{8{v0UpdateVec_7_bits_mask[1]}}, {8{v0UpdateVec_7_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_39 = {{8{v0UpdateVec_7_bits_mask[3]}}, {8{v0UpdateVec_7_bits_mask[2]}}};
  wire [31:0]       maskExt_39 = {maskExt_hi_39, maskExt_lo_39};
  wire [15:0]       maskExt_lo_40 = {{8{v0UpdateVec_8_bits_mask[1]}}, {8{v0UpdateVec_8_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_40 = {{8{v0UpdateVec_8_bits_mask[3]}}, {8{v0UpdateVec_8_bits_mask[2]}}};
  wire [31:0]       maskExt_40 = {maskExt_hi_40, maskExt_lo_40};
  wire [15:0]       maskExt_lo_41 = {{8{v0UpdateVec_9_bits_mask[1]}}, {8{v0UpdateVec_9_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_41 = {{8{v0UpdateVec_9_bits_mask[3]}}, {8{v0UpdateVec_9_bits_mask[2]}}};
  wire [31:0]       maskExt_41 = {maskExt_hi_41, maskExt_lo_41};
  wire [15:0]       maskExt_lo_42 = {{8{v0UpdateVec_10_bits_mask[1]}}, {8{v0UpdateVec_10_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_42 = {{8{v0UpdateVec_10_bits_mask[3]}}, {8{v0UpdateVec_10_bits_mask[2]}}};
  wire [31:0]       maskExt_42 = {maskExt_hi_42, maskExt_lo_42};
  wire [15:0]       maskExt_lo_43 = {{8{v0UpdateVec_11_bits_mask[1]}}, {8{v0UpdateVec_11_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_43 = {{8{v0UpdateVec_11_bits_mask[3]}}, {8{v0UpdateVec_11_bits_mask[2]}}};
  wire [31:0]       maskExt_43 = {maskExt_hi_43, maskExt_lo_43};
  wire [15:0]       maskExt_lo_44 = {{8{v0UpdateVec_12_bits_mask[1]}}, {8{v0UpdateVec_12_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_44 = {{8{v0UpdateVec_12_bits_mask[3]}}, {8{v0UpdateVec_12_bits_mask[2]}}};
  wire [31:0]       maskExt_44 = {maskExt_hi_44, maskExt_lo_44};
  wire [15:0]       maskExt_lo_45 = {{8{v0UpdateVec_13_bits_mask[1]}}, {8{v0UpdateVec_13_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_45 = {{8{v0UpdateVec_13_bits_mask[3]}}, {8{v0UpdateVec_13_bits_mask[2]}}};
  wire [31:0]       maskExt_45 = {maskExt_hi_45, maskExt_lo_45};
  wire [15:0]       maskExt_lo_46 = {{8{v0UpdateVec_14_bits_mask[1]}}, {8{v0UpdateVec_14_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_46 = {{8{v0UpdateVec_14_bits_mask[3]}}, {8{v0UpdateVec_14_bits_mask[2]}}};
  wire [31:0]       maskExt_46 = {maskExt_hi_46, maskExt_lo_46};
  wire [15:0]       maskExt_lo_47 = {{8{v0UpdateVec_15_bits_mask[1]}}, {8{v0UpdateVec_15_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_47 = {{8{v0UpdateVec_15_bits_mask[3]}}, {8{v0UpdateVec_15_bits_mask[2]}}};
  wire [31:0]       maskExt_47 = {maskExt_hi_47, maskExt_lo_47};
  wire [15:0]       maskExt_lo_48 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_48 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]       maskExt_48 = {maskExt_hi_48, maskExt_lo_48};
  wire [15:0]       maskExt_lo_49 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_49 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]       maskExt_49 = {maskExt_hi_49, maskExt_lo_49};
  wire [15:0]       maskExt_lo_50 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_50 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]       maskExt_50 = {maskExt_hi_50, maskExt_lo_50};
  wire [15:0]       maskExt_lo_51 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_51 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]       maskExt_51 = {maskExt_hi_51, maskExt_lo_51};
  wire [15:0]       maskExt_lo_52 = {{8{v0UpdateVec_4_bits_mask[1]}}, {8{v0UpdateVec_4_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_52 = {{8{v0UpdateVec_4_bits_mask[3]}}, {8{v0UpdateVec_4_bits_mask[2]}}};
  wire [31:0]       maskExt_52 = {maskExt_hi_52, maskExt_lo_52};
  wire [15:0]       maskExt_lo_53 = {{8{v0UpdateVec_5_bits_mask[1]}}, {8{v0UpdateVec_5_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_53 = {{8{v0UpdateVec_5_bits_mask[3]}}, {8{v0UpdateVec_5_bits_mask[2]}}};
  wire [31:0]       maskExt_53 = {maskExt_hi_53, maskExt_lo_53};
  wire [15:0]       maskExt_lo_54 = {{8{v0UpdateVec_6_bits_mask[1]}}, {8{v0UpdateVec_6_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_54 = {{8{v0UpdateVec_6_bits_mask[3]}}, {8{v0UpdateVec_6_bits_mask[2]}}};
  wire [31:0]       maskExt_54 = {maskExt_hi_54, maskExt_lo_54};
  wire [15:0]       maskExt_lo_55 = {{8{v0UpdateVec_7_bits_mask[1]}}, {8{v0UpdateVec_7_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_55 = {{8{v0UpdateVec_7_bits_mask[3]}}, {8{v0UpdateVec_7_bits_mask[2]}}};
  wire [31:0]       maskExt_55 = {maskExt_hi_55, maskExt_lo_55};
  wire [15:0]       maskExt_lo_56 = {{8{v0UpdateVec_8_bits_mask[1]}}, {8{v0UpdateVec_8_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_56 = {{8{v0UpdateVec_8_bits_mask[3]}}, {8{v0UpdateVec_8_bits_mask[2]}}};
  wire [31:0]       maskExt_56 = {maskExt_hi_56, maskExt_lo_56};
  wire [15:0]       maskExt_lo_57 = {{8{v0UpdateVec_9_bits_mask[1]}}, {8{v0UpdateVec_9_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_57 = {{8{v0UpdateVec_9_bits_mask[3]}}, {8{v0UpdateVec_9_bits_mask[2]}}};
  wire [31:0]       maskExt_57 = {maskExt_hi_57, maskExt_lo_57};
  wire [15:0]       maskExt_lo_58 = {{8{v0UpdateVec_10_bits_mask[1]}}, {8{v0UpdateVec_10_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_58 = {{8{v0UpdateVec_10_bits_mask[3]}}, {8{v0UpdateVec_10_bits_mask[2]}}};
  wire [31:0]       maskExt_58 = {maskExt_hi_58, maskExt_lo_58};
  wire [15:0]       maskExt_lo_59 = {{8{v0UpdateVec_11_bits_mask[1]}}, {8{v0UpdateVec_11_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_59 = {{8{v0UpdateVec_11_bits_mask[3]}}, {8{v0UpdateVec_11_bits_mask[2]}}};
  wire [31:0]       maskExt_59 = {maskExt_hi_59, maskExt_lo_59};
  wire [15:0]       maskExt_lo_60 = {{8{v0UpdateVec_12_bits_mask[1]}}, {8{v0UpdateVec_12_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_60 = {{8{v0UpdateVec_12_bits_mask[3]}}, {8{v0UpdateVec_12_bits_mask[2]}}};
  wire [31:0]       maskExt_60 = {maskExt_hi_60, maskExt_lo_60};
  wire [15:0]       maskExt_lo_61 = {{8{v0UpdateVec_13_bits_mask[1]}}, {8{v0UpdateVec_13_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_61 = {{8{v0UpdateVec_13_bits_mask[3]}}, {8{v0UpdateVec_13_bits_mask[2]}}};
  wire [31:0]       maskExt_61 = {maskExt_hi_61, maskExt_lo_61};
  wire [15:0]       maskExt_lo_62 = {{8{v0UpdateVec_14_bits_mask[1]}}, {8{v0UpdateVec_14_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_62 = {{8{v0UpdateVec_14_bits_mask[3]}}, {8{v0UpdateVec_14_bits_mask[2]}}};
  wire [31:0]       maskExt_62 = {maskExt_hi_62, maskExt_lo_62};
  wire [15:0]       maskExt_lo_63 = {{8{v0UpdateVec_15_bits_mask[1]}}, {8{v0UpdateVec_15_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_63 = {{8{v0UpdateVec_15_bits_mask[3]}}, {8{v0UpdateVec_15_bits_mask[2]}}};
  wire [31:0]       maskExt_63 = {maskExt_hi_63, maskExt_lo_63};
  wire              alwaysMerge = {request_bits_instructionInformation_mop_0, request_bits_instructionInformation_lumop_0[2:0], request_bits_instructionInformation_lumop_0[4]} == 6'h0;
  wire              useLoadUnit = alwaysMerge & ~request_bits_instructionInformation_isStore_0;
  wire              useStoreUnit = alwaysMerge & request_bits_instructionInformation_isStore_0;
  wire              useOtherUnit = ~alwaysMerge;
  wire              addressCheck = _otherUnit_status_idle & (~useOtherUnit | _loadUnit_status_idle & _storeUnit_status_idle);
  wire              unitReady = useLoadUnit & _loadUnit_status_idle | useStoreUnit & _storeUnit_status_idle | useOtherUnit & _otherUnit_status_idle;
  wire              request_ready_0 = unitReady & addressCheck;
  wire              requestFire = request_ready_0 & request_valid_0;
  wire              reqEnq_0 = useLoadUnit & requestFire;
  wire              reqEnq_1 = useStoreUnit & requestFire;
  wire              reqEnq_2 = useOtherUnit & requestFire;
  wire [4:0]        maskSelect = _loadUnit_maskSelect_valid ? _loadUnit_maskSelect_bits : 5'h0;
  wire [63:0]       _GEN = {v0_1, v0_0};
  wire [63:0]       loadUnit_maskInput_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]       storeUnit_maskInput_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]       otherUnit_maskInput_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]       _GEN_0 = {v0_3, v0_2};
  wire [63:0]       loadUnit_maskInput_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi = _GEN_0;
  wire [63:0]       storeUnit_maskInput_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi = _GEN_0;
  wire [63:0]       otherUnit_maskInput_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi = _GEN_0;
  wire [127:0]      loadUnit_maskInput_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo};
  wire [63:0]       _GEN_1 = {v0_5, v0_4};
  wire [63:0]       loadUnit_maskInput_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]       storeUnit_maskInput_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]       otherUnit_maskInput_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]       _GEN_2 = {v0_7, v0_6};
  wire [63:0]       loadUnit_maskInput_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi = _GEN_2;
  wire [63:0]       storeUnit_maskInput_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi = _GEN_2;
  wire [63:0]       otherUnit_maskInput_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi = _GEN_2;
  wire [127:0]      loadUnit_maskInput_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo};
  wire [255:0]      loadUnit_maskInput_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo};
  wire [63:0]       _GEN_3 = {v0_9, v0_8};
  wire [63:0]       loadUnit_maskInput_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]       storeUnit_maskInput_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]       otherUnit_maskInput_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]       _GEN_4 = {v0_11, v0_10};
  wire [63:0]       loadUnit_maskInput_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi = _GEN_4;
  wire [63:0]       storeUnit_maskInput_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi = _GEN_4;
  wire [63:0]       otherUnit_maskInput_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi = _GEN_4;
  wire [127:0]      loadUnit_maskInput_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo};
  wire [63:0]       _GEN_5 = {v0_13, v0_12};
  wire [63:0]       loadUnit_maskInput_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]       storeUnit_maskInput_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]       otherUnit_maskInput_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]       _GEN_6 = {v0_15, v0_14};
  wire [63:0]       loadUnit_maskInput_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi = _GEN_6;
  wire [63:0]       storeUnit_maskInput_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi = _GEN_6;
  wire [63:0]       otherUnit_maskInput_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi = _GEN_6;
  wire [127:0]      loadUnit_maskInput_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo};
  wire [255:0]      loadUnit_maskInput_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo};
  wire [511:0]      loadUnit_maskInput_lo_lo = {loadUnit_maskInput_lo_lo_hi, loadUnit_maskInput_lo_lo_lo};
  wire [63:0]       _GEN_7 = {v0_17, v0_16};
  wire [63:0]       loadUnit_maskInput_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]       storeUnit_maskInput_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]       otherUnit_maskInput_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]       _GEN_8 = {v0_19, v0_18};
  wire [63:0]       loadUnit_maskInput_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi = _GEN_8;
  wire [63:0]       storeUnit_maskInput_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi = _GEN_8;
  wire [63:0]       otherUnit_maskInput_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi = _GEN_8;
  wire [127:0]      loadUnit_maskInput_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo};
  wire [63:0]       _GEN_9 = {v0_21, v0_20};
  wire [63:0]       loadUnit_maskInput_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]       storeUnit_maskInput_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]       otherUnit_maskInput_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]       _GEN_10 = {v0_23, v0_22};
  wire [63:0]       loadUnit_maskInput_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi = _GEN_10;
  wire [63:0]       storeUnit_maskInput_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi = _GEN_10;
  wire [63:0]       otherUnit_maskInput_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi = _GEN_10;
  wire [127:0]      loadUnit_maskInput_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo};
  wire [255:0]      loadUnit_maskInput_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo};
  wire [63:0]       _GEN_11 = {v0_25, v0_24};
  wire [63:0]       loadUnit_maskInput_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]       storeUnit_maskInput_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]       otherUnit_maskInput_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]       _GEN_12 = {v0_27, v0_26};
  wire [63:0]       loadUnit_maskInput_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi = _GEN_12;
  wire [63:0]       storeUnit_maskInput_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi = _GEN_12;
  wire [63:0]       otherUnit_maskInput_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi = _GEN_12;
  wire [127:0]      loadUnit_maskInput_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo};
  wire [63:0]       _GEN_13 = {v0_29, v0_28};
  wire [63:0]       loadUnit_maskInput_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]       storeUnit_maskInput_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]       otherUnit_maskInput_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]       _GEN_14 = {v0_31, v0_30};
  wire [63:0]       loadUnit_maskInput_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi = _GEN_14;
  wire [63:0]       storeUnit_maskInput_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi = _GEN_14;
  wire [63:0]       otherUnit_maskInput_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi = _GEN_14;
  wire [127:0]      loadUnit_maskInput_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo};
  wire [255:0]      loadUnit_maskInput_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo};
  wire [511:0]      loadUnit_maskInput_lo_hi = {loadUnit_maskInput_lo_hi_hi, loadUnit_maskInput_lo_hi_lo};
  wire [1023:0]     loadUnit_maskInput_lo = {loadUnit_maskInput_lo_hi, loadUnit_maskInput_lo_lo};
  wire [63:0]       _GEN_15 = {v0_33, v0_32};
  wire [63:0]       loadUnit_maskInput_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]       storeUnit_maskInput_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]       otherUnit_maskInput_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]       _GEN_16 = {v0_35, v0_34};
  wire [63:0]       loadUnit_maskInput_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi = _GEN_16;
  wire [63:0]       storeUnit_maskInput_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi = _GEN_16;
  wire [63:0]       otherUnit_maskInput_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi = _GEN_16;
  wire [127:0]      loadUnit_maskInput_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo};
  wire [63:0]       _GEN_17 = {v0_37, v0_36};
  wire [63:0]       loadUnit_maskInput_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]       storeUnit_maskInput_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]       otherUnit_maskInput_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]       _GEN_18 = {v0_39, v0_38};
  wire [63:0]       loadUnit_maskInput_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi = _GEN_18;
  wire [63:0]       storeUnit_maskInput_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi = _GEN_18;
  wire [63:0]       otherUnit_maskInput_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi = _GEN_18;
  wire [127:0]      loadUnit_maskInput_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo};
  wire [255:0]      loadUnit_maskInput_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo};
  wire [63:0]       _GEN_19 = {v0_41, v0_40};
  wire [63:0]       loadUnit_maskInput_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]       storeUnit_maskInput_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]       otherUnit_maskInput_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]       _GEN_20 = {v0_43, v0_42};
  wire [63:0]       loadUnit_maskInput_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi = _GEN_20;
  wire [63:0]       storeUnit_maskInput_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi = _GEN_20;
  wire [63:0]       otherUnit_maskInput_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi = _GEN_20;
  wire [127:0]      loadUnit_maskInput_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo};
  wire [63:0]       _GEN_21 = {v0_45, v0_44};
  wire [63:0]       loadUnit_maskInput_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]       storeUnit_maskInput_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]       otherUnit_maskInput_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]       _GEN_22 = {v0_47, v0_46};
  wire [63:0]       loadUnit_maskInput_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi = _GEN_22;
  wire [63:0]       storeUnit_maskInput_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi = _GEN_22;
  wire [63:0]       otherUnit_maskInput_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi = _GEN_22;
  wire [127:0]      loadUnit_maskInput_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo};
  wire [255:0]      loadUnit_maskInput_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo};
  wire [511:0]      loadUnit_maskInput_hi_lo = {loadUnit_maskInput_hi_lo_hi, loadUnit_maskInput_hi_lo_lo};
  wire [63:0]       _GEN_23 = {v0_49, v0_48};
  wire [63:0]       loadUnit_maskInput_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]       storeUnit_maskInput_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]       otherUnit_maskInput_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]       _GEN_24 = {v0_51, v0_50};
  wire [63:0]       loadUnit_maskInput_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi = _GEN_24;
  wire [63:0]       storeUnit_maskInput_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi = _GEN_24;
  wire [63:0]       otherUnit_maskInput_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi = _GEN_24;
  wire [127:0]      loadUnit_maskInput_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo};
  wire [63:0]       _GEN_25 = {v0_53, v0_52};
  wire [63:0]       loadUnit_maskInput_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]       storeUnit_maskInput_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]       otherUnit_maskInput_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]       _GEN_26 = {v0_55, v0_54};
  wire [63:0]       loadUnit_maskInput_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi = _GEN_26;
  wire [63:0]       storeUnit_maskInput_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi = _GEN_26;
  wire [63:0]       otherUnit_maskInput_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi = _GEN_26;
  wire [127:0]      loadUnit_maskInput_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo};
  wire [255:0]      loadUnit_maskInput_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo};
  wire [63:0]       _GEN_27 = {v0_57, v0_56};
  wire [63:0]       loadUnit_maskInput_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]       storeUnit_maskInput_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]       otherUnit_maskInput_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]       _GEN_28 = {v0_59, v0_58};
  wire [63:0]       loadUnit_maskInput_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi = _GEN_28;
  wire [63:0]       storeUnit_maskInput_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi = _GEN_28;
  wire [63:0]       otherUnit_maskInput_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi = _GEN_28;
  wire [127:0]      loadUnit_maskInput_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo};
  wire [63:0]       _GEN_29 = {v0_61, v0_60};
  wire [63:0]       loadUnit_maskInput_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]       storeUnit_maskInput_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]       otherUnit_maskInput_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]       _GEN_30 = {v0_63, v0_62};
  wire [63:0]       loadUnit_maskInput_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi = _GEN_30;
  wire [63:0]       storeUnit_maskInput_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi = _GEN_30;
  wire [63:0]       otherUnit_maskInput_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi = _GEN_30;
  wire [127:0]      loadUnit_maskInput_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo};
  wire [255:0]      loadUnit_maskInput_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo};
  wire [511:0]      loadUnit_maskInput_hi_hi = {loadUnit_maskInput_hi_hi_hi, loadUnit_maskInput_hi_hi_lo};
  wire [1023:0]     loadUnit_maskInput_hi = {loadUnit_maskInput_hi_hi, loadUnit_maskInput_hi_lo};
  wire [31:0][63:0] _GEN_31 =
    {{loadUnit_maskInput_hi[1023:960]},
     {loadUnit_maskInput_hi[959:896]},
     {loadUnit_maskInput_hi[895:832]},
     {loadUnit_maskInput_hi[831:768]},
     {loadUnit_maskInput_hi[767:704]},
     {loadUnit_maskInput_hi[703:640]},
     {loadUnit_maskInput_hi[639:576]},
     {loadUnit_maskInput_hi[575:512]},
     {loadUnit_maskInput_hi[511:448]},
     {loadUnit_maskInput_hi[447:384]},
     {loadUnit_maskInput_hi[383:320]},
     {loadUnit_maskInput_hi[319:256]},
     {loadUnit_maskInput_hi[255:192]},
     {loadUnit_maskInput_hi[191:128]},
     {loadUnit_maskInput_hi[127:64]},
     {loadUnit_maskInput_hi[63:0]},
     {loadUnit_maskInput_lo[1023:960]},
     {loadUnit_maskInput_lo[959:896]},
     {loadUnit_maskInput_lo[895:832]},
     {loadUnit_maskInput_lo[831:768]},
     {loadUnit_maskInput_lo[767:704]},
     {loadUnit_maskInput_lo[703:640]},
     {loadUnit_maskInput_lo[639:576]},
     {loadUnit_maskInput_lo[575:512]},
     {loadUnit_maskInput_lo[511:448]},
     {loadUnit_maskInput_lo[447:384]},
     {loadUnit_maskInput_lo[383:320]},
     {loadUnit_maskInput_lo[319:256]},
     {loadUnit_maskInput_lo[255:192]},
     {loadUnit_maskInput_lo[191:128]},
     {loadUnit_maskInput_lo[127:64]},
     {loadUnit_maskInput_lo[63:0]}};
  wire [4:0]        maskSelect_1 = _storeUnit_maskSelect_valid ? _storeUnit_maskSelect_bits : 5'h0;
  wire [127:0]      storeUnit_maskInput_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo};
  wire [127:0]      storeUnit_maskInput_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo};
  wire [255:0]      storeUnit_maskInput_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo};
  wire [127:0]      storeUnit_maskInput_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo};
  wire [127:0]      storeUnit_maskInput_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo};
  wire [255:0]      storeUnit_maskInput_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo};
  wire [511:0]      storeUnit_maskInput_lo_lo = {storeUnit_maskInput_lo_lo_hi, storeUnit_maskInput_lo_lo_lo};
  wire [127:0]      storeUnit_maskInput_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo};
  wire [127:0]      storeUnit_maskInput_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo};
  wire [255:0]      storeUnit_maskInput_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo};
  wire [127:0]      storeUnit_maskInput_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo};
  wire [127:0]      storeUnit_maskInput_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo};
  wire [255:0]      storeUnit_maskInput_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo};
  wire [511:0]      storeUnit_maskInput_lo_hi = {storeUnit_maskInput_lo_hi_hi, storeUnit_maskInput_lo_hi_lo};
  wire [1023:0]     storeUnit_maskInput_lo = {storeUnit_maskInput_lo_hi, storeUnit_maskInput_lo_lo};
  wire [127:0]      storeUnit_maskInput_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo};
  wire [127:0]      storeUnit_maskInput_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo};
  wire [255:0]      storeUnit_maskInput_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo};
  wire [127:0]      storeUnit_maskInput_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo};
  wire [127:0]      storeUnit_maskInput_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo};
  wire [255:0]      storeUnit_maskInput_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo};
  wire [511:0]      storeUnit_maskInput_hi_lo = {storeUnit_maskInput_hi_lo_hi, storeUnit_maskInput_hi_lo_lo};
  wire [127:0]      storeUnit_maskInput_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo};
  wire [127:0]      storeUnit_maskInput_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo};
  wire [255:0]      storeUnit_maskInput_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo};
  wire [127:0]      storeUnit_maskInput_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo};
  wire [127:0]      storeUnit_maskInput_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo};
  wire [255:0]      storeUnit_maskInput_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo};
  wire [511:0]      storeUnit_maskInput_hi_hi = {storeUnit_maskInput_hi_hi_hi, storeUnit_maskInput_hi_hi_lo};
  wire [1023:0]     storeUnit_maskInput_hi = {storeUnit_maskInput_hi_hi, storeUnit_maskInput_hi_lo};
  wire [31:0][63:0] _GEN_32 =
    {{storeUnit_maskInput_hi[1023:960]},
     {storeUnit_maskInput_hi[959:896]},
     {storeUnit_maskInput_hi[895:832]},
     {storeUnit_maskInput_hi[831:768]},
     {storeUnit_maskInput_hi[767:704]},
     {storeUnit_maskInput_hi[703:640]},
     {storeUnit_maskInput_hi[639:576]},
     {storeUnit_maskInput_hi[575:512]},
     {storeUnit_maskInput_hi[511:448]},
     {storeUnit_maskInput_hi[447:384]},
     {storeUnit_maskInput_hi[383:320]},
     {storeUnit_maskInput_hi[319:256]},
     {storeUnit_maskInput_hi[255:192]},
     {storeUnit_maskInput_hi[191:128]},
     {storeUnit_maskInput_hi[127:64]},
     {storeUnit_maskInput_hi[63:0]},
     {storeUnit_maskInput_lo[1023:960]},
     {storeUnit_maskInput_lo[959:896]},
     {storeUnit_maskInput_lo[895:832]},
     {storeUnit_maskInput_lo[831:768]},
     {storeUnit_maskInput_lo[767:704]},
     {storeUnit_maskInput_lo[703:640]},
     {storeUnit_maskInput_lo[639:576]},
     {storeUnit_maskInput_lo[575:512]},
     {storeUnit_maskInput_lo[511:448]},
     {storeUnit_maskInput_lo[447:384]},
     {storeUnit_maskInput_lo[383:320]},
     {storeUnit_maskInput_lo[319:256]},
     {storeUnit_maskInput_lo[255:192]},
     {storeUnit_maskInput_lo[191:128]},
     {storeUnit_maskInput_lo[127:64]},
     {storeUnit_maskInput_lo[63:0]}};
  wire [4:0]        maskSelect_2 = _otherUnit_maskSelect_valid ? _otherUnit_maskSelect_bits : 5'h0;
  wire [127:0]      otherUnit_maskInput_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo};
  wire [127:0]      otherUnit_maskInput_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo};
  wire [255:0]      otherUnit_maskInput_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo};
  wire [127:0]      otherUnit_maskInput_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo};
  wire [127:0]      otherUnit_maskInput_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo};
  wire [255:0]      otherUnit_maskInput_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo};
  wire [511:0]      otherUnit_maskInput_lo_lo = {otherUnit_maskInput_lo_lo_hi, otherUnit_maskInput_lo_lo_lo};
  wire [127:0]      otherUnit_maskInput_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo};
  wire [127:0]      otherUnit_maskInput_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo};
  wire [255:0]      otherUnit_maskInput_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo};
  wire [127:0]      otherUnit_maskInput_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo};
  wire [127:0]      otherUnit_maskInput_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo};
  wire [255:0]      otherUnit_maskInput_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo};
  wire [511:0]      otherUnit_maskInput_lo_hi = {otherUnit_maskInput_lo_hi_hi, otherUnit_maskInput_lo_hi_lo};
  wire [1023:0]     otherUnit_maskInput_lo = {otherUnit_maskInput_lo_hi, otherUnit_maskInput_lo_lo};
  wire [127:0]      otherUnit_maskInput_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo};
  wire [127:0]      otherUnit_maskInput_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo};
  wire [255:0]      otherUnit_maskInput_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo};
  wire [127:0]      otherUnit_maskInput_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo};
  wire [127:0]      otherUnit_maskInput_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo};
  wire [255:0]      otherUnit_maskInput_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo};
  wire [511:0]      otherUnit_maskInput_hi_lo = {otherUnit_maskInput_hi_lo_hi, otherUnit_maskInput_hi_lo_lo};
  wire [127:0]      otherUnit_maskInput_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo};
  wire [127:0]      otherUnit_maskInput_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo};
  wire [255:0]      otherUnit_maskInput_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo};
  wire [127:0]      otherUnit_maskInput_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo};
  wire [127:0]      otherUnit_maskInput_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo};
  wire [255:0]      otherUnit_maskInput_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo};
  wire [511:0]      otherUnit_maskInput_hi_hi = {otherUnit_maskInput_hi_hi_hi, otherUnit_maskInput_hi_hi_lo};
  wire [1023:0]     otherUnit_maskInput_hi = {otherUnit_maskInput_hi_hi, otherUnit_maskInput_hi_lo};
  wire [31:0][63:0] _GEN_33 =
    {{otherUnit_maskInput_hi[1023:960]},
     {otherUnit_maskInput_hi[959:896]},
     {otherUnit_maskInput_hi[895:832]},
     {otherUnit_maskInput_hi[831:768]},
     {otherUnit_maskInput_hi[767:704]},
     {otherUnit_maskInput_hi[703:640]},
     {otherUnit_maskInput_hi[639:576]},
     {otherUnit_maskInput_hi[575:512]},
     {otherUnit_maskInput_hi[511:448]},
     {otherUnit_maskInput_hi[447:384]},
     {otherUnit_maskInput_hi[383:320]},
     {otherUnit_maskInput_hi[319:256]},
     {otherUnit_maskInput_hi[255:192]},
     {otherUnit_maskInput_hi[191:128]},
     {otherUnit_maskInput_hi[127:64]},
     {otherUnit_maskInput_hi[63:0]},
     {otherUnit_maskInput_lo[1023:960]},
     {otherUnit_maskInput_lo[959:896]},
     {otherUnit_maskInput_lo[895:832]},
     {otherUnit_maskInput_lo[831:768]},
     {otherUnit_maskInput_lo[767:704]},
     {otherUnit_maskInput_lo[703:640]},
     {otherUnit_maskInput_lo[639:576]},
     {otherUnit_maskInput_lo[575:512]},
     {otherUnit_maskInput_lo[511:448]},
     {otherUnit_maskInput_lo[447:384]},
     {otherUnit_maskInput_lo[383:320]},
     {otherUnit_maskInput_lo[319:256]},
     {otherUnit_maskInput_lo[255:192]},
     {otherUnit_maskInput_lo[191:128]},
     {otherUnit_maskInput_lo[127:64]},
     {otherUnit_maskInput_lo[63:0]}};
  wire              vrfWritePort_0_valid_0 = writeQueueVec_0_deq_valid;
  wire [4:0]        vrfWritePort_0_bits_vd_0 = writeQueueVec_0_deq_bits_data_vd;
  wire [1:0]        vrfWritePort_0_bits_offset_0 = writeQueueVec_0_deq_bits_data_offset;
  wire [3:0]        vrfWritePort_0_bits_mask_0 = writeQueueVec_0_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_0_bits_data_0 = writeQueueVec_0_deq_bits_data_data;
  wire              vrfWritePort_0_bits_last_0 = writeQueueVec_0_deq_bits_data_last;
  wire [2:0]        vrfWritePort_0_bits_instructionIndex_0 = writeQueueVec_0_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_enq_bits = writeQueueVec_0_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_0_enq_bits_data_data;
  wire              writeQueueVec_0_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi = {writeQueueVec_0_enq_bits_data_data, writeQueueVec_0_enq_bits_data_last};
  wire [2:0]        writeQueueVec_0_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo = {writeQueueVec_dataIn_lo_hi, writeQueueVec_0_enq_bits_data_instructionIndex};
  wire [4:0]        writeQueueVec_0_enq_bits_data_vd;
  wire [1:0]        writeQueueVec_0_enq_bits_data_offset;
  wire [6:0]        writeQueueVec_dataIn_hi_hi = {writeQueueVec_0_enq_bits_data_vd, writeQueueVec_0_enq_bits_data_offset};
  wire [3:0]        writeQueueVec_0_enq_bits_data_mask;
  wire [10:0]       writeQueueVec_dataIn_hi = {writeQueueVec_dataIn_hi_hi, writeQueueVec_0_enq_bits_data_mask};
  wire [62:0]       writeQueueVec_dataIn = {writeQueueVec_dataIn_hi, writeQueueVec_dataIn_lo, 16'h1};
  wire [15:0]       writeQueueVec_dataOut_targetLane = _writeQueueVec_fifo_data_out[15:0];
  wire [2:0]        writeQueueVec_dataOut_data_instructionIndex = _writeQueueVec_fifo_data_out[18:16];
  wire              writeQueueVec_dataOut_data_last = _writeQueueVec_fifo_data_out[19];
  wire [31:0]       writeQueueVec_dataOut_data_data = _writeQueueVec_fifo_data_out[51:20];
  wire [3:0]        writeQueueVec_dataOut_data_mask = _writeQueueVec_fifo_data_out[55:52];
  wire [1:0]        writeQueueVec_dataOut_data_offset = _writeQueueVec_fifo_data_out[57:56];
  wire [4:0]        writeQueueVec_dataOut_data_vd = _writeQueueVec_fifo_data_out[62:58];
  wire              writeQueueVec_0_enq_ready = ~_writeQueueVec_fifo_full;
  wire              writeQueueVec_0_enq_valid;
  wire              _probeWire_slots_0_writeValid_T = writeQueueVec_0_enq_ready & writeQueueVec_0_enq_valid;
  assign writeQueueVec_0_deq_valid = ~_writeQueueVec_fifo_empty | writeQueueVec_0_enq_valid;
  assign writeQueueVec_0_deq_bits_data_vd = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_vd : writeQueueVec_dataOut_data_vd;
  assign writeQueueVec_0_deq_bits_data_offset = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_offset : writeQueueVec_dataOut_data_offset;
  assign writeQueueVec_0_deq_bits_data_mask = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_mask : writeQueueVec_dataOut_data_mask;
  assign writeQueueVec_0_deq_bits_data_data = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_data : writeQueueVec_dataOut_data_data;
  assign writeQueueVec_0_deq_bits_data_last = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_last : writeQueueVec_dataOut_data_last;
  assign writeQueueVec_0_deq_bits_data_instructionIndex = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_instructionIndex : writeQueueVec_dataOut_data_instructionIndex;
  wire [15:0]       writeQueueVec_0_deq_bits_targetLane = _writeQueueVec_fifo_empty ? 16'h1 : writeQueueVec_dataOut_targetLane;
  wire              vrfWritePort_1_valid_0 = writeQueueVec_1_deq_valid;
  wire [4:0]        vrfWritePort_1_bits_vd_0 = writeQueueVec_1_deq_bits_data_vd;
  wire [1:0]        vrfWritePort_1_bits_offset_0 = writeQueueVec_1_deq_bits_data_offset;
  wire [3:0]        vrfWritePort_1_bits_mask_0 = writeQueueVec_1_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_1_bits_data_0 = writeQueueVec_1_deq_bits_data_data;
  wire              vrfWritePort_1_bits_last_0 = writeQueueVec_1_deq_bits_data_last;
  wire [2:0]        vrfWritePort_1_bits_instructionIndex_0 = writeQueueVec_1_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_1_enq_bits = writeQueueVec_1_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_1_enq_bits_data_data;
  wire              writeQueueVec_1_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_1 = {writeQueueVec_1_enq_bits_data_data, writeQueueVec_1_enq_bits_data_last};
  wire [2:0]        writeQueueVec_1_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_1 = {writeQueueVec_dataIn_lo_hi_1, writeQueueVec_1_enq_bits_data_instructionIndex};
  wire [4:0]        writeQueueVec_1_enq_bits_data_vd;
  wire [1:0]        writeQueueVec_1_enq_bits_data_offset;
  wire [6:0]        writeQueueVec_dataIn_hi_hi_1 = {writeQueueVec_1_enq_bits_data_vd, writeQueueVec_1_enq_bits_data_offset};
  wire [3:0]        writeQueueVec_1_enq_bits_data_mask;
  wire [10:0]       writeQueueVec_dataIn_hi_1 = {writeQueueVec_dataIn_hi_hi_1, writeQueueVec_1_enq_bits_data_mask};
  wire [62:0]       writeQueueVec_dataIn_1 = {writeQueueVec_dataIn_hi_1, writeQueueVec_dataIn_lo_1, 16'h2};
  wire [15:0]       writeQueueVec_dataOut_1_targetLane = _writeQueueVec_fifo_1_data_out[15:0];
  wire [2:0]        writeQueueVec_dataOut_1_data_instructionIndex = _writeQueueVec_fifo_1_data_out[18:16];
  wire              writeQueueVec_dataOut_1_data_last = _writeQueueVec_fifo_1_data_out[19];
  wire [31:0]       writeQueueVec_dataOut_1_data_data = _writeQueueVec_fifo_1_data_out[51:20];
  wire [3:0]        writeQueueVec_dataOut_1_data_mask = _writeQueueVec_fifo_1_data_out[55:52];
  wire [1:0]        writeQueueVec_dataOut_1_data_offset = _writeQueueVec_fifo_1_data_out[57:56];
  wire [4:0]        writeQueueVec_dataOut_1_data_vd = _writeQueueVec_fifo_1_data_out[62:58];
  wire              writeQueueVec_1_enq_ready = ~_writeQueueVec_fifo_1_full;
  wire              writeQueueVec_1_enq_valid;
  wire              _probeWire_slots_1_writeValid_T = writeQueueVec_1_enq_ready & writeQueueVec_1_enq_valid;
  assign writeQueueVec_1_deq_valid = ~_writeQueueVec_fifo_1_empty | writeQueueVec_1_enq_valid;
  assign writeQueueVec_1_deq_bits_data_vd = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_vd : writeQueueVec_dataOut_1_data_vd;
  assign writeQueueVec_1_deq_bits_data_offset = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_offset : writeQueueVec_dataOut_1_data_offset;
  assign writeQueueVec_1_deq_bits_data_mask = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_mask : writeQueueVec_dataOut_1_data_mask;
  assign writeQueueVec_1_deq_bits_data_data = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_data : writeQueueVec_dataOut_1_data_data;
  assign writeQueueVec_1_deq_bits_data_last = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_last : writeQueueVec_dataOut_1_data_last;
  assign writeQueueVec_1_deq_bits_data_instructionIndex = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_instructionIndex : writeQueueVec_dataOut_1_data_instructionIndex;
  wire [15:0]       writeQueueVec_1_deq_bits_targetLane = _writeQueueVec_fifo_1_empty ? 16'h2 : writeQueueVec_dataOut_1_targetLane;
  wire              vrfWritePort_2_valid_0 = writeQueueVec_2_deq_valid;
  wire [4:0]        vrfWritePort_2_bits_vd_0 = writeQueueVec_2_deq_bits_data_vd;
  wire [1:0]        vrfWritePort_2_bits_offset_0 = writeQueueVec_2_deq_bits_data_offset;
  wire [3:0]        vrfWritePort_2_bits_mask_0 = writeQueueVec_2_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_2_bits_data_0 = writeQueueVec_2_deq_bits_data_data;
  wire              vrfWritePort_2_bits_last_0 = writeQueueVec_2_deq_bits_data_last;
  wire [2:0]        vrfWritePort_2_bits_instructionIndex_0 = writeQueueVec_2_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_2_enq_bits = writeQueueVec_2_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_2_enq_bits_data_data;
  wire              writeQueueVec_2_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_2 = {writeQueueVec_2_enq_bits_data_data, writeQueueVec_2_enq_bits_data_last};
  wire [2:0]        writeQueueVec_2_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_2 = {writeQueueVec_dataIn_lo_hi_2, writeQueueVec_2_enq_bits_data_instructionIndex};
  wire [4:0]        writeQueueVec_2_enq_bits_data_vd;
  wire [1:0]        writeQueueVec_2_enq_bits_data_offset;
  wire [6:0]        writeQueueVec_dataIn_hi_hi_2 = {writeQueueVec_2_enq_bits_data_vd, writeQueueVec_2_enq_bits_data_offset};
  wire [3:0]        writeQueueVec_2_enq_bits_data_mask;
  wire [10:0]       writeQueueVec_dataIn_hi_2 = {writeQueueVec_dataIn_hi_hi_2, writeQueueVec_2_enq_bits_data_mask};
  wire [62:0]       writeQueueVec_dataIn_2 = {writeQueueVec_dataIn_hi_2, writeQueueVec_dataIn_lo_2, 16'h4};
  wire [15:0]       writeQueueVec_dataOut_2_targetLane = _writeQueueVec_fifo_2_data_out[15:0];
  wire [2:0]        writeQueueVec_dataOut_2_data_instructionIndex = _writeQueueVec_fifo_2_data_out[18:16];
  wire              writeQueueVec_dataOut_2_data_last = _writeQueueVec_fifo_2_data_out[19];
  wire [31:0]       writeQueueVec_dataOut_2_data_data = _writeQueueVec_fifo_2_data_out[51:20];
  wire [3:0]        writeQueueVec_dataOut_2_data_mask = _writeQueueVec_fifo_2_data_out[55:52];
  wire [1:0]        writeQueueVec_dataOut_2_data_offset = _writeQueueVec_fifo_2_data_out[57:56];
  wire [4:0]        writeQueueVec_dataOut_2_data_vd = _writeQueueVec_fifo_2_data_out[62:58];
  wire              writeQueueVec_2_enq_ready = ~_writeQueueVec_fifo_2_full;
  wire              writeQueueVec_2_enq_valid;
  wire              _probeWire_slots_2_writeValid_T = writeQueueVec_2_enq_ready & writeQueueVec_2_enq_valid;
  assign writeQueueVec_2_deq_valid = ~_writeQueueVec_fifo_2_empty | writeQueueVec_2_enq_valid;
  assign writeQueueVec_2_deq_bits_data_vd = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_vd : writeQueueVec_dataOut_2_data_vd;
  assign writeQueueVec_2_deq_bits_data_offset = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_offset : writeQueueVec_dataOut_2_data_offset;
  assign writeQueueVec_2_deq_bits_data_mask = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_mask : writeQueueVec_dataOut_2_data_mask;
  assign writeQueueVec_2_deq_bits_data_data = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_data : writeQueueVec_dataOut_2_data_data;
  assign writeQueueVec_2_deq_bits_data_last = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_last : writeQueueVec_dataOut_2_data_last;
  assign writeQueueVec_2_deq_bits_data_instructionIndex = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_instructionIndex : writeQueueVec_dataOut_2_data_instructionIndex;
  wire [15:0]       writeQueueVec_2_deq_bits_targetLane = _writeQueueVec_fifo_2_empty ? 16'h4 : writeQueueVec_dataOut_2_targetLane;
  wire              vrfWritePort_3_valid_0 = writeQueueVec_3_deq_valid;
  wire [4:0]        vrfWritePort_3_bits_vd_0 = writeQueueVec_3_deq_bits_data_vd;
  wire [1:0]        vrfWritePort_3_bits_offset_0 = writeQueueVec_3_deq_bits_data_offset;
  wire [3:0]        vrfWritePort_3_bits_mask_0 = writeQueueVec_3_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_3_bits_data_0 = writeQueueVec_3_deq_bits_data_data;
  wire              vrfWritePort_3_bits_last_0 = writeQueueVec_3_deq_bits_data_last;
  wire [2:0]        vrfWritePort_3_bits_instructionIndex_0 = writeQueueVec_3_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_3_enq_bits = writeQueueVec_3_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_3_enq_bits_data_data;
  wire              writeQueueVec_3_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_3 = {writeQueueVec_3_enq_bits_data_data, writeQueueVec_3_enq_bits_data_last};
  wire [2:0]        writeQueueVec_3_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_3 = {writeQueueVec_dataIn_lo_hi_3, writeQueueVec_3_enq_bits_data_instructionIndex};
  wire [4:0]        writeQueueVec_3_enq_bits_data_vd;
  wire [1:0]        writeQueueVec_3_enq_bits_data_offset;
  wire [6:0]        writeQueueVec_dataIn_hi_hi_3 = {writeQueueVec_3_enq_bits_data_vd, writeQueueVec_3_enq_bits_data_offset};
  wire [3:0]        writeQueueVec_3_enq_bits_data_mask;
  wire [10:0]       writeQueueVec_dataIn_hi_3 = {writeQueueVec_dataIn_hi_hi_3, writeQueueVec_3_enq_bits_data_mask};
  wire [62:0]       writeQueueVec_dataIn_3 = {writeQueueVec_dataIn_hi_3, writeQueueVec_dataIn_lo_3, 16'h8};
  wire [15:0]       writeQueueVec_dataOut_3_targetLane = _writeQueueVec_fifo_3_data_out[15:0];
  wire [2:0]        writeQueueVec_dataOut_3_data_instructionIndex = _writeQueueVec_fifo_3_data_out[18:16];
  wire              writeQueueVec_dataOut_3_data_last = _writeQueueVec_fifo_3_data_out[19];
  wire [31:0]       writeQueueVec_dataOut_3_data_data = _writeQueueVec_fifo_3_data_out[51:20];
  wire [3:0]        writeQueueVec_dataOut_3_data_mask = _writeQueueVec_fifo_3_data_out[55:52];
  wire [1:0]        writeQueueVec_dataOut_3_data_offset = _writeQueueVec_fifo_3_data_out[57:56];
  wire [4:0]        writeQueueVec_dataOut_3_data_vd = _writeQueueVec_fifo_3_data_out[62:58];
  wire              writeQueueVec_3_enq_ready = ~_writeQueueVec_fifo_3_full;
  wire              writeQueueVec_3_enq_valid;
  wire              _probeWire_slots_3_writeValid_T = writeQueueVec_3_enq_ready & writeQueueVec_3_enq_valid;
  assign writeQueueVec_3_deq_valid = ~_writeQueueVec_fifo_3_empty | writeQueueVec_3_enq_valid;
  assign writeQueueVec_3_deq_bits_data_vd = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_vd : writeQueueVec_dataOut_3_data_vd;
  assign writeQueueVec_3_deq_bits_data_offset = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_offset : writeQueueVec_dataOut_3_data_offset;
  assign writeQueueVec_3_deq_bits_data_mask = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_mask : writeQueueVec_dataOut_3_data_mask;
  assign writeQueueVec_3_deq_bits_data_data = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_data : writeQueueVec_dataOut_3_data_data;
  assign writeQueueVec_3_deq_bits_data_last = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_last : writeQueueVec_dataOut_3_data_last;
  assign writeQueueVec_3_deq_bits_data_instructionIndex = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_instructionIndex : writeQueueVec_dataOut_3_data_instructionIndex;
  wire [15:0]       writeQueueVec_3_deq_bits_targetLane = _writeQueueVec_fifo_3_empty ? 16'h8 : writeQueueVec_dataOut_3_targetLane;
  wire              vrfWritePort_4_valid_0 = writeQueueVec_4_deq_valid;
  wire [4:0]        vrfWritePort_4_bits_vd_0 = writeQueueVec_4_deq_bits_data_vd;
  wire [1:0]        vrfWritePort_4_bits_offset_0 = writeQueueVec_4_deq_bits_data_offset;
  wire [3:0]        vrfWritePort_4_bits_mask_0 = writeQueueVec_4_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_4_bits_data_0 = writeQueueVec_4_deq_bits_data_data;
  wire              vrfWritePort_4_bits_last_0 = writeQueueVec_4_deq_bits_data_last;
  wire [2:0]        vrfWritePort_4_bits_instructionIndex_0 = writeQueueVec_4_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_4_enq_bits = writeQueueVec_4_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_4_enq_bits_data_data;
  wire              writeQueueVec_4_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_4 = {writeQueueVec_4_enq_bits_data_data, writeQueueVec_4_enq_bits_data_last};
  wire [2:0]        writeQueueVec_4_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_4 = {writeQueueVec_dataIn_lo_hi_4, writeQueueVec_4_enq_bits_data_instructionIndex};
  wire [4:0]        writeQueueVec_4_enq_bits_data_vd;
  wire [1:0]        writeQueueVec_4_enq_bits_data_offset;
  wire [6:0]        writeQueueVec_dataIn_hi_hi_4 = {writeQueueVec_4_enq_bits_data_vd, writeQueueVec_4_enq_bits_data_offset};
  wire [3:0]        writeQueueVec_4_enq_bits_data_mask;
  wire [10:0]       writeQueueVec_dataIn_hi_4 = {writeQueueVec_dataIn_hi_hi_4, writeQueueVec_4_enq_bits_data_mask};
  wire [62:0]       writeQueueVec_dataIn_4 = {writeQueueVec_dataIn_hi_4, writeQueueVec_dataIn_lo_4, 16'h10};
  wire [15:0]       writeQueueVec_dataOut_4_targetLane = _writeQueueVec_fifo_4_data_out[15:0];
  wire [2:0]        writeQueueVec_dataOut_4_data_instructionIndex = _writeQueueVec_fifo_4_data_out[18:16];
  wire              writeQueueVec_dataOut_4_data_last = _writeQueueVec_fifo_4_data_out[19];
  wire [31:0]       writeQueueVec_dataOut_4_data_data = _writeQueueVec_fifo_4_data_out[51:20];
  wire [3:0]        writeQueueVec_dataOut_4_data_mask = _writeQueueVec_fifo_4_data_out[55:52];
  wire [1:0]        writeQueueVec_dataOut_4_data_offset = _writeQueueVec_fifo_4_data_out[57:56];
  wire [4:0]        writeQueueVec_dataOut_4_data_vd = _writeQueueVec_fifo_4_data_out[62:58];
  wire              writeQueueVec_4_enq_ready = ~_writeQueueVec_fifo_4_full;
  wire              writeQueueVec_4_enq_valid;
  wire              _probeWire_slots_4_writeValid_T = writeQueueVec_4_enq_ready & writeQueueVec_4_enq_valid;
  assign writeQueueVec_4_deq_valid = ~_writeQueueVec_fifo_4_empty | writeQueueVec_4_enq_valid;
  assign writeQueueVec_4_deq_bits_data_vd = _writeQueueVec_fifo_4_empty ? writeQueueVec_4_enq_bits_data_vd : writeQueueVec_dataOut_4_data_vd;
  assign writeQueueVec_4_deq_bits_data_offset = _writeQueueVec_fifo_4_empty ? writeQueueVec_4_enq_bits_data_offset : writeQueueVec_dataOut_4_data_offset;
  assign writeQueueVec_4_deq_bits_data_mask = _writeQueueVec_fifo_4_empty ? writeQueueVec_4_enq_bits_data_mask : writeQueueVec_dataOut_4_data_mask;
  assign writeQueueVec_4_deq_bits_data_data = _writeQueueVec_fifo_4_empty ? writeQueueVec_4_enq_bits_data_data : writeQueueVec_dataOut_4_data_data;
  assign writeQueueVec_4_deq_bits_data_last = _writeQueueVec_fifo_4_empty ? writeQueueVec_4_enq_bits_data_last : writeQueueVec_dataOut_4_data_last;
  assign writeQueueVec_4_deq_bits_data_instructionIndex = _writeQueueVec_fifo_4_empty ? writeQueueVec_4_enq_bits_data_instructionIndex : writeQueueVec_dataOut_4_data_instructionIndex;
  wire [15:0]       writeQueueVec_4_deq_bits_targetLane = _writeQueueVec_fifo_4_empty ? 16'h10 : writeQueueVec_dataOut_4_targetLane;
  wire              vrfWritePort_5_valid_0 = writeQueueVec_5_deq_valid;
  wire [4:0]        vrfWritePort_5_bits_vd_0 = writeQueueVec_5_deq_bits_data_vd;
  wire [1:0]        vrfWritePort_5_bits_offset_0 = writeQueueVec_5_deq_bits_data_offset;
  wire [3:0]        vrfWritePort_5_bits_mask_0 = writeQueueVec_5_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_5_bits_data_0 = writeQueueVec_5_deq_bits_data_data;
  wire              vrfWritePort_5_bits_last_0 = writeQueueVec_5_deq_bits_data_last;
  wire [2:0]        vrfWritePort_5_bits_instructionIndex_0 = writeQueueVec_5_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_5_enq_bits = writeQueueVec_5_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_5_enq_bits_data_data;
  wire              writeQueueVec_5_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_5 = {writeQueueVec_5_enq_bits_data_data, writeQueueVec_5_enq_bits_data_last};
  wire [2:0]        writeQueueVec_5_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_5 = {writeQueueVec_dataIn_lo_hi_5, writeQueueVec_5_enq_bits_data_instructionIndex};
  wire [4:0]        writeQueueVec_5_enq_bits_data_vd;
  wire [1:0]        writeQueueVec_5_enq_bits_data_offset;
  wire [6:0]        writeQueueVec_dataIn_hi_hi_5 = {writeQueueVec_5_enq_bits_data_vd, writeQueueVec_5_enq_bits_data_offset};
  wire [3:0]        writeQueueVec_5_enq_bits_data_mask;
  wire [10:0]       writeQueueVec_dataIn_hi_5 = {writeQueueVec_dataIn_hi_hi_5, writeQueueVec_5_enq_bits_data_mask};
  wire [62:0]       writeQueueVec_dataIn_5 = {writeQueueVec_dataIn_hi_5, writeQueueVec_dataIn_lo_5, 16'h20};
  wire [15:0]       writeQueueVec_dataOut_5_targetLane = _writeQueueVec_fifo_5_data_out[15:0];
  wire [2:0]        writeQueueVec_dataOut_5_data_instructionIndex = _writeQueueVec_fifo_5_data_out[18:16];
  wire              writeQueueVec_dataOut_5_data_last = _writeQueueVec_fifo_5_data_out[19];
  wire [31:0]       writeQueueVec_dataOut_5_data_data = _writeQueueVec_fifo_5_data_out[51:20];
  wire [3:0]        writeQueueVec_dataOut_5_data_mask = _writeQueueVec_fifo_5_data_out[55:52];
  wire [1:0]        writeQueueVec_dataOut_5_data_offset = _writeQueueVec_fifo_5_data_out[57:56];
  wire [4:0]        writeQueueVec_dataOut_5_data_vd = _writeQueueVec_fifo_5_data_out[62:58];
  wire              writeQueueVec_5_enq_ready = ~_writeQueueVec_fifo_5_full;
  wire              writeQueueVec_5_enq_valid;
  wire              _probeWire_slots_5_writeValid_T = writeQueueVec_5_enq_ready & writeQueueVec_5_enq_valid;
  assign writeQueueVec_5_deq_valid = ~_writeQueueVec_fifo_5_empty | writeQueueVec_5_enq_valid;
  assign writeQueueVec_5_deq_bits_data_vd = _writeQueueVec_fifo_5_empty ? writeQueueVec_5_enq_bits_data_vd : writeQueueVec_dataOut_5_data_vd;
  assign writeQueueVec_5_deq_bits_data_offset = _writeQueueVec_fifo_5_empty ? writeQueueVec_5_enq_bits_data_offset : writeQueueVec_dataOut_5_data_offset;
  assign writeQueueVec_5_deq_bits_data_mask = _writeQueueVec_fifo_5_empty ? writeQueueVec_5_enq_bits_data_mask : writeQueueVec_dataOut_5_data_mask;
  assign writeQueueVec_5_deq_bits_data_data = _writeQueueVec_fifo_5_empty ? writeQueueVec_5_enq_bits_data_data : writeQueueVec_dataOut_5_data_data;
  assign writeQueueVec_5_deq_bits_data_last = _writeQueueVec_fifo_5_empty ? writeQueueVec_5_enq_bits_data_last : writeQueueVec_dataOut_5_data_last;
  assign writeQueueVec_5_deq_bits_data_instructionIndex = _writeQueueVec_fifo_5_empty ? writeQueueVec_5_enq_bits_data_instructionIndex : writeQueueVec_dataOut_5_data_instructionIndex;
  wire [15:0]       writeQueueVec_5_deq_bits_targetLane = _writeQueueVec_fifo_5_empty ? 16'h20 : writeQueueVec_dataOut_5_targetLane;
  wire              vrfWritePort_6_valid_0 = writeQueueVec_6_deq_valid;
  wire [4:0]        vrfWritePort_6_bits_vd_0 = writeQueueVec_6_deq_bits_data_vd;
  wire [1:0]        vrfWritePort_6_bits_offset_0 = writeQueueVec_6_deq_bits_data_offset;
  wire [3:0]        vrfWritePort_6_bits_mask_0 = writeQueueVec_6_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_6_bits_data_0 = writeQueueVec_6_deq_bits_data_data;
  wire              vrfWritePort_6_bits_last_0 = writeQueueVec_6_deq_bits_data_last;
  wire [2:0]        vrfWritePort_6_bits_instructionIndex_0 = writeQueueVec_6_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_6_enq_bits = writeQueueVec_6_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_6_enq_bits_data_data;
  wire              writeQueueVec_6_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_6 = {writeQueueVec_6_enq_bits_data_data, writeQueueVec_6_enq_bits_data_last};
  wire [2:0]        writeQueueVec_6_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_6 = {writeQueueVec_dataIn_lo_hi_6, writeQueueVec_6_enq_bits_data_instructionIndex};
  wire [4:0]        writeQueueVec_6_enq_bits_data_vd;
  wire [1:0]        writeQueueVec_6_enq_bits_data_offset;
  wire [6:0]        writeQueueVec_dataIn_hi_hi_6 = {writeQueueVec_6_enq_bits_data_vd, writeQueueVec_6_enq_bits_data_offset};
  wire [3:0]        writeQueueVec_6_enq_bits_data_mask;
  wire [10:0]       writeQueueVec_dataIn_hi_6 = {writeQueueVec_dataIn_hi_hi_6, writeQueueVec_6_enq_bits_data_mask};
  wire [62:0]       writeQueueVec_dataIn_6 = {writeQueueVec_dataIn_hi_6, writeQueueVec_dataIn_lo_6, 16'h40};
  wire [15:0]       writeQueueVec_dataOut_6_targetLane = _writeQueueVec_fifo_6_data_out[15:0];
  wire [2:0]        writeQueueVec_dataOut_6_data_instructionIndex = _writeQueueVec_fifo_6_data_out[18:16];
  wire              writeQueueVec_dataOut_6_data_last = _writeQueueVec_fifo_6_data_out[19];
  wire [31:0]       writeQueueVec_dataOut_6_data_data = _writeQueueVec_fifo_6_data_out[51:20];
  wire [3:0]        writeQueueVec_dataOut_6_data_mask = _writeQueueVec_fifo_6_data_out[55:52];
  wire [1:0]        writeQueueVec_dataOut_6_data_offset = _writeQueueVec_fifo_6_data_out[57:56];
  wire [4:0]        writeQueueVec_dataOut_6_data_vd = _writeQueueVec_fifo_6_data_out[62:58];
  wire              writeQueueVec_6_enq_ready = ~_writeQueueVec_fifo_6_full;
  wire              writeQueueVec_6_enq_valid;
  wire              _probeWire_slots_6_writeValid_T = writeQueueVec_6_enq_ready & writeQueueVec_6_enq_valid;
  assign writeQueueVec_6_deq_valid = ~_writeQueueVec_fifo_6_empty | writeQueueVec_6_enq_valid;
  assign writeQueueVec_6_deq_bits_data_vd = _writeQueueVec_fifo_6_empty ? writeQueueVec_6_enq_bits_data_vd : writeQueueVec_dataOut_6_data_vd;
  assign writeQueueVec_6_deq_bits_data_offset = _writeQueueVec_fifo_6_empty ? writeQueueVec_6_enq_bits_data_offset : writeQueueVec_dataOut_6_data_offset;
  assign writeQueueVec_6_deq_bits_data_mask = _writeQueueVec_fifo_6_empty ? writeQueueVec_6_enq_bits_data_mask : writeQueueVec_dataOut_6_data_mask;
  assign writeQueueVec_6_deq_bits_data_data = _writeQueueVec_fifo_6_empty ? writeQueueVec_6_enq_bits_data_data : writeQueueVec_dataOut_6_data_data;
  assign writeQueueVec_6_deq_bits_data_last = _writeQueueVec_fifo_6_empty ? writeQueueVec_6_enq_bits_data_last : writeQueueVec_dataOut_6_data_last;
  assign writeQueueVec_6_deq_bits_data_instructionIndex = _writeQueueVec_fifo_6_empty ? writeQueueVec_6_enq_bits_data_instructionIndex : writeQueueVec_dataOut_6_data_instructionIndex;
  wire [15:0]       writeQueueVec_6_deq_bits_targetLane = _writeQueueVec_fifo_6_empty ? 16'h40 : writeQueueVec_dataOut_6_targetLane;
  wire              vrfWritePort_7_valid_0 = writeQueueVec_7_deq_valid;
  wire [4:0]        vrfWritePort_7_bits_vd_0 = writeQueueVec_7_deq_bits_data_vd;
  wire [1:0]        vrfWritePort_7_bits_offset_0 = writeQueueVec_7_deq_bits_data_offset;
  wire [3:0]        vrfWritePort_7_bits_mask_0 = writeQueueVec_7_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_7_bits_data_0 = writeQueueVec_7_deq_bits_data_data;
  wire              vrfWritePort_7_bits_last_0 = writeQueueVec_7_deq_bits_data_last;
  wire [2:0]        vrfWritePort_7_bits_instructionIndex_0 = writeQueueVec_7_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_7_enq_bits = writeQueueVec_7_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_7_enq_bits_data_data;
  wire              writeQueueVec_7_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_7 = {writeQueueVec_7_enq_bits_data_data, writeQueueVec_7_enq_bits_data_last};
  wire [2:0]        writeQueueVec_7_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_7 = {writeQueueVec_dataIn_lo_hi_7, writeQueueVec_7_enq_bits_data_instructionIndex};
  wire [4:0]        writeQueueVec_7_enq_bits_data_vd;
  wire [1:0]        writeQueueVec_7_enq_bits_data_offset;
  wire [6:0]        writeQueueVec_dataIn_hi_hi_7 = {writeQueueVec_7_enq_bits_data_vd, writeQueueVec_7_enq_bits_data_offset};
  wire [3:0]        writeQueueVec_7_enq_bits_data_mask;
  wire [10:0]       writeQueueVec_dataIn_hi_7 = {writeQueueVec_dataIn_hi_hi_7, writeQueueVec_7_enq_bits_data_mask};
  wire [62:0]       writeQueueVec_dataIn_7 = {writeQueueVec_dataIn_hi_7, writeQueueVec_dataIn_lo_7, 16'h80};
  wire [15:0]       writeQueueVec_dataOut_7_targetLane = _writeQueueVec_fifo_7_data_out[15:0];
  wire [2:0]        writeQueueVec_dataOut_7_data_instructionIndex = _writeQueueVec_fifo_7_data_out[18:16];
  wire              writeQueueVec_dataOut_7_data_last = _writeQueueVec_fifo_7_data_out[19];
  wire [31:0]       writeQueueVec_dataOut_7_data_data = _writeQueueVec_fifo_7_data_out[51:20];
  wire [3:0]        writeQueueVec_dataOut_7_data_mask = _writeQueueVec_fifo_7_data_out[55:52];
  wire [1:0]        writeQueueVec_dataOut_7_data_offset = _writeQueueVec_fifo_7_data_out[57:56];
  wire [4:0]        writeQueueVec_dataOut_7_data_vd = _writeQueueVec_fifo_7_data_out[62:58];
  wire              writeQueueVec_7_enq_ready = ~_writeQueueVec_fifo_7_full;
  wire              writeQueueVec_7_enq_valid;
  wire              _probeWire_slots_7_writeValid_T = writeQueueVec_7_enq_ready & writeQueueVec_7_enq_valid;
  assign writeQueueVec_7_deq_valid = ~_writeQueueVec_fifo_7_empty | writeQueueVec_7_enq_valid;
  assign writeQueueVec_7_deq_bits_data_vd = _writeQueueVec_fifo_7_empty ? writeQueueVec_7_enq_bits_data_vd : writeQueueVec_dataOut_7_data_vd;
  assign writeQueueVec_7_deq_bits_data_offset = _writeQueueVec_fifo_7_empty ? writeQueueVec_7_enq_bits_data_offset : writeQueueVec_dataOut_7_data_offset;
  assign writeQueueVec_7_deq_bits_data_mask = _writeQueueVec_fifo_7_empty ? writeQueueVec_7_enq_bits_data_mask : writeQueueVec_dataOut_7_data_mask;
  assign writeQueueVec_7_deq_bits_data_data = _writeQueueVec_fifo_7_empty ? writeQueueVec_7_enq_bits_data_data : writeQueueVec_dataOut_7_data_data;
  assign writeQueueVec_7_deq_bits_data_last = _writeQueueVec_fifo_7_empty ? writeQueueVec_7_enq_bits_data_last : writeQueueVec_dataOut_7_data_last;
  assign writeQueueVec_7_deq_bits_data_instructionIndex = _writeQueueVec_fifo_7_empty ? writeQueueVec_7_enq_bits_data_instructionIndex : writeQueueVec_dataOut_7_data_instructionIndex;
  wire [15:0]       writeQueueVec_7_deq_bits_targetLane = _writeQueueVec_fifo_7_empty ? 16'h80 : writeQueueVec_dataOut_7_targetLane;
  wire              vrfWritePort_8_valid_0 = writeQueueVec_8_deq_valid;
  wire [4:0]        vrfWritePort_8_bits_vd_0 = writeQueueVec_8_deq_bits_data_vd;
  wire [1:0]        vrfWritePort_8_bits_offset_0 = writeQueueVec_8_deq_bits_data_offset;
  wire [3:0]        vrfWritePort_8_bits_mask_0 = writeQueueVec_8_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_8_bits_data_0 = writeQueueVec_8_deq_bits_data_data;
  wire              vrfWritePort_8_bits_last_0 = writeQueueVec_8_deq_bits_data_last;
  wire [2:0]        vrfWritePort_8_bits_instructionIndex_0 = writeQueueVec_8_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_8_enq_bits = writeQueueVec_8_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_8_enq_bits_data_data;
  wire              writeQueueVec_8_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_8 = {writeQueueVec_8_enq_bits_data_data, writeQueueVec_8_enq_bits_data_last};
  wire [2:0]        writeQueueVec_8_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_8 = {writeQueueVec_dataIn_lo_hi_8, writeQueueVec_8_enq_bits_data_instructionIndex};
  wire [4:0]        writeQueueVec_8_enq_bits_data_vd;
  wire [1:0]        writeQueueVec_8_enq_bits_data_offset;
  wire [6:0]        writeQueueVec_dataIn_hi_hi_8 = {writeQueueVec_8_enq_bits_data_vd, writeQueueVec_8_enq_bits_data_offset};
  wire [3:0]        writeQueueVec_8_enq_bits_data_mask;
  wire [10:0]       writeQueueVec_dataIn_hi_8 = {writeQueueVec_dataIn_hi_hi_8, writeQueueVec_8_enq_bits_data_mask};
  wire [62:0]       writeQueueVec_dataIn_8 = {writeQueueVec_dataIn_hi_8, writeQueueVec_dataIn_lo_8, 16'h100};
  wire [15:0]       writeQueueVec_dataOut_8_targetLane = _writeQueueVec_fifo_8_data_out[15:0];
  wire [2:0]        writeQueueVec_dataOut_8_data_instructionIndex = _writeQueueVec_fifo_8_data_out[18:16];
  wire              writeQueueVec_dataOut_8_data_last = _writeQueueVec_fifo_8_data_out[19];
  wire [31:0]       writeQueueVec_dataOut_8_data_data = _writeQueueVec_fifo_8_data_out[51:20];
  wire [3:0]        writeQueueVec_dataOut_8_data_mask = _writeQueueVec_fifo_8_data_out[55:52];
  wire [1:0]        writeQueueVec_dataOut_8_data_offset = _writeQueueVec_fifo_8_data_out[57:56];
  wire [4:0]        writeQueueVec_dataOut_8_data_vd = _writeQueueVec_fifo_8_data_out[62:58];
  wire              writeQueueVec_8_enq_ready = ~_writeQueueVec_fifo_8_full;
  wire              writeQueueVec_8_enq_valid;
  wire              _probeWire_slots_8_writeValid_T = writeQueueVec_8_enq_ready & writeQueueVec_8_enq_valid;
  assign writeQueueVec_8_deq_valid = ~_writeQueueVec_fifo_8_empty | writeQueueVec_8_enq_valid;
  assign writeQueueVec_8_deq_bits_data_vd = _writeQueueVec_fifo_8_empty ? writeQueueVec_8_enq_bits_data_vd : writeQueueVec_dataOut_8_data_vd;
  assign writeQueueVec_8_deq_bits_data_offset = _writeQueueVec_fifo_8_empty ? writeQueueVec_8_enq_bits_data_offset : writeQueueVec_dataOut_8_data_offset;
  assign writeQueueVec_8_deq_bits_data_mask = _writeQueueVec_fifo_8_empty ? writeQueueVec_8_enq_bits_data_mask : writeQueueVec_dataOut_8_data_mask;
  assign writeQueueVec_8_deq_bits_data_data = _writeQueueVec_fifo_8_empty ? writeQueueVec_8_enq_bits_data_data : writeQueueVec_dataOut_8_data_data;
  assign writeQueueVec_8_deq_bits_data_last = _writeQueueVec_fifo_8_empty ? writeQueueVec_8_enq_bits_data_last : writeQueueVec_dataOut_8_data_last;
  assign writeQueueVec_8_deq_bits_data_instructionIndex = _writeQueueVec_fifo_8_empty ? writeQueueVec_8_enq_bits_data_instructionIndex : writeQueueVec_dataOut_8_data_instructionIndex;
  wire [15:0]       writeQueueVec_8_deq_bits_targetLane = _writeQueueVec_fifo_8_empty ? 16'h100 : writeQueueVec_dataOut_8_targetLane;
  wire              vrfWritePort_9_valid_0 = writeQueueVec_9_deq_valid;
  wire [4:0]        vrfWritePort_9_bits_vd_0 = writeQueueVec_9_deq_bits_data_vd;
  wire [1:0]        vrfWritePort_9_bits_offset_0 = writeQueueVec_9_deq_bits_data_offset;
  wire [3:0]        vrfWritePort_9_bits_mask_0 = writeQueueVec_9_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_9_bits_data_0 = writeQueueVec_9_deq_bits_data_data;
  wire              vrfWritePort_9_bits_last_0 = writeQueueVec_9_deq_bits_data_last;
  wire [2:0]        vrfWritePort_9_bits_instructionIndex_0 = writeQueueVec_9_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_9_enq_bits = writeQueueVec_9_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_9_enq_bits_data_data;
  wire              writeQueueVec_9_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_9 = {writeQueueVec_9_enq_bits_data_data, writeQueueVec_9_enq_bits_data_last};
  wire [2:0]        writeQueueVec_9_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_9 = {writeQueueVec_dataIn_lo_hi_9, writeQueueVec_9_enq_bits_data_instructionIndex};
  wire [4:0]        writeQueueVec_9_enq_bits_data_vd;
  wire [1:0]        writeQueueVec_9_enq_bits_data_offset;
  wire [6:0]        writeQueueVec_dataIn_hi_hi_9 = {writeQueueVec_9_enq_bits_data_vd, writeQueueVec_9_enq_bits_data_offset};
  wire [3:0]        writeQueueVec_9_enq_bits_data_mask;
  wire [10:0]       writeQueueVec_dataIn_hi_9 = {writeQueueVec_dataIn_hi_hi_9, writeQueueVec_9_enq_bits_data_mask};
  wire [62:0]       writeQueueVec_dataIn_9 = {writeQueueVec_dataIn_hi_9, writeQueueVec_dataIn_lo_9, 16'h200};
  wire [15:0]       writeQueueVec_dataOut_9_targetLane = _writeQueueVec_fifo_9_data_out[15:0];
  wire [2:0]        writeQueueVec_dataOut_9_data_instructionIndex = _writeQueueVec_fifo_9_data_out[18:16];
  wire              writeQueueVec_dataOut_9_data_last = _writeQueueVec_fifo_9_data_out[19];
  wire [31:0]       writeQueueVec_dataOut_9_data_data = _writeQueueVec_fifo_9_data_out[51:20];
  wire [3:0]        writeQueueVec_dataOut_9_data_mask = _writeQueueVec_fifo_9_data_out[55:52];
  wire [1:0]        writeQueueVec_dataOut_9_data_offset = _writeQueueVec_fifo_9_data_out[57:56];
  wire [4:0]        writeQueueVec_dataOut_9_data_vd = _writeQueueVec_fifo_9_data_out[62:58];
  wire              writeQueueVec_9_enq_ready = ~_writeQueueVec_fifo_9_full;
  wire              writeQueueVec_9_enq_valid;
  wire              _probeWire_slots_9_writeValid_T = writeQueueVec_9_enq_ready & writeQueueVec_9_enq_valid;
  assign writeQueueVec_9_deq_valid = ~_writeQueueVec_fifo_9_empty | writeQueueVec_9_enq_valid;
  assign writeQueueVec_9_deq_bits_data_vd = _writeQueueVec_fifo_9_empty ? writeQueueVec_9_enq_bits_data_vd : writeQueueVec_dataOut_9_data_vd;
  assign writeQueueVec_9_deq_bits_data_offset = _writeQueueVec_fifo_9_empty ? writeQueueVec_9_enq_bits_data_offset : writeQueueVec_dataOut_9_data_offset;
  assign writeQueueVec_9_deq_bits_data_mask = _writeQueueVec_fifo_9_empty ? writeQueueVec_9_enq_bits_data_mask : writeQueueVec_dataOut_9_data_mask;
  assign writeQueueVec_9_deq_bits_data_data = _writeQueueVec_fifo_9_empty ? writeQueueVec_9_enq_bits_data_data : writeQueueVec_dataOut_9_data_data;
  assign writeQueueVec_9_deq_bits_data_last = _writeQueueVec_fifo_9_empty ? writeQueueVec_9_enq_bits_data_last : writeQueueVec_dataOut_9_data_last;
  assign writeQueueVec_9_deq_bits_data_instructionIndex = _writeQueueVec_fifo_9_empty ? writeQueueVec_9_enq_bits_data_instructionIndex : writeQueueVec_dataOut_9_data_instructionIndex;
  wire [15:0]       writeQueueVec_9_deq_bits_targetLane = _writeQueueVec_fifo_9_empty ? 16'h200 : writeQueueVec_dataOut_9_targetLane;
  wire              vrfWritePort_10_valid_0 = writeQueueVec_10_deq_valid;
  wire [4:0]        vrfWritePort_10_bits_vd_0 = writeQueueVec_10_deq_bits_data_vd;
  wire [1:0]        vrfWritePort_10_bits_offset_0 = writeQueueVec_10_deq_bits_data_offset;
  wire [3:0]        vrfWritePort_10_bits_mask_0 = writeQueueVec_10_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_10_bits_data_0 = writeQueueVec_10_deq_bits_data_data;
  wire              vrfWritePort_10_bits_last_0 = writeQueueVec_10_deq_bits_data_last;
  wire [2:0]        vrfWritePort_10_bits_instructionIndex_0 = writeQueueVec_10_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_10_enq_bits = writeQueueVec_10_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_10_enq_bits_data_data;
  wire              writeQueueVec_10_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_10 = {writeQueueVec_10_enq_bits_data_data, writeQueueVec_10_enq_bits_data_last};
  wire [2:0]        writeQueueVec_10_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_10 = {writeQueueVec_dataIn_lo_hi_10, writeQueueVec_10_enq_bits_data_instructionIndex};
  wire [4:0]        writeQueueVec_10_enq_bits_data_vd;
  wire [1:0]        writeQueueVec_10_enq_bits_data_offset;
  wire [6:0]        writeQueueVec_dataIn_hi_hi_10 = {writeQueueVec_10_enq_bits_data_vd, writeQueueVec_10_enq_bits_data_offset};
  wire [3:0]        writeQueueVec_10_enq_bits_data_mask;
  wire [10:0]       writeQueueVec_dataIn_hi_10 = {writeQueueVec_dataIn_hi_hi_10, writeQueueVec_10_enq_bits_data_mask};
  wire [62:0]       writeQueueVec_dataIn_10 = {writeQueueVec_dataIn_hi_10, writeQueueVec_dataIn_lo_10, 16'h400};
  wire [15:0]       writeQueueVec_dataOut_10_targetLane = _writeQueueVec_fifo_10_data_out[15:0];
  wire [2:0]        writeQueueVec_dataOut_10_data_instructionIndex = _writeQueueVec_fifo_10_data_out[18:16];
  wire              writeQueueVec_dataOut_10_data_last = _writeQueueVec_fifo_10_data_out[19];
  wire [31:0]       writeQueueVec_dataOut_10_data_data = _writeQueueVec_fifo_10_data_out[51:20];
  wire [3:0]        writeQueueVec_dataOut_10_data_mask = _writeQueueVec_fifo_10_data_out[55:52];
  wire [1:0]        writeQueueVec_dataOut_10_data_offset = _writeQueueVec_fifo_10_data_out[57:56];
  wire [4:0]        writeQueueVec_dataOut_10_data_vd = _writeQueueVec_fifo_10_data_out[62:58];
  wire              writeQueueVec_10_enq_ready = ~_writeQueueVec_fifo_10_full;
  wire              writeQueueVec_10_enq_valid;
  wire              _probeWire_slots_10_writeValid_T = writeQueueVec_10_enq_ready & writeQueueVec_10_enq_valid;
  assign writeQueueVec_10_deq_valid = ~_writeQueueVec_fifo_10_empty | writeQueueVec_10_enq_valid;
  assign writeQueueVec_10_deq_bits_data_vd = _writeQueueVec_fifo_10_empty ? writeQueueVec_10_enq_bits_data_vd : writeQueueVec_dataOut_10_data_vd;
  assign writeQueueVec_10_deq_bits_data_offset = _writeQueueVec_fifo_10_empty ? writeQueueVec_10_enq_bits_data_offset : writeQueueVec_dataOut_10_data_offset;
  assign writeQueueVec_10_deq_bits_data_mask = _writeQueueVec_fifo_10_empty ? writeQueueVec_10_enq_bits_data_mask : writeQueueVec_dataOut_10_data_mask;
  assign writeQueueVec_10_deq_bits_data_data = _writeQueueVec_fifo_10_empty ? writeQueueVec_10_enq_bits_data_data : writeQueueVec_dataOut_10_data_data;
  assign writeQueueVec_10_deq_bits_data_last = _writeQueueVec_fifo_10_empty ? writeQueueVec_10_enq_bits_data_last : writeQueueVec_dataOut_10_data_last;
  assign writeQueueVec_10_deq_bits_data_instructionIndex = _writeQueueVec_fifo_10_empty ? writeQueueVec_10_enq_bits_data_instructionIndex : writeQueueVec_dataOut_10_data_instructionIndex;
  wire [15:0]       writeQueueVec_10_deq_bits_targetLane = _writeQueueVec_fifo_10_empty ? 16'h400 : writeQueueVec_dataOut_10_targetLane;
  wire              vrfWritePort_11_valid_0 = writeQueueVec_11_deq_valid;
  wire [4:0]        vrfWritePort_11_bits_vd_0 = writeQueueVec_11_deq_bits_data_vd;
  wire [1:0]        vrfWritePort_11_bits_offset_0 = writeQueueVec_11_deq_bits_data_offset;
  wire [3:0]        vrfWritePort_11_bits_mask_0 = writeQueueVec_11_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_11_bits_data_0 = writeQueueVec_11_deq_bits_data_data;
  wire              vrfWritePort_11_bits_last_0 = writeQueueVec_11_deq_bits_data_last;
  wire [2:0]        vrfWritePort_11_bits_instructionIndex_0 = writeQueueVec_11_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_11_enq_bits = writeQueueVec_11_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_11_enq_bits_data_data;
  wire              writeQueueVec_11_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_11 = {writeQueueVec_11_enq_bits_data_data, writeQueueVec_11_enq_bits_data_last};
  wire [2:0]        writeQueueVec_11_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_11 = {writeQueueVec_dataIn_lo_hi_11, writeQueueVec_11_enq_bits_data_instructionIndex};
  wire [4:0]        writeQueueVec_11_enq_bits_data_vd;
  wire [1:0]        writeQueueVec_11_enq_bits_data_offset;
  wire [6:0]        writeQueueVec_dataIn_hi_hi_11 = {writeQueueVec_11_enq_bits_data_vd, writeQueueVec_11_enq_bits_data_offset};
  wire [3:0]        writeQueueVec_11_enq_bits_data_mask;
  wire [10:0]       writeQueueVec_dataIn_hi_11 = {writeQueueVec_dataIn_hi_hi_11, writeQueueVec_11_enq_bits_data_mask};
  wire [62:0]       writeQueueVec_dataIn_11 = {writeQueueVec_dataIn_hi_11, writeQueueVec_dataIn_lo_11, 16'h800};
  wire [15:0]       writeQueueVec_dataOut_11_targetLane = _writeQueueVec_fifo_11_data_out[15:0];
  wire [2:0]        writeQueueVec_dataOut_11_data_instructionIndex = _writeQueueVec_fifo_11_data_out[18:16];
  wire              writeQueueVec_dataOut_11_data_last = _writeQueueVec_fifo_11_data_out[19];
  wire [31:0]       writeQueueVec_dataOut_11_data_data = _writeQueueVec_fifo_11_data_out[51:20];
  wire [3:0]        writeQueueVec_dataOut_11_data_mask = _writeQueueVec_fifo_11_data_out[55:52];
  wire [1:0]        writeQueueVec_dataOut_11_data_offset = _writeQueueVec_fifo_11_data_out[57:56];
  wire [4:0]        writeQueueVec_dataOut_11_data_vd = _writeQueueVec_fifo_11_data_out[62:58];
  wire              writeQueueVec_11_enq_ready = ~_writeQueueVec_fifo_11_full;
  wire              writeQueueVec_11_enq_valid;
  wire              _probeWire_slots_11_writeValid_T = writeQueueVec_11_enq_ready & writeQueueVec_11_enq_valid;
  assign writeQueueVec_11_deq_valid = ~_writeQueueVec_fifo_11_empty | writeQueueVec_11_enq_valid;
  assign writeQueueVec_11_deq_bits_data_vd = _writeQueueVec_fifo_11_empty ? writeQueueVec_11_enq_bits_data_vd : writeQueueVec_dataOut_11_data_vd;
  assign writeQueueVec_11_deq_bits_data_offset = _writeQueueVec_fifo_11_empty ? writeQueueVec_11_enq_bits_data_offset : writeQueueVec_dataOut_11_data_offset;
  assign writeQueueVec_11_deq_bits_data_mask = _writeQueueVec_fifo_11_empty ? writeQueueVec_11_enq_bits_data_mask : writeQueueVec_dataOut_11_data_mask;
  assign writeQueueVec_11_deq_bits_data_data = _writeQueueVec_fifo_11_empty ? writeQueueVec_11_enq_bits_data_data : writeQueueVec_dataOut_11_data_data;
  assign writeQueueVec_11_deq_bits_data_last = _writeQueueVec_fifo_11_empty ? writeQueueVec_11_enq_bits_data_last : writeQueueVec_dataOut_11_data_last;
  assign writeQueueVec_11_deq_bits_data_instructionIndex = _writeQueueVec_fifo_11_empty ? writeQueueVec_11_enq_bits_data_instructionIndex : writeQueueVec_dataOut_11_data_instructionIndex;
  wire [15:0]       writeQueueVec_11_deq_bits_targetLane = _writeQueueVec_fifo_11_empty ? 16'h800 : writeQueueVec_dataOut_11_targetLane;
  wire              vrfWritePort_12_valid_0 = writeQueueVec_12_deq_valid;
  wire [4:0]        vrfWritePort_12_bits_vd_0 = writeQueueVec_12_deq_bits_data_vd;
  wire [1:0]        vrfWritePort_12_bits_offset_0 = writeQueueVec_12_deq_bits_data_offset;
  wire [3:0]        vrfWritePort_12_bits_mask_0 = writeQueueVec_12_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_12_bits_data_0 = writeQueueVec_12_deq_bits_data_data;
  wire              vrfWritePort_12_bits_last_0 = writeQueueVec_12_deq_bits_data_last;
  wire [2:0]        vrfWritePort_12_bits_instructionIndex_0 = writeQueueVec_12_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_12_enq_bits = writeQueueVec_12_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_12_enq_bits_data_data;
  wire              writeQueueVec_12_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_12 = {writeQueueVec_12_enq_bits_data_data, writeQueueVec_12_enq_bits_data_last};
  wire [2:0]        writeQueueVec_12_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_12 = {writeQueueVec_dataIn_lo_hi_12, writeQueueVec_12_enq_bits_data_instructionIndex};
  wire [4:0]        writeQueueVec_12_enq_bits_data_vd;
  wire [1:0]        writeQueueVec_12_enq_bits_data_offset;
  wire [6:0]        writeQueueVec_dataIn_hi_hi_12 = {writeQueueVec_12_enq_bits_data_vd, writeQueueVec_12_enq_bits_data_offset};
  wire [3:0]        writeQueueVec_12_enq_bits_data_mask;
  wire [10:0]       writeQueueVec_dataIn_hi_12 = {writeQueueVec_dataIn_hi_hi_12, writeQueueVec_12_enq_bits_data_mask};
  wire [62:0]       writeQueueVec_dataIn_12 = {writeQueueVec_dataIn_hi_12, writeQueueVec_dataIn_lo_12, 16'h1000};
  wire [15:0]       writeQueueVec_dataOut_12_targetLane = _writeQueueVec_fifo_12_data_out[15:0];
  wire [2:0]        writeQueueVec_dataOut_12_data_instructionIndex = _writeQueueVec_fifo_12_data_out[18:16];
  wire              writeQueueVec_dataOut_12_data_last = _writeQueueVec_fifo_12_data_out[19];
  wire [31:0]       writeQueueVec_dataOut_12_data_data = _writeQueueVec_fifo_12_data_out[51:20];
  wire [3:0]        writeQueueVec_dataOut_12_data_mask = _writeQueueVec_fifo_12_data_out[55:52];
  wire [1:0]        writeQueueVec_dataOut_12_data_offset = _writeQueueVec_fifo_12_data_out[57:56];
  wire [4:0]        writeQueueVec_dataOut_12_data_vd = _writeQueueVec_fifo_12_data_out[62:58];
  wire              writeQueueVec_12_enq_ready = ~_writeQueueVec_fifo_12_full;
  wire              writeQueueVec_12_enq_valid;
  wire              _probeWire_slots_12_writeValid_T = writeQueueVec_12_enq_ready & writeQueueVec_12_enq_valid;
  assign writeQueueVec_12_deq_valid = ~_writeQueueVec_fifo_12_empty | writeQueueVec_12_enq_valid;
  assign writeQueueVec_12_deq_bits_data_vd = _writeQueueVec_fifo_12_empty ? writeQueueVec_12_enq_bits_data_vd : writeQueueVec_dataOut_12_data_vd;
  assign writeQueueVec_12_deq_bits_data_offset = _writeQueueVec_fifo_12_empty ? writeQueueVec_12_enq_bits_data_offset : writeQueueVec_dataOut_12_data_offset;
  assign writeQueueVec_12_deq_bits_data_mask = _writeQueueVec_fifo_12_empty ? writeQueueVec_12_enq_bits_data_mask : writeQueueVec_dataOut_12_data_mask;
  assign writeQueueVec_12_deq_bits_data_data = _writeQueueVec_fifo_12_empty ? writeQueueVec_12_enq_bits_data_data : writeQueueVec_dataOut_12_data_data;
  assign writeQueueVec_12_deq_bits_data_last = _writeQueueVec_fifo_12_empty ? writeQueueVec_12_enq_bits_data_last : writeQueueVec_dataOut_12_data_last;
  assign writeQueueVec_12_deq_bits_data_instructionIndex = _writeQueueVec_fifo_12_empty ? writeQueueVec_12_enq_bits_data_instructionIndex : writeQueueVec_dataOut_12_data_instructionIndex;
  wire [15:0]       writeQueueVec_12_deq_bits_targetLane = _writeQueueVec_fifo_12_empty ? 16'h1000 : writeQueueVec_dataOut_12_targetLane;
  wire              vrfWritePort_13_valid_0 = writeQueueVec_13_deq_valid;
  wire [4:0]        vrfWritePort_13_bits_vd_0 = writeQueueVec_13_deq_bits_data_vd;
  wire [1:0]        vrfWritePort_13_bits_offset_0 = writeQueueVec_13_deq_bits_data_offset;
  wire [3:0]        vrfWritePort_13_bits_mask_0 = writeQueueVec_13_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_13_bits_data_0 = writeQueueVec_13_deq_bits_data_data;
  wire              vrfWritePort_13_bits_last_0 = writeQueueVec_13_deq_bits_data_last;
  wire [2:0]        vrfWritePort_13_bits_instructionIndex_0 = writeQueueVec_13_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_13_enq_bits = writeQueueVec_13_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_13_enq_bits_data_data;
  wire              writeQueueVec_13_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_13 = {writeQueueVec_13_enq_bits_data_data, writeQueueVec_13_enq_bits_data_last};
  wire [2:0]        writeQueueVec_13_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_13 = {writeQueueVec_dataIn_lo_hi_13, writeQueueVec_13_enq_bits_data_instructionIndex};
  wire [4:0]        writeQueueVec_13_enq_bits_data_vd;
  wire [1:0]        writeQueueVec_13_enq_bits_data_offset;
  wire [6:0]        writeQueueVec_dataIn_hi_hi_13 = {writeQueueVec_13_enq_bits_data_vd, writeQueueVec_13_enq_bits_data_offset};
  wire [3:0]        writeQueueVec_13_enq_bits_data_mask;
  wire [10:0]       writeQueueVec_dataIn_hi_13 = {writeQueueVec_dataIn_hi_hi_13, writeQueueVec_13_enq_bits_data_mask};
  wire [62:0]       writeQueueVec_dataIn_13 = {writeQueueVec_dataIn_hi_13, writeQueueVec_dataIn_lo_13, 16'h2000};
  wire [15:0]       writeQueueVec_dataOut_13_targetLane = _writeQueueVec_fifo_13_data_out[15:0];
  wire [2:0]        writeQueueVec_dataOut_13_data_instructionIndex = _writeQueueVec_fifo_13_data_out[18:16];
  wire              writeQueueVec_dataOut_13_data_last = _writeQueueVec_fifo_13_data_out[19];
  wire [31:0]       writeQueueVec_dataOut_13_data_data = _writeQueueVec_fifo_13_data_out[51:20];
  wire [3:0]        writeQueueVec_dataOut_13_data_mask = _writeQueueVec_fifo_13_data_out[55:52];
  wire [1:0]        writeQueueVec_dataOut_13_data_offset = _writeQueueVec_fifo_13_data_out[57:56];
  wire [4:0]        writeQueueVec_dataOut_13_data_vd = _writeQueueVec_fifo_13_data_out[62:58];
  wire              writeQueueVec_13_enq_ready = ~_writeQueueVec_fifo_13_full;
  wire              writeQueueVec_13_enq_valid;
  wire              _probeWire_slots_13_writeValid_T = writeQueueVec_13_enq_ready & writeQueueVec_13_enq_valid;
  assign writeQueueVec_13_deq_valid = ~_writeQueueVec_fifo_13_empty | writeQueueVec_13_enq_valid;
  assign writeQueueVec_13_deq_bits_data_vd = _writeQueueVec_fifo_13_empty ? writeQueueVec_13_enq_bits_data_vd : writeQueueVec_dataOut_13_data_vd;
  assign writeQueueVec_13_deq_bits_data_offset = _writeQueueVec_fifo_13_empty ? writeQueueVec_13_enq_bits_data_offset : writeQueueVec_dataOut_13_data_offset;
  assign writeQueueVec_13_deq_bits_data_mask = _writeQueueVec_fifo_13_empty ? writeQueueVec_13_enq_bits_data_mask : writeQueueVec_dataOut_13_data_mask;
  assign writeQueueVec_13_deq_bits_data_data = _writeQueueVec_fifo_13_empty ? writeQueueVec_13_enq_bits_data_data : writeQueueVec_dataOut_13_data_data;
  assign writeQueueVec_13_deq_bits_data_last = _writeQueueVec_fifo_13_empty ? writeQueueVec_13_enq_bits_data_last : writeQueueVec_dataOut_13_data_last;
  assign writeQueueVec_13_deq_bits_data_instructionIndex = _writeQueueVec_fifo_13_empty ? writeQueueVec_13_enq_bits_data_instructionIndex : writeQueueVec_dataOut_13_data_instructionIndex;
  wire [15:0]       writeQueueVec_13_deq_bits_targetLane = _writeQueueVec_fifo_13_empty ? 16'h2000 : writeQueueVec_dataOut_13_targetLane;
  wire              vrfWritePort_14_valid_0 = writeQueueVec_14_deq_valid;
  wire [4:0]        vrfWritePort_14_bits_vd_0 = writeQueueVec_14_deq_bits_data_vd;
  wire [1:0]        vrfWritePort_14_bits_offset_0 = writeQueueVec_14_deq_bits_data_offset;
  wire [3:0]        vrfWritePort_14_bits_mask_0 = writeQueueVec_14_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_14_bits_data_0 = writeQueueVec_14_deq_bits_data_data;
  wire              vrfWritePort_14_bits_last_0 = writeQueueVec_14_deq_bits_data_last;
  wire [2:0]        vrfWritePort_14_bits_instructionIndex_0 = writeQueueVec_14_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_14_enq_bits = writeQueueVec_14_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_14_enq_bits_data_data;
  wire              writeQueueVec_14_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_14 = {writeQueueVec_14_enq_bits_data_data, writeQueueVec_14_enq_bits_data_last};
  wire [2:0]        writeQueueVec_14_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_14 = {writeQueueVec_dataIn_lo_hi_14, writeQueueVec_14_enq_bits_data_instructionIndex};
  wire [4:0]        writeQueueVec_14_enq_bits_data_vd;
  wire [1:0]        writeQueueVec_14_enq_bits_data_offset;
  wire [6:0]        writeQueueVec_dataIn_hi_hi_14 = {writeQueueVec_14_enq_bits_data_vd, writeQueueVec_14_enq_bits_data_offset};
  wire [3:0]        writeQueueVec_14_enq_bits_data_mask;
  wire [10:0]       writeQueueVec_dataIn_hi_14 = {writeQueueVec_dataIn_hi_hi_14, writeQueueVec_14_enq_bits_data_mask};
  wire [62:0]       writeQueueVec_dataIn_14 = {writeQueueVec_dataIn_hi_14, writeQueueVec_dataIn_lo_14, 16'h4000};
  wire [15:0]       writeQueueVec_dataOut_14_targetLane = _writeQueueVec_fifo_14_data_out[15:0];
  wire [2:0]        writeQueueVec_dataOut_14_data_instructionIndex = _writeQueueVec_fifo_14_data_out[18:16];
  wire              writeQueueVec_dataOut_14_data_last = _writeQueueVec_fifo_14_data_out[19];
  wire [31:0]       writeQueueVec_dataOut_14_data_data = _writeQueueVec_fifo_14_data_out[51:20];
  wire [3:0]        writeQueueVec_dataOut_14_data_mask = _writeQueueVec_fifo_14_data_out[55:52];
  wire [1:0]        writeQueueVec_dataOut_14_data_offset = _writeQueueVec_fifo_14_data_out[57:56];
  wire [4:0]        writeQueueVec_dataOut_14_data_vd = _writeQueueVec_fifo_14_data_out[62:58];
  wire              writeQueueVec_14_enq_ready = ~_writeQueueVec_fifo_14_full;
  wire              writeQueueVec_14_enq_valid;
  wire              _probeWire_slots_14_writeValid_T = writeQueueVec_14_enq_ready & writeQueueVec_14_enq_valid;
  assign writeQueueVec_14_deq_valid = ~_writeQueueVec_fifo_14_empty | writeQueueVec_14_enq_valid;
  assign writeQueueVec_14_deq_bits_data_vd = _writeQueueVec_fifo_14_empty ? writeQueueVec_14_enq_bits_data_vd : writeQueueVec_dataOut_14_data_vd;
  assign writeQueueVec_14_deq_bits_data_offset = _writeQueueVec_fifo_14_empty ? writeQueueVec_14_enq_bits_data_offset : writeQueueVec_dataOut_14_data_offset;
  assign writeQueueVec_14_deq_bits_data_mask = _writeQueueVec_fifo_14_empty ? writeQueueVec_14_enq_bits_data_mask : writeQueueVec_dataOut_14_data_mask;
  assign writeQueueVec_14_deq_bits_data_data = _writeQueueVec_fifo_14_empty ? writeQueueVec_14_enq_bits_data_data : writeQueueVec_dataOut_14_data_data;
  assign writeQueueVec_14_deq_bits_data_last = _writeQueueVec_fifo_14_empty ? writeQueueVec_14_enq_bits_data_last : writeQueueVec_dataOut_14_data_last;
  assign writeQueueVec_14_deq_bits_data_instructionIndex = _writeQueueVec_fifo_14_empty ? writeQueueVec_14_enq_bits_data_instructionIndex : writeQueueVec_dataOut_14_data_instructionIndex;
  wire [15:0]       writeQueueVec_14_deq_bits_targetLane = _writeQueueVec_fifo_14_empty ? 16'h4000 : writeQueueVec_dataOut_14_targetLane;
  wire              vrfWritePort_15_valid_0 = writeQueueVec_15_deq_valid;
  wire [4:0]        vrfWritePort_15_bits_vd_0 = writeQueueVec_15_deq_bits_data_vd;
  wire [1:0]        vrfWritePort_15_bits_offset_0 = writeQueueVec_15_deq_bits_data_offset;
  wire [3:0]        vrfWritePort_15_bits_mask_0 = writeQueueVec_15_deq_bits_data_mask;
  wire [31:0]       vrfWritePort_15_bits_data_0 = writeQueueVec_15_deq_bits_data_data;
  wire              vrfWritePort_15_bits_last_0 = writeQueueVec_15_deq_bits_data_last;
  wire [2:0]        vrfWritePort_15_bits_instructionIndex_0 = writeQueueVec_15_deq_bits_data_instructionIndex;
  wire [2:0]        writeIndexQueue_15_enq_bits = writeQueueVec_15_deq_bits_data_instructionIndex;
  wire [31:0]       writeQueueVec_15_enq_bits_data_data;
  wire              writeQueueVec_15_enq_bits_data_last;
  wire [32:0]       writeQueueVec_dataIn_lo_hi_15 = {writeQueueVec_15_enq_bits_data_data, writeQueueVec_15_enq_bits_data_last};
  wire [2:0]        writeQueueVec_15_enq_bits_data_instructionIndex;
  wire [35:0]       writeQueueVec_dataIn_lo_15 = {writeQueueVec_dataIn_lo_hi_15, writeQueueVec_15_enq_bits_data_instructionIndex};
  wire [4:0]        writeQueueVec_15_enq_bits_data_vd;
  wire [1:0]        writeQueueVec_15_enq_bits_data_offset;
  wire [6:0]        writeQueueVec_dataIn_hi_hi_15 = {writeQueueVec_15_enq_bits_data_vd, writeQueueVec_15_enq_bits_data_offset};
  wire [3:0]        writeQueueVec_15_enq_bits_data_mask;
  wire [10:0]       writeQueueVec_dataIn_hi_15 = {writeQueueVec_dataIn_hi_hi_15, writeQueueVec_15_enq_bits_data_mask};
  wire [62:0]       writeQueueVec_dataIn_15 = {writeQueueVec_dataIn_hi_15, writeQueueVec_dataIn_lo_15, 16'h8000};
  wire [15:0]       writeQueueVec_dataOut_15_targetLane = _writeQueueVec_fifo_15_data_out[15:0];
  wire [2:0]        writeQueueVec_dataOut_15_data_instructionIndex = _writeQueueVec_fifo_15_data_out[18:16];
  wire              writeQueueVec_dataOut_15_data_last = _writeQueueVec_fifo_15_data_out[19];
  wire [31:0]       writeQueueVec_dataOut_15_data_data = _writeQueueVec_fifo_15_data_out[51:20];
  wire [3:0]        writeQueueVec_dataOut_15_data_mask = _writeQueueVec_fifo_15_data_out[55:52];
  wire [1:0]        writeQueueVec_dataOut_15_data_offset = _writeQueueVec_fifo_15_data_out[57:56];
  wire [4:0]        writeQueueVec_dataOut_15_data_vd = _writeQueueVec_fifo_15_data_out[62:58];
  wire              writeQueueVec_15_enq_ready = ~_writeQueueVec_fifo_15_full;
  wire              writeQueueVec_15_enq_valid;
  wire              _probeWire_slots_15_writeValid_T = writeQueueVec_15_enq_ready & writeQueueVec_15_enq_valid;
  assign writeQueueVec_15_deq_valid = ~_writeQueueVec_fifo_15_empty | writeQueueVec_15_enq_valid;
  assign writeQueueVec_15_deq_bits_data_vd = _writeQueueVec_fifo_15_empty ? writeQueueVec_15_enq_bits_data_vd : writeQueueVec_dataOut_15_data_vd;
  assign writeQueueVec_15_deq_bits_data_offset = _writeQueueVec_fifo_15_empty ? writeQueueVec_15_enq_bits_data_offset : writeQueueVec_dataOut_15_data_offset;
  assign writeQueueVec_15_deq_bits_data_mask = _writeQueueVec_fifo_15_empty ? writeQueueVec_15_enq_bits_data_mask : writeQueueVec_dataOut_15_data_mask;
  assign writeQueueVec_15_deq_bits_data_data = _writeQueueVec_fifo_15_empty ? writeQueueVec_15_enq_bits_data_data : writeQueueVec_dataOut_15_data_data;
  assign writeQueueVec_15_deq_bits_data_last = _writeQueueVec_fifo_15_empty ? writeQueueVec_15_enq_bits_data_last : writeQueueVec_dataOut_15_data_last;
  assign writeQueueVec_15_deq_bits_data_instructionIndex = _writeQueueVec_fifo_15_empty ? writeQueueVec_15_enq_bits_data_instructionIndex : writeQueueVec_dataOut_15_data_instructionIndex;
  wire [15:0]       writeQueueVec_15_deq_bits_targetLane = _writeQueueVec_fifo_15_empty ? 16'h8000 : writeQueueVec_dataOut_15_targetLane;
  wire              otherUnitTargetQueue_deq_valid;
  assign otherUnitTargetQueue_deq_valid = ~_otherUnitTargetQueue_fifo_empty;
  wire              otherUnitTargetQueue_deq_ready;
  wire              otherUnitTargetQueue_enq_ready = ~_otherUnitTargetQueue_fifo_full | otherUnitTargetQueue_deq_ready;
  wire              otherUnitTargetQueue_enq_valid;
  wire              otherUnitDataQueueVec_0_enq_ready = ~_otherUnitDataQueueVec_fifo_full;
  wire              otherUnitDataQueueVec_0_deq_ready;
  wire              otherUnitDataQueueVec_0_enq_valid;
  wire              otherUnitDataQueueVec_0_deq_valid = ~_otherUnitDataQueueVec_fifo_empty | otherUnitDataQueueVec_0_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_0_deq_bits = _otherUnitDataQueueVec_fifo_empty ? otherUnitDataQueueVec_0_enq_bits : _otherUnitDataQueueVec_fifo_data_out;
  wire              otherUnitDataQueueVec_1_enq_ready = ~_otherUnitDataQueueVec_fifo_1_full;
  wire              otherUnitDataQueueVec_1_deq_ready;
  wire              otherUnitDataQueueVec_1_enq_valid;
  wire              otherUnitDataQueueVec_1_deq_valid = ~_otherUnitDataQueueVec_fifo_1_empty | otherUnitDataQueueVec_1_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_1_deq_bits = _otherUnitDataQueueVec_fifo_1_empty ? otherUnitDataQueueVec_1_enq_bits : _otherUnitDataQueueVec_fifo_1_data_out;
  wire              otherUnitDataQueueVec_2_enq_ready = ~_otherUnitDataQueueVec_fifo_2_full;
  wire              otherUnitDataQueueVec_2_deq_ready;
  wire              otherUnitDataQueueVec_2_enq_valid;
  wire              otherUnitDataQueueVec_2_deq_valid = ~_otherUnitDataQueueVec_fifo_2_empty | otherUnitDataQueueVec_2_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_2_deq_bits = _otherUnitDataQueueVec_fifo_2_empty ? otherUnitDataQueueVec_2_enq_bits : _otherUnitDataQueueVec_fifo_2_data_out;
  wire              otherUnitDataQueueVec_3_enq_ready = ~_otherUnitDataQueueVec_fifo_3_full;
  wire              otherUnitDataQueueVec_3_deq_ready;
  wire              otherUnitDataQueueVec_3_enq_valid;
  wire              otherUnitDataQueueVec_3_deq_valid = ~_otherUnitDataQueueVec_fifo_3_empty | otherUnitDataQueueVec_3_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_3_deq_bits = _otherUnitDataQueueVec_fifo_3_empty ? otherUnitDataQueueVec_3_enq_bits : _otherUnitDataQueueVec_fifo_3_data_out;
  wire              otherUnitDataQueueVec_4_enq_ready = ~_otherUnitDataQueueVec_fifo_4_full;
  wire              otherUnitDataQueueVec_4_deq_ready;
  wire              otherUnitDataQueueVec_4_enq_valid;
  wire              otherUnitDataQueueVec_4_deq_valid = ~_otherUnitDataQueueVec_fifo_4_empty | otherUnitDataQueueVec_4_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_4_deq_bits = _otherUnitDataQueueVec_fifo_4_empty ? otherUnitDataQueueVec_4_enq_bits : _otherUnitDataQueueVec_fifo_4_data_out;
  wire              otherUnitDataQueueVec_5_enq_ready = ~_otherUnitDataQueueVec_fifo_5_full;
  wire              otherUnitDataQueueVec_5_deq_ready;
  wire              otherUnitDataQueueVec_5_enq_valid;
  wire              otherUnitDataQueueVec_5_deq_valid = ~_otherUnitDataQueueVec_fifo_5_empty | otherUnitDataQueueVec_5_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_5_deq_bits = _otherUnitDataQueueVec_fifo_5_empty ? otherUnitDataQueueVec_5_enq_bits : _otherUnitDataQueueVec_fifo_5_data_out;
  wire              otherUnitDataQueueVec_6_enq_ready = ~_otherUnitDataQueueVec_fifo_6_full;
  wire              otherUnitDataQueueVec_6_deq_ready;
  wire              otherUnitDataQueueVec_6_enq_valid;
  wire              otherUnitDataQueueVec_6_deq_valid = ~_otherUnitDataQueueVec_fifo_6_empty | otherUnitDataQueueVec_6_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_6_deq_bits = _otherUnitDataQueueVec_fifo_6_empty ? otherUnitDataQueueVec_6_enq_bits : _otherUnitDataQueueVec_fifo_6_data_out;
  wire              otherUnitDataQueueVec_7_enq_ready = ~_otherUnitDataQueueVec_fifo_7_full;
  wire              otherUnitDataQueueVec_7_deq_ready;
  wire              otherUnitDataQueueVec_7_enq_valid;
  wire              otherUnitDataQueueVec_7_deq_valid = ~_otherUnitDataQueueVec_fifo_7_empty | otherUnitDataQueueVec_7_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_7_deq_bits = _otherUnitDataQueueVec_fifo_7_empty ? otherUnitDataQueueVec_7_enq_bits : _otherUnitDataQueueVec_fifo_7_data_out;
  wire              otherUnitDataQueueVec_8_enq_ready = ~_otherUnitDataQueueVec_fifo_8_full;
  wire              otherUnitDataQueueVec_8_deq_ready;
  wire              otherUnitDataQueueVec_8_enq_valid;
  wire              otherUnitDataQueueVec_8_deq_valid = ~_otherUnitDataQueueVec_fifo_8_empty | otherUnitDataQueueVec_8_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_8_deq_bits = _otherUnitDataQueueVec_fifo_8_empty ? otherUnitDataQueueVec_8_enq_bits : _otherUnitDataQueueVec_fifo_8_data_out;
  wire              otherUnitDataQueueVec_9_enq_ready = ~_otherUnitDataQueueVec_fifo_9_full;
  wire              otherUnitDataQueueVec_9_deq_ready;
  wire              otherUnitDataQueueVec_9_enq_valid;
  wire              otherUnitDataQueueVec_9_deq_valid = ~_otherUnitDataQueueVec_fifo_9_empty | otherUnitDataQueueVec_9_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_9_deq_bits = _otherUnitDataQueueVec_fifo_9_empty ? otherUnitDataQueueVec_9_enq_bits : _otherUnitDataQueueVec_fifo_9_data_out;
  wire              otherUnitDataQueueVec_10_enq_ready = ~_otherUnitDataQueueVec_fifo_10_full;
  wire              otherUnitDataQueueVec_10_deq_ready;
  wire              otherUnitDataQueueVec_10_enq_valid;
  wire              otherUnitDataQueueVec_10_deq_valid = ~_otherUnitDataQueueVec_fifo_10_empty | otherUnitDataQueueVec_10_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_10_deq_bits = _otherUnitDataQueueVec_fifo_10_empty ? otherUnitDataQueueVec_10_enq_bits : _otherUnitDataQueueVec_fifo_10_data_out;
  wire              otherUnitDataQueueVec_11_enq_ready = ~_otherUnitDataQueueVec_fifo_11_full;
  wire              otherUnitDataQueueVec_11_deq_ready;
  wire              otherUnitDataQueueVec_11_enq_valid;
  wire              otherUnitDataQueueVec_11_deq_valid = ~_otherUnitDataQueueVec_fifo_11_empty | otherUnitDataQueueVec_11_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_11_deq_bits = _otherUnitDataQueueVec_fifo_11_empty ? otherUnitDataQueueVec_11_enq_bits : _otherUnitDataQueueVec_fifo_11_data_out;
  wire              otherUnitDataQueueVec_12_enq_ready = ~_otherUnitDataQueueVec_fifo_12_full;
  wire              otherUnitDataQueueVec_12_deq_ready;
  wire              otherUnitDataQueueVec_12_enq_valid;
  wire              otherUnitDataQueueVec_12_deq_valid = ~_otherUnitDataQueueVec_fifo_12_empty | otherUnitDataQueueVec_12_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_12_deq_bits = _otherUnitDataQueueVec_fifo_12_empty ? otherUnitDataQueueVec_12_enq_bits : _otherUnitDataQueueVec_fifo_12_data_out;
  wire              otherUnitDataQueueVec_13_enq_ready = ~_otherUnitDataQueueVec_fifo_13_full;
  wire              otherUnitDataQueueVec_13_deq_ready;
  wire              otherUnitDataQueueVec_13_enq_valid;
  wire              otherUnitDataQueueVec_13_deq_valid = ~_otherUnitDataQueueVec_fifo_13_empty | otherUnitDataQueueVec_13_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_13_deq_bits = _otherUnitDataQueueVec_fifo_13_empty ? otherUnitDataQueueVec_13_enq_bits : _otherUnitDataQueueVec_fifo_13_data_out;
  wire              otherUnitDataQueueVec_14_enq_ready = ~_otherUnitDataQueueVec_fifo_14_full;
  wire              otherUnitDataQueueVec_14_deq_ready;
  wire              otherUnitDataQueueVec_14_enq_valid;
  wire              otherUnitDataQueueVec_14_deq_valid = ~_otherUnitDataQueueVec_fifo_14_empty | otherUnitDataQueueVec_14_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_14_deq_bits = _otherUnitDataQueueVec_fifo_14_empty ? otherUnitDataQueueVec_14_enq_bits : _otherUnitDataQueueVec_fifo_14_data_out;
  wire              otherUnitDataQueueVec_15_enq_ready = ~_otherUnitDataQueueVec_fifo_15_full;
  wire              otherUnitDataQueueVec_15_deq_ready;
  wire              otherUnitDataQueueVec_15_enq_valid;
  wire              otherUnitDataQueueVec_15_deq_valid = ~_otherUnitDataQueueVec_fifo_15_empty | otherUnitDataQueueVec_15_enq_valid;
  wire [31:0]       otherUnitDataQueueVec_15_deq_bits = _otherUnitDataQueueVec_fifo_15_empty ? otherUnitDataQueueVec_15_enq_bits : _otherUnitDataQueueVec_fifo_15_data_out;
  wire [15:0]       otherTryReadVrf = _otherUnit_vrfReadDataPorts_valid ? _otherUnit_status_targetLane : 16'h0;
  wire              vrfReadDataPorts_0_valid_0 = otherTryReadVrf[0] | _storeUnit_vrfReadDataPorts_0_valid;
  wire [4:0]        vrfReadDataPorts_0_bits_vs_0 = otherTryReadVrf[0] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_0_bits_vs;
  wire [1:0]        vrfReadDataPorts_0_bits_offset_0 = otherTryReadVrf[0] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_0_bits_offset;
  wire [2:0]        vrfReadDataPorts_0_bits_instructionIndex_0 = otherTryReadVrf[0] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_0_bits_instructionIndex;
  wire              otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_0_enq_valid = vrfReadResults_0_valid & ~otherUnitTargetQueue_empty;
  wire [15:0]       dataDeqFire;
  assign otherUnitDataQueueVec_0_deq_ready = dataDeqFire[0];
  wire              vrfReadDataPorts_1_valid_0 = otherTryReadVrf[1] | _storeUnit_vrfReadDataPorts_1_valid;
  wire [4:0]        vrfReadDataPorts_1_bits_vs_0 = otherTryReadVrf[1] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_1_bits_vs;
  wire [1:0]        vrfReadDataPorts_1_bits_offset_0 = otherTryReadVrf[1] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_1_bits_offset;
  wire [2:0]        vrfReadDataPorts_1_bits_instructionIndex_0 = otherTryReadVrf[1] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_1_bits_instructionIndex;
  assign otherUnitDataQueueVec_1_enq_valid = vrfReadResults_1_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_1_deq_ready = dataDeqFire[1];
  wire              vrfReadDataPorts_2_valid_0 = otherTryReadVrf[2] | _storeUnit_vrfReadDataPorts_2_valid;
  wire [4:0]        vrfReadDataPorts_2_bits_vs_0 = otherTryReadVrf[2] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_2_bits_vs;
  wire [1:0]        vrfReadDataPorts_2_bits_offset_0 = otherTryReadVrf[2] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_2_bits_offset;
  wire [2:0]        vrfReadDataPorts_2_bits_instructionIndex_0 = otherTryReadVrf[2] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_2_bits_instructionIndex;
  assign otherUnitDataQueueVec_2_enq_valid = vrfReadResults_2_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_2_deq_ready = dataDeqFire[2];
  wire              vrfReadDataPorts_3_valid_0 = otherTryReadVrf[3] | _storeUnit_vrfReadDataPorts_3_valid;
  wire [4:0]        vrfReadDataPorts_3_bits_vs_0 = otherTryReadVrf[3] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_3_bits_vs;
  wire [1:0]        vrfReadDataPorts_3_bits_offset_0 = otherTryReadVrf[3] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_3_bits_offset;
  wire [2:0]        vrfReadDataPorts_3_bits_instructionIndex_0 = otherTryReadVrf[3] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_3_bits_instructionIndex;
  assign otherUnitDataQueueVec_3_enq_valid = vrfReadResults_3_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_3_deq_ready = dataDeqFire[3];
  wire              vrfReadDataPorts_4_valid_0 = otherTryReadVrf[4] | _storeUnit_vrfReadDataPorts_4_valid;
  wire [4:0]        vrfReadDataPorts_4_bits_vs_0 = otherTryReadVrf[4] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_4_bits_vs;
  wire [1:0]        vrfReadDataPorts_4_bits_offset_0 = otherTryReadVrf[4] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_4_bits_offset;
  wire [2:0]        vrfReadDataPorts_4_bits_instructionIndex_0 = otherTryReadVrf[4] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_4_bits_instructionIndex;
  assign otherUnitDataQueueVec_4_enq_valid = vrfReadResults_4_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_4_deq_ready = dataDeqFire[4];
  wire              vrfReadDataPorts_5_valid_0 = otherTryReadVrf[5] | _storeUnit_vrfReadDataPorts_5_valid;
  wire [4:0]        vrfReadDataPorts_5_bits_vs_0 = otherTryReadVrf[5] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_5_bits_vs;
  wire [1:0]        vrfReadDataPorts_5_bits_offset_0 = otherTryReadVrf[5] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_5_bits_offset;
  wire [2:0]        vrfReadDataPorts_5_bits_instructionIndex_0 = otherTryReadVrf[5] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_5_bits_instructionIndex;
  assign otherUnitDataQueueVec_5_enq_valid = vrfReadResults_5_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_5_deq_ready = dataDeqFire[5];
  wire              vrfReadDataPorts_6_valid_0 = otherTryReadVrf[6] | _storeUnit_vrfReadDataPorts_6_valid;
  wire [4:0]        vrfReadDataPorts_6_bits_vs_0 = otherTryReadVrf[6] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_6_bits_vs;
  wire [1:0]        vrfReadDataPorts_6_bits_offset_0 = otherTryReadVrf[6] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_6_bits_offset;
  wire [2:0]        vrfReadDataPorts_6_bits_instructionIndex_0 = otherTryReadVrf[6] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_6_bits_instructionIndex;
  assign otherUnitDataQueueVec_6_enq_valid = vrfReadResults_6_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_6_deq_ready = dataDeqFire[6];
  wire              vrfReadDataPorts_7_valid_0 = otherTryReadVrf[7] | _storeUnit_vrfReadDataPorts_7_valid;
  wire [4:0]        vrfReadDataPorts_7_bits_vs_0 = otherTryReadVrf[7] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_7_bits_vs;
  wire [1:0]        vrfReadDataPorts_7_bits_offset_0 = otherTryReadVrf[7] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_7_bits_offset;
  wire [2:0]        vrfReadDataPorts_7_bits_instructionIndex_0 = otherTryReadVrf[7] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_7_bits_instructionIndex;
  assign otherUnitDataQueueVec_7_enq_valid = vrfReadResults_7_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_7_deq_ready = dataDeqFire[7];
  wire              vrfReadDataPorts_8_valid_0 = otherTryReadVrf[8] | _storeUnit_vrfReadDataPorts_8_valid;
  wire [4:0]        vrfReadDataPorts_8_bits_vs_0 = otherTryReadVrf[8] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_8_bits_vs;
  wire [1:0]        vrfReadDataPorts_8_bits_offset_0 = otherTryReadVrf[8] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_8_bits_offset;
  wire [2:0]        vrfReadDataPorts_8_bits_instructionIndex_0 = otherTryReadVrf[8] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_8_bits_instructionIndex;
  assign otherUnitDataQueueVec_8_enq_valid = vrfReadResults_8_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_8_deq_ready = dataDeqFire[8];
  wire              vrfReadDataPorts_9_valid_0 = otherTryReadVrf[9] | _storeUnit_vrfReadDataPorts_9_valid;
  wire [4:0]        vrfReadDataPorts_9_bits_vs_0 = otherTryReadVrf[9] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_9_bits_vs;
  wire [1:0]        vrfReadDataPorts_9_bits_offset_0 = otherTryReadVrf[9] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_9_bits_offset;
  wire [2:0]        vrfReadDataPorts_9_bits_instructionIndex_0 = otherTryReadVrf[9] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_9_bits_instructionIndex;
  assign otherUnitDataQueueVec_9_enq_valid = vrfReadResults_9_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_9_deq_ready = dataDeqFire[9];
  wire              vrfReadDataPorts_10_valid_0 = otherTryReadVrf[10] | _storeUnit_vrfReadDataPorts_10_valid;
  wire [4:0]        vrfReadDataPorts_10_bits_vs_0 = otherTryReadVrf[10] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_10_bits_vs;
  wire [1:0]        vrfReadDataPorts_10_bits_offset_0 = otherTryReadVrf[10] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_10_bits_offset;
  wire [2:0]        vrfReadDataPorts_10_bits_instructionIndex_0 = otherTryReadVrf[10] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_10_bits_instructionIndex;
  assign otherUnitDataQueueVec_10_enq_valid = vrfReadResults_10_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_10_deq_ready = dataDeqFire[10];
  wire              vrfReadDataPorts_11_valid_0 = otherTryReadVrf[11] | _storeUnit_vrfReadDataPorts_11_valid;
  wire [4:0]        vrfReadDataPorts_11_bits_vs_0 = otherTryReadVrf[11] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_11_bits_vs;
  wire [1:0]        vrfReadDataPorts_11_bits_offset_0 = otherTryReadVrf[11] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_11_bits_offset;
  wire [2:0]        vrfReadDataPorts_11_bits_instructionIndex_0 = otherTryReadVrf[11] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_11_bits_instructionIndex;
  assign otherUnitDataQueueVec_11_enq_valid = vrfReadResults_11_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_11_deq_ready = dataDeqFire[11];
  wire              vrfReadDataPorts_12_valid_0 = otherTryReadVrf[12] | _storeUnit_vrfReadDataPorts_12_valid;
  wire [4:0]        vrfReadDataPorts_12_bits_vs_0 = otherTryReadVrf[12] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_12_bits_vs;
  wire [1:0]        vrfReadDataPorts_12_bits_offset_0 = otherTryReadVrf[12] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_12_bits_offset;
  wire [2:0]        vrfReadDataPorts_12_bits_instructionIndex_0 = otherTryReadVrf[12] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_12_bits_instructionIndex;
  assign otherUnitDataQueueVec_12_enq_valid = vrfReadResults_12_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_12_deq_ready = dataDeqFire[12];
  wire              vrfReadDataPorts_13_valid_0 = otherTryReadVrf[13] | _storeUnit_vrfReadDataPorts_13_valid;
  wire [4:0]        vrfReadDataPorts_13_bits_vs_0 = otherTryReadVrf[13] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_13_bits_vs;
  wire [1:0]        vrfReadDataPorts_13_bits_offset_0 = otherTryReadVrf[13] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_13_bits_offset;
  wire [2:0]        vrfReadDataPorts_13_bits_instructionIndex_0 = otherTryReadVrf[13] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_13_bits_instructionIndex;
  assign otherUnitDataQueueVec_13_enq_valid = vrfReadResults_13_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_13_deq_ready = dataDeqFire[13];
  wire              vrfReadDataPorts_14_valid_0 = otherTryReadVrf[14] | _storeUnit_vrfReadDataPorts_14_valid;
  wire [4:0]        vrfReadDataPorts_14_bits_vs_0 = otherTryReadVrf[14] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_14_bits_vs;
  wire [1:0]        vrfReadDataPorts_14_bits_offset_0 = otherTryReadVrf[14] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_14_bits_offset;
  wire [2:0]        vrfReadDataPorts_14_bits_instructionIndex_0 = otherTryReadVrf[14] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_14_bits_instructionIndex;
  assign otherUnitDataQueueVec_14_enq_valid = vrfReadResults_14_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_14_deq_ready = dataDeqFire[14];
  wire              vrfReadDataPorts_15_valid_0 = otherTryReadVrf[15] | _storeUnit_vrfReadDataPorts_15_valid;
  wire [4:0]        vrfReadDataPorts_15_bits_vs_0 = otherTryReadVrf[15] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_15_bits_vs;
  wire [1:0]        vrfReadDataPorts_15_bits_offset_0 = otherTryReadVrf[15] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_15_bits_offset;
  wire [2:0]        vrfReadDataPorts_15_bits_instructionIndex_0 = otherTryReadVrf[15] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_15_bits_instructionIndex;
  assign otherUnitDataQueueVec_15_enq_valid = vrfReadResults_15_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_15_deq_ready = dataDeqFire[15];
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_lo_lo_lo = {vrfReadDataPorts_1_ready_0, vrfReadDataPorts_0_ready_0};
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_lo_lo_hi = {vrfReadDataPorts_3_ready_0, vrfReadDataPorts_2_ready_0};
  wire [3:0]        otherUnit_vrfReadDataPorts_ready_lo_lo = {otherUnit_vrfReadDataPorts_ready_lo_lo_hi, otherUnit_vrfReadDataPorts_ready_lo_lo_lo};
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_lo_hi_lo = {vrfReadDataPorts_5_ready_0, vrfReadDataPorts_4_ready_0};
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_lo_hi_hi = {vrfReadDataPorts_7_ready_0, vrfReadDataPorts_6_ready_0};
  wire [3:0]        otherUnit_vrfReadDataPorts_ready_lo_hi = {otherUnit_vrfReadDataPorts_ready_lo_hi_hi, otherUnit_vrfReadDataPorts_ready_lo_hi_lo};
  wire [7:0]        otherUnit_vrfReadDataPorts_ready_lo = {otherUnit_vrfReadDataPorts_ready_lo_hi, otherUnit_vrfReadDataPorts_ready_lo_lo};
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_hi_lo_lo = {vrfReadDataPorts_9_ready_0, vrfReadDataPorts_8_ready_0};
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_hi_lo_hi = {vrfReadDataPorts_11_ready_0, vrfReadDataPorts_10_ready_0};
  wire [3:0]        otherUnit_vrfReadDataPorts_ready_hi_lo = {otherUnit_vrfReadDataPorts_ready_hi_lo_hi, otherUnit_vrfReadDataPorts_ready_hi_lo_lo};
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_hi_hi_lo = {vrfReadDataPorts_13_ready_0, vrfReadDataPorts_12_ready_0};
  wire [1:0]        otherUnit_vrfReadDataPorts_ready_hi_hi_hi = {vrfReadDataPorts_15_ready_0, vrfReadDataPorts_14_ready_0};
  wire [3:0]        otherUnit_vrfReadDataPorts_ready_hi_hi = {otherUnit_vrfReadDataPorts_ready_hi_hi_hi, otherUnit_vrfReadDataPorts_ready_hi_hi_lo};
  wire [7:0]        otherUnit_vrfReadDataPorts_ready_hi = {otherUnit_vrfReadDataPorts_ready_hi_hi, otherUnit_vrfReadDataPorts_ready_hi_lo};
  wire              otherUnit_vrfReadDataPorts_ready = (|(otherTryReadVrf & {otherUnit_vrfReadDataPorts_ready_hi, otherUnit_vrfReadDataPorts_ready_lo})) & otherUnitTargetQueue_enq_ready;
  assign otherUnitTargetQueue_enq_valid = otherUnit_vrfReadDataPorts_ready & _otherUnit_vrfReadDataPorts_valid;
  wire [15:0]       otherUnitTargetQueue_deq_bits;
  wire [1:0]        otherUnit_vrfReadResults_valid_lo_lo_lo = {otherUnitDataQueueVec_1_deq_valid, otherUnitDataQueueVec_0_deq_valid};
  wire [1:0]        otherUnit_vrfReadResults_valid_lo_lo_hi = {otherUnitDataQueueVec_3_deq_valid, otherUnitDataQueueVec_2_deq_valid};
  wire [3:0]        otherUnit_vrfReadResults_valid_lo_lo = {otherUnit_vrfReadResults_valid_lo_lo_hi, otherUnit_vrfReadResults_valid_lo_lo_lo};
  wire [1:0]        otherUnit_vrfReadResults_valid_lo_hi_lo = {otherUnitDataQueueVec_5_deq_valid, otherUnitDataQueueVec_4_deq_valid};
  wire [1:0]        otherUnit_vrfReadResults_valid_lo_hi_hi = {otherUnitDataQueueVec_7_deq_valid, otherUnitDataQueueVec_6_deq_valid};
  wire [3:0]        otherUnit_vrfReadResults_valid_lo_hi = {otherUnit_vrfReadResults_valid_lo_hi_hi, otherUnit_vrfReadResults_valid_lo_hi_lo};
  wire [7:0]        otherUnit_vrfReadResults_valid_lo = {otherUnit_vrfReadResults_valid_lo_hi, otherUnit_vrfReadResults_valid_lo_lo};
  wire [1:0]        otherUnit_vrfReadResults_valid_hi_lo_lo = {otherUnitDataQueueVec_9_deq_valid, otherUnitDataQueueVec_8_deq_valid};
  wire [1:0]        otherUnit_vrfReadResults_valid_hi_lo_hi = {otherUnitDataQueueVec_11_deq_valid, otherUnitDataQueueVec_10_deq_valid};
  wire [3:0]        otherUnit_vrfReadResults_valid_hi_lo = {otherUnit_vrfReadResults_valid_hi_lo_hi, otherUnit_vrfReadResults_valid_hi_lo_lo};
  wire [1:0]        otherUnit_vrfReadResults_valid_hi_hi_lo = {otherUnitDataQueueVec_13_deq_valid, otherUnitDataQueueVec_12_deq_valid};
  wire [1:0]        otherUnit_vrfReadResults_valid_hi_hi_hi = {otherUnitDataQueueVec_15_deq_valid, otherUnitDataQueueVec_14_deq_valid};
  wire [3:0]        otherUnit_vrfReadResults_valid_hi_hi = {otherUnit_vrfReadResults_valid_hi_hi_hi, otherUnit_vrfReadResults_valid_hi_hi_lo};
  wire [7:0]        otherUnit_vrfReadResults_valid_hi = {otherUnit_vrfReadResults_valid_hi_hi, otherUnit_vrfReadResults_valid_hi_lo};
  assign otherUnitTargetQueue_deq_ready = otherUnitTargetQueue_deq_valid & (|(otherUnitTargetQueue_deq_bits & {otherUnit_vrfReadResults_valid_hi, otherUnit_vrfReadResults_valid_lo}));
  assign dataDeqFire = otherUnitTargetQueue_deq_ready ? otherUnitTargetQueue_deq_bits : 16'h0;
  wire [15:0]       otherTryToWrite = _otherUnit_vrfWritePort_valid ? _otherUnit_status_targetLane : 16'h0;
  wire [1:0]        otherUnit_vrfWritePort_ready_lo_lo_lo = {writeQueueVec_1_enq_ready, writeQueueVec_0_enq_ready};
  wire [1:0]        otherUnit_vrfWritePort_ready_lo_lo_hi = {writeQueueVec_3_enq_ready, writeQueueVec_2_enq_ready};
  wire [3:0]        otherUnit_vrfWritePort_ready_lo_lo = {otherUnit_vrfWritePort_ready_lo_lo_hi, otherUnit_vrfWritePort_ready_lo_lo_lo};
  wire [1:0]        otherUnit_vrfWritePort_ready_lo_hi_lo = {writeQueueVec_5_enq_ready, writeQueueVec_4_enq_ready};
  wire [1:0]        otherUnit_vrfWritePort_ready_lo_hi_hi = {writeQueueVec_7_enq_ready, writeQueueVec_6_enq_ready};
  wire [3:0]        otherUnit_vrfWritePort_ready_lo_hi = {otherUnit_vrfWritePort_ready_lo_hi_hi, otherUnit_vrfWritePort_ready_lo_hi_lo};
  wire [7:0]        otherUnit_vrfWritePort_ready_lo = {otherUnit_vrfWritePort_ready_lo_hi, otherUnit_vrfWritePort_ready_lo_lo};
  wire [1:0]        otherUnit_vrfWritePort_ready_hi_lo_lo = {writeQueueVec_9_enq_ready, writeQueueVec_8_enq_ready};
  wire [1:0]        otherUnit_vrfWritePort_ready_hi_lo_hi = {writeQueueVec_11_enq_ready, writeQueueVec_10_enq_ready};
  wire [3:0]        otherUnit_vrfWritePort_ready_hi_lo = {otherUnit_vrfWritePort_ready_hi_lo_hi, otherUnit_vrfWritePort_ready_hi_lo_lo};
  wire [1:0]        otherUnit_vrfWritePort_ready_hi_hi_lo = {writeQueueVec_13_enq_ready, writeQueueVec_12_enq_ready};
  wire [1:0]        otherUnit_vrfWritePort_ready_hi_hi_hi = {writeQueueVec_15_enq_ready, writeQueueVec_14_enq_ready};
  wire [3:0]        otherUnit_vrfWritePort_ready_hi_hi = {otherUnit_vrfWritePort_ready_hi_hi_hi, otherUnit_vrfWritePort_ready_hi_hi_lo};
  wire [7:0]        otherUnit_vrfWritePort_ready_hi = {otherUnit_vrfWritePort_ready_hi_hi, otherUnit_vrfWritePort_ready_hi_lo};
  assign writeQueueVec_0_enq_valid = otherTryToWrite[0] | _loadUnit_vrfWritePort_0_valid;
  assign writeQueueVec_0_enq_bits_data_vd = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_0_bits_vd;
  assign writeQueueVec_0_enq_bits_data_offset = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_0_bits_offset;
  assign writeQueueVec_0_enq_bits_data_mask = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_0_bits_mask;
  assign writeQueueVec_0_enq_bits_data_data = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_0_bits_data;
  assign writeQueueVec_0_enq_bits_data_last = otherTryToWrite[0] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_0_enq_bits_data_instructionIndex = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_0_bits_instructionIndex;
  assign writeQueueVec_1_enq_valid = otherTryToWrite[1] | _loadUnit_vrfWritePort_1_valid;
  assign writeQueueVec_1_enq_bits_data_vd = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_1_bits_vd;
  assign writeQueueVec_1_enq_bits_data_offset = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_1_bits_offset;
  assign writeQueueVec_1_enq_bits_data_mask = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_1_bits_mask;
  assign writeQueueVec_1_enq_bits_data_data = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_1_bits_data;
  assign writeQueueVec_1_enq_bits_data_last = otherTryToWrite[1] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_1_enq_bits_data_instructionIndex = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_1_bits_instructionIndex;
  assign writeQueueVec_2_enq_valid = otherTryToWrite[2] | _loadUnit_vrfWritePort_2_valid;
  assign writeQueueVec_2_enq_bits_data_vd = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_2_bits_vd;
  assign writeQueueVec_2_enq_bits_data_offset = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_2_bits_offset;
  assign writeQueueVec_2_enq_bits_data_mask = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_2_bits_mask;
  assign writeQueueVec_2_enq_bits_data_data = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_2_bits_data;
  assign writeQueueVec_2_enq_bits_data_last = otherTryToWrite[2] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_2_enq_bits_data_instructionIndex = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_2_bits_instructionIndex;
  assign writeQueueVec_3_enq_valid = otherTryToWrite[3] | _loadUnit_vrfWritePort_3_valid;
  assign writeQueueVec_3_enq_bits_data_vd = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_3_bits_vd;
  assign writeQueueVec_3_enq_bits_data_offset = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_3_bits_offset;
  assign writeQueueVec_3_enq_bits_data_mask = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_3_bits_mask;
  assign writeQueueVec_3_enq_bits_data_data = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_3_bits_data;
  assign writeQueueVec_3_enq_bits_data_last = otherTryToWrite[3] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_3_enq_bits_data_instructionIndex = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_3_bits_instructionIndex;
  assign writeQueueVec_4_enq_valid = otherTryToWrite[4] | _loadUnit_vrfWritePort_4_valid;
  assign writeQueueVec_4_enq_bits_data_vd = otherTryToWrite[4] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_4_bits_vd;
  assign writeQueueVec_4_enq_bits_data_offset = otherTryToWrite[4] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_4_bits_offset;
  assign writeQueueVec_4_enq_bits_data_mask = otherTryToWrite[4] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_4_bits_mask;
  assign writeQueueVec_4_enq_bits_data_data = otherTryToWrite[4] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_4_bits_data;
  assign writeQueueVec_4_enq_bits_data_last = otherTryToWrite[4] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_4_enq_bits_data_instructionIndex = otherTryToWrite[4] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_4_bits_instructionIndex;
  assign writeQueueVec_5_enq_valid = otherTryToWrite[5] | _loadUnit_vrfWritePort_5_valid;
  assign writeQueueVec_5_enq_bits_data_vd = otherTryToWrite[5] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_5_bits_vd;
  assign writeQueueVec_5_enq_bits_data_offset = otherTryToWrite[5] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_5_bits_offset;
  assign writeQueueVec_5_enq_bits_data_mask = otherTryToWrite[5] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_5_bits_mask;
  assign writeQueueVec_5_enq_bits_data_data = otherTryToWrite[5] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_5_bits_data;
  assign writeQueueVec_5_enq_bits_data_last = otherTryToWrite[5] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_5_enq_bits_data_instructionIndex = otherTryToWrite[5] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_5_bits_instructionIndex;
  assign writeQueueVec_6_enq_valid = otherTryToWrite[6] | _loadUnit_vrfWritePort_6_valid;
  assign writeQueueVec_6_enq_bits_data_vd = otherTryToWrite[6] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_6_bits_vd;
  assign writeQueueVec_6_enq_bits_data_offset = otherTryToWrite[6] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_6_bits_offset;
  assign writeQueueVec_6_enq_bits_data_mask = otherTryToWrite[6] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_6_bits_mask;
  assign writeQueueVec_6_enq_bits_data_data = otherTryToWrite[6] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_6_bits_data;
  assign writeQueueVec_6_enq_bits_data_last = otherTryToWrite[6] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_6_enq_bits_data_instructionIndex = otherTryToWrite[6] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_6_bits_instructionIndex;
  assign writeQueueVec_7_enq_valid = otherTryToWrite[7] | _loadUnit_vrfWritePort_7_valid;
  assign writeQueueVec_7_enq_bits_data_vd = otherTryToWrite[7] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_7_bits_vd;
  assign writeQueueVec_7_enq_bits_data_offset = otherTryToWrite[7] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_7_bits_offset;
  assign writeQueueVec_7_enq_bits_data_mask = otherTryToWrite[7] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_7_bits_mask;
  assign writeQueueVec_7_enq_bits_data_data = otherTryToWrite[7] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_7_bits_data;
  assign writeQueueVec_7_enq_bits_data_last = otherTryToWrite[7] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_7_enq_bits_data_instructionIndex = otherTryToWrite[7] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_7_bits_instructionIndex;
  assign writeQueueVec_8_enq_valid = otherTryToWrite[8] | _loadUnit_vrfWritePort_8_valid;
  assign writeQueueVec_8_enq_bits_data_vd = otherTryToWrite[8] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_8_bits_vd;
  assign writeQueueVec_8_enq_bits_data_offset = otherTryToWrite[8] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_8_bits_offset;
  assign writeQueueVec_8_enq_bits_data_mask = otherTryToWrite[8] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_8_bits_mask;
  assign writeQueueVec_8_enq_bits_data_data = otherTryToWrite[8] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_8_bits_data;
  assign writeQueueVec_8_enq_bits_data_last = otherTryToWrite[8] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_8_enq_bits_data_instructionIndex = otherTryToWrite[8] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_8_bits_instructionIndex;
  assign writeQueueVec_9_enq_valid = otherTryToWrite[9] | _loadUnit_vrfWritePort_9_valid;
  assign writeQueueVec_9_enq_bits_data_vd = otherTryToWrite[9] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_9_bits_vd;
  assign writeQueueVec_9_enq_bits_data_offset = otherTryToWrite[9] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_9_bits_offset;
  assign writeQueueVec_9_enq_bits_data_mask = otherTryToWrite[9] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_9_bits_mask;
  assign writeQueueVec_9_enq_bits_data_data = otherTryToWrite[9] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_9_bits_data;
  assign writeQueueVec_9_enq_bits_data_last = otherTryToWrite[9] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_9_enq_bits_data_instructionIndex = otherTryToWrite[9] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_9_bits_instructionIndex;
  assign writeQueueVec_10_enq_valid = otherTryToWrite[10] | _loadUnit_vrfWritePort_10_valid;
  assign writeQueueVec_10_enq_bits_data_vd = otherTryToWrite[10] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_10_bits_vd;
  assign writeQueueVec_10_enq_bits_data_offset = otherTryToWrite[10] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_10_bits_offset;
  assign writeQueueVec_10_enq_bits_data_mask = otherTryToWrite[10] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_10_bits_mask;
  assign writeQueueVec_10_enq_bits_data_data = otherTryToWrite[10] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_10_bits_data;
  assign writeQueueVec_10_enq_bits_data_last = otherTryToWrite[10] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_10_enq_bits_data_instructionIndex = otherTryToWrite[10] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_10_bits_instructionIndex;
  assign writeQueueVec_11_enq_valid = otherTryToWrite[11] | _loadUnit_vrfWritePort_11_valid;
  assign writeQueueVec_11_enq_bits_data_vd = otherTryToWrite[11] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_11_bits_vd;
  assign writeQueueVec_11_enq_bits_data_offset = otherTryToWrite[11] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_11_bits_offset;
  assign writeQueueVec_11_enq_bits_data_mask = otherTryToWrite[11] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_11_bits_mask;
  assign writeQueueVec_11_enq_bits_data_data = otherTryToWrite[11] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_11_bits_data;
  assign writeQueueVec_11_enq_bits_data_last = otherTryToWrite[11] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_11_enq_bits_data_instructionIndex = otherTryToWrite[11] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_11_bits_instructionIndex;
  assign writeQueueVec_12_enq_valid = otherTryToWrite[12] | _loadUnit_vrfWritePort_12_valid;
  assign writeQueueVec_12_enq_bits_data_vd = otherTryToWrite[12] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_12_bits_vd;
  assign writeQueueVec_12_enq_bits_data_offset = otherTryToWrite[12] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_12_bits_offset;
  assign writeQueueVec_12_enq_bits_data_mask = otherTryToWrite[12] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_12_bits_mask;
  assign writeQueueVec_12_enq_bits_data_data = otherTryToWrite[12] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_12_bits_data;
  assign writeQueueVec_12_enq_bits_data_last = otherTryToWrite[12] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_12_enq_bits_data_instructionIndex = otherTryToWrite[12] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_12_bits_instructionIndex;
  assign writeQueueVec_13_enq_valid = otherTryToWrite[13] | _loadUnit_vrfWritePort_13_valid;
  assign writeQueueVec_13_enq_bits_data_vd = otherTryToWrite[13] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_13_bits_vd;
  assign writeQueueVec_13_enq_bits_data_offset = otherTryToWrite[13] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_13_bits_offset;
  assign writeQueueVec_13_enq_bits_data_mask = otherTryToWrite[13] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_13_bits_mask;
  assign writeQueueVec_13_enq_bits_data_data = otherTryToWrite[13] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_13_bits_data;
  assign writeQueueVec_13_enq_bits_data_last = otherTryToWrite[13] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_13_enq_bits_data_instructionIndex = otherTryToWrite[13] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_13_bits_instructionIndex;
  assign writeQueueVec_14_enq_valid = otherTryToWrite[14] | _loadUnit_vrfWritePort_14_valid;
  assign writeQueueVec_14_enq_bits_data_vd = otherTryToWrite[14] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_14_bits_vd;
  assign writeQueueVec_14_enq_bits_data_offset = otherTryToWrite[14] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_14_bits_offset;
  assign writeQueueVec_14_enq_bits_data_mask = otherTryToWrite[14] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_14_bits_mask;
  assign writeQueueVec_14_enq_bits_data_data = otherTryToWrite[14] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_14_bits_data;
  assign writeQueueVec_14_enq_bits_data_last = otherTryToWrite[14] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_14_enq_bits_data_instructionIndex = otherTryToWrite[14] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_14_bits_instructionIndex;
  assign writeQueueVec_15_enq_valid = otherTryToWrite[15] | _loadUnit_vrfWritePort_15_valid;
  assign writeQueueVec_15_enq_bits_data_vd = otherTryToWrite[15] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_15_bits_vd;
  assign writeQueueVec_15_enq_bits_data_offset = otherTryToWrite[15] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_15_bits_offset;
  assign writeQueueVec_15_enq_bits_data_mask = otherTryToWrite[15] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_15_bits_mask;
  assign writeQueueVec_15_enq_bits_data_data = otherTryToWrite[15] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_15_bits_data;
  assign writeQueueVec_15_enq_bits_data_last = otherTryToWrite[15] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_15_enq_bits_data_instructionIndex = otherTryToWrite[15] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_15_bits_instructionIndex;
  wire [7:0]        _GEN_34 = {5'h0, _loadUnit_status_instructionIndex};
  wire [7:0]        _GEN_35 = {5'h0, _otherUnit_status_instructionIndex};
  wire [7:0]        dataInMSHR = (_loadUnit_status_idle ? 8'h0 : 8'h1 << _GEN_34) | (_otherUnit_status_idle | _otherUnit_status_isStore ? 8'h0 : 8'h1 << _GEN_35);
  reg  [6:0]        queueCount_0;
  reg  [6:0]        queueCount_1;
  reg  [6:0]        queueCount_2;
  reg  [6:0]        queueCount_3;
  reg  [6:0]        queueCount_4;
  reg  [6:0]        queueCount_5;
  reg  [6:0]        queueCount_6;
  reg  [6:0]        queueCount_7;
  wire [7:0]        enqOH = 8'h1 << writeQueueVec_0_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq = _probeWire_slots_0_writeValid_T ? enqOH : 8'h0;
  wire              writeIndexQueue_deq_valid;
  assign writeIndexQueue_deq_valid = ~_writeIndexQueue_fifo_empty;
  wire              writeIndexQueue_enq_ready = ~_writeIndexQueue_fifo_full;
  wire              writeIndexQueue_enq_valid;
  assign writeIndexQueue_enq_valid = writeQueueVec_0_deq_ready & writeQueueVec_0_deq_valid;
  wire [2:0]        writeIndexQueue_deq_bits;
  wire [7:0]        queueDeq = writeIndexQueue_deq_ready & writeIndexQueue_deq_valid ? 8'h1 << writeIndexQueue_deq_bits : 8'h0;
  wire [6:0]        counterUpdate = queueEnq[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_1 = queueEnq[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_2 = queueEnq[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_3 = queueEnq[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_4 = queueEnq[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_5 = queueEnq[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_6 = queueEnq[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_7 = queueEnq[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_0_lo_lo = {|queueCount_1, |queueCount_0};
  wire [1:0]        dataInWriteQueue_0_lo_hi = {|queueCount_3, |queueCount_2};
  wire [3:0]        dataInWriteQueue_0_lo = {dataInWriteQueue_0_lo_hi, dataInWriteQueue_0_lo_lo};
  wire [1:0]        dataInWriteQueue_0_hi_lo = {|queueCount_5, |queueCount_4};
  wire [1:0]        dataInWriteQueue_0_hi_hi = {|queueCount_7, |queueCount_6};
  wire [3:0]        dataInWriteQueue_0_hi = {dataInWriteQueue_0_hi_hi, dataInWriteQueue_0_hi_lo};
  reg  [6:0]        queueCount_0_1;
  reg  [6:0]        queueCount_1_1;
  reg  [6:0]        queueCount_2_1;
  reg  [6:0]        queueCount_3_1;
  reg  [6:0]        queueCount_4_1;
  reg  [6:0]        queueCount_5_1;
  reg  [6:0]        queueCount_6_1;
  reg  [6:0]        queueCount_7_1;
  wire [7:0]        enqOH_1 = 8'h1 << writeQueueVec_1_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_1 = _probeWire_slots_1_writeValid_T ? enqOH_1 : 8'h0;
  wire              writeIndexQueue_1_deq_valid;
  assign writeIndexQueue_1_deq_valid = ~_writeIndexQueue_fifo_1_empty;
  wire              writeIndexQueue_1_enq_ready = ~_writeIndexQueue_fifo_1_full;
  wire              writeIndexQueue_1_enq_valid;
  assign writeIndexQueue_1_enq_valid = writeQueueVec_1_deq_ready & writeQueueVec_1_deq_valid;
  wire [2:0]        writeIndexQueue_1_deq_bits;
  wire [7:0]        queueDeq_1 = writeIndexQueue_1_deq_ready & writeIndexQueue_1_deq_valid ? 8'h1 << writeIndexQueue_1_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_8 = queueEnq_1[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_9 = queueEnq_1[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_10 = queueEnq_1[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_11 = queueEnq_1[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_12 = queueEnq_1[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_13 = queueEnq_1[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_14 = queueEnq_1[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_15 = queueEnq_1[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_1_lo_lo = {|queueCount_1_1, |queueCount_0_1};
  wire [1:0]        dataInWriteQueue_1_lo_hi = {|queueCount_3_1, |queueCount_2_1};
  wire [3:0]        dataInWriteQueue_1_lo = {dataInWriteQueue_1_lo_hi, dataInWriteQueue_1_lo_lo};
  wire [1:0]        dataInWriteQueue_1_hi_lo = {|queueCount_5_1, |queueCount_4_1};
  wire [1:0]        dataInWriteQueue_1_hi_hi = {|queueCount_7_1, |queueCount_6_1};
  wire [3:0]        dataInWriteQueue_1_hi = {dataInWriteQueue_1_hi_hi, dataInWriteQueue_1_hi_lo};
  reg  [6:0]        queueCount_0_2;
  reg  [6:0]        queueCount_1_2;
  reg  [6:0]        queueCount_2_2;
  reg  [6:0]        queueCount_3_2;
  reg  [6:0]        queueCount_4_2;
  reg  [6:0]        queueCount_5_2;
  reg  [6:0]        queueCount_6_2;
  reg  [6:0]        queueCount_7_2;
  wire [7:0]        enqOH_2 = 8'h1 << writeQueueVec_2_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_2 = _probeWire_slots_2_writeValid_T ? enqOH_2 : 8'h0;
  wire              writeIndexQueue_2_deq_valid;
  assign writeIndexQueue_2_deq_valid = ~_writeIndexQueue_fifo_2_empty;
  wire              writeIndexQueue_2_enq_ready = ~_writeIndexQueue_fifo_2_full;
  wire              writeIndexQueue_2_enq_valid;
  assign writeIndexQueue_2_enq_valid = writeQueueVec_2_deq_ready & writeQueueVec_2_deq_valid;
  wire [2:0]        writeIndexQueue_2_deq_bits;
  wire [7:0]        queueDeq_2 = writeIndexQueue_2_deq_ready & writeIndexQueue_2_deq_valid ? 8'h1 << writeIndexQueue_2_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_16 = queueEnq_2[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_17 = queueEnq_2[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_18 = queueEnq_2[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_19 = queueEnq_2[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_20 = queueEnq_2[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_21 = queueEnq_2[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_22 = queueEnq_2[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_23 = queueEnq_2[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_2_lo_lo = {|queueCount_1_2, |queueCount_0_2};
  wire [1:0]        dataInWriteQueue_2_lo_hi = {|queueCount_3_2, |queueCount_2_2};
  wire [3:0]        dataInWriteQueue_2_lo = {dataInWriteQueue_2_lo_hi, dataInWriteQueue_2_lo_lo};
  wire [1:0]        dataInWriteQueue_2_hi_lo = {|queueCount_5_2, |queueCount_4_2};
  wire [1:0]        dataInWriteQueue_2_hi_hi = {|queueCount_7_2, |queueCount_6_2};
  wire [3:0]        dataInWriteQueue_2_hi = {dataInWriteQueue_2_hi_hi, dataInWriteQueue_2_hi_lo};
  reg  [6:0]        queueCount_0_3;
  reg  [6:0]        queueCount_1_3;
  reg  [6:0]        queueCount_2_3;
  reg  [6:0]        queueCount_3_3;
  reg  [6:0]        queueCount_4_3;
  reg  [6:0]        queueCount_5_3;
  reg  [6:0]        queueCount_6_3;
  reg  [6:0]        queueCount_7_3;
  wire [7:0]        enqOH_3 = 8'h1 << writeQueueVec_3_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_3 = _probeWire_slots_3_writeValid_T ? enqOH_3 : 8'h0;
  wire              writeIndexQueue_3_deq_valid;
  assign writeIndexQueue_3_deq_valid = ~_writeIndexQueue_fifo_3_empty;
  wire              writeIndexQueue_3_enq_ready = ~_writeIndexQueue_fifo_3_full;
  wire              writeIndexQueue_3_enq_valid;
  assign writeIndexQueue_3_enq_valid = writeQueueVec_3_deq_ready & writeQueueVec_3_deq_valid;
  wire [2:0]        writeIndexQueue_3_deq_bits;
  wire [7:0]        queueDeq_3 = writeIndexQueue_3_deq_ready & writeIndexQueue_3_deq_valid ? 8'h1 << writeIndexQueue_3_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_24 = queueEnq_3[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_25 = queueEnq_3[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_26 = queueEnq_3[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_27 = queueEnq_3[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_28 = queueEnq_3[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_29 = queueEnq_3[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_30 = queueEnq_3[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_31 = queueEnq_3[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_3_lo_lo = {|queueCount_1_3, |queueCount_0_3};
  wire [1:0]        dataInWriteQueue_3_lo_hi = {|queueCount_3_3, |queueCount_2_3};
  wire [3:0]        dataInWriteQueue_3_lo = {dataInWriteQueue_3_lo_hi, dataInWriteQueue_3_lo_lo};
  wire [1:0]        dataInWriteQueue_3_hi_lo = {|queueCount_5_3, |queueCount_4_3};
  wire [1:0]        dataInWriteQueue_3_hi_hi = {|queueCount_7_3, |queueCount_6_3};
  wire [3:0]        dataInWriteQueue_3_hi = {dataInWriteQueue_3_hi_hi, dataInWriteQueue_3_hi_lo};
  reg  [6:0]        queueCount_0_4;
  reg  [6:0]        queueCount_1_4;
  reg  [6:0]        queueCount_2_4;
  reg  [6:0]        queueCount_3_4;
  reg  [6:0]        queueCount_4_4;
  reg  [6:0]        queueCount_5_4;
  reg  [6:0]        queueCount_6_4;
  reg  [6:0]        queueCount_7_4;
  wire [7:0]        enqOH_4 = 8'h1 << writeQueueVec_4_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_4 = _probeWire_slots_4_writeValid_T ? enqOH_4 : 8'h0;
  wire              writeIndexQueue_4_deq_valid;
  assign writeIndexQueue_4_deq_valid = ~_writeIndexQueue_fifo_4_empty;
  wire              writeIndexQueue_4_enq_ready = ~_writeIndexQueue_fifo_4_full;
  wire              writeIndexQueue_4_enq_valid;
  assign writeIndexQueue_4_enq_valid = writeQueueVec_4_deq_ready & writeQueueVec_4_deq_valid;
  wire [2:0]        writeIndexQueue_4_deq_bits;
  wire [7:0]        queueDeq_4 = writeIndexQueue_4_deq_ready & writeIndexQueue_4_deq_valid ? 8'h1 << writeIndexQueue_4_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_32 = queueEnq_4[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_33 = queueEnq_4[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_34 = queueEnq_4[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_35 = queueEnq_4[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_36 = queueEnq_4[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_37 = queueEnq_4[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_38 = queueEnq_4[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_39 = queueEnq_4[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_4_lo_lo = {|queueCount_1_4, |queueCount_0_4};
  wire [1:0]        dataInWriteQueue_4_lo_hi = {|queueCount_3_4, |queueCount_2_4};
  wire [3:0]        dataInWriteQueue_4_lo = {dataInWriteQueue_4_lo_hi, dataInWriteQueue_4_lo_lo};
  wire [1:0]        dataInWriteQueue_4_hi_lo = {|queueCount_5_4, |queueCount_4_4};
  wire [1:0]        dataInWriteQueue_4_hi_hi = {|queueCount_7_4, |queueCount_6_4};
  wire [3:0]        dataInWriteQueue_4_hi = {dataInWriteQueue_4_hi_hi, dataInWriteQueue_4_hi_lo};
  reg  [6:0]        queueCount_0_5;
  reg  [6:0]        queueCount_1_5;
  reg  [6:0]        queueCount_2_5;
  reg  [6:0]        queueCount_3_5;
  reg  [6:0]        queueCount_4_5;
  reg  [6:0]        queueCount_5_5;
  reg  [6:0]        queueCount_6_5;
  reg  [6:0]        queueCount_7_5;
  wire [7:0]        enqOH_5 = 8'h1 << writeQueueVec_5_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_5 = _probeWire_slots_5_writeValid_T ? enqOH_5 : 8'h0;
  wire              writeIndexQueue_5_deq_valid;
  assign writeIndexQueue_5_deq_valid = ~_writeIndexQueue_fifo_5_empty;
  wire              writeIndexQueue_5_enq_ready = ~_writeIndexQueue_fifo_5_full;
  wire              writeIndexQueue_5_enq_valid;
  assign writeIndexQueue_5_enq_valid = writeQueueVec_5_deq_ready & writeQueueVec_5_deq_valid;
  wire [2:0]        writeIndexQueue_5_deq_bits;
  wire [7:0]        queueDeq_5 = writeIndexQueue_5_deq_ready & writeIndexQueue_5_deq_valid ? 8'h1 << writeIndexQueue_5_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_40 = queueEnq_5[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_41 = queueEnq_5[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_42 = queueEnq_5[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_43 = queueEnq_5[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_44 = queueEnq_5[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_45 = queueEnq_5[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_46 = queueEnq_5[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_47 = queueEnq_5[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_5_lo_lo = {|queueCount_1_5, |queueCount_0_5};
  wire [1:0]        dataInWriteQueue_5_lo_hi = {|queueCount_3_5, |queueCount_2_5};
  wire [3:0]        dataInWriteQueue_5_lo = {dataInWriteQueue_5_lo_hi, dataInWriteQueue_5_lo_lo};
  wire [1:0]        dataInWriteQueue_5_hi_lo = {|queueCount_5_5, |queueCount_4_5};
  wire [1:0]        dataInWriteQueue_5_hi_hi = {|queueCount_7_5, |queueCount_6_5};
  wire [3:0]        dataInWriteQueue_5_hi = {dataInWriteQueue_5_hi_hi, dataInWriteQueue_5_hi_lo};
  reg  [6:0]        queueCount_0_6;
  reg  [6:0]        queueCount_1_6;
  reg  [6:0]        queueCount_2_6;
  reg  [6:0]        queueCount_3_6;
  reg  [6:0]        queueCount_4_6;
  reg  [6:0]        queueCount_5_6;
  reg  [6:0]        queueCount_6_6;
  reg  [6:0]        queueCount_7_6;
  wire [7:0]        enqOH_6 = 8'h1 << writeQueueVec_6_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_6 = _probeWire_slots_6_writeValid_T ? enqOH_6 : 8'h0;
  wire              writeIndexQueue_6_deq_valid;
  assign writeIndexQueue_6_deq_valid = ~_writeIndexQueue_fifo_6_empty;
  wire              writeIndexQueue_6_enq_ready = ~_writeIndexQueue_fifo_6_full;
  wire              writeIndexQueue_6_enq_valid;
  assign writeIndexQueue_6_enq_valid = writeQueueVec_6_deq_ready & writeQueueVec_6_deq_valid;
  wire [2:0]        writeIndexQueue_6_deq_bits;
  wire [7:0]        queueDeq_6 = writeIndexQueue_6_deq_ready & writeIndexQueue_6_deq_valid ? 8'h1 << writeIndexQueue_6_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_48 = queueEnq_6[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_49 = queueEnq_6[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_50 = queueEnq_6[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_51 = queueEnq_6[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_52 = queueEnq_6[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_53 = queueEnq_6[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_54 = queueEnq_6[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_55 = queueEnq_6[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_6_lo_lo = {|queueCount_1_6, |queueCount_0_6};
  wire [1:0]        dataInWriteQueue_6_lo_hi = {|queueCount_3_6, |queueCount_2_6};
  wire [3:0]        dataInWriteQueue_6_lo = {dataInWriteQueue_6_lo_hi, dataInWriteQueue_6_lo_lo};
  wire [1:0]        dataInWriteQueue_6_hi_lo = {|queueCount_5_6, |queueCount_4_6};
  wire [1:0]        dataInWriteQueue_6_hi_hi = {|queueCount_7_6, |queueCount_6_6};
  wire [3:0]        dataInWriteQueue_6_hi = {dataInWriteQueue_6_hi_hi, dataInWriteQueue_6_hi_lo};
  reg  [6:0]        queueCount_0_7;
  reg  [6:0]        queueCount_1_7;
  reg  [6:0]        queueCount_2_7;
  reg  [6:0]        queueCount_3_7;
  reg  [6:0]        queueCount_4_7;
  reg  [6:0]        queueCount_5_7;
  reg  [6:0]        queueCount_6_7;
  reg  [6:0]        queueCount_7_7;
  wire [7:0]        enqOH_7 = 8'h1 << writeQueueVec_7_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_7 = _probeWire_slots_7_writeValid_T ? enqOH_7 : 8'h0;
  wire              writeIndexQueue_7_deq_valid;
  assign writeIndexQueue_7_deq_valid = ~_writeIndexQueue_fifo_7_empty;
  wire              writeIndexQueue_7_enq_ready = ~_writeIndexQueue_fifo_7_full;
  wire              writeIndexQueue_7_enq_valid;
  assign writeIndexQueue_7_enq_valid = writeQueueVec_7_deq_ready & writeQueueVec_7_deq_valid;
  wire [2:0]        writeIndexQueue_7_deq_bits;
  wire [7:0]        queueDeq_7 = writeIndexQueue_7_deq_ready & writeIndexQueue_7_deq_valid ? 8'h1 << writeIndexQueue_7_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_56 = queueEnq_7[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_57 = queueEnq_7[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_58 = queueEnq_7[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_59 = queueEnq_7[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_60 = queueEnq_7[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_61 = queueEnq_7[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_62 = queueEnq_7[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_63 = queueEnq_7[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_7_lo_lo = {|queueCount_1_7, |queueCount_0_7};
  wire [1:0]        dataInWriteQueue_7_lo_hi = {|queueCount_3_7, |queueCount_2_7};
  wire [3:0]        dataInWriteQueue_7_lo = {dataInWriteQueue_7_lo_hi, dataInWriteQueue_7_lo_lo};
  wire [1:0]        dataInWriteQueue_7_hi_lo = {|queueCount_5_7, |queueCount_4_7};
  wire [1:0]        dataInWriteQueue_7_hi_hi = {|queueCount_7_7, |queueCount_6_7};
  wire [3:0]        dataInWriteQueue_7_hi = {dataInWriteQueue_7_hi_hi, dataInWriteQueue_7_hi_lo};
  reg  [6:0]        queueCount_0_8;
  reg  [6:0]        queueCount_1_8;
  reg  [6:0]        queueCount_2_8;
  reg  [6:0]        queueCount_3_8;
  reg  [6:0]        queueCount_4_8;
  reg  [6:0]        queueCount_5_8;
  reg  [6:0]        queueCount_6_8;
  reg  [6:0]        queueCount_7_8;
  wire [7:0]        enqOH_8 = 8'h1 << writeQueueVec_8_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_8 = _probeWire_slots_8_writeValid_T ? enqOH_8 : 8'h0;
  wire              writeIndexQueue_8_deq_valid;
  assign writeIndexQueue_8_deq_valid = ~_writeIndexQueue_fifo_8_empty;
  wire              writeIndexQueue_8_enq_ready = ~_writeIndexQueue_fifo_8_full;
  wire              writeIndexQueue_8_enq_valid;
  assign writeIndexQueue_8_enq_valid = writeQueueVec_8_deq_ready & writeQueueVec_8_deq_valid;
  wire [2:0]        writeIndexQueue_8_deq_bits;
  wire [7:0]        queueDeq_8 = writeIndexQueue_8_deq_ready & writeIndexQueue_8_deq_valid ? 8'h1 << writeIndexQueue_8_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_64 = queueEnq_8[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_65 = queueEnq_8[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_66 = queueEnq_8[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_67 = queueEnq_8[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_68 = queueEnq_8[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_69 = queueEnq_8[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_70 = queueEnq_8[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_71 = queueEnq_8[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_8_lo_lo = {|queueCount_1_8, |queueCount_0_8};
  wire [1:0]        dataInWriteQueue_8_lo_hi = {|queueCount_3_8, |queueCount_2_8};
  wire [3:0]        dataInWriteQueue_8_lo = {dataInWriteQueue_8_lo_hi, dataInWriteQueue_8_lo_lo};
  wire [1:0]        dataInWriteQueue_8_hi_lo = {|queueCount_5_8, |queueCount_4_8};
  wire [1:0]        dataInWriteQueue_8_hi_hi = {|queueCount_7_8, |queueCount_6_8};
  wire [3:0]        dataInWriteQueue_8_hi = {dataInWriteQueue_8_hi_hi, dataInWriteQueue_8_hi_lo};
  reg  [6:0]        queueCount_0_9;
  reg  [6:0]        queueCount_1_9;
  reg  [6:0]        queueCount_2_9;
  reg  [6:0]        queueCount_3_9;
  reg  [6:0]        queueCount_4_9;
  reg  [6:0]        queueCount_5_9;
  reg  [6:0]        queueCount_6_9;
  reg  [6:0]        queueCount_7_9;
  wire [7:0]        enqOH_9 = 8'h1 << writeQueueVec_9_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_9 = _probeWire_slots_9_writeValid_T ? enqOH_9 : 8'h0;
  wire              writeIndexQueue_9_deq_valid;
  assign writeIndexQueue_9_deq_valid = ~_writeIndexQueue_fifo_9_empty;
  wire              writeIndexQueue_9_enq_ready = ~_writeIndexQueue_fifo_9_full;
  wire              writeIndexQueue_9_enq_valid;
  assign writeIndexQueue_9_enq_valid = writeQueueVec_9_deq_ready & writeQueueVec_9_deq_valid;
  wire [2:0]        writeIndexQueue_9_deq_bits;
  wire [7:0]        queueDeq_9 = writeIndexQueue_9_deq_ready & writeIndexQueue_9_deq_valid ? 8'h1 << writeIndexQueue_9_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_72 = queueEnq_9[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_73 = queueEnq_9[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_74 = queueEnq_9[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_75 = queueEnq_9[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_76 = queueEnq_9[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_77 = queueEnq_9[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_78 = queueEnq_9[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_79 = queueEnq_9[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_9_lo_lo = {|queueCount_1_9, |queueCount_0_9};
  wire [1:0]        dataInWriteQueue_9_lo_hi = {|queueCount_3_9, |queueCount_2_9};
  wire [3:0]        dataInWriteQueue_9_lo = {dataInWriteQueue_9_lo_hi, dataInWriteQueue_9_lo_lo};
  wire [1:0]        dataInWriteQueue_9_hi_lo = {|queueCount_5_9, |queueCount_4_9};
  wire [1:0]        dataInWriteQueue_9_hi_hi = {|queueCount_7_9, |queueCount_6_9};
  wire [3:0]        dataInWriteQueue_9_hi = {dataInWriteQueue_9_hi_hi, dataInWriteQueue_9_hi_lo};
  reg  [6:0]        queueCount_0_10;
  reg  [6:0]        queueCount_1_10;
  reg  [6:0]        queueCount_2_10;
  reg  [6:0]        queueCount_3_10;
  reg  [6:0]        queueCount_4_10;
  reg  [6:0]        queueCount_5_10;
  reg  [6:0]        queueCount_6_10;
  reg  [6:0]        queueCount_7_10;
  wire [7:0]        enqOH_10 = 8'h1 << writeQueueVec_10_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_10 = _probeWire_slots_10_writeValid_T ? enqOH_10 : 8'h0;
  wire              writeIndexQueue_10_deq_valid;
  assign writeIndexQueue_10_deq_valid = ~_writeIndexQueue_fifo_10_empty;
  wire              writeIndexQueue_10_enq_ready = ~_writeIndexQueue_fifo_10_full;
  wire              writeIndexQueue_10_enq_valid;
  assign writeIndexQueue_10_enq_valid = writeQueueVec_10_deq_ready & writeQueueVec_10_deq_valid;
  wire [2:0]        writeIndexQueue_10_deq_bits;
  wire [7:0]        queueDeq_10 = writeIndexQueue_10_deq_ready & writeIndexQueue_10_deq_valid ? 8'h1 << writeIndexQueue_10_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_80 = queueEnq_10[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_81 = queueEnq_10[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_82 = queueEnq_10[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_83 = queueEnq_10[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_84 = queueEnq_10[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_85 = queueEnq_10[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_86 = queueEnq_10[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_87 = queueEnq_10[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_10_lo_lo = {|queueCount_1_10, |queueCount_0_10};
  wire [1:0]        dataInWriteQueue_10_lo_hi = {|queueCount_3_10, |queueCount_2_10};
  wire [3:0]        dataInWriteQueue_10_lo = {dataInWriteQueue_10_lo_hi, dataInWriteQueue_10_lo_lo};
  wire [1:0]        dataInWriteQueue_10_hi_lo = {|queueCount_5_10, |queueCount_4_10};
  wire [1:0]        dataInWriteQueue_10_hi_hi = {|queueCount_7_10, |queueCount_6_10};
  wire [3:0]        dataInWriteQueue_10_hi = {dataInWriteQueue_10_hi_hi, dataInWriteQueue_10_hi_lo};
  reg  [6:0]        queueCount_0_11;
  reg  [6:0]        queueCount_1_11;
  reg  [6:0]        queueCount_2_11;
  reg  [6:0]        queueCount_3_11;
  reg  [6:0]        queueCount_4_11;
  reg  [6:0]        queueCount_5_11;
  reg  [6:0]        queueCount_6_11;
  reg  [6:0]        queueCount_7_11;
  wire [7:0]        enqOH_11 = 8'h1 << writeQueueVec_11_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_11 = _probeWire_slots_11_writeValid_T ? enqOH_11 : 8'h0;
  wire              writeIndexQueue_11_deq_valid;
  assign writeIndexQueue_11_deq_valid = ~_writeIndexQueue_fifo_11_empty;
  wire              writeIndexQueue_11_enq_ready = ~_writeIndexQueue_fifo_11_full;
  wire              writeIndexQueue_11_enq_valid;
  assign writeIndexQueue_11_enq_valid = writeQueueVec_11_deq_ready & writeQueueVec_11_deq_valid;
  wire [2:0]        writeIndexQueue_11_deq_bits;
  wire [7:0]        queueDeq_11 = writeIndexQueue_11_deq_ready & writeIndexQueue_11_deq_valid ? 8'h1 << writeIndexQueue_11_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_88 = queueEnq_11[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_89 = queueEnq_11[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_90 = queueEnq_11[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_91 = queueEnq_11[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_92 = queueEnq_11[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_93 = queueEnq_11[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_94 = queueEnq_11[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_95 = queueEnq_11[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_11_lo_lo = {|queueCount_1_11, |queueCount_0_11};
  wire [1:0]        dataInWriteQueue_11_lo_hi = {|queueCount_3_11, |queueCount_2_11};
  wire [3:0]        dataInWriteQueue_11_lo = {dataInWriteQueue_11_lo_hi, dataInWriteQueue_11_lo_lo};
  wire [1:0]        dataInWriteQueue_11_hi_lo = {|queueCount_5_11, |queueCount_4_11};
  wire [1:0]        dataInWriteQueue_11_hi_hi = {|queueCount_7_11, |queueCount_6_11};
  wire [3:0]        dataInWriteQueue_11_hi = {dataInWriteQueue_11_hi_hi, dataInWriteQueue_11_hi_lo};
  reg  [6:0]        queueCount_0_12;
  reg  [6:0]        queueCount_1_12;
  reg  [6:0]        queueCount_2_12;
  reg  [6:0]        queueCount_3_12;
  reg  [6:0]        queueCount_4_12;
  reg  [6:0]        queueCount_5_12;
  reg  [6:0]        queueCount_6_12;
  reg  [6:0]        queueCount_7_12;
  wire [7:0]        enqOH_12 = 8'h1 << writeQueueVec_12_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_12 = _probeWire_slots_12_writeValid_T ? enqOH_12 : 8'h0;
  wire              writeIndexQueue_12_deq_valid;
  assign writeIndexQueue_12_deq_valid = ~_writeIndexQueue_fifo_12_empty;
  wire              writeIndexQueue_12_enq_ready = ~_writeIndexQueue_fifo_12_full;
  wire              writeIndexQueue_12_enq_valid;
  assign writeIndexQueue_12_enq_valid = writeQueueVec_12_deq_ready & writeQueueVec_12_deq_valid;
  wire [2:0]        writeIndexQueue_12_deq_bits;
  wire [7:0]        queueDeq_12 = writeIndexQueue_12_deq_ready & writeIndexQueue_12_deq_valid ? 8'h1 << writeIndexQueue_12_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_96 = queueEnq_12[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_97 = queueEnq_12[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_98 = queueEnq_12[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_99 = queueEnq_12[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_100 = queueEnq_12[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_101 = queueEnq_12[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_102 = queueEnq_12[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_103 = queueEnq_12[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_12_lo_lo = {|queueCount_1_12, |queueCount_0_12};
  wire [1:0]        dataInWriteQueue_12_lo_hi = {|queueCount_3_12, |queueCount_2_12};
  wire [3:0]        dataInWriteQueue_12_lo = {dataInWriteQueue_12_lo_hi, dataInWriteQueue_12_lo_lo};
  wire [1:0]        dataInWriteQueue_12_hi_lo = {|queueCount_5_12, |queueCount_4_12};
  wire [1:0]        dataInWriteQueue_12_hi_hi = {|queueCount_7_12, |queueCount_6_12};
  wire [3:0]        dataInWriteQueue_12_hi = {dataInWriteQueue_12_hi_hi, dataInWriteQueue_12_hi_lo};
  reg  [6:0]        queueCount_0_13;
  reg  [6:0]        queueCount_1_13;
  reg  [6:0]        queueCount_2_13;
  reg  [6:0]        queueCount_3_13;
  reg  [6:0]        queueCount_4_13;
  reg  [6:0]        queueCount_5_13;
  reg  [6:0]        queueCount_6_13;
  reg  [6:0]        queueCount_7_13;
  wire [7:0]        enqOH_13 = 8'h1 << writeQueueVec_13_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_13 = _probeWire_slots_13_writeValid_T ? enqOH_13 : 8'h0;
  wire              writeIndexQueue_13_deq_valid;
  assign writeIndexQueue_13_deq_valid = ~_writeIndexQueue_fifo_13_empty;
  wire              writeIndexQueue_13_enq_ready = ~_writeIndexQueue_fifo_13_full;
  wire              writeIndexQueue_13_enq_valid;
  assign writeIndexQueue_13_enq_valid = writeQueueVec_13_deq_ready & writeQueueVec_13_deq_valid;
  wire [2:0]        writeIndexQueue_13_deq_bits;
  wire [7:0]        queueDeq_13 = writeIndexQueue_13_deq_ready & writeIndexQueue_13_deq_valid ? 8'h1 << writeIndexQueue_13_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_104 = queueEnq_13[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_105 = queueEnq_13[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_106 = queueEnq_13[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_107 = queueEnq_13[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_108 = queueEnq_13[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_109 = queueEnq_13[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_110 = queueEnq_13[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_111 = queueEnq_13[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_13_lo_lo = {|queueCount_1_13, |queueCount_0_13};
  wire [1:0]        dataInWriteQueue_13_lo_hi = {|queueCount_3_13, |queueCount_2_13};
  wire [3:0]        dataInWriteQueue_13_lo = {dataInWriteQueue_13_lo_hi, dataInWriteQueue_13_lo_lo};
  wire [1:0]        dataInWriteQueue_13_hi_lo = {|queueCount_5_13, |queueCount_4_13};
  wire [1:0]        dataInWriteQueue_13_hi_hi = {|queueCount_7_13, |queueCount_6_13};
  wire [3:0]        dataInWriteQueue_13_hi = {dataInWriteQueue_13_hi_hi, dataInWriteQueue_13_hi_lo};
  reg  [6:0]        queueCount_0_14;
  reg  [6:0]        queueCount_1_14;
  reg  [6:0]        queueCount_2_14;
  reg  [6:0]        queueCount_3_14;
  reg  [6:0]        queueCount_4_14;
  reg  [6:0]        queueCount_5_14;
  reg  [6:0]        queueCount_6_14;
  reg  [6:0]        queueCount_7_14;
  wire [7:0]        enqOH_14 = 8'h1 << writeQueueVec_14_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_14 = _probeWire_slots_14_writeValid_T ? enqOH_14 : 8'h0;
  wire              writeIndexQueue_14_deq_valid;
  assign writeIndexQueue_14_deq_valid = ~_writeIndexQueue_fifo_14_empty;
  wire              writeIndexQueue_14_enq_ready = ~_writeIndexQueue_fifo_14_full;
  wire              writeIndexQueue_14_enq_valid;
  assign writeIndexQueue_14_enq_valid = writeQueueVec_14_deq_ready & writeQueueVec_14_deq_valid;
  wire [2:0]        writeIndexQueue_14_deq_bits;
  wire [7:0]        queueDeq_14 = writeIndexQueue_14_deq_ready & writeIndexQueue_14_deq_valid ? 8'h1 << writeIndexQueue_14_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_112 = queueEnq_14[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_113 = queueEnq_14[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_114 = queueEnq_14[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_115 = queueEnq_14[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_116 = queueEnq_14[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_117 = queueEnq_14[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_118 = queueEnq_14[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_119 = queueEnq_14[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_14_lo_lo = {|queueCount_1_14, |queueCount_0_14};
  wire [1:0]        dataInWriteQueue_14_lo_hi = {|queueCount_3_14, |queueCount_2_14};
  wire [3:0]        dataInWriteQueue_14_lo = {dataInWriteQueue_14_lo_hi, dataInWriteQueue_14_lo_lo};
  wire [1:0]        dataInWriteQueue_14_hi_lo = {|queueCount_5_14, |queueCount_4_14};
  wire [1:0]        dataInWriteQueue_14_hi_hi = {|queueCount_7_14, |queueCount_6_14};
  wire [3:0]        dataInWriteQueue_14_hi = {dataInWriteQueue_14_hi_hi, dataInWriteQueue_14_hi_lo};
  reg  [6:0]        queueCount_0_15;
  reg  [6:0]        queueCount_1_15;
  reg  [6:0]        queueCount_2_15;
  reg  [6:0]        queueCount_3_15;
  reg  [6:0]        queueCount_4_15;
  reg  [6:0]        queueCount_5_15;
  reg  [6:0]        queueCount_6_15;
  reg  [6:0]        queueCount_7_15;
  wire [7:0]        enqOH_15 = 8'h1 << writeQueueVec_15_enq_bits_data_instructionIndex;
  wire [7:0]        queueEnq_15 = _probeWire_slots_15_writeValid_T ? enqOH_15 : 8'h0;
  wire              writeIndexQueue_15_deq_valid;
  assign writeIndexQueue_15_deq_valid = ~_writeIndexQueue_fifo_15_empty;
  wire              writeIndexQueue_15_enq_ready = ~_writeIndexQueue_fifo_15_full;
  wire              writeIndexQueue_15_enq_valid;
  assign writeIndexQueue_15_enq_valid = writeQueueVec_15_deq_ready & writeQueueVec_15_deq_valid;
  wire [2:0]        writeIndexQueue_15_deq_bits;
  wire [7:0]        queueDeq_15 = writeIndexQueue_15_deq_ready & writeIndexQueue_15_deq_valid ? 8'h1 << writeIndexQueue_15_deq_bits : 8'h0;
  wire [6:0]        counterUpdate_120 = queueEnq_15[0] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_121 = queueEnq_15[1] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_122 = queueEnq_15[2] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_123 = queueEnq_15[3] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_124 = queueEnq_15[4] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_125 = queueEnq_15[5] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_126 = queueEnq_15[6] ? 7'h1 : 7'h7F;
  wire [6:0]        counterUpdate_127 = queueEnq_15[7] ? 7'h1 : 7'h7F;
  wire [1:0]        dataInWriteQueue_15_lo_lo = {|queueCount_1_15, |queueCount_0_15};
  wire [1:0]        dataInWriteQueue_15_lo_hi = {|queueCount_3_15, |queueCount_2_15};
  wire [3:0]        dataInWriteQueue_15_lo = {dataInWriteQueue_15_lo_hi, dataInWriteQueue_15_lo_lo};
  wire [1:0]        dataInWriteQueue_15_hi_lo = {|queueCount_5_15, |queueCount_4_15};
  wire [1:0]        dataInWriteQueue_15_hi_hi = {|queueCount_7_15, |queueCount_6_15};
  wire [3:0]        dataInWriteQueue_15_hi = {dataInWriteQueue_15_hi_hi, dataInWriteQueue_15_hi_lo};
  wire              sourceQueue_deq_valid;
  assign sourceQueue_deq_valid = ~_sourceQueue_fifo_empty;
  wire              sourceQueue_enq_ready = ~_sourceQueue_fifo_full;
  wire              sourceQueue_enq_valid;
  wire              sourceQueue_deq_ready;
  wire              axi4Port_ar_valid_0 = _loadUnit_memRequest_valid & sourceQueue_enq_ready;
  wire              axi4Port_r_ready_0;
  assign sourceQueue_enq_valid = _loadUnit_memRequest_valid & axi4Port_ar_ready_0;
  assign sourceQueue_deq_ready = axi4Port_r_ready_0 & axi4Port_r_valid_0;
  assign dataQueue_deq_valid = ~_dataQueue_fifo_empty;
  wire              axi4Port_w_valid_0 = dataQueue_deq_valid;
  wire [511:0]      dataQueue_dataOut_data;
  wire [511:0]      axi4Port_w_bits_data_0 = dataQueue_deq_bits_data;
  wire [63:0]       dataQueue_dataOut_mask;
  wire [63:0]       axi4Port_w_bits_strb_0 = dataQueue_deq_bits_mask;
  wire [5:0]        dataQueue_dataOut_index;
  wire [31:0]       dataQueue_dataOut_address;
  wire [5:0]        dataQueue_enq_bits_index;
  wire [31:0]       dataQueue_enq_bits_address;
  wire [37:0]       dataQueue_dataIn_lo = {dataQueue_enq_bits_index, dataQueue_enq_bits_address};
  wire [511:0]      dataQueue_enq_bits_data;
  wire [63:0]       dataQueue_enq_bits_mask;
  wire [575:0]      dataQueue_dataIn_hi = {dataQueue_enq_bits_data, dataQueue_enq_bits_mask};
  wire [613:0]      dataQueue_dataIn = {dataQueue_dataIn_hi, dataQueue_dataIn_lo};
  assign dataQueue_dataOut_address = _dataQueue_fifo_data_out[31:0];
  assign dataQueue_dataOut_index = _dataQueue_fifo_data_out[37:32];
  assign dataQueue_dataOut_mask = _dataQueue_fifo_data_out[101:38];
  assign dataQueue_dataOut_data = _dataQueue_fifo_data_out[613:102];
  assign dataQueue_deq_bits_data = dataQueue_dataOut_data;
  assign dataQueue_deq_bits_mask = dataQueue_dataOut_mask;
  wire [5:0]        dataQueue_deq_bits_index = dataQueue_dataOut_index;
  wire [31:0]       dataQueue_deq_bits_address = dataQueue_dataOut_address;
  wire              dataQueue_enq_ready = ~_dataQueue_fifo_full;
  wire              dataQueue_enq_valid;
  wire              axi4Port_aw_valid_0 = _storeUnit_memRequest_valid & dataQueue_enq_ready;
  wire [1:0]        axi4Port_aw_bits_id_0 = _storeUnit_memRequest_bits_index[1:0];
  assign dataQueue_enq_valid = _storeUnit_memRequest_valid & axi4Port_aw_ready_0;
  wire              simpleSourceQueue_deq_valid;
  assign simpleSourceQueue_deq_valid = ~_simpleSourceQueue_fifo_empty;
  wire              simpleSourceQueue_enq_ready = ~_simpleSourceQueue_fifo_full;
  wire              simpleSourceQueue_enq_valid;
  wire              simpleSourceQueue_deq_ready;
  wire              simpleAccessPorts_ar_valid_0 = _otherUnit_memReadRequest_valid & simpleSourceQueue_enq_ready;
  wire              simpleAccessPorts_r_ready_0;
  assign simpleSourceQueue_enq_valid = _otherUnit_memReadRequest_valid & simpleAccessPorts_ar_ready_0;
  assign simpleSourceQueue_deq_ready = simpleAccessPorts_r_ready_0 & simpleAccessPorts_r_valid_0;
  assign simpleDataQueue_deq_valid = ~_simpleDataQueue_fifo_empty;
  wire              simpleAccessPorts_w_valid_0 = simpleDataQueue_deq_valid;
  wire [31:0]       simpleDataQueue_dataOut_data;
  wire [31:0]       simpleAccessPorts_w_bits_data_0 = simpleDataQueue_deq_bits_data;
  wire [3:0]        simpleDataQueue_dataOut_mask;
  wire [3:0]        simpleAccessPorts_w_bits_strb_0 = simpleDataQueue_deq_bits_mask;
  wire [7:0]        simpleDataQueue_dataOut_source;
  wire [31:0]       simpleDataQueue_dataOut_address;
  wire [1:0]        simpleDataQueue_dataOut_size;
  wire [31:0]       simpleDataQueue_enq_bits_address;
  wire [1:0]        simpleDataQueue_enq_bits_size;
  wire [33:0]       simpleDataQueue_dataIn_lo = {simpleDataQueue_enq_bits_address, simpleDataQueue_enq_bits_size};
  wire [31:0]       simpleDataQueue_enq_bits_data;
  wire [3:0]        simpleDataQueue_enq_bits_mask;
  wire [35:0]       simpleDataQueue_dataIn_hi_hi = {simpleDataQueue_enq_bits_data, simpleDataQueue_enq_bits_mask};
  wire [7:0]        simpleDataQueue_enq_bits_source;
  wire [43:0]       simpleDataQueue_dataIn_hi = {simpleDataQueue_dataIn_hi_hi, simpleDataQueue_enq_bits_source};
  wire [77:0]       simpleDataQueue_dataIn = {simpleDataQueue_dataIn_hi, simpleDataQueue_dataIn_lo};
  assign simpleDataQueue_dataOut_size = _simpleDataQueue_fifo_data_out[1:0];
  assign simpleDataQueue_dataOut_address = _simpleDataQueue_fifo_data_out[33:2];
  assign simpleDataQueue_dataOut_source = _simpleDataQueue_fifo_data_out[41:34];
  assign simpleDataQueue_dataOut_mask = _simpleDataQueue_fifo_data_out[45:42];
  assign simpleDataQueue_dataOut_data = _simpleDataQueue_fifo_data_out[77:46];
  assign simpleDataQueue_deq_bits_data = simpleDataQueue_dataOut_data;
  assign simpleDataQueue_deq_bits_mask = simpleDataQueue_dataOut_mask;
  wire [7:0]        simpleDataQueue_deq_bits_source = simpleDataQueue_dataOut_source;
  wire [31:0]       simpleDataQueue_deq_bits_address = simpleDataQueue_dataOut_address;
  wire [1:0]        simpleDataQueue_deq_bits_size = simpleDataQueue_dataOut_size;
  wire              simpleDataQueue_enq_ready = ~_simpleDataQueue_fifo_full;
  wire              simpleDataQueue_enq_valid;
  wire              simpleAccessPorts_aw_valid_0 = _otherUnit_memWriteRequest_valid & dataQueue_enq_ready;
  wire [2:0]        simpleAccessPorts_aw_bits_size_0 = {1'h0, _otherUnit_memWriteRequest_bits_size};
  wire [1:0]        simpleAccessPorts_aw_bits_id_0 = _otherUnit_memWriteRequest_bits_source[1:0];
  assign simpleDataQueue_enq_valid = _otherUnit_memWriteRequest_valid & simpleAccessPorts_aw_ready_0;
  wire [1:0]        tokenIO_offsetGroupRelease_lo_lo_lo = {_otherUnit_offsetRelease_1, _otherUnit_offsetRelease_0};
  wire [1:0]        tokenIO_offsetGroupRelease_lo_lo_hi = {_otherUnit_offsetRelease_3, _otherUnit_offsetRelease_2};
  wire [3:0]        tokenIO_offsetGroupRelease_lo_lo = {tokenIO_offsetGroupRelease_lo_lo_hi, tokenIO_offsetGroupRelease_lo_lo_lo};
  wire [1:0]        tokenIO_offsetGroupRelease_lo_hi_lo = {_otherUnit_offsetRelease_5, _otherUnit_offsetRelease_4};
  wire [1:0]        tokenIO_offsetGroupRelease_lo_hi_hi = {_otherUnit_offsetRelease_7, _otherUnit_offsetRelease_6};
  wire [3:0]        tokenIO_offsetGroupRelease_lo_hi = {tokenIO_offsetGroupRelease_lo_hi_hi, tokenIO_offsetGroupRelease_lo_hi_lo};
  wire [7:0]        tokenIO_offsetGroupRelease_lo = {tokenIO_offsetGroupRelease_lo_hi, tokenIO_offsetGroupRelease_lo_lo};
  wire [1:0]        tokenIO_offsetGroupRelease_hi_lo_lo = {_otherUnit_offsetRelease_9, _otherUnit_offsetRelease_8};
  wire [1:0]        tokenIO_offsetGroupRelease_hi_lo_hi = {_otherUnit_offsetRelease_11, _otherUnit_offsetRelease_10};
  wire [3:0]        tokenIO_offsetGroupRelease_hi_lo = {tokenIO_offsetGroupRelease_hi_lo_hi, tokenIO_offsetGroupRelease_hi_lo_lo};
  wire [1:0]        tokenIO_offsetGroupRelease_hi_hi_lo = {_otherUnit_offsetRelease_13, _otherUnit_offsetRelease_12};
  wire [1:0]        tokenIO_offsetGroupRelease_hi_hi_hi = {_otherUnit_offsetRelease_15, _otherUnit_offsetRelease_14};
  wire [3:0]        tokenIO_offsetGroupRelease_hi_hi = {tokenIO_offsetGroupRelease_hi_hi_hi, tokenIO_offsetGroupRelease_hi_hi_lo};
  wire [7:0]        tokenIO_offsetGroupRelease_hi = {tokenIO_offsetGroupRelease_hi_hi, tokenIO_offsetGroupRelease_hi_lo};
  wire              unitOrder =
    _loadUnit_status_instructionIndex == _storeUnit_status_instructionIndex | _loadUnit_status_instructionIndex[1:0] < _storeUnit_status_instructionIndex[1:0] ^ _loadUnit_status_instructionIndex[2] ^ _storeUnit_status_instructionIndex[2];
  wire              loadAddressConflict = _loadUnit_status_startAddress >= _storeUnit_status_startAddress & _loadUnit_status_startAddress <= _storeUnit_status_endAddress;
  wire              storeAddressConflict = _storeUnit_status_startAddress >= _loadUnit_status_startAddress & _storeUnit_status_startAddress <= _loadUnit_status_endAddress;
  wire              stallLoad = ~unitOrder & loadAddressConflict & ~_storeUnit_status_idle;
  wire              stallStore = unitOrder & storeAddressConflict & ~_loadUnit_status_idle;
  always @(posedge clock) begin
    if (reset) begin
      v0_0 <= 32'h0;
      v0_1 <= 32'h0;
      v0_2 <= 32'h0;
      v0_3 <= 32'h0;
      v0_4 <= 32'h0;
      v0_5 <= 32'h0;
      v0_6 <= 32'h0;
      v0_7 <= 32'h0;
      v0_8 <= 32'h0;
      v0_9 <= 32'h0;
      v0_10 <= 32'h0;
      v0_11 <= 32'h0;
      v0_12 <= 32'h0;
      v0_13 <= 32'h0;
      v0_14 <= 32'h0;
      v0_15 <= 32'h0;
      v0_16 <= 32'h0;
      v0_17 <= 32'h0;
      v0_18 <= 32'h0;
      v0_19 <= 32'h0;
      v0_20 <= 32'h0;
      v0_21 <= 32'h0;
      v0_22 <= 32'h0;
      v0_23 <= 32'h0;
      v0_24 <= 32'h0;
      v0_25 <= 32'h0;
      v0_26 <= 32'h0;
      v0_27 <= 32'h0;
      v0_28 <= 32'h0;
      v0_29 <= 32'h0;
      v0_30 <= 32'h0;
      v0_31 <= 32'h0;
      v0_32 <= 32'h0;
      v0_33 <= 32'h0;
      v0_34 <= 32'h0;
      v0_35 <= 32'h0;
      v0_36 <= 32'h0;
      v0_37 <= 32'h0;
      v0_38 <= 32'h0;
      v0_39 <= 32'h0;
      v0_40 <= 32'h0;
      v0_41 <= 32'h0;
      v0_42 <= 32'h0;
      v0_43 <= 32'h0;
      v0_44 <= 32'h0;
      v0_45 <= 32'h0;
      v0_46 <= 32'h0;
      v0_47 <= 32'h0;
      v0_48 <= 32'h0;
      v0_49 <= 32'h0;
      v0_50 <= 32'h0;
      v0_51 <= 32'h0;
      v0_52 <= 32'h0;
      v0_53 <= 32'h0;
      v0_54 <= 32'h0;
      v0_55 <= 32'h0;
      v0_56 <= 32'h0;
      v0_57 <= 32'h0;
      v0_58 <= 32'h0;
      v0_59 <= 32'h0;
      v0_60 <= 32'h0;
      v0_61 <= 32'h0;
      v0_62 <= 32'h0;
      v0_63 <= 32'h0;
      queueCount_0 <= 7'h0;
      queueCount_1 <= 7'h0;
      queueCount_2 <= 7'h0;
      queueCount_3 <= 7'h0;
      queueCount_4 <= 7'h0;
      queueCount_5 <= 7'h0;
      queueCount_6 <= 7'h0;
      queueCount_7 <= 7'h0;
      queueCount_0_1 <= 7'h0;
      queueCount_1_1 <= 7'h0;
      queueCount_2_1 <= 7'h0;
      queueCount_3_1 <= 7'h0;
      queueCount_4_1 <= 7'h0;
      queueCount_5_1 <= 7'h0;
      queueCount_6_1 <= 7'h0;
      queueCount_7_1 <= 7'h0;
      queueCount_0_2 <= 7'h0;
      queueCount_1_2 <= 7'h0;
      queueCount_2_2 <= 7'h0;
      queueCount_3_2 <= 7'h0;
      queueCount_4_2 <= 7'h0;
      queueCount_5_2 <= 7'h0;
      queueCount_6_2 <= 7'h0;
      queueCount_7_2 <= 7'h0;
      queueCount_0_3 <= 7'h0;
      queueCount_1_3 <= 7'h0;
      queueCount_2_3 <= 7'h0;
      queueCount_3_3 <= 7'h0;
      queueCount_4_3 <= 7'h0;
      queueCount_5_3 <= 7'h0;
      queueCount_6_3 <= 7'h0;
      queueCount_7_3 <= 7'h0;
      queueCount_0_4 <= 7'h0;
      queueCount_1_4 <= 7'h0;
      queueCount_2_4 <= 7'h0;
      queueCount_3_4 <= 7'h0;
      queueCount_4_4 <= 7'h0;
      queueCount_5_4 <= 7'h0;
      queueCount_6_4 <= 7'h0;
      queueCount_7_4 <= 7'h0;
      queueCount_0_5 <= 7'h0;
      queueCount_1_5 <= 7'h0;
      queueCount_2_5 <= 7'h0;
      queueCount_3_5 <= 7'h0;
      queueCount_4_5 <= 7'h0;
      queueCount_5_5 <= 7'h0;
      queueCount_6_5 <= 7'h0;
      queueCount_7_5 <= 7'h0;
      queueCount_0_6 <= 7'h0;
      queueCount_1_6 <= 7'h0;
      queueCount_2_6 <= 7'h0;
      queueCount_3_6 <= 7'h0;
      queueCount_4_6 <= 7'h0;
      queueCount_5_6 <= 7'h0;
      queueCount_6_6 <= 7'h0;
      queueCount_7_6 <= 7'h0;
      queueCount_0_7 <= 7'h0;
      queueCount_1_7 <= 7'h0;
      queueCount_2_7 <= 7'h0;
      queueCount_3_7 <= 7'h0;
      queueCount_4_7 <= 7'h0;
      queueCount_5_7 <= 7'h0;
      queueCount_6_7 <= 7'h0;
      queueCount_7_7 <= 7'h0;
      queueCount_0_8 <= 7'h0;
      queueCount_1_8 <= 7'h0;
      queueCount_2_8 <= 7'h0;
      queueCount_3_8 <= 7'h0;
      queueCount_4_8 <= 7'h0;
      queueCount_5_8 <= 7'h0;
      queueCount_6_8 <= 7'h0;
      queueCount_7_8 <= 7'h0;
      queueCount_0_9 <= 7'h0;
      queueCount_1_9 <= 7'h0;
      queueCount_2_9 <= 7'h0;
      queueCount_3_9 <= 7'h0;
      queueCount_4_9 <= 7'h0;
      queueCount_5_9 <= 7'h0;
      queueCount_6_9 <= 7'h0;
      queueCount_7_9 <= 7'h0;
      queueCount_0_10 <= 7'h0;
      queueCount_1_10 <= 7'h0;
      queueCount_2_10 <= 7'h0;
      queueCount_3_10 <= 7'h0;
      queueCount_4_10 <= 7'h0;
      queueCount_5_10 <= 7'h0;
      queueCount_6_10 <= 7'h0;
      queueCount_7_10 <= 7'h0;
      queueCount_0_11 <= 7'h0;
      queueCount_1_11 <= 7'h0;
      queueCount_2_11 <= 7'h0;
      queueCount_3_11 <= 7'h0;
      queueCount_4_11 <= 7'h0;
      queueCount_5_11 <= 7'h0;
      queueCount_6_11 <= 7'h0;
      queueCount_7_11 <= 7'h0;
      queueCount_0_12 <= 7'h0;
      queueCount_1_12 <= 7'h0;
      queueCount_2_12 <= 7'h0;
      queueCount_3_12 <= 7'h0;
      queueCount_4_12 <= 7'h0;
      queueCount_5_12 <= 7'h0;
      queueCount_6_12 <= 7'h0;
      queueCount_7_12 <= 7'h0;
      queueCount_0_13 <= 7'h0;
      queueCount_1_13 <= 7'h0;
      queueCount_2_13 <= 7'h0;
      queueCount_3_13 <= 7'h0;
      queueCount_4_13 <= 7'h0;
      queueCount_5_13 <= 7'h0;
      queueCount_6_13 <= 7'h0;
      queueCount_7_13 <= 7'h0;
      queueCount_0_14 <= 7'h0;
      queueCount_1_14 <= 7'h0;
      queueCount_2_14 <= 7'h0;
      queueCount_3_14 <= 7'h0;
      queueCount_4_14 <= 7'h0;
      queueCount_5_14 <= 7'h0;
      queueCount_6_14 <= 7'h0;
      queueCount_7_14 <= 7'h0;
      queueCount_0_15 <= 7'h0;
      queueCount_1_15 <= 7'h0;
      queueCount_2_15 <= 7'h0;
      queueCount_3_15 <= 7'h0;
      queueCount_4_15 <= 7'h0;
      queueCount_5_15 <= 7'h0;
      queueCount_6_15 <= 7'h0;
      queueCount_7_15 <= 7'h0;
    end
    else begin
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 2'h0)
        v0_0 <= v0_0 & ~maskExt | maskExt & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 2'h0)
        v0_1 <= v0_1 & ~maskExt_1 | maskExt_1 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 2'h0)
        v0_2 <= v0_2 & ~maskExt_2 | maskExt_2 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 2'h0)
        v0_3 <= v0_3 & ~maskExt_3 | maskExt_3 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_4_valid & v0UpdateVec_4_bits_offset == 2'h0)
        v0_4 <= v0_4 & ~maskExt_4 | maskExt_4 & v0UpdateVec_4_bits_data;
      if (v0UpdateVec_5_valid & v0UpdateVec_5_bits_offset == 2'h0)
        v0_5 <= v0_5 & ~maskExt_5 | maskExt_5 & v0UpdateVec_5_bits_data;
      if (v0UpdateVec_6_valid & v0UpdateVec_6_bits_offset == 2'h0)
        v0_6 <= v0_6 & ~maskExt_6 | maskExt_6 & v0UpdateVec_6_bits_data;
      if (v0UpdateVec_7_valid & v0UpdateVec_7_bits_offset == 2'h0)
        v0_7 <= v0_7 & ~maskExt_7 | maskExt_7 & v0UpdateVec_7_bits_data;
      if (v0UpdateVec_8_valid & v0UpdateVec_8_bits_offset == 2'h0)
        v0_8 <= v0_8 & ~maskExt_8 | maskExt_8 & v0UpdateVec_8_bits_data;
      if (v0UpdateVec_9_valid & v0UpdateVec_9_bits_offset == 2'h0)
        v0_9 <= v0_9 & ~maskExt_9 | maskExt_9 & v0UpdateVec_9_bits_data;
      if (v0UpdateVec_10_valid & v0UpdateVec_10_bits_offset == 2'h0)
        v0_10 <= v0_10 & ~maskExt_10 | maskExt_10 & v0UpdateVec_10_bits_data;
      if (v0UpdateVec_11_valid & v0UpdateVec_11_bits_offset == 2'h0)
        v0_11 <= v0_11 & ~maskExt_11 | maskExt_11 & v0UpdateVec_11_bits_data;
      if (v0UpdateVec_12_valid & v0UpdateVec_12_bits_offset == 2'h0)
        v0_12 <= v0_12 & ~maskExt_12 | maskExt_12 & v0UpdateVec_12_bits_data;
      if (v0UpdateVec_13_valid & v0UpdateVec_13_bits_offset == 2'h0)
        v0_13 <= v0_13 & ~maskExt_13 | maskExt_13 & v0UpdateVec_13_bits_data;
      if (v0UpdateVec_14_valid & v0UpdateVec_14_bits_offset == 2'h0)
        v0_14 <= v0_14 & ~maskExt_14 | maskExt_14 & v0UpdateVec_14_bits_data;
      if (v0UpdateVec_15_valid & v0UpdateVec_15_bits_offset == 2'h0)
        v0_15 <= v0_15 & ~maskExt_15 | maskExt_15 & v0UpdateVec_15_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 2'h1)
        v0_16 <= v0_16 & ~maskExt_16 | maskExt_16 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 2'h1)
        v0_17 <= v0_17 & ~maskExt_17 | maskExt_17 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 2'h1)
        v0_18 <= v0_18 & ~maskExt_18 | maskExt_18 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 2'h1)
        v0_19 <= v0_19 & ~maskExt_19 | maskExt_19 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_4_valid & v0UpdateVec_4_bits_offset == 2'h1)
        v0_20 <= v0_20 & ~maskExt_20 | maskExt_20 & v0UpdateVec_4_bits_data;
      if (v0UpdateVec_5_valid & v0UpdateVec_5_bits_offset == 2'h1)
        v0_21 <= v0_21 & ~maskExt_21 | maskExt_21 & v0UpdateVec_5_bits_data;
      if (v0UpdateVec_6_valid & v0UpdateVec_6_bits_offset == 2'h1)
        v0_22 <= v0_22 & ~maskExt_22 | maskExt_22 & v0UpdateVec_6_bits_data;
      if (v0UpdateVec_7_valid & v0UpdateVec_7_bits_offset == 2'h1)
        v0_23 <= v0_23 & ~maskExt_23 | maskExt_23 & v0UpdateVec_7_bits_data;
      if (v0UpdateVec_8_valid & v0UpdateVec_8_bits_offset == 2'h1)
        v0_24 <= v0_24 & ~maskExt_24 | maskExt_24 & v0UpdateVec_8_bits_data;
      if (v0UpdateVec_9_valid & v0UpdateVec_9_bits_offset == 2'h1)
        v0_25 <= v0_25 & ~maskExt_25 | maskExt_25 & v0UpdateVec_9_bits_data;
      if (v0UpdateVec_10_valid & v0UpdateVec_10_bits_offset == 2'h1)
        v0_26 <= v0_26 & ~maskExt_26 | maskExt_26 & v0UpdateVec_10_bits_data;
      if (v0UpdateVec_11_valid & v0UpdateVec_11_bits_offset == 2'h1)
        v0_27 <= v0_27 & ~maskExt_27 | maskExt_27 & v0UpdateVec_11_bits_data;
      if (v0UpdateVec_12_valid & v0UpdateVec_12_bits_offset == 2'h1)
        v0_28 <= v0_28 & ~maskExt_28 | maskExt_28 & v0UpdateVec_12_bits_data;
      if (v0UpdateVec_13_valid & v0UpdateVec_13_bits_offset == 2'h1)
        v0_29 <= v0_29 & ~maskExt_29 | maskExt_29 & v0UpdateVec_13_bits_data;
      if (v0UpdateVec_14_valid & v0UpdateVec_14_bits_offset == 2'h1)
        v0_30 <= v0_30 & ~maskExt_30 | maskExt_30 & v0UpdateVec_14_bits_data;
      if (v0UpdateVec_15_valid & v0UpdateVec_15_bits_offset == 2'h1)
        v0_31 <= v0_31 & ~maskExt_31 | maskExt_31 & v0UpdateVec_15_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 2'h2)
        v0_32 <= v0_32 & ~maskExt_32 | maskExt_32 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 2'h2)
        v0_33 <= v0_33 & ~maskExt_33 | maskExt_33 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 2'h2)
        v0_34 <= v0_34 & ~maskExt_34 | maskExt_34 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 2'h2)
        v0_35 <= v0_35 & ~maskExt_35 | maskExt_35 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_4_valid & v0UpdateVec_4_bits_offset == 2'h2)
        v0_36 <= v0_36 & ~maskExt_36 | maskExt_36 & v0UpdateVec_4_bits_data;
      if (v0UpdateVec_5_valid & v0UpdateVec_5_bits_offset == 2'h2)
        v0_37 <= v0_37 & ~maskExt_37 | maskExt_37 & v0UpdateVec_5_bits_data;
      if (v0UpdateVec_6_valid & v0UpdateVec_6_bits_offset == 2'h2)
        v0_38 <= v0_38 & ~maskExt_38 | maskExt_38 & v0UpdateVec_6_bits_data;
      if (v0UpdateVec_7_valid & v0UpdateVec_7_bits_offset == 2'h2)
        v0_39 <= v0_39 & ~maskExt_39 | maskExt_39 & v0UpdateVec_7_bits_data;
      if (v0UpdateVec_8_valid & v0UpdateVec_8_bits_offset == 2'h2)
        v0_40 <= v0_40 & ~maskExt_40 | maskExt_40 & v0UpdateVec_8_bits_data;
      if (v0UpdateVec_9_valid & v0UpdateVec_9_bits_offset == 2'h2)
        v0_41 <= v0_41 & ~maskExt_41 | maskExt_41 & v0UpdateVec_9_bits_data;
      if (v0UpdateVec_10_valid & v0UpdateVec_10_bits_offset == 2'h2)
        v0_42 <= v0_42 & ~maskExt_42 | maskExt_42 & v0UpdateVec_10_bits_data;
      if (v0UpdateVec_11_valid & v0UpdateVec_11_bits_offset == 2'h2)
        v0_43 <= v0_43 & ~maskExt_43 | maskExt_43 & v0UpdateVec_11_bits_data;
      if (v0UpdateVec_12_valid & v0UpdateVec_12_bits_offset == 2'h2)
        v0_44 <= v0_44 & ~maskExt_44 | maskExt_44 & v0UpdateVec_12_bits_data;
      if (v0UpdateVec_13_valid & v0UpdateVec_13_bits_offset == 2'h2)
        v0_45 <= v0_45 & ~maskExt_45 | maskExt_45 & v0UpdateVec_13_bits_data;
      if (v0UpdateVec_14_valid & v0UpdateVec_14_bits_offset == 2'h2)
        v0_46 <= v0_46 & ~maskExt_46 | maskExt_46 & v0UpdateVec_14_bits_data;
      if (v0UpdateVec_15_valid & v0UpdateVec_15_bits_offset == 2'h2)
        v0_47 <= v0_47 & ~maskExt_47 | maskExt_47 & v0UpdateVec_15_bits_data;
      if (v0UpdateVec_0_valid & (&v0UpdateVec_0_bits_offset))
        v0_48 <= v0_48 & ~maskExt_48 | maskExt_48 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & (&v0UpdateVec_1_bits_offset))
        v0_49 <= v0_49 & ~maskExt_49 | maskExt_49 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & (&v0UpdateVec_2_bits_offset))
        v0_50 <= v0_50 & ~maskExt_50 | maskExt_50 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & (&v0UpdateVec_3_bits_offset))
        v0_51 <= v0_51 & ~maskExt_51 | maskExt_51 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_4_valid & (&v0UpdateVec_4_bits_offset))
        v0_52 <= v0_52 & ~maskExt_52 | maskExt_52 & v0UpdateVec_4_bits_data;
      if (v0UpdateVec_5_valid & (&v0UpdateVec_5_bits_offset))
        v0_53 <= v0_53 & ~maskExt_53 | maskExt_53 & v0UpdateVec_5_bits_data;
      if (v0UpdateVec_6_valid & (&v0UpdateVec_6_bits_offset))
        v0_54 <= v0_54 & ~maskExt_54 | maskExt_54 & v0UpdateVec_6_bits_data;
      if (v0UpdateVec_7_valid & (&v0UpdateVec_7_bits_offset))
        v0_55 <= v0_55 & ~maskExt_55 | maskExt_55 & v0UpdateVec_7_bits_data;
      if (v0UpdateVec_8_valid & (&v0UpdateVec_8_bits_offset))
        v0_56 <= v0_56 & ~maskExt_56 | maskExt_56 & v0UpdateVec_8_bits_data;
      if (v0UpdateVec_9_valid & (&v0UpdateVec_9_bits_offset))
        v0_57 <= v0_57 & ~maskExt_57 | maskExt_57 & v0UpdateVec_9_bits_data;
      if (v0UpdateVec_10_valid & (&v0UpdateVec_10_bits_offset))
        v0_58 <= v0_58 & ~maskExt_58 | maskExt_58 & v0UpdateVec_10_bits_data;
      if (v0UpdateVec_11_valid & (&v0UpdateVec_11_bits_offset))
        v0_59 <= v0_59 & ~maskExt_59 | maskExt_59 & v0UpdateVec_11_bits_data;
      if (v0UpdateVec_12_valid & (&v0UpdateVec_12_bits_offset))
        v0_60 <= v0_60 & ~maskExt_60 | maskExt_60 & v0UpdateVec_12_bits_data;
      if (v0UpdateVec_13_valid & (&v0UpdateVec_13_bits_offset))
        v0_61 <= v0_61 & ~maskExt_61 | maskExt_61 & v0UpdateVec_13_bits_data;
      if (v0UpdateVec_14_valid & (&v0UpdateVec_14_bits_offset))
        v0_62 <= v0_62 & ~maskExt_62 | maskExt_62 & v0UpdateVec_14_bits_data;
      if (v0UpdateVec_15_valid & (&v0UpdateVec_15_bits_offset))
        v0_63 <= v0_63 & ~maskExt_63 | maskExt_63 & v0UpdateVec_15_bits_data;
      if (queueEnq[0] ^ queueDeq[0])
        queueCount_0 <= queueCount_0 + counterUpdate;
      if (queueEnq[1] ^ queueDeq[1])
        queueCount_1 <= queueCount_1 + counterUpdate_1;
      if (queueEnq[2] ^ queueDeq[2])
        queueCount_2 <= queueCount_2 + counterUpdate_2;
      if (queueEnq[3] ^ queueDeq[3])
        queueCount_3 <= queueCount_3 + counterUpdate_3;
      if (queueEnq[4] ^ queueDeq[4])
        queueCount_4 <= queueCount_4 + counterUpdate_4;
      if (queueEnq[5] ^ queueDeq[5])
        queueCount_5 <= queueCount_5 + counterUpdate_5;
      if (queueEnq[6] ^ queueDeq[6])
        queueCount_6 <= queueCount_6 + counterUpdate_6;
      if (queueEnq[7] ^ queueDeq[7])
        queueCount_7 <= queueCount_7 + counterUpdate_7;
      if (queueEnq_1[0] ^ queueDeq_1[0])
        queueCount_0_1 <= queueCount_0_1 + counterUpdate_8;
      if (queueEnq_1[1] ^ queueDeq_1[1])
        queueCount_1_1 <= queueCount_1_1 + counterUpdate_9;
      if (queueEnq_1[2] ^ queueDeq_1[2])
        queueCount_2_1 <= queueCount_2_1 + counterUpdate_10;
      if (queueEnq_1[3] ^ queueDeq_1[3])
        queueCount_3_1 <= queueCount_3_1 + counterUpdate_11;
      if (queueEnq_1[4] ^ queueDeq_1[4])
        queueCount_4_1 <= queueCount_4_1 + counterUpdate_12;
      if (queueEnq_1[5] ^ queueDeq_1[5])
        queueCount_5_1 <= queueCount_5_1 + counterUpdate_13;
      if (queueEnq_1[6] ^ queueDeq_1[6])
        queueCount_6_1 <= queueCount_6_1 + counterUpdate_14;
      if (queueEnq_1[7] ^ queueDeq_1[7])
        queueCount_7_1 <= queueCount_7_1 + counterUpdate_15;
      if (queueEnq_2[0] ^ queueDeq_2[0])
        queueCount_0_2 <= queueCount_0_2 + counterUpdate_16;
      if (queueEnq_2[1] ^ queueDeq_2[1])
        queueCount_1_2 <= queueCount_1_2 + counterUpdate_17;
      if (queueEnq_2[2] ^ queueDeq_2[2])
        queueCount_2_2 <= queueCount_2_2 + counterUpdate_18;
      if (queueEnq_2[3] ^ queueDeq_2[3])
        queueCount_3_2 <= queueCount_3_2 + counterUpdate_19;
      if (queueEnq_2[4] ^ queueDeq_2[4])
        queueCount_4_2 <= queueCount_4_2 + counterUpdate_20;
      if (queueEnq_2[5] ^ queueDeq_2[5])
        queueCount_5_2 <= queueCount_5_2 + counterUpdate_21;
      if (queueEnq_2[6] ^ queueDeq_2[6])
        queueCount_6_2 <= queueCount_6_2 + counterUpdate_22;
      if (queueEnq_2[7] ^ queueDeq_2[7])
        queueCount_7_2 <= queueCount_7_2 + counterUpdate_23;
      if (queueEnq_3[0] ^ queueDeq_3[0])
        queueCount_0_3 <= queueCount_0_3 + counterUpdate_24;
      if (queueEnq_3[1] ^ queueDeq_3[1])
        queueCount_1_3 <= queueCount_1_3 + counterUpdate_25;
      if (queueEnq_3[2] ^ queueDeq_3[2])
        queueCount_2_3 <= queueCount_2_3 + counterUpdate_26;
      if (queueEnq_3[3] ^ queueDeq_3[3])
        queueCount_3_3 <= queueCount_3_3 + counterUpdate_27;
      if (queueEnq_3[4] ^ queueDeq_3[4])
        queueCount_4_3 <= queueCount_4_3 + counterUpdate_28;
      if (queueEnq_3[5] ^ queueDeq_3[5])
        queueCount_5_3 <= queueCount_5_3 + counterUpdate_29;
      if (queueEnq_3[6] ^ queueDeq_3[6])
        queueCount_6_3 <= queueCount_6_3 + counterUpdate_30;
      if (queueEnq_3[7] ^ queueDeq_3[7])
        queueCount_7_3 <= queueCount_7_3 + counterUpdate_31;
      if (queueEnq_4[0] ^ queueDeq_4[0])
        queueCount_0_4 <= queueCount_0_4 + counterUpdate_32;
      if (queueEnq_4[1] ^ queueDeq_4[1])
        queueCount_1_4 <= queueCount_1_4 + counterUpdate_33;
      if (queueEnq_4[2] ^ queueDeq_4[2])
        queueCount_2_4 <= queueCount_2_4 + counterUpdate_34;
      if (queueEnq_4[3] ^ queueDeq_4[3])
        queueCount_3_4 <= queueCount_3_4 + counterUpdate_35;
      if (queueEnq_4[4] ^ queueDeq_4[4])
        queueCount_4_4 <= queueCount_4_4 + counterUpdate_36;
      if (queueEnq_4[5] ^ queueDeq_4[5])
        queueCount_5_4 <= queueCount_5_4 + counterUpdate_37;
      if (queueEnq_4[6] ^ queueDeq_4[6])
        queueCount_6_4 <= queueCount_6_4 + counterUpdate_38;
      if (queueEnq_4[7] ^ queueDeq_4[7])
        queueCount_7_4 <= queueCount_7_4 + counterUpdate_39;
      if (queueEnq_5[0] ^ queueDeq_5[0])
        queueCount_0_5 <= queueCount_0_5 + counterUpdate_40;
      if (queueEnq_5[1] ^ queueDeq_5[1])
        queueCount_1_5 <= queueCount_1_5 + counterUpdate_41;
      if (queueEnq_5[2] ^ queueDeq_5[2])
        queueCount_2_5 <= queueCount_2_5 + counterUpdate_42;
      if (queueEnq_5[3] ^ queueDeq_5[3])
        queueCount_3_5 <= queueCount_3_5 + counterUpdate_43;
      if (queueEnq_5[4] ^ queueDeq_5[4])
        queueCount_4_5 <= queueCount_4_5 + counterUpdate_44;
      if (queueEnq_5[5] ^ queueDeq_5[5])
        queueCount_5_5 <= queueCount_5_5 + counterUpdate_45;
      if (queueEnq_5[6] ^ queueDeq_5[6])
        queueCount_6_5 <= queueCount_6_5 + counterUpdate_46;
      if (queueEnq_5[7] ^ queueDeq_5[7])
        queueCount_7_5 <= queueCount_7_5 + counterUpdate_47;
      if (queueEnq_6[0] ^ queueDeq_6[0])
        queueCount_0_6 <= queueCount_0_6 + counterUpdate_48;
      if (queueEnq_6[1] ^ queueDeq_6[1])
        queueCount_1_6 <= queueCount_1_6 + counterUpdate_49;
      if (queueEnq_6[2] ^ queueDeq_6[2])
        queueCount_2_6 <= queueCount_2_6 + counterUpdate_50;
      if (queueEnq_6[3] ^ queueDeq_6[3])
        queueCount_3_6 <= queueCount_3_6 + counterUpdate_51;
      if (queueEnq_6[4] ^ queueDeq_6[4])
        queueCount_4_6 <= queueCount_4_6 + counterUpdate_52;
      if (queueEnq_6[5] ^ queueDeq_6[5])
        queueCount_5_6 <= queueCount_5_6 + counterUpdate_53;
      if (queueEnq_6[6] ^ queueDeq_6[6])
        queueCount_6_6 <= queueCount_6_6 + counterUpdate_54;
      if (queueEnq_6[7] ^ queueDeq_6[7])
        queueCount_7_6 <= queueCount_7_6 + counterUpdate_55;
      if (queueEnq_7[0] ^ queueDeq_7[0])
        queueCount_0_7 <= queueCount_0_7 + counterUpdate_56;
      if (queueEnq_7[1] ^ queueDeq_7[1])
        queueCount_1_7 <= queueCount_1_7 + counterUpdate_57;
      if (queueEnq_7[2] ^ queueDeq_7[2])
        queueCount_2_7 <= queueCount_2_7 + counterUpdate_58;
      if (queueEnq_7[3] ^ queueDeq_7[3])
        queueCount_3_7 <= queueCount_3_7 + counterUpdate_59;
      if (queueEnq_7[4] ^ queueDeq_7[4])
        queueCount_4_7 <= queueCount_4_7 + counterUpdate_60;
      if (queueEnq_7[5] ^ queueDeq_7[5])
        queueCount_5_7 <= queueCount_5_7 + counterUpdate_61;
      if (queueEnq_7[6] ^ queueDeq_7[6])
        queueCount_6_7 <= queueCount_6_7 + counterUpdate_62;
      if (queueEnq_7[7] ^ queueDeq_7[7])
        queueCount_7_7 <= queueCount_7_7 + counterUpdate_63;
      if (queueEnq_8[0] ^ queueDeq_8[0])
        queueCount_0_8 <= queueCount_0_8 + counterUpdate_64;
      if (queueEnq_8[1] ^ queueDeq_8[1])
        queueCount_1_8 <= queueCount_1_8 + counterUpdate_65;
      if (queueEnq_8[2] ^ queueDeq_8[2])
        queueCount_2_8 <= queueCount_2_8 + counterUpdate_66;
      if (queueEnq_8[3] ^ queueDeq_8[3])
        queueCount_3_8 <= queueCount_3_8 + counterUpdate_67;
      if (queueEnq_8[4] ^ queueDeq_8[4])
        queueCount_4_8 <= queueCount_4_8 + counterUpdate_68;
      if (queueEnq_8[5] ^ queueDeq_8[5])
        queueCount_5_8 <= queueCount_5_8 + counterUpdate_69;
      if (queueEnq_8[6] ^ queueDeq_8[6])
        queueCount_6_8 <= queueCount_6_8 + counterUpdate_70;
      if (queueEnq_8[7] ^ queueDeq_8[7])
        queueCount_7_8 <= queueCount_7_8 + counterUpdate_71;
      if (queueEnq_9[0] ^ queueDeq_9[0])
        queueCount_0_9 <= queueCount_0_9 + counterUpdate_72;
      if (queueEnq_9[1] ^ queueDeq_9[1])
        queueCount_1_9 <= queueCount_1_9 + counterUpdate_73;
      if (queueEnq_9[2] ^ queueDeq_9[2])
        queueCount_2_9 <= queueCount_2_9 + counterUpdate_74;
      if (queueEnq_9[3] ^ queueDeq_9[3])
        queueCount_3_9 <= queueCount_3_9 + counterUpdate_75;
      if (queueEnq_9[4] ^ queueDeq_9[4])
        queueCount_4_9 <= queueCount_4_9 + counterUpdate_76;
      if (queueEnq_9[5] ^ queueDeq_9[5])
        queueCount_5_9 <= queueCount_5_9 + counterUpdate_77;
      if (queueEnq_9[6] ^ queueDeq_9[6])
        queueCount_6_9 <= queueCount_6_9 + counterUpdate_78;
      if (queueEnq_9[7] ^ queueDeq_9[7])
        queueCount_7_9 <= queueCount_7_9 + counterUpdate_79;
      if (queueEnq_10[0] ^ queueDeq_10[0])
        queueCount_0_10 <= queueCount_0_10 + counterUpdate_80;
      if (queueEnq_10[1] ^ queueDeq_10[1])
        queueCount_1_10 <= queueCount_1_10 + counterUpdate_81;
      if (queueEnq_10[2] ^ queueDeq_10[2])
        queueCount_2_10 <= queueCount_2_10 + counterUpdate_82;
      if (queueEnq_10[3] ^ queueDeq_10[3])
        queueCount_3_10 <= queueCount_3_10 + counterUpdate_83;
      if (queueEnq_10[4] ^ queueDeq_10[4])
        queueCount_4_10 <= queueCount_4_10 + counterUpdate_84;
      if (queueEnq_10[5] ^ queueDeq_10[5])
        queueCount_5_10 <= queueCount_5_10 + counterUpdate_85;
      if (queueEnq_10[6] ^ queueDeq_10[6])
        queueCount_6_10 <= queueCount_6_10 + counterUpdate_86;
      if (queueEnq_10[7] ^ queueDeq_10[7])
        queueCount_7_10 <= queueCount_7_10 + counterUpdate_87;
      if (queueEnq_11[0] ^ queueDeq_11[0])
        queueCount_0_11 <= queueCount_0_11 + counterUpdate_88;
      if (queueEnq_11[1] ^ queueDeq_11[1])
        queueCount_1_11 <= queueCount_1_11 + counterUpdate_89;
      if (queueEnq_11[2] ^ queueDeq_11[2])
        queueCount_2_11 <= queueCount_2_11 + counterUpdate_90;
      if (queueEnq_11[3] ^ queueDeq_11[3])
        queueCount_3_11 <= queueCount_3_11 + counterUpdate_91;
      if (queueEnq_11[4] ^ queueDeq_11[4])
        queueCount_4_11 <= queueCount_4_11 + counterUpdate_92;
      if (queueEnq_11[5] ^ queueDeq_11[5])
        queueCount_5_11 <= queueCount_5_11 + counterUpdate_93;
      if (queueEnq_11[6] ^ queueDeq_11[6])
        queueCount_6_11 <= queueCount_6_11 + counterUpdate_94;
      if (queueEnq_11[7] ^ queueDeq_11[7])
        queueCount_7_11 <= queueCount_7_11 + counterUpdate_95;
      if (queueEnq_12[0] ^ queueDeq_12[0])
        queueCount_0_12 <= queueCount_0_12 + counterUpdate_96;
      if (queueEnq_12[1] ^ queueDeq_12[1])
        queueCount_1_12 <= queueCount_1_12 + counterUpdate_97;
      if (queueEnq_12[2] ^ queueDeq_12[2])
        queueCount_2_12 <= queueCount_2_12 + counterUpdate_98;
      if (queueEnq_12[3] ^ queueDeq_12[3])
        queueCount_3_12 <= queueCount_3_12 + counterUpdate_99;
      if (queueEnq_12[4] ^ queueDeq_12[4])
        queueCount_4_12 <= queueCount_4_12 + counterUpdate_100;
      if (queueEnq_12[5] ^ queueDeq_12[5])
        queueCount_5_12 <= queueCount_5_12 + counterUpdate_101;
      if (queueEnq_12[6] ^ queueDeq_12[6])
        queueCount_6_12 <= queueCount_6_12 + counterUpdate_102;
      if (queueEnq_12[7] ^ queueDeq_12[7])
        queueCount_7_12 <= queueCount_7_12 + counterUpdate_103;
      if (queueEnq_13[0] ^ queueDeq_13[0])
        queueCount_0_13 <= queueCount_0_13 + counterUpdate_104;
      if (queueEnq_13[1] ^ queueDeq_13[1])
        queueCount_1_13 <= queueCount_1_13 + counterUpdate_105;
      if (queueEnq_13[2] ^ queueDeq_13[2])
        queueCount_2_13 <= queueCount_2_13 + counterUpdate_106;
      if (queueEnq_13[3] ^ queueDeq_13[3])
        queueCount_3_13 <= queueCount_3_13 + counterUpdate_107;
      if (queueEnq_13[4] ^ queueDeq_13[4])
        queueCount_4_13 <= queueCount_4_13 + counterUpdate_108;
      if (queueEnq_13[5] ^ queueDeq_13[5])
        queueCount_5_13 <= queueCount_5_13 + counterUpdate_109;
      if (queueEnq_13[6] ^ queueDeq_13[6])
        queueCount_6_13 <= queueCount_6_13 + counterUpdate_110;
      if (queueEnq_13[7] ^ queueDeq_13[7])
        queueCount_7_13 <= queueCount_7_13 + counterUpdate_111;
      if (queueEnq_14[0] ^ queueDeq_14[0])
        queueCount_0_14 <= queueCount_0_14 + counterUpdate_112;
      if (queueEnq_14[1] ^ queueDeq_14[1])
        queueCount_1_14 <= queueCount_1_14 + counterUpdate_113;
      if (queueEnq_14[2] ^ queueDeq_14[2])
        queueCount_2_14 <= queueCount_2_14 + counterUpdate_114;
      if (queueEnq_14[3] ^ queueDeq_14[3])
        queueCount_3_14 <= queueCount_3_14 + counterUpdate_115;
      if (queueEnq_14[4] ^ queueDeq_14[4])
        queueCount_4_14 <= queueCount_4_14 + counterUpdate_116;
      if (queueEnq_14[5] ^ queueDeq_14[5])
        queueCount_5_14 <= queueCount_5_14 + counterUpdate_117;
      if (queueEnq_14[6] ^ queueDeq_14[6])
        queueCount_6_14 <= queueCount_6_14 + counterUpdate_118;
      if (queueEnq_14[7] ^ queueDeq_14[7])
        queueCount_7_14 <= queueCount_7_14 + counterUpdate_119;
      if (queueEnq_15[0] ^ queueDeq_15[0])
        queueCount_0_15 <= queueCount_0_15 + counterUpdate_120;
      if (queueEnq_15[1] ^ queueDeq_15[1])
        queueCount_1_15 <= queueCount_1_15 + counterUpdate_121;
      if (queueEnq_15[2] ^ queueDeq_15[2])
        queueCount_2_15 <= queueCount_2_15 + counterUpdate_122;
      if (queueEnq_15[3] ^ queueDeq_15[3])
        queueCount_3_15 <= queueCount_3_15 + counterUpdate_123;
      if (queueEnq_15[4] ^ queueDeq_15[4])
        queueCount_4_15 <= queueCount_4_15 + counterUpdate_124;
      if (queueEnq_15[5] ^ queueDeq_15[5])
        queueCount_5_15 <= queueCount_5_15 + counterUpdate_125;
      if (queueEnq_15[6] ^ queueDeq_15[6])
        queueCount_6_15 <= queueCount_6_15 + counterUpdate_126;
      if (queueEnq_15[7] ^ queueDeq_15[7])
        queueCount_7_15 <= queueCount_7_15 + counterUpdate_127;
    end
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:91];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [6:0] i = 7'h0; i < 7'h5C; i += 7'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        v0_0 = _RANDOM[7'h0];
        v0_1 = _RANDOM[7'h1];
        v0_2 = _RANDOM[7'h2];
        v0_3 = _RANDOM[7'h3];
        v0_4 = _RANDOM[7'h4];
        v0_5 = _RANDOM[7'h5];
        v0_6 = _RANDOM[7'h6];
        v0_7 = _RANDOM[7'h7];
        v0_8 = _RANDOM[7'h8];
        v0_9 = _RANDOM[7'h9];
        v0_10 = _RANDOM[7'hA];
        v0_11 = _RANDOM[7'hB];
        v0_12 = _RANDOM[7'hC];
        v0_13 = _RANDOM[7'hD];
        v0_14 = _RANDOM[7'hE];
        v0_15 = _RANDOM[7'hF];
        v0_16 = _RANDOM[7'h10];
        v0_17 = _RANDOM[7'h11];
        v0_18 = _RANDOM[7'h12];
        v0_19 = _RANDOM[7'h13];
        v0_20 = _RANDOM[7'h14];
        v0_21 = _RANDOM[7'h15];
        v0_22 = _RANDOM[7'h16];
        v0_23 = _RANDOM[7'h17];
        v0_24 = _RANDOM[7'h18];
        v0_25 = _RANDOM[7'h19];
        v0_26 = _RANDOM[7'h1A];
        v0_27 = _RANDOM[7'h1B];
        v0_28 = _RANDOM[7'h1C];
        v0_29 = _RANDOM[7'h1D];
        v0_30 = _RANDOM[7'h1E];
        v0_31 = _RANDOM[7'h1F];
        v0_32 = _RANDOM[7'h20];
        v0_33 = _RANDOM[7'h21];
        v0_34 = _RANDOM[7'h22];
        v0_35 = _RANDOM[7'h23];
        v0_36 = _RANDOM[7'h24];
        v0_37 = _RANDOM[7'h25];
        v0_38 = _RANDOM[7'h26];
        v0_39 = _RANDOM[7'h27];
        v0_40 = _RANDOM[7'h28];
        v0_41 = _RANDOM[7'h29];
        v0_42 = _RANDOM[7'h2A];
        v0_43 = _RANDOM[7'h2B];
        v0_44 = _RANDOM[7'h2C];
        v0_45 = _RANDOM[7'h2D];
        v0_46 = _RANDOM[7'h2E];
        v0_47 = _RANDOM[7'h2F];
        v0_48 = _RANDOM[7'h30];
        v0_49 = _RANDOM[7'h31];
        v0_50 = _RANDOM[7'h32];
        v0_51 = _RANDOM[7'h33];
        v0_52 = _RANDOM[7'h34];
        v0_53 = _RANDOM[7'h35];
        v0_54 = _RANDOM[7'h36];
        v0_55 = _RANDOM[7'h37];
        v0_56 = _RANDOM[7'h38];
        v0_57 = _RANDOM[7'h39];
        v0_58 = _RANDOM[7'h3A];
        v0_59 = _RANDOM[7'h3B];
        v0_60 = _RANDOM[7'h3C];
        v0_61 = _RANDOM[7'h3D];
        v0_62 = _RANDOM[7'h3E];
        v0_63 = _RANDOM[7'h3F];
        queueCount_0 = _RANDOM[7'h40][6:0];
        queueCount_1 = _RANDOM[7'h40][13:7];
        queueCount_2 = _RANDOM[7'h40][20:14];
        queueCount_3 = _RANDOM[7'h40][27:21];
        queueCount_4 = {_RANDOM[7'h40][31:28], _RANDOM[7'h41][2:0]};
        queueCount_5 = _RANDOM[7'h41][9:3];
        queueCount_6 = _RANDOM[7'h41][16:10];
        queueCount_7 = _RANDOM[7'h41][23:17];
        queueCount_0_1 = _RANDOM[7'h41][30:24];
        queueCount_1_1 = {_RANDOM[7'h41][31], _RANDOM[7'h42][5:0]};
        queueCount_2_1 = _RANDOM[7'h42][12:6];
        queueCount_3_1 = _RANDOM[7'h42][19:13];
        queueCount_4_1 = _RANDOM[7'h42][26:20];
        queueCount_5_1 = {_RANDOM[7'h42][31:27], _RANDOM[7'h43][1:0]};
        queueCount_6_1 = _RANDOM[7'h43][8:2];
        queueCount_7_1 = _RANDOM[7'h43][15:9];
        queueCount_0_2 = _RANDOM[7'h43][22:16];
        queueCount_1_2 = _RANDOM[7'h43][29:23];
        queueCount_2_2 = {_RANDOM[7'h43][31:30], _RANDOM[7'h44][4:0]};
        queueCount_3_2 = _RANDOM[7'h44][11:5];
        queueCount_4_2 = _RANDOM[7'h44][18:12];
        queueCount_5_2 = _RANDOM[7'h44][25:19];
        queueCount_6_2 = {_RANDOM[7'h44][31:26], _RANDOM[7'h45][0]};
        queueCount_7_2 = _RANDOM[7'h45][7:1];
        queueCount_0_3 = _RANDOM[7'h45][14:8];
        queueCount_1_3 = _RANDOM[7'h45][21:15];
        queueCount_2_3 = _RANDOM[7'h45][28:22];
        queueCount_3_3 = {_RANDOM[7'h45][31:29], _RANDOM[7'h46][3:0]};
        queueCount_4_3 = _RANDOM[7'h46][10:4];
        queueCount_5_3 = _RANDOM[7'h46][17:11];
        queueCount_6_3 = _RANDOM[7'h46][24:18];
        queueCount_7_3 = _RANDOM[7'h46][31:25];
        queueCount_0_4 = _RANDOM[7'h47][6:0];
        queueCount_1_4 = _RANDOM[7'h47][13:7];
        queueCount_2_4 = _RANDOM[7'h47][20:14];
        queueCount_3_4 = _RANDOM[7'h47][27:21];
        queueCount_4_4 = {_RANDOM[7'h47][31:28], _RANDOM[7'h48][2:0]};
        queueCount_5_4 = _RANDOM[7'h48][9:3];
        queueCount_6_4 = _RANDOM[7'h48][16:10];
        queueCount_7_4 = _RANDOM[7'h48][23:17];
        queueCount_0_5 = _RANDOM[7'h48][30:24];
        queueCount_1_5 = {_RANDOM[7'h48][31], _RANDOM[7'h49][5:0]};
        queueCount_2_5 = _RANDOM[7'h49][12:6];
        queueCount_3_5 = _RANDOM[7'h49][19:13];
        queueCount_4_5 = _RANDOM[7'h49][26:20];
        queueCount_5_5 = {_RANDOM[7'h49][31:27], _RANDOM[7'h4A][1:0]};
        queueCount_6_5 = _RANDOM[7'h4A][8:2];
        queueCount_7_5 = _RANDOM[7'h4A][15:9];
        queueCount_0_6 = _RANDOM[7'h4A][22:16];
        queueCount_1_6 = _RANDOM[7'h4A][29:23];
        queueCount_2_6 = {_RANDOM[7'h4A][31:30], _RANDOM[7'h4B][4:0]};
        queueCount_3_6 = _RANDOM[7'h4B][11:5];
        queueCount_4_6 = _RANDOM[7'h4B][18:12];
        queueCount_5_6 = _RANDOM[7'h4B][25:19];
        queueCount_6_6 = {_RANDOM[7'h4B][31:26], _RANDOM[7'h4C][0]};
        queueCount_7_6 = _RANDOM[7'h4C][7:1];
        queueCount_0_7 = _RANDOM[7'h4C][14:8];
        queueCount_1_7 = _RANDOM[7'h4C][21:15];
        queueCount_2_7 = _RANDOM[7'h4C][28:22];
        queueCount_3_7 = {_RANDOM[7'h4C][31:29], _RANDOM[7'h4D][3:0]};
        queueCount_4_7 = _RANDOM[7'h4D][10:4];
        queueCount_5_7 = _RANDOM[7'h4D][17:11];
        queueCount_6_7 = _RANDOM[7'h4D][24:18];
        queueCount_7_7 = _RANDOM[7'h4D][31:25];
        queueCount_0_8 = _RANDOM[7'h4E][6:0];
        queueCount_1_8 = _RANDOM[7'h4E][13:7];
        queueCount_2_8 = _RANDOM[7'h4E][20:14];
        queueCount_3_8 = _RANDOM[7'h4E][27:21];
        queueCount_4_8 = {_RANDOM[7'h4E][31:28], _RANDOM[7'h4F][2:0]};
        queueCount_5_8 = _RANDOM[7'h4F][9:3];
        queueCount_6_8 = _RANDOM[7'h4F][16:10];
        queueCount_7_8 = _RANDOM[7'h4F][23:17];
        queueCount_0_9 = _RANDOM[7'h4F][30:24];
        queueCount_1_9 = {_RANDOM[7'h4F][31], _RANDOM[7'h50][5:0]};
        queueCount_2_9 = _RANDOM[7'h50][12:6];
        queueCount_3_9 = _RANDOM[7'h50][19:13];
        queueCount_4_9 = _RANDOM[7'h50][26:20];
        queueCount_5_9 = {_RANDOM[7'h50][31:27], _RANDOM[7'h51][1:0]};
        queueCount_6_9 = _RANDOM[7'h51][8:2];
        queueCount_7_9 = _RANDOM[7'h51][15:9];
        queueCount_0_10 = _RANDOM[7'h51][22:16];
        queueCount_1_10 = _RANDOM[7'h51][29:23];
        queueCount_2_10 = {_RANDOM[7'h51][31:30], _RANDOM[7'h52][4:0]};
        queueCount_3_10 = _RANDOM[7'h52][11:5];
        queueCount_4_10 = _RANDOM[7'h52][18:12];
        queueCount_5_10 = _RANDOM[7'h52][25:19];
        queueCount_6_10 = {_RANDOM[7'h52][31:26], _RANDOM[7'h53][0]};
        queueCount_7_10 = _RANDOM[7'h53][7:1];
        queueCount_0_11 = _RANDOM[7'h53][14:8];
        queueCount_1_11 = _RANDOM[7'h53][21:15];
        queueCount_2_11 = _RANDOM[7'h53][28:22];
        queueCount_3_11 = {_RANDOM[7'h53][31:29], _RANDOM[7'h54][3:0]};
        queueCount_4_11 = _RANDOM[7'h54][10:4];
        queueCount_5_11 = _RANDOM[7'h54][17:11];
        queueCount_6_11 = _RANDOM[7'h54][24:18];
        queueCount_7_11 = _RANDOM[7'h54][31:25];
        queueCount_0_12 = _RANDOM[7'h55][6:0];
        queueCount_1_12 = _RANDOM[7'h55][13:7];
        queueCount_2_12 = _RANDOM[7'h55][20:14];
        queueCount_3_12 = _RANDOM[7'h55][27:21];
        queueCount_4_12 = {_RANDOM[7'h55][31:28], _RANDOM[7'h56][2:0]};
        queueCount_5_12 = _RANDOM[7'h56][9:3];
        queueCount_6_12 = _RANDOM[7'h56][16:10];
        queueCount_7_12 = _RANDOM[7'h56][23:17];
        queueCount_0_13 = _RANDOM[7'h56][30:24];
        queueCount_1_13 = {_RANDOM[7'h56][31], _RANDOM[7'h57][5:0]};
        queueCount_2_13 = _RANDOM[7'h57][12:6];
        queueCount_3_13 = _RANDOM[7'h57][19:13];
        queueCount_4_13 = _RANDOM[7'h57][26:20];
        queueCount_5_13 = {_RANDOM[7'h57][31:27], _RANDOM[7'h58][1:0]};
        queueCount_6_13 = _RANDOM[7'h58][8:2];
        queueCount_7_13 = _RANDOM[7'h58][15:9];
        queueCount_0_14 = _RANDOM[7'h58][22:16];
        queueCount_1_14 = _RANDOM[7'h58][29:23];
        queueCount_2_14 = {_RANDOM[7'h58][31:30], _RANDOM[7'h59][4:0]};
        queueCount_3_14 = _RANDOM[7'h59][11:5];
        queueCount_4_14 = _RANDOM[7'h59][18:12];
        queueCount_5_14 = _RANDOM[7'h59][25:19];
        queueCount_6_14 = {_RANDOM[7'h59][31:26], _RANDOM[7'h5A][0]};
        queueCount_7_14 = _RANDOM[7'h5A][7:1];
        queueCount_0_15 = _RANDOM[7'h5A][14:8];
        queueCount_1_15 = _RANDOM[7'h5A][21:15];
        queueCount_2_15 = _RANDOM[7'h5A][28:22];
        queueCount_3_15 = {_RANDOM[7'h5A][31:29], _RANDOM[7'h5B][3:0]};
        queueCount_4_15 = _RANDOM[7'h5B][10:4];
        queueCount_5_15 = _RANDOM[7'h5B][17:11];
        queueCount_6_15 = _RANDOM[7'h5B][24:18];
        queueCount_7_15 = _RANDOM[7'h5B][31:25];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  wire [5:0]        sourceQueue_deq_bits;
  wire [31:0]       axi4Port_aw_bits_addr_0;
  assign axi4Port_aw_bits_addr_0 = _storeUnit_memRequest_bits_address;
  assign dataQueue_enq_bits_index = _storeUnit_memRequest_bits_index;
  assign dataQueue_enq_bits_address = _storeUnit_memRequest_bits_address;
  wire [8:0]        simpleSourceQueue_deq_bits;
  wire [31:0]       simpleAccessPorts_aw_bits_addr_0;
  assign simpleAccessPorts_aw_bits_addr_0 = _otherUnit_memWriteRequest_bits_address;
  wire [15:0]       otherUnitTargetQueue_enq_bits;
  assign otherUnitTargetQueue_enq_bits = _otherUnit_status_targetLane;
  assign simpleDataQueue_enq_bits_source = _otherUnit_memWriteRequest_bits_source;
  assign simpleDataQueue_enq_bits_address = _otherUnit_memWriteRequest_bits_address;
  assign simpleDataQueue_enq_bits_size = _otherUnit_memWriteRequest_bits_size;
  wire              writeQueueVec_0_empty;
  assign writeQueueVec_0_empty = _writeQueueVec_fifo_empty;
  wire              writeQueueVec_0_full;
  assign writeQueueVec_0_full = _writeQueueVec_fifo_full;
  wire              writeQueueVec_1_empty;
  assign writeQueueVec_1_empty = _writeQueueVec_fifo_1_empty;
  wire              writeQueueVec_1_full;
  assign writeQueueVec_1_full = _writeQueueVec_fifo_1_full;
  wire              writeQueueVec_2_empty;
  assign writeQueueVec_2_empty = _writeQueueVec_fifo_2_empty;
  wire              writeQueueVec_2_full;
  assign writeQueueVec_2_full = _writeQueueVec_fifo_2_full;
  wire              writeQueueVec_3_empty;
  assign writeQueueVec_3_empty = _writeQueueVec_fifo_3_empty;
  wire              writeQueueVec_3_full;
  assign writeQueueVec_3_full = _writeQueueVec_fifo_3_full;
  wire              writeQueueVec_4_empty;
  assign writeQueueVec_4_empty = _writeQueueVec_fifo_4_empty;
  wire              writeQueueVec_4_full;
  assign writeQueueVec_4_full = _writeQueueVec_fifo_4_full;
  wire              writeQueueVec_5_empty;
  assign writeQueueVec_5_empty = _writeQueueVec_fifo_5_empty;
  wire              writeQueueVec_5_full;
  assign writeQueueVec_5_full = _writeQueueVec_fifo_5_full;
  wire              writeQueueVec_6_empty;
  assign writeQueueVec_6_empty = _writeQueueVec_fifo_6_empty;
  wire              writeQueueVec_6_full;
  assign writeQueueVec_6_full = _writeQueueVec_fifo_6_full;
  wire              writeQueueVec_7_empty;
  assign writeQueueVec_7_empty = _writeQueueVec_fifo_7_empty;
  wire              writeQueueVec_7_full;
  assign writeQueueVec_7_full = _writeQueueVec_fifo_7_full;
  wire              writeQueueVec_8_empty;
  assign writeQueueVec_8_empty = _writeQueueVec_fifo_8_empty;
  wire              writeQueueVec_8_full;
  assign writeQueueVec_8_full = _writeQueueVec_fifo_8_full;
  wire              writeQueueVec_9_empty;
  assign writeQueueVec_9_empty = _writeQueueVec_fifo_9_empty;
  wire              writeQueueVec_9_full;
  assign writeQueueVec_9_full = _writeQueueVec_fifo_9_full;
  wire              writeQueueVec_10_empty;
  assign writeQueueVec_10_empty = _writeQueueVec_fifo_10_empty;
  wire              writeQueueVec_10_full;
  assign writeQueueVec_10_full = _writeQueueVec_fifo_10_full;
  wire              writeQueueVec_11_empty;
  assign writeQueueVec_11_empty = _writeQueueVec_fifo_11_empty;
  wire              writeQueueVec_11_full;
  assign writeQueueVec_11_full = _writeQueueVec_fifo_11_full;
  wire              writeQueueVec_12_empty;
  assign writeQueueVec_12_empty = _writeQueueVec_fifo_12_empty;
  wire              writeQueueVec_12_full;
  assign writeQueueVec_12_full = _writeQueueVec_fifo_12_full;
  wire              writeQueueVec_13_empty;
  assign writeQueueVec_13_empty = _writeQueueVec_fifo_13_empty;
  wire              writeQueueVec_13_full;
  assign writeQueueVec_13_full = _writeQueueVec_fifo_13_full;
  wire              writeQueueVec_14_empty;
  assign writeQueueVec_14_empty = _writeQueueVec_fifo_14_empty;
  wire              writeQueueVec_14_full;
  assign writeQueueVec_14_full = _writeQueueVec_fifo_14_full;
  wire              writeQueueVec_15_empty;
  assign writeQueueVec_15_empty = _writeQueueVec_fifo_15_empty;
  wire              writeQueueVec_15_full;
  assign writeQueueVec_15_full = _writeQueueVec_fifo_15_full;
  assign otherUnitTargetQueue_empty = _otherUnitTargetQueue_fifo_empty;
  wire              otherUnitTargetQueue_full;
  assign otherUnitTargetQueue_full = _otherUnitTargetQueue_fifo_full;
  wire              otherUnitDataQueueVec_0_empty;
  assign otherUnitDataQueueVec_0_empty = _otherUnitDataQueueVec_fifo_empty;
  wire              otherUnitDataQueueVec_0_full;
  assign otherUnitDataQueueVec_0_full = _otherUnitDataQueueVec_fifo_full;
  wire              otherUnitDataQueueVec_1_empty;
  assign otherUnitDataQueueVec_1_empty = _otherUnitDataQueueVec_fifo_1_empty;
  wire              otherUnitDataQueueVec_1_full;
  assign otherUnitDataQueueVec_1_full = _otherUnitDataQueueVec_fifo_1_full;
  wire              otherUnitDataQueueVec_2_empty;
  assign otherUnitDataQueueVec_2_empty = _otherUnitDataQueueVec_fifo_2_empty;
  wire              otherUnitDataQueueVec_2_full;
  assign otherUnitDataQueueVec_2_full = _otherUnitDataQueueVec_fifo_2_full;
  wire              otherUnitDataQueueVec_3_empty;
  assign otherUnitDataQueueVec_3_empty = _otherUnitDataQueueVec_fifo_3_empty;
  wire              otherUnitDataQueueVec_3_full;
  assign otherUnitDataQueueVec_3_full = _otherUnitDataQueueVec_fifo_3_full;
  wire              otherUnitDataQueueVec_4_empty;
  assign otherUnitDataQueueVec_4_empty = _otherUnitDataQueueVec_fifo_4_empty;
  wire              otherUnitDataQueueVec_4_full;
  assign otherUnitDataQueueVec_4_full = _otherUnitDataQueueVec_fifo_4_full;
  wire              otherUnitDataQueueVec_5_empty;
  assign otherUnitDataQueueVec_5_empty = _otherUnitDataQueueVec_fifo_5_empty;
  wire              otherUnitDataQueueVec_5_full;
  assign otherUnitDataQueueVec_5_full = _otherUnitDataQueueVec_fifo_5_full;
  wire              otherUnitDataQueueVec_6_empty;
  assign otherUnitDataQueueVec_6_empty = _otherUnitDataQueueVec_fifo_6_empty;
  wire              otherUnitDataQueueVec_6_full;
  assign otherUnitDataQueueVec_6_full = _otherUnitDataQueueVec_fifo_6_full;
  wire              otherUnitDataQueueVec_7_empty;
  assign otherUnitDataQueueVec_7_empty = _otherUnitDataQueueVec_fifo_7_empty;
  wire              otherUnitDataQueueVec_7_full;
  assign otherUnitDataQueueVec_7_full = _otherUnitDataQueueVec_fifo_7_full;
  wire              otherUnitDataQueueVec_8_empty;
  assign otherUnitDataQueueVec_8_empty = _otherUnitDataQueueVec_fifo_8_empty;
  wire              otherUnitDataQueueVec_8_full;
  assign otherUnitDataQueueVec_8_full = _otherUnitDataQueueVec_fifo_8_full;
  wire              otherUnitDataQueueVec_9_empty;
  assign otherUnitDataQueueVec_9_empty = _otherUnitDataQueueVec_fifo_9_empty;
  wire              otherUnitDataQueueVec_9_full;
  assign otherUnitDataQueueVec_9_full = _otherUnitDataQueueVec_fifo_9_full;
  wire              otherUnitDataQueueVec_10_empty;
  assign otherUnitDataQueueVec_10_empty = _otherUnitDataQueueVec_fifo_10_empty;
  wire              otherUnitDataQueueVec_10_full;
  assign otherUnitDataQueueVec_10_full = _otherUnitDataQueueVec_fifo_10_full;
  wire              otherUnitDataQueueVec_11_empty;
  assign otherUnitDataQueueVec_11_empty = _otherUnitDataQueueVec_fifo_11_empty;
  wire              otherUnitDataQueueVec_11_full;
  assign otherUnitDataQueueVec_11_full = _otherUnitDataQueueVec_fifo_11_full;
  wire              otherUnitDataQueueVec_12_empty;
  assign otherUnitDataQueueVec_12_empty = _otherUnitDataQueueVec_fifo_12_empty;
  wire              otherUnitDataQueueVec_12_full;
  assign otherUnitDataQueueVec_12_full = _otherUnitDataQueueVec_fifo_12_full;
  wire              otherUnitDataQueueVec_13_empty;
  assign otherUnitDataQueueVec_13_empty = _otherUnitDataQueueVec_fifo_13_empty;
  wire              otherUnitDataQueueVec_13_full;
  assign otherUnitDataQueueVec_13_full = _otherUnitDataQueueVec_fifo_13_full;
  wire              otherUnitDataQueueVec_14_empty;
  assign otherUnitDataQueueVec_14_empty = _otherUnitDataQueueVec_fifo_14_empty;
  wire              otherUnitDataQueueVec_14_full;
  assign otherUnitDataQueueVec_14_full = _otherUnitDataQueueVec_fifo_14_full;
  wire              otherUnitDataQueueVec_15_empty;
  assign otherUnitDataQueueVec_15_empty = _otherUnitDataQueueVec_fifo_15_empty;
  wire              otherUnitDataQueueVec_15_full;
  assign otherUnitDataQueueVec_15_full = _otherUnitDataQueueVec_fifo_15_full;
  wire              writeIndexQueue_empty;
  assign writeIndexQueue_empty = _writeIndexQueue_fifo_empty;
  wire              writeIndexQueue_full;
  assign writeIndexQueue_full = _writeIndexQueue_fifo_full;
  wire              writeIndexQueue_1_empty;
  assign writeIndexQueue_1_empty = _writeIndexQueue_fifo_1_empty;
  wire              writeIndexQueue_1_full;
  assign writeIndexQueue_1_full = _writeIndexQueue_fifo_1_full;
  wire              writeIndexQueue_2_empty;
  assign writeIndexQueue_2_empty = _writeIndexQueue_fifo_2_empty;
  wire              writeIndexQueue_2_full;
  assign writeIndexQueue_2_full = _writeIndexQueue_fifo_2_full;
  wire              writeIndexQueue_3_empty;
  assign writeIndexQueue_3_empty = _writeIndexQueue_fifo_3_empty;
  wire              writeIndexQueue_3_full;
  assign writeIndexQueue_3_full = _writeIndexQueue_fifo_3_full;
  wire              writeIndexQueue_4_empty;
  assign writeIndexQueue_4_empty = _writeIndexQueue_fifo_4_empty;
  wire              writeIndexQueue_4_full;
  assign writeIndexQueue_4_full = _writeIndexQueue_fifo_4_full;
  wire              writeIndexQueue_5_empty;
  assign writeIndexQueue_5_empty = _writeIndexQueue_fifo_5_empty;
  wire              writeIndexQueue_5_full;
  assign writeIndexQueue_5_full = _writeIndexQueue_fifo_5_full;
  wire              writeIndexQueue_6_empty;
  assign writeIndexQueue_6_empty = _writeIndexQueue_fifo_6_empty;
  wire              writeIndexQueue_6_full;
  assign writeIndexQueue_6_full = _writeIndexQueue_fifo_6_full;
  wire              writeIndexQueue_7_empty;
  assign writeIndexQueue_7_empty = _writeIndexQueue_fifo_7_empty;
  wire              writeIndexQueue_7_full;
  assign writeIndexQueue_7_full = _writeIndexQueue_fifo_7_full;
  wire              writeIndexQueue_8_empty;
  assign writeIndexQueue_8_empty = _writeIndexQueue_fifo_8_empty;
  wire              writeIndexQueue_8_full;
  assign writeIndexQueue_8_full = _writeIndexQueue_fifo_8_full;
  wire              writeIndexQueue_9_empty;
  assign writeIndexQueue_9_empty = _writeIndexQueue_fifo_9_empty;
  wire              writeIndexQueue_9_full;
  assign writeIndexQueue_9_full = _writeIndexQueue_fifo_9_full;
  wire              writeIndexQueue_10_empty;
  assign writeIndexQueue_10_empty = _writeIndexQueue_fifo_10_empty;
  wire              writeIndexQueue_10_full;
  assign writeIndexQueue_10_full = _writeIndexQueue_fifo_10_full;
  wire              writeIndexQueue_11_empty;
  assign writeIndexQueue_11_empty = _writeIndexQueue_fifo_11_empty;
  wire              writeIndexQueue_11_full;
  assign writeIndexQueue_11_full = _writeIndexQueue_fifo_11_full;
  wire              writeIndexQueue_12_empty;
  assign writeIndexQueue_12_empty = _writeIndexQueue_fifo_12_empty;
  wire              writeIndexQueue_12_full;
  assign writeIndexQueue_12_full = _writeIndexQueue_fifo_12_full;
  wire              writeIndexQueue_13_empty;
  assign writeIndexQueue_13_empty = _writeIndexQueue_fifo_13_empty;
  wire              writeIndexQueue_13_full;
  assign writeIndexQueue_13_full = _writeIndexQueue_fifo_13_full;
  wire              writeIndexQueue_14_empty;
  assign writeIndexQueue_14_empty = _writeIndexQueue_fifo_14_empty;
  wire              writeIndexQueue_14_full;
  assign writeIndexQueue_14_full = _writeIndexQueue_fifo_14_full;
  wire              writeIndexQueue_15_empty;
  assign writeIndexQueue_15_empty = _writeIndexQueue_fifo_15_empty;
  wire              writeIndexQueue_15_full;
  assign writeIndexQueue_15_full = _writeIndexQueue_fifo_15_full;
  wire              sourceQueue_empty;
  assign sourceQueue_empty = _sourceQueue_fifo_empty;
  wire              sourceQueue_full;
  assign sourceQueue_full = _sourceQueue_fifo_full;
  wire              dataQueue_empty;
  assign dataQueue_empty = _dataQueue_fifo_empty;
  wire              dataQueue_full;
  assign dataQueue_full = _dataQueue_fifo_full;
  wire              simpleSourceQueue_empty;
  assign simpleSourceQueue_empty = _simpleSourceQueue_fifo_empty;
  wire              simpleSourceQueue_full;
  assign simpleSourceQueue_full = _simpleSourceQueue_fifo_full;
  wire              simpleDataQueue_empty;
  assign simpleDataQueue_empty = _simpleDataQueue_fifo_empty;
  wire              simpleDataQueue_full;
  assign simpleDataQueue_full = _simpleDataQueue_fifo_full;
  LoadUnit loadUnit (
    .clock                                                  (clock),
    .reset                                                  (reset),
    .lsuRequest_valid                                       (reqEnq_0),
    .lsuRequest_bits_instructionInformation_nf              (request_bits_instructionInformation_nf_0),
    .lsuRequest_bits_instructionInformation_mew             (request_bits_instructionInformation_mew_0),
    .lsuRequest_bits_instructionInformation_mop             (request_bits_instructionInformation_mop_0),
    .lsuRequest_bits_instructionInformation_lumop           (request_bits_instructionInformation_lumop_0),
    .lsuRequest_bits_instructionInformation_eew             (request_bits_instructionInformation_eew_0),
    .lsuRequest_bits_instructionInformation_vs3             (request_bits_instructionInformation_vs3_0),
    .lsuRequest_bits_instructionInformation_isStore         (request_bits_instructionInformation_isStore_0),
    .lsuRequest_bits_instructionInformation_maskedLoadStore (request_bits_instructionInformation_maskedLoadStore_0),
    .lsuRequest_bits_rs1Data                                (request_bits_rs1Data_0),
    .lsuRequest_bits_rs2Data                                (request_bits_rs2Data_0),
    .lsuRequest_bits_instructionIndex                       (request_bits_instructionIndex_0),
    .csrInterface_vl                                        (csrInterface_vl),
    .csrInterface_vStart                                    (csrInterface_vStart),
    .csrInterface_vlmul                                     (csrInterface_vlmul),
    .csrInterface_vSew                                      (csrInterface_vSew),
    .csrInterface_vxrm                                      (csrInterface_vxrm),
    .csrInterface_vta                                       (csrInterface_vta),
    .csrInterface_vma                                       (csrInterface_vma),
    .maskInput                                              (_GEN_31[maskSelect]),
    .maskSelect_valid                                       (_loadUnit_maskSelect_valid),
    .maskSelect_bits                                        (_loadUnit_maskSelect_bits),
    .addressConflict                                        (stallLoad),
    .memRequest_ready                                       (sourceQueue_enq_ready & axi4Port_ar_ready_0),
    .memRequest_valid                                       (_loadUnit_memRequest_valid),
    .memRequest_bits_src                                    (sourceQueue_enq_bits),
    .memRequest_bits_address                                (axi4Port_ar_bits_addr_0),
    .memResponse_ready                                      (axi4Port_r_ready_0),
    .memResponse_valid                                      (axi4Port_r_valid_0),
    .memResponse_bits_data                                  (axi4Port_r_bits_data_0),
    .memResponse_bits_index                                 (sourceQueue_deq_bits),
    .status_idle                                            (_loadUnit_status_idle),
    .status_last                                            (_loadUnit_status_last),
    .status_instructionIndex                                (_loadUnit_status_instructionIndex),
    .status_changeMaskGroup                                 (/* unused */),
    .status_startAddress                                    (_loadUnit_status_startAddress),
    .status_endAddress                                      (_loadUnit_status_endAddress),
    .vrfWritePort_0_ready                                   (writeQueueVec_0_enq_ready & ~(otherTryToWrite[0])),
    .vrfWritePort_0_valid                                   (_loadUnit_vrfWritePort_0_valid),
    .vrfWritePort_0_bits_vd                                 (_loadUnit_vrfWritePort_0_bits_vd),
    .vrfWritePort_0_bits_offset                             (_loadUnit_vrfWritePort_0_bits_offset),
    .vrfWritePort_0_bits_mask                               (_loadUnit_vrfWritePort_0_bits_mask),
    .vrfWritePort_0_bits_data                               (_loadUnit_vrfWritePort_0_bits_data),
    .vrfWritePort_0_bits_instructionIndex                   (_loadUnit_vrfWritePort_0_bits_instructionIndex),
    .vrfWritePort_1_ready                                   (writeQueueVec_1_enq_ready & ~(otherTryToWrite[1])),
    .vrfWritePort_1_valid                                   (_loadUnit_vrfWritePort_1_valid),
    .vrfWritePort_1_bits_vd                                 (_loadUnit_vrfWritePort_1_bits_vd),
    .vrfWritePort_1_bits_offset                             (_loadUnit_vrfWritePort_1_bits_offset),
    .vrfWritePort_1_bits_mask                               (_loadUnit_vrfWritePort_1_bits_mask),
    .vrfWritePort_1_bits_data                               (_loadUnit_vrfWritePort_1_bits_data),
    .vrfWritePort_1_bits_instructionIndex                   (_loadUnit_vrfWritePort_1_bits_instructionIndex),
    .vrfWritePort_2_ready                                   (writeQueueVec_2_enq_ready & ~(otherTryToWrite[2])),
    .vrfWritePort_2_valid                                   (_loadUnit_vrfWritePort_2_valid),
    .vrfWritePort_2_bits_vd                                 (_loadUnit_vrfWritePort_2_bits_vd),
    .vrfWritePort_2_bits_offset                             (_loadUnit_vrfWritePort_2_bits_offset),
    .vrfWritePort_2_bits_mask                               (_loadUnit_vrfWritePort_2_bits_mask),
    .vrfWritePort_2_bits_data                               (_loadUnit_vrfWritePort_2_bits_data),
    .vrfWritePort_2_bits_instructionIndex                   (_loadUnit_vrfWritePort_2_bits_instructionIndex),
    .vrfWritePort_3_ready                                   (writeQueueVec_3_enq_ready & ~(otherTryToWrite[3])),
    .vrfWritePort_3_valid                                   (_loadUnit_vrfWritePort_3_valid),
    .vrfWritePort_3_bits_vd                                 (_loadUnit_vrfWritePort_3_bits_vd),
    .vrfWritePort_3_bits_offset                             (_loadUnit_vrfWritePort_3_bits_offset),
    .vrfWritePort_3_bits_mask                               (_loadUnit_vrfWritePort_3_bits_mask),
    .vrfWritePort_3_bits_data                               (_loadUnit_vrfWritePort_3_bits_data),
    .vrfWritePort_3_bits_instructionIndex                   (_loadUnit_vrfWritePort_3_bits_instructionIndex),
    .vrfWritePort_4_ready                                   (writeQueueVec_4_enq_ready & ~(otherTryToWrite[4])),
    .vrfWritePort_4_valid                                   (_loadUnit_vrfWritePort_4_valid),
    .vrfWritePort_4_bits_vd                                 (_loadUnit_vrfWritePort_4_bits_vd),
    .vrfWritePort_4_bits_offset                             (_loadUnit_vrfWritePort_4_bits_offset),
    .vrfWritePort_4_bits_mask                               (_loadUnit_vrfWritePort_4_bits_mask),
    .vrfWritePort_4_bits_data                               (_loadUnit_vrfWritePort_4_bits_data),
    .vrfWritePort_4_bits_instructionIndex                   (_loadUnit_vrfWritePort_4_bits_instructionIndex),
    .vrfWritePort_5_ready                                   (writeQueueVec_5_enq_ready & ~(otherTryToWrite[5])),
    .vrfWritePort_5_valid                                   (_loadUnit_vrfWritePort_5_valid),
    .vrfWritePort_5_bits_vd                                 (_loadUnit_vrfWritePort_5_bits_vd),
    .vrfWritePort_5_bits_offset                             (_loadUnit_vrfWritePort_5_bits_offset),
    .vrfWritePort_5_bits_mask                               (_loadUnit_vrfWritePort_5_bits_mask),
    .vrfWritePort_5_bits_data                               (_loadUnit_vrfWritePort_5_bits_data),
    .vrfWritePort_5_bits_instructionIndex                   (_loadUnit_vrfWritePort_5_bits_instructionIndex),
    .vrfWritePort_6_ready                                   (writeQueueVec_6_enq_ready & ~(otherTryToWrite[6])),
    .vrfWritePort_6_valid                                   (_loadUnit_vrfWritePort_6_valid),
    .vrfWritePort_6_bits_vd                                 (_loadUnit_vrfWritePort_6_bits_vd),
    .vrfWritePort_6_bits_offset                             (_loadUnit_vrfWritePort_6_bits_offset),
    .vrfWritePort_6_bits_mask                               (_loadUnit_vrfWritePort_6_bits_mask),
    .vrfWritePort_6_bits_data                               (_loadUnit_vrfWritePort_6_bits_data),
    .vrfWritePort_6_bits_instructionIndex                   (_loadUnit_vrfWritePort_6_bits_instructionIndex),
    .vrfWritePort_7_ready                                   (writeQueueVec_7_enq_ready & ~(otherTryToWrite[7])),
    .vrfWritePort_7_valid                                   (_loadUnit_vrfWritePort_7_valid),
    .vrfWritePort_7_bits_vd                                 (_loadUnit_vrfWritePort_7_bits_vd),
    .vrfWritePort_7_bits_offset                             (_loadUnit_vrfWritePort_7_bits_offset),
    .vrfWritePort_7_bits_mask                               (_loadUnit_vrfWritePort_7_bits_mask),
    .vrfWritePort_7_bits_data                               (_loadUnit_vrfWritePort_7_bits_data),
    .vrfWritePort_7_bits_instructionIndex                   (_loadUnit_vrfWritePort_7_bits_instructionIndex),
    .vrfWritePort_8_ready                                   (writeQueueVec_8_enq_ready & ~(otherTryToWrite[8])),
    .vrfWritePort_8_valid                                   (_loadUnit_vrfWritePort_8_valid),
    .vrfWritePort_8_bits_vd                                 (_loadUnit_vrfWritePort_8_bits_vd),
    .vrfWritePort_8_bits_offset                             (_loadUnit_vrfWritePort_8_bits_offset),
    .vrfWritePort_8_bits_mask                               (_loadUnit_vrfWritePort_8_bits_mask),
    .vrfWritePort_8_bits_data                               (_loadUnit_vrfWritePort_8_bits_data),
    .vrfWritePort_8_bits_instructionIndex                   (_loadUnit_vrfWritePort_8_bits_instructionIndex),
    .vrfWritePort_9_ready                                   (writeQueueVec_9_enq_ready & ~(otherTryToWrite[9])),
    .vrfWritePort_9_valid                                   (_loadUnit_vrfWritePort_9_valid),
    .vrfWritePort_9_bits_vd                                 (_loadUnit_vrfWritePort_9_bits_vd),
    .vrfWritePort_9_bits_offset                             (_loadUnit_vrfWritePort_9_bits_offset),
    .vrfWritePort_9_bits_mask                               (_loadUnit_vrfWritePort_9_bits_mask),
    .vrfWritePort_9_bits_data                               (_loadUnit_vrfWritePort_9_bits_data),
    .vrfWritePort_9_bits_instructionIndex                   (_loadUnit_vrfWritePort_9_bits_instructionIndex),
    .vrfWritePort_10_ready                                  (writeQueueVec_10_enq_ready & ~(otherTryToWrite[10])),
    .vrfWritePort_10_valid                                  (_loadUnit_vrfWritePort_10_valid),
    .vrfWritePort_10_bits_vd                                (_loadUnit_vrfWritePort_10_bits_vd),
    .vrfWritePort_10_bits_offset                            (_loadUnit_vrfWritePort_10_bits_offset),
    .vrfWritePort_10_bits_mask                              (_loadUnit_vrfWritePort_10_bits_mask),
    .vrfWritePort_10_bits_data                              (_loadUnit_vrfWritePort_10_bits_data),
    .vrfWritePort_10_bits_instructionIndex                  (_loadUnit_vrfWritePort_10_bits_instructionIndex),
    .vrfWritePort_11_ready                                  (writeQueueVec_11_enq_ready & ~(otherTryToWrite[11])),
    .vrfWritePort_11_valid                                  (_loadUnit_vrfWritePort_11_valid),
    .vrfWritePort_11_bits_vd                                (_loadUnit_vrfWritePort_11_bits_vd),
    .vrfWritePort_11_bits_offset                            (_loadUnit_vrfWritePort_11_bits_offset),
    .vrfWritePort_11_bits_mask                              (_loadUnit_vrfWritePort_11_bits_mask),
    .vrfWritePort_11_bits_data                              (_loadUnit_vrfWritePort_11_bits_data),
    .vrfWritePort_11_bits_instructionIndex                  (_loadUnit_vrfWritePort_11_bits_instructionIndex),
    .vrfWritePort_12_ready                                  (writeQueueVec_12_enq_ready & ~(otherTryToWrite[12])),
    .vrfWritePort_12_valid                                  (_loadUnit_vrfWritePort_12_valid),
    .vrfWritePort_12_bits_vd                                (_loadUnit_vrfWritePort_12_bits_vd),
    .vrfWritePort_12_bits_offset                            (_loadUnit_vrfWritePort_12_bits_offset),
    .vrfWritePort_12_bits_mask                              (_loadUnit_vrfWritePort_12_bits_mask),
    .vrfWritePort_12_bits_data                              (_loadUnit_vrfWritePort_12_bits_data),
    .vrfWritePort_12_bits_instructionIndex                  (_loadUnit_vrfWritePort_12_bits_instructionIndex),
    .vrfWritePort_13_ready                                  (writeQueueVec_13_enq_ready & ~(otherTryToWrite[13])),
    .vrfWritePort_13_valid                                  (_loadUnit_vrfWritePort_13_valid),
    .vrfWritePort_13_bits_vd                                (_loadUnit_vrfWritePort_13_bits_vd),
    .vrfWritePort_13_bits_offset                            (_loadUnit_vrfWritePort_13_bits_offset),
    .vrfWritePort_13_bits_mask                              (_loadUnit_vrfWritePort_13_bits_mask),
    .vrfWritePort_13_bits_data                              (_loadUnit_vrfWritePort_13_bits_data),
    .vrfWritePort_13_bits_instructionIndex                  (_loadUnit_vrfWritePort_13_bits_instructionIndex),
    .vrfWritePort_14_ready                                  (writeQueueVec_14_enq_ready & ~(otherTryToWrite[14])),
    .vrfWritePort_14_valid                                  (_loadUnit_vrfWritePort_14_valid),
    .vrfWritePort_14_bits_vd                                (_loadUnit_vrfWritePort_14_bits_vd),
    .vrfWritePort_14_bits_offset                            (_loadUnit_vrfWritePort_14_bits_offset),
    .vrfWritePort_14_bits_mask                              (_loadUnit_vrfWritePort_14_bits_mask),
    .vrfWritePort_14_bits_data                              (_loadUnit_vrfWritePort_14_bits_data),
    .vrfWritePort_14_bits_instructionIndex                  (_loadUnit_vrfWritePort_14_bits_instructionIndex),
    .vrfWritePort_15_ready                                  (writeQueueVec_15_enq_ready & ~(otherTryToWrite[15])),
    .vrfWritePort_15_valid                                  (_loadUnit_vrfWritePort_15_valid),
    .vrfWritePort_15_bits_vd                                (_loadUnit_vrfWritePort_15_bits_vd),
    .vrfWritePort_15_bits_offset                            (_loadUnit_vrfWritePort_15_bits_offset),
    .vrfWritePort_15_bits_mask                              (_loadUnit_vrfWritePort_15_bits_mask),
    .vrfWritePort_15_bits_data                              (_loadUnit_vrfWritePort_15_bits_data),
    .vrfWritePort_15_bits_instructionIndex                  (_loadUnit_vrfWritePort_15_bits_instructionIndex)
  );
  StoreUnit storeUnit (
    .clock                                                  (clock),
    .reset                                                  (reset),
    .lsuRequest_valid                                       (reqEnq_1),
    .lsuRequest_bits_instructionInformation_nf              (request_bits_instructionInformation_nf_0),
    .lsuRequest_bits_instructionInformation_mew             (request_bits_instructionInformation_mew_0),
    .lsuRequest_bits_instructionInformation_mop             (request_bits_instructionInformation_mop_0),
    .lsuRequest_bits_instructionInformation_lumop           (request_bits_instructionInformation_lumop_0),
    .lsuRequest_bits_instructionInformation_eew             (request_bits_instructionInformation_eew_0),
    .lsuRequest_bits_instructionInformation_vs3             (request_bits_instructionInformation_vs3_0),
    .lsuRequest_bits_instructionInformation_isStore         (request_bits_instructionInformation_isStore_0),
    .lsuRequest_bits_instructionInformation_maskedLoadStore (request_bits_instructionInformation_maskedLoadStore_0),
    .lsuRequest_bits_rs1Data                                (request_bits_rs1Data_0),
    .lsuRequest_bits_rs2Data                                (request_bits_rs2Data_0),
    .lsuRequest_bits_instructionIndex                       (request_bits_instructionIndex_0),
    .csrInterface_vl                                        (csrInterface_vl),
    .csrInterface_vStart                                    (csrInterface_vStart),
    .csrInterface_vlmul                                     (csrInterface_vlmul),
    .csrInterface_vSew                                      (csrInterface_vSew),
    .csrInterface_vxrm                                      (csrInterface_vxrm),
    .csrInterface_vta                                       (csrInterface_vta),
    .csrInterface_vma                                       (csrInterface_vma),
    .maskInput                                              (_GEN_32[maskSelect_1]),
    .maskSelect_valid                                       (_storeUnit_maskSelect_valid),
    .maskSelect_bits                                        (_storeUnit_maskSelect_bits),
    .memRequest_ready                                       (axi4Port_aw_ready_0 & dataQueue_enq_ready),
    .memRequest_valid                                       (_storeUnit_memRequest_valid),
    .memRequest_bits_data                                   (dataQueue_enq_bits_data),
    .memRequest_bits_mask                                   (dataQueue_enq_bits_mask),
    .memRequest_bits_index                                  (_storeUnit_memRequest_bits_index),
    .memRequest_bits_address                                (_storeUnit_memRequest_bits_address),
    .status_idle                                            (_storeUnit_status_idle),
    .status_last                                            (_storeUnit_status_last),
    .status_instructionIndex                                (_storeUnit_status_instructionIndex),
    .status_changeMaskGroup                                 (/* unused */),
    .status_startAddress                                    (_storeUnit_status_startAddress),
    .status_endAddress                                      (_storeUnit_status_endAddress),
    .vrfReadDataPorts_0_ready                               (vrfReadDataPorts_0_ready_0 & ~(otherTryReadVrf[0])),
    .vrfReadDataPorts_0_valid                               (_storeUnit_vrfReadDataPorts_0_valid),
    .vrfReadDataPorts_0_bits_vs                             (_storeUnit_vrfReadDataPorts_0_bits_vs),
    .vrfReadDataPorts_0_bits_offset                         (_storeUnit_vrfReadDataPorts_0_bits_offset),
    .vrfReadDataPorts_0_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_0_bits_instructionIndex),
    .vrfReadDataPorts_1_ready                               (vrfReadDataPorts_1_ready_0 & ~(otherTryReadVrf[1])),
    .vrfReadDataPorts_1_valid                               (_storeUnit_vrfReadDataPorts_1_valid),
    .vrfReadDataPorts_1_bits_vs                             (_storeUnit_vrfReadDataPorts_1_bits_vs),
    .vrfReadDataPorts_1_bits_offset                         (_storeUnit_vrfReadDataPorts_1_bits_offset),
    .vrfReadDataPorts_1_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_1_bits_instructionIndex),
    .vrfReadDataPorts_2_ready                               (vrfReadDataPorts_2_ready_0 & ~(otherTryReadVrf[2])),
    .vrfReadDataPorts_2_valid                               (_storeUnit_vrfReadDataPorts_2_valid),
    .vrfReadDataPorts_2_bits_vs                             (_storeUnit_vrfReadDataPorts_2_bits_vs),
    .vrfReadDataPorts_2_bits_offset                         (_storeUnit_vrfReadDataPorts_2_bits_offset),
    .vrfReadDataPorts_2_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_2_bits_instructionIndex),
    .vrfReadDataPorts_3_ready                               (vrfReadDataPorts_3_ready_0 & ~(otherTryReadVrf[3])),
    .vrfReadDataPorts_3_valid                               (_storeUnit_vrfReadDataPorts_3_valid),
    .vrfReadDataPorts_3_bits_vs                             (_storeUnit_vrfReadDataPorts_3_bits_vs),
    .vrfReadDataPorts_3_bits_offset                         (_storeUnit_vrfReadDataPorts_3_bits_offset),
    .vrfReadDataPorts_3_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_3_bits_instructionIndex),
    .vrfReadDataPorts_4_ready                               (vrfReadDataPorts_4_ready_0 & ~(otherTryReadVrf[4])),
    .vrfReadDataPorts_4_valid                               (_storeUnit_vrfReadDataPorts_4_valid),
    .vrfReadDataPorts_4_bits_vs                             (_storeUnit_vrfReadDataPorts_4_bits_vs),
    .vrfReadDataPorts_4_bits_offset                         (_storeUnit_vrfReadDataPorts_4_bits_offset),
    .vrfReadDataPorts_4_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_4_bits_instructionIndex),
    .vrfReadDataPorts_5_ready                               (vrfReadDataPorts_5_ready_0 & ~(otherTryReadVrf[5])),
    .vrfReadDataPorts_5_valid                               (_storeUnit_vrfReadDataPorts_5_valid),
    .vrfReadDataPorts_5_bits_vs                             (_storeUnit_vrfReadDataPorts_5_bits_vs),
    .vrfReadDataPorts_5_bits_offset                         (_storeUnit_vrfReadDataPorts_5_bits_offset),
    .vrfReadDataPorts_5_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_5_bits_instructionIndex),
    .vrfReadDataPorts_6_ready                               (vrfReadDataPorts_6_ready_0 & ~(otherTryReadVrf[6])),
    .vrfReadDataPorts_6_valid                               (_storeUnit_vrfReadDataPorts_6_valid),
    .vrfReadDataPorts_6_bits_vs                             (_storeUnit_vrfReadDataPorts_6_bits_vs),
    .vrfReadDataPorts_6_bits_offset                         (_storeUnit_vrfReadDataPorts_6_bits_offset),
    .vrfReadDataPorts_6_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_6_bits_instructionIndex),
    .vrfReadDataPorts_7_ready                               (vrfReadDataPorts_7_ready_0 & ~(otherTryReadVrf[7])),
    .vrfReadDataPorts_7_valid                               (_storeUnit_vrfReadDataPorts_7_valid),
    .vrfReadDataPorts_7_bits_vs                             (_storeUnit_vrfReadDataPorts_7_bits_vs),
    .vrfReadDataPorts_7_bits_offset                         (_storeUnit_vrfReadDataPorts_7_bits_offset),
    .vrfReadDataPorts_7_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_7_bits_instructionIndex),
    .vrfReadDataPorts_8_ready                               (vrfReadDataPorts_8_ready_0 & ~(otherTryReadVrf[8])),
    .vrfReadDataPorts_8_valid                               (_storeUnit_vrfReadDataPorts_8_valid),
    .vrfReadDataPorts_8_bits_vs                             (_storeUnit_vrfReadDataPorts_8_bits_vs),
    .vrfReadDataPorts_8_bits_offset                         (_storeUnit_vrfReadDataPorts_8_bits_offset),
    .vrfReadDataPorts_8_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_8_bits_instructionIndex),
    .vrfReadDataPorts_9_ready                               (vrfReadDataPorts_9_ready_0 & ~(otherTryReadVrf[9])),
    .vrfReadDataPorts_9_valid                               (_storeUnit_vrfReadDataPorts_9_valid),
    .vrfReadDataPorts_9_bits_vs                             (_storeUnit_vrfReadDataPorts_9_bits_vs),
    .vrfReadDataPorts_9_bits_offset                         (_storeUnit_vrfReadDataPorts_9_bits_offset),
    .vrfReadDataPorts_9_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_9_bits_instructionIndex),
    .vrfReadDataPorts_10_ready                              (vrfReadDataPorts_10_ready_0 & ~(otherTryReadVrf[10])),
    .vrfReadDataPorts_10_valid                              (_storeUnit_vrfReadDataPorts_10_valid),
    .vrfReadDataPorts_10_bits_vs                            (_storeUnit_vrfReadDataPorts_10_bits_vs),
    .vrfReadDataPorts_10_bits_offset                        (_storeUnit_vrfReadDataPorts_10_bits_offset),
    .vrfReadDataPorts_10_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_10_bits_instructionIndex),
    .vrfReadDataPorts_11_ready                              (vrfReadDataPorts_11_ready_0 & ~(otherTryReadVrf[11])),
    .vrfReadDataPorts_11_valid                              (_storeUnit_vrfReadDataPorts_11_valid),
    .vrfReadDataPorts_11_bits_vs                            (_storeUnit_vrfReadDataPorts_11_bits_vs),
    .vrfReadDataPorts_11_bits_offset                        (_storeUnit_vrfReadDataPorts_11_bits_offset),
    .vrfReadDataPorts_11_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_11_bits_instructionIndex),
    .vrfReadDataPorts_12_ready                              (vrfReadDataPorts_12_ready_0 & ~(otherTryReadVrf[12])),
    .vrfReadDataPorts_12_valid                              (_storeUnit_vrfReadDataPorts_12_valid),
    .vrfReadDataPorts_12_bits_vs                            (_storeUnit_vrfReadDataPorts_12_bits_vs),
    .vrfReadDataPorts_12_bits_offset                        (_storeUnit_vrfReadDataPorts_12_bits_offset),
    .vrfReadDataPorts_12_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_12_bits_instructionIndex),
    .vrfReadDataPorts_13_ready                              (vrfReadDataPorts_13_ready_0 & ~(otherTryReadVrf[13])),
    .vrfReadDataPorts_13_valid                              (_storeUnit_vrfReadDataPorts_13_valid),
    .vrfReadDataPorts_13_bits_vs                            (_storeUnit_vrfReadDataPorts_13_bits_vs),
    .vrfReadDataPorts_13_bits_offset                        (_storeUnit_vrfReadDataPorts_13_bits_offset),
    .vrfReadDataPorts_13_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_13_bits_instructionIndex),
    .vrfReadDataPorts_14_ready                              (vrfReadDataPorts_14_ready_0 & ~(otherTryReadVrf[14])),
    .vrfReadDataPorts_14_valid                              (_storeUnit_vrfReadDataPorts_14_valid),
    .vrfReadDataPorts_14_bits_vs                            (_storeUnit_vrfReadDataPorts_14_bits_vs),
    .vrfReadDataPorts_14_bits_offset                        (_storeUnit_vrfReadDataPorts_14_bits_offset),
    .vrfReadDataPorts_14_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_14_bits_instructionIndex),
    .vrfReadDataPorts_15_ready                              (vrfReadDataPorts_15_ready_0 & ~(otherTryReadVrf[15])),
    .vrfReadDataPorts_15_valid                              (_storeUnit_vrfReadDataPorts_15_valid),
    .vrfReadDataPorts_15_bits_vs                            (_storeUnit_vrfReadDataPorts_15_bits_vs),
    .vrfReadDataPorts_15_bits_offset                        (_storeUnit_vrfReadDataPorts_15_bits_offset),
    .vrfReadDataPorts_15_bits_instructionIndex              (_storeUnit_vrfReadDataPorts_15_bits_instructionIndex),
    .vrfReadResults_0_valid                                 (vrfReadResults_0_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_0_bits                                  (vrfReadResults_0_bits),
    .vrfReadResults_1_valid                                 (vrfReadResults_1_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_1_bits                                  (vrfReadResults_1_bits),
    .vrfReadResults_2_valid                                 (vrfReadResults_2_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_2_bits                                  (vrfReadResults_2_bits),
    .vrfReadResults_3_valid                                 (vrfReadResults_3_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_3_bits                                  (vrfReadResults_3_bits),
    .vrfReadResults_4_valid                                 (vrfReadResults_4_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_4_bits                                  (vrfReadResults_4_bits),
    .vrfReadResults_5_valid                                 (vrfReadResults_5_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_5_bits                                  (vrfReadResults_5_bits),
    .vrfReadResults_6_valid                                 (vrfReadResults_6_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_6_bits                                  (vrfReadResults_6_bits),
    .vrfReadResults_7_valid                                 (vrfReadResults_7_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_7_bits                                  (vrfReadResults_7_bits),
    .vrfReadResults_8_valid                                 (vrfReadResults_8_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_8_bits                                  (vrfReadResults_8_bits),
    .vrfReadResults_9_valid                                 (vrfReadResults_9_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_9_bits                                  (vrfReadResults_9_bits),
    .vrfReadResults_10_valid                                (vrfReadResults_10_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_10_bits                                 (vrfReadResults_10_bits),
    .vrfReadResults_11_valid                                (vrfReadResults_11_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_11_bits                                 (vrfReadResults_11_bits),
    .vrfReadResults_12_valid                                (vrfReadResults_12_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_12_bits                                 (vrfReadResults_12_bits),
    .vrfReadResults_13_valid                                (vrfReadResults_13_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_13_bits                                 (vrfReadResults_13_bits),
    .vrfReadResults_14_valid                                (vrfReadResults_14_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_14_bits                                 (vrfReadResults_14_bits),
    .vrfReadResults_15_valid                                (vrfReadResults_15_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_15_bits                                 (vrfReadResults_15_bits),
    .storeResponse                                          (axi4Port_b_valid_0)
  );
  SimpleAccessUnit otherUnit (
    .clock                                                  (clock),
    .reset                                                  (reset),
    .lsuRequest_valid                                       (reqEnq_2),
    .lsuRequest_bits_instructionInformation_nf              (request_bits_instructionInformation_nf_0),
    .lsuRequest_bits_instructionInformation_mew             (request_bits_instructionInformation_mew_0),
    .lsuRequest_bits_instructionInformation_mop             (request_bits_instructionInformation_mop_0),
    .lsuRequest_bits_instructionInformation_lumop           (request_bits_instructionInformation_lumop_0),
    .lsuRequest_bits_instructionInformation_eew             (request_bits_instructionInformation_eew_0),
    .lsuRequest_bits_instructionInformation_vs3             (request_bits_instructionInformation_vs3_0),
    .lsuRequest_bits_instructionInformation_isStore         (request_bits_instructionInformation_isStore_0),
    .lsuRequest_bits_instructionInformation_maskedLoadStore (request_bits_instructionInformation_maskedLoadStore_0),
    .lsuRequest_bits_rs1Data                                (request_bits_rs1Data_0),
    .lsuRequest_bits_rs2Data                                (request_bits_rs2Data_0),
    .lsuRequest_bits_instructionIndex                       (request_bits_instructionIndex_0),
    .vrfReadDataPorts_ready                                 (otherUnit_vrfReadDataPorts_ready),
    .vrfReadDataPorts_valid                                 (_otherUnit_vrfReadDataPorts_valid),
    .vrfReadDataPorts_bits_vs                               (_otherUnit_vrfReadDataPorts_bits_vs),
    .vrfReadDataPorts_bits_offset                           (_otherUnit_vrfReadDataPorts_bits_offset),
    .vrfReadDataPorts_bits_instructionIndex                 (_otherUnit_vrfReadDataPorts_bits_instructionIndex),
    .vrfReadResults_valid                                   (otherUnitTargetQueue_deq_ready),
    .vrfReadResults_bits
      ((otherUnitTargetQueue_deq_bits[0] ? otherUnitDataQueueVec_0_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[1] ? otherUnitDataQueueVec_1_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[2] ? otherUnitDataQueueVec_2_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[3] ? otherUnitDataQueueVec_3_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[4] ? otherUnitDataQueueVec_4_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[5] ? otherUnitDataQueueVec_5_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[6] ? otherUnitDataQueueVec_6_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[7] ? otherUnitDataQueueVec_7_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[8] ? otherUnitDataQueueVec_8_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[9] ? otherUnitDataQueueVec_9_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[10] ? otherUnitDataQueueVec_10_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[11] ? otherUnitDataQueueVec_11_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[12] ? otherUnitDataQueueVec_12_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[13] ? otherUnitDataQueueVec_13_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[14] ? otherUnitDataQueueVec_14_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[15] ? otherUnitDataQueueVec_15_deq_bits : 32'h0)),
    .offsetReadResult_0_valid                               (offsetReadResult_0_valid),
    .offsetReadResult_0_bits                                (offsetReadResult_0_bits),
    .offsetReadResult_1_valid                               (offsetReadResult_1_valid),
    .offsetReadResult_1_bits                                (offsetReadResult_1_bits),
    .offsetReadResult_2_valid                               (offsetReadResult_2_valid),
    .offsetReadResult_2_bits                                (offsetReadResult_2_bits),
    .offsetReadResult_3_valid                               (offsetReadResult_3_valid),
    .offsetReadResult_3_bits                                (offsetReadResult_3_bits),
    .offsetReadResult_4_valid                               (offsetReadResult_4_valid),
    .offsetReadResult_4_bits                                (offsetReadResult_4_bits),
    .offsetReadResult_5_valid                               (offsetReadResult_5_valid),
    .offsetReadResult_5_bits                                (offsetReadResult_5_bits),
    .offsetReadResult_6_valid                               (offsetReadResult_6_valid),
    .offsetReadResult_6_bits                                (offsetReadResult_6_bits),
    .offsetReadResult_7_valid                               (offsetReadResult_7_valid),
    .offsetReadResult_7_bits                                (offsetReadResult_7_bits),
    .offsetReadResult_8_valid                               (offsetReadResult_8_valid),
    .offsetReadResult_8_bits                                (offsetReadResult_8_bits),
    .offsetReadResult_9_valid                               (offsetReadResult_9_valid),
    .offsetReadResult_9_bits                                (offsetReadResult_9_bits),
    .offsetReadResult_10_valid                              (offsetReadResult_10_valid),
    .offsetReadResult_10_bits                               (offsetReadResult_10_bits),
    .offsetReadResult_11_valid                              (offsetReadResult_11_valid),
    .offsetReadResult_11_bits                               (offsetReadResult_11_bits),
    .offsetReadResult_12_valid                              (offsetReadResult_12_valid),
    .offsetReadResult_12_bits                               (offsetReadResult_12_bits),
    .offsetReadResult_13_valid                              (offsetReadResult_13_valid),
    .offsetReadResult_13_bits                               (offsetReadResult_13_bits),
    .offsetReadResult_14_valid                              (offsetReadResult_14_valid),
    .offsetReadResult_14_bits                               (offsetReadResult_14_bits),
    .offsetReadResult_15_valid                              (offsetReadResult_15_valid),
    .offsetReadResult_15_bits                               (offsetReadResult_15_bits),
    .maskInput                                              (_GEN_33[maskSelect_2]),
    .maskSelect_valid                                       (_otherUnit_maskSelect_valid),
    .maskSelect_bits                                        (_otherUnit_maskSelect_bits),
    .memReadRequest_ready                                   (simpleSourceQueue_enq_ready & simpleAccessPorts_ar_ready_0),
    .memReadRequest_valid                                   (_otherUnit_memReadRequest_valid),
    .memReadRequest_bits_address                            (simpleAccessPorts_ar_bits_addr_0),
    .memReadRequest_bits_source                             (simpleSourceQueue_enq_bits),
    .memReadResponse_ready                                  (simpleAccessPorts_r_ready_0),
    .memReadResponse_valid                                  (simpleAccessPorts_r_valid_0),
    .memReadResponse_bits_data                              (simpleAccessPorts_r_bits_data_0),
    .memReadResponse_bits_source                            (simpleSourceQueue_deq_bits),
    .memWriteRequest_ready                                  (simpleAccessPorts_aw_ready_0 & simpleDataQueue_enq_ready),
    .memWriteRequest_valid                                  (_otherUnit_memWriteRequest_valid),
    .memWriteRequest_bits_data                              (simpleDataQueue_enq_bits_data),
    .memWriteRequest_bits_mask                              (simpleDataQueue_enq_bits_mask),
    .memWriteRequest_bits_source                            (_otherUnit_memWriteRequest_bits_source),
    .memWriteRequest_bits_address                           (_otherUnit_memWriteRequest_bits_address),
    .memWriteRequest_bits_size                              (_otherUnit_memWriteRequest_bits_size),
    .vrfWritePort_ready                                     (|(_otherUnit_status_targetLane & {otherUnit_vrfWritePort_ready_hi, otherUnit_vrfWritePort_ready_lo})),
    .vrfWritePort_valid                                     (_otherUnit_vrfWritePort_valid),
    .vrfWritePort_bits_vd                                   (_otherUnit_vrfWritePort_bits_vd),
    .vrfWritePort_bits_offset                               (_otherUnit_vrfWritePort_bits_offset),
    .vrfWritePort_bits_mask                                 (_otherUnit_vrfWritePort_bits_mask),
    .vrfWritePort_bits_data                                 (_otherUnit_vrfWritePort_bits_data),
    .vrfWritePort_bits_last                                 (_otherUnit_vrfWritePort_bits_last),
    .vrfWritePort_bits_instructionIndex                     (_otherUnit_vrfWritePort_bits_instructionIndex),
    .csrInterface_vl                                        (csrInterface_vl),
    .csrInterface_vStart                                    (csrInterface_vStart),
    .csrInterface_vlmul                                     (csrInterface_vlmul),
    .csrInterface_vSew                                      (csrInterface_vSew),
    .csrInterface_vxrm                                      (csrInterface_vxrm),
    .csrInterface_vta                                       (csrInterface_vta),
    .csrInterface_vma                                       (csrInterface_vma),
    .status_idle                                            (_otherUnit_status_idle),
    .status_last                                            (_otherUnit_status_last),
    .status_instructionIndex                                (_otherUnit_status_instructionIndex),
    .status_targetLane                                      (_otherUnit_status_targetLane),
    .status_isStore                                         (_otherUnit_status_isStore),
    .offsetRelease_0                                        (_otherUnit_offsetRelease_0),
    .offsetRelease_1                                        (_otherUnit_offsetRelease_1),
    .offsetRelease_2                                        (_otherUnit_offsetRelease_2),
    .offsetRelease_3                                        (_otherUnit_offsetRelease_3),
    .offsetRelease_4                                        (_otherUnit_offsetRelease_4),
    .offsetRelease_5                                        (_otherUnit_offsetRelease_5),
    .offsetRelease_6                                        (_otherUnit_offsetRelease_6),
    .offsetRelease_7                                        (_otherUnit_offsetRelease_7),
    .offsetRelease_8                                        (_otherUnit_offsetRelease_8),
    .offsetRelease_9                                        (_otherUnit_offsetRelease_9),
    .offsetRelease_10                                       (_otherUnit_offsetRelease_10),
    .offsetRelease_11                                       (_otherUnit_offsetRelease_11),
    .offsetRelease_12                                       (_otherUnit_offsetRelease_12),
    .offsetRelease_13                                       (_otherUnit_offsetRelease_13),
    .offsetRelease_14                                       (_otherUnit_offsetRelease_14),
    .offsetRelease_15                                       (_otherUnit_offsetRelease_15)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(63)
  ) writeQueueVec_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_0_writeValid_T & ~(_writeQueueVec_fifo_empty & writeQueueVec_0_deq_ready))),
    .pop_req_n    (~(writeQueueVec_0_deq_ready & ~_writeQueueVec_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn),
    .empty        (_writeQueueVec_fifo_empty),
    .almost_empty (writeQueueVec_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_0_almostFull),
    .full         (_writeQueueVec_fifo_full),
    .error        (_writeQueueVec_fifo_error),
    .data_out     (_writeQueueVec_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(63)
  ) writeQueueVec_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_1_writeValid_T & ~(_writeQueueVec_fifo_1_empty & writeQueueVec_1_deq_ready))),
    .pop_req_n    (~(writeQueueVec_1_deq_ready & ~_writeQueueVec_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_1),
    .empty        (_writeQueueVec_fifo_1_empty),
    .almost_empty (writeQueueVec_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_1_almostFull),
    .full         (_writeQueueVec_fifo_1_full),
    .error        (_writeQueueVec_fifo_1_error),
    .data_out     (_writeQueueVec_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(63)
  ) writeQueueVec_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_2_writeValid_T & ~(_writeQueueVec_fifo_2_empty & writeQueueVec_2_deq_ready))),
    .pop_req_n    (~(writeQueueVec_2_deq_ready & ~_writeQueueVec_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_2),
    .empty        (_writeQueueVec_fifo_2_empty),
    .almost_empty (writeQueueVec_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_2_almostFull),
    .full         (_writeQueueVec_fifo_2_full),
    .error        (_writeQueueVec_fifo_2_error),
    .data_out     (_writeQueueVec_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(63)
  ) writeQueueVec_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_3_writeValid_T & ~(_writeQueueVec_fifo_3_empty & writeQueueVec_3_deq_ready))),
    .pop_req_n    (~(writeQueueVec_3_deq_ready & ~_writeQueueVec_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_3),
    .empty        (_writeQueueVec_fifo_3_empty),
    .almost_empty (writeQueueVec_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_3_almostFull),
    .full         (_writeQueueVec_fifo_3_full),
    .error        (_writeQueueVec_fifo_3_error),
    .data_out     (_writeQueueVec_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(63)
  ) writeQueueVec_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_4_writeValid_T & ~(_writeQueueVec_fifo_4_empty & writeQueueVec_4_deq_ready))),
    .pop_req_n    (~(writeQueueVec_4_deq_ready & ~_writeQueueVec_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_4),
    .empty        (_writeQueueVec_fifo_4_empty),
    .almost_empty (writeQueueVec_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_4_almostFull),
    .full         (_writeQueueVec_fifo_4_full),
    .error        (_writeQueueVec_fifo_4_error),
    .data_out     (_writeQueueVec_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(63)
  ) writeQueueVec_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_5_writeValid_T & ~(_writeQueueVec_fifo_5_empty & writeQueueVec_5_deq_ready))),
    .pop_req_n    (~(writeQueueVec_5_deq_ready & ~_writeQueueVec_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_5),
    .empty        (_writeQueueVec_fifo_5_empty),
    .almost_empty (writeQueueVec_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_5_almostFull),
    .full         (_writeQueueVec_fifo_5_full),
    .error        (_writeQueueVec_fifo_5_error),
    .data_out     (_writeQueueVec_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(63)
  ) writeQueueVec_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_6_writeValid_T & ~(_writeQueueVec_fifo_6_empty & writeQueueVec_6_deq_ready))),
    .pop_req_n    (~(writeQueueVec_6_deq_ready & ~_writeQueueVec_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_6),
    .empty        (_writeQueueVec_fifo_6_empty),
    .almost_empty (writeQueueVec_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_6_almostFull),
    .full         (_writeQueueVec_fifo_6_full),
    .error        (_writeQueueVec_fifo_6_error),
    .data_out     (_writeQueueVec_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(63)
  ) writeQueueVec_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_7_writeValid_T & ~(_writeQueueVec_fifo_7_empty & writeQueueVec_7_deq_ready))),
    .pop_req_n    (~(writeQueueVec_7_deq_ready & ~_writeQueueVec_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_7),
    .empty        (_writeQueueVec_fifo_7_empty),
    .almost_empty (writeQueueVec_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_7_almostFull),
    .full         (_writeQueueVec_fifo_7_full),
    .error        (_writeQueueVec_fifo_7_error),
    .data_out     (_writeQueueVec_fifo_7_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(63)
  ) writeQueueVec_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_8_writeValid_T & ~(_writeQueueVec_fifo_8_empty & writeQueueVec_8_deq_ready))),
    .pop_req_n    (~(writeQueueVec_8_deq_ready & ~_writeQueueVec_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_8),
    .empty        (_writeQueueVec_fifo_8_empty),
    .almost_empty (writeQueueVec_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_8_almostFull),
    .full         (_writeQueueVec_fifo_8_full),
    .error        (_writeQueueVec_fifo_8_error),
    .data_out     (_writeQueueVec_fifo_8_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(63)
  ) writeQueueVec_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_9_writeValid_T & ~(_writeQueueVec_fifo_9_empty & writeQueueVec_9_deq_ready))),
    .pop_req_n    (~(writeQueueVec_9_deq_ready & ~_writeQueueVec_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_9),
    .empty        (_writeQueueVec_fifo_9_empty),
    .almost_empty (writeQueueVec_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_9_almostFull),
    .full         (_writeQueueVec_fifo_9_full),
    .error        (_writeQueueVec_fifo_9_error),
    .data_out     (_writeQueueVec_fifo_9_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(63)
  ) writeQueueVec_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_10_writeValid_T & ~(_writeQueueVec_fifo_10_empty & writeQueueVec_10_deq_ready))),
    .pop_req_n    (~(writeQueueVec_10_deq_ready & ~_writeQueueVec_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_10),
    .empty        (_writeQueueVec_fifo_10_empty),
    .almost_empty (writeQueueVec_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_10_almostFull),
    .full         (_writeQueueVec_fifo_10_full),
    .error        (_writeQueueVec_fifo_10_error),
    .data_out     (_writeQueueVec_fifo_10_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(63)
  ) writeQueueVec_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_11_writeValid_T & ~(_writeQueueVec_fifo_11_empty & writeQueueVec_11_deq_ready))),
    .pop_req_n    (~(writeQueueVec_11_deq_ready & ~_writeQueueVec_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_11),
    .empty        (_writeQueueVec_fifo_11_empty),
    .almost_empty (writeQueueVec_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_11_almostFull),
    .full         (_writeQueueVec_fifo_11_full),
    .error        (_writeQueueVec_fifo_11_error),
    .data_out     (_writeQueueVec_fifo_11_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(63)
  ) writeQueueVec_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_12_writeValid_T & ~(_writeQueueVec_fifo_12_empty & writeQueueVec_12_deq_ready))),
    .pop_req_n    (~(writeQueueVec_12_deq_ready & ~_writeQueueVec_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_12),
    .empty        (_writeQueueVec_fifo_12_empty),
    .almost_empty (writeQueueVec_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_12_almostFull),
    .full         (_writeQueueVec_fifo_12_full),
    .error        (_writeQueueVec_fifo_12_error),
    .data_out     (_writeQueueVec_fifo_12_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(63)
  ) writeQueueVec_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_13_writeValid_T & ~(_writeQueueVec_fifo_13_empty & writeQueueVec_13_deq_ready))),
    .pop_req_n    (~(writeQueueVec_13_deq_ready & ~_writeQueueVec_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_13),
    .empty        (_writeQueueVec_fifo_13_empty),
    .almost_empty (writeQueueVec_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_13_almostFull),
    .full         (_writeQueueVec_fifo_13_full),
    .error        (_writeQueueVec_fifo_13_error),
    .data_out     (_writeQueueVec_fifo_13_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(63)
  ) writeQueueVec_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_14_writeValid_T & ~(_writeQueueVec_fifo_14_empty & writeQueueVec_14_deq_ready))),
    .pop_req_n    (~(writeQueueVec_14_deq_ready & ~_writeQueueVec_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_14),
    .empty        (_writeQueueVec_fifo_14_empty),
    .almost_empty (writeQueueVec_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_14_almostFull),
    .full         (_writeQueueVec_fifo_14_full),
    .error        (_writeQueueVec_fifo_14_error),
    .data_out     (_writeQueueVec_fifo_14_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(63)
  ) writeQueueVec_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_15_writeValid_T & ~(_writeQueueVec_fifo_15_empty & writeQueueVec_15_deq_ready))),
    .pop_req_n    (~(writeQueueVec_15_deq_ready & ~_writeQueueVec_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_15),
    .empty        (_writeQueueVec_fifo_15_empty),
    .almost_empty (writeQueueVec_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_15_almostFull),
    .full         (_writeQueueVec_fifo_15_full),
    .error        (_writeQueueVec_fifo_15_error),
    .data_out     (_writeQueueVec_fifo_15_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(16)
  ) otherUnitTargetQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitTargetQueue_enq_ready & otherUnitTargetQueue_enq_valid)),
    .pop_req_n    (~(otherUnitTargetQueue_deq_ready & ~_otherUnitTargetQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitTargetQueue_enq_bits),
    .empty        (_otherUnitTargetQueue_fifo_empty),
    .almost_empty (otherUnitTargetQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitTargetQueue_almostFull),
    .full         (_otherUnitTargetQueue_fifo_full),
    .error        (_otherUnitTargetQueue_fifo_error),
    .data_out     (otherUnitTargetQueue_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_0_enq_ready & otherUnitDataQueueVec_0_enq_valid & ~(_otherUnitDataQueueVec_fifo_empty & otherUnitDataQueueVec_0_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_0_deq_ready & ~_otherUnitDataQueueVec_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_0_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_empty),
    .almost_empty (otherUnitDataQueueVec_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_0_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_full),
    .error        (_otherUnitDataQueueVec_fifo_error),
    .data_out     (_otherUnitDataQueueVec_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_1_enq_ready & otherUnitDataQueueVec_1_enq_valid & ~(_otherUnitDataQueueVec_fifo_1_empty & otherUnitDataQueueVec_1_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_1_deq_ready & ~_otherUnitDataQueueVec_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_1_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_1_empty),
    .almost_empty (otherUnitDataQueueVec_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_1_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_1_full),
    .error        (_otherUnitDataQueueVec_fifo_1_error),
    .data_out     (_otherUnitDataQueueVec_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_2_enq_ready & otherUnitDataQueueVec_2_enq_valid & ~(_otherUnitDataQueueVec_fifo_2_empty & otherUnitDataQueueVec_2_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_2_deq_ready & ~_otherUnitDataQueueVec_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_2_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_2_empty),
    .almost_empty (otherUnitDataQueueVec_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_2_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_2_full),
    .error        (_otherUnitDataQueueVec_fifo_2_error),
    .data_out     (_otherUnitDataQueueVec_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_3_enq_ready & otherUnitDataQueueVec_3_enq_valid & ~(_otherUnitDataQueueVec_fifo_3_empty & otherUnitDataQueueVec_3_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_3_deq_ready & ~_otherUnitDataQueueVec_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_3_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_3_empty),
    .almost_empty (otherUnitDataQueueVec_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_3_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_3_full),
    .error        (_otherUnitDataQueueVec_fifo_3_error),
    .data_out     (_otherUnitDataQueueVec_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_4_enq_ready & otherUnitDataQueueVec_4_enq_valid & ~(_otherUnitDataQueueVec_fifo_4_empty & otherUnitDataQueueVec_4_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_4_deq_ready & ~_otherUnitDataQueueVec_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_4_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_4_empty),
    .almost_empty (otherUnitDataQueueVec_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_4_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_4_full),
    .error        (_otherUnitDataQueueVec_fifo_4_error),
    .data_out     (_otherUnitDataQueueVec_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_5_enq_ready & otherUnitDataQueueVec_5_enq_valid & ~(_otherUnitDataQueueVec_fifo_5_empty & otherUnitDataQueueVec_5_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_5_deq_ready & ~_otherUnitDataQueueVec_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_5_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_5_empty),
    .almost_empty (otherUnitDataQueueVec_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_5_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_5_full),
    .error        (_otherUnitDataQueueVec_fifo_5_error),
    .data_out     (_otherUnitDataQueueVec_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_6_enq_ready & otherUnitDataQueueVec_6_enq_valid & ~(_otherUnitDataQueueVec_fifo_6_empty & otherUnitDataQueueVec_6_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_6_deq_ready & ~_otherUnitDataQueueVec_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_6_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_6_empty),
    .almost_empty (otherUnitDataQueueVec_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_6_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_6_full),
    .error        (_otherUnitDataQueueVec_fifo_6_error),
    .data_out     (_otherUnitDataQueueVec_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_7_enq_ready & otherUnitDataQueueVec_7_enq_valid & ~(_otherUnitDataQueueVec_fifo_7_empty & otherUnitDataQueueVec_7_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_7_deq_ready & ~_otherUnitDataQueueVec_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_7_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_7_empty),
    .almost_empty (otherUnitDataQueueVec_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_7_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_7_full),
    .error        (_otherUnitDataQueueVec_fifo_7_error),
    .data_out     (_otherUnitDataQueueVec_fifo_7_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_8_enq_ready & otherUnitDataQueueVec_8_enq_valid & ~(_otherUnitDataQueueVec_fifo_8_empty & otherUnitDataQueueVec_8_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_8_deq_ready & ~_otherUnitDataQueueVec_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_8_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_8_empty),
    .almost_empty (otherUnitDataQueueVec_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_8_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_8_full),
    .error        (_otherUnitDataQueueVec_fifo_8_error),
    .data_out     (_otherUnitDataQueueVec_fifo_8_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_9_enq_ready & otherUnitDataQueueVec_9_enq_valid & ~(_otherUnitDataQueueVec_fifo_9_empty & otherUnitDataQueueVec_9_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_9_deq_ready & ~_otherUnitDataQueueVec_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_9_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_9_empty),
    .almost_empty (otherUnitDataQueueVec_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_9_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_9_full),
    .error        (_otherUnitDataQueueVec_fifo_9_error),
    .data_out     (_otherUnitDataQueueVec_fifo_9_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_10_enq_ready & otherUnitDataQueueVec_10_enq_valid & ~(_otherUnitDataQueueVec_fifo_10_empty & otherUnitDataQueueVec_10_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_10_deq_ready & ~_otherUnitDataQueueVec_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_10_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_10_empty),
    .almost_empty (otherUnitDataQueueVec_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_10_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_10_full),
    .error        (_otherUnitDataQueueVec_fifo_10_error),
    .data_out     (_otherUnitDataQueueVec_fifo_10_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_11_enq_ready & otherUnitDataQueueVec_11_enq_valid & ~(_otherUnitDataQueueVec_fifo_11_empty & otherUnitDataQueueVec_11_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_11_deq_ready & ~_otherUnitDataQueueVec_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_11_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_11_empty),
    .almost_empty (otherUnitDataQueueVec_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_11_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_11_full),
    .error        (_otherUnitDataQueueVec_fifo_11_error),
    .data_out     (_otherUnitDataQueueVec_fifo_11_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_12_enq_ready & otherUnitDataQueueVec_12_enq_valid & ~(_otherUnitDataQueueVec_fifo_12_empty & otherUnitDataQueueVec_12_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_12_deq_ready & ~_otherUnitDataQueueVec_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_12_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_12_empty),
    .almost_empty (otherUnitDataQueueVec_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_12_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_12_full),
    .error        (_otherUnitDataQueueVec_fifo_12_error),
    .data_out     (_otherUnitDataQueueVec_fifo_12_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_13_enq_ready & otherUnitDataQueueVec_13_enq_valid & ~(_otherUnitDataQueueVec_fifo_13_empty & otherUnitDataQueueVec_13_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_13_deq_ready & ~_otherUnitDataQueueVec_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_13_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_13_empty),
    .almost_empty (otherUnitDataQueueVec_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_13_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_13_full),
    .error        (_otherUnitDataQueueVec_fifo_13_error),
    .data_out     (_otherUnitDataQueueVec_fifo_13_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_14_enq_ready & otherUnitDataQueueVec_14_enq_valid & ~(_otherUnitDataQueueVec_fifo_14_empty & otherUnitDataQueueVec_14_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_14_deq_ready & ~_otherUnitDataQueueVec_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_14_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_14_empty),
    .almost_empty (otherUnitDataQueueVec_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_14_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_14_full),
    .error        (_otherUnitDataQueueVec_fifo_14_error),
    .data_out     (_otherUnitDataQueueVec_fifo_14_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_15_enq_ready & otherUnitDataQueueVec_15_enq_valid & ~(_otherUnitDataQueueVec_fifo_15_empty & otherUnitDataQueueVec_15_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_15_deq_ready & ~_otherUnitDataQueueVec_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_15_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_15_empty),
    .almost_empty (otherUnitDataQueueVec_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_15_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_15_full),
    .error        (_otherUnitDataQueueVec_fifo_15_error),
    .data_out     (_otherUnitDataQueueVec_fifo_15_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_enq_ready & writeIndexQueue_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_deq_ready & ~_writeIndexQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_enq_bits),
    .empty        (_writeIndexQueue_fifo_empty),
    .almost_empty (writeIndexQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_almostFull),
    .full         (_writeIndexQueue_fifo_full),
    .error        (_writeIndexQueue_fifo_error),
    .data_out     (writeIndexQueue_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_1_enq_ready & writeIndexQueue_1_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_1_deq_ready & ~_writeIndexQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_1_enq_bits),
    .empty        (_writeIndexQueue_fifo_1_empty),
    .almost_empty (writeIndexQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_1_almostFull),
    .full         (_writeIndexQueue_fifo_1_full),
    .error        (_writeIndexQueue_fifo_1_error),
    .data_out     (writeIndexQueue_1_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_2_enq_ready & writeIndexQueue_2_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_2_deq_ready & ~_writeIndexQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_2_enq_bits),
    .empty        (_writeIndexQueue_fifo_2_empty),
    .almost_empty (writeIndexQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_2_almostFull),
    .full         (_writeIndexQueue_fifo_2_full),
    .error        (_writeIndexQueue_fifo_2_error),
    .data_out     (writeIndexQueue_2_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_3_enq_ready & writeIndexQueue_3_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_3_deq_ready & ~_writeIndexQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_3_enq_bits),
    .empty        (_writeIndexQueue_fifo_3_empty),
    .almost_empty (writeIndexQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_3_almostFull),
    .full         (_writeIndexQueue_fifo_3_full),
    .error        (_writeIndexQueue_fifo_3_error),
    .data_out     (writeIndexQueue_3_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_4_enq_ready & writeIndexQueue_4_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_4_deq_ready & ~_writeIndexQueue_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_4_enq_bits),
    .empty        (_writeIndexQueue_fifo_4_empty),
    .almost_empty (writeIndexQueue_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_4_almostFull),
    .full         (_writeIndexQueue_fifo_4_full),
    .error        (_writeIndexQueue_fifo_4_error),
    .data_out     (writeIndexQueue_4_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_5_enq_ready & writeIndexQueue_5_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_5_deq_ready & ~_writeIndexQueue_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_5_enq_bits),
    .empty        (_writeIndexQueue_fifo_5_empty),
    .almost_empty (writeIndexQueue_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_5_almostFull),
    .full         (_writeIndexQueue_fifo_5_full),
    .error        (_writeIndexQueue_fifo_5_error),
    .data_out     (writeIndexQueue_5_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_6_enq_ready & writeIndexQueue_6_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_6_deq_ready & ~_writeIndexQueue_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_6_enq_bits),
    .empty        (_writeIndexQueue_fifo_6_empty),
    .almost_empty (writeIndexQueue_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_6_almostFull),
    .full         (_writeIndexQueue_fifo_6_full),
    .error        (_writeIndexQueue_fifo_6_error),
    .data_out     (writeIndexQueue_6_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_7_enq_ready & writeIndexQueue_7_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_7_deq_ready & ~_writeIndexQueue_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_7_enq_bits),
    .empty        (_writeIndexQueue_fifo_7_empty),
    .almost_empty (writeIndexQueue_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_7_almostFull),
    .full         (_writeIndexQueue_fifo_7_full),
    .error        (_writeIndexQueue_fifo_7_error),
    .data_out     (writeIndexQueue_7_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_8_enq_ready & writeIndexQueue_8_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_8_deq_ready & ~_writeIndexQueue_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_8_enq_bits),
    .empty        (_writeIndexQueue_fifo_8_empty),
    .almost_empty (writeIndexQueue_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_8_almostFull),
    .full         (_writeIndexQueue_fifo_8_full),
    .error        (_writeIndexQueue_fifo_8_error),
    .data_out     (writeIndexQueue_8_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_9_enq_ready & writeIndexQueue_9_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_9_deq_ready & ~_writeIndexQueue_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_9_enq_bits),
    .empty        (_writeIndexQueue_fifo_9_empty),
    .almost_empty (writeIndexQueue_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_9_almostFull),
    .full         (_writeIndexQueue_fifo_9_full),
    .error        (_writeIndexQueue_fifo_9_error),
    .data_out     (writeIndexQueue_9_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_10_enq_ready & writeIndexQueue_10_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_10_deq_ready & ~_writeIndexQueue_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_10_enq_bits),
    .empty        (_writeIndexQueue_fifo_10_empty),
    .almost_empty (writeIndexQueue_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_10_almostFull),
    .full         (_writeIndexQueue_fifo_10_full),
    .error        (_writeIndexQueue_fifo_10_error),
    .data_out     (writeIndexQueue_10_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_11_enq_ready & writeIndexQueue_11_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_11_deq_ready & ~_writeIndexQueue_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_11_enq_bits),
    .empty        (_writeIndexQueue_fifo_11_empty),
    .almost_empty (writeIndexQueue_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_11_almostFull),
    .full         (_writeIndexQueue_fifo_11_full),
    .error        (_writeIndexQueue_fifo_11_error),
    .data_out     (writeIndexQueue_11_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_12_enq_ready & writeIndexQueue_12_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_12_deq_ready & ~_writeIndexQueue_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_12_enq_bits),
    .empty        (_writeIndexQueue_fifo_12_empty),
    .almost_empty (writeIndexQueue_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_12_almostFull),
    .full         (_writeIndexQueue_fifo_12_full),
    .error        (_writeIndexQueue_fifo_12_error),
    .data_out     (writeIndexQueue_12_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_13_enq_ready & writeIndexQueue_13_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_13_deq_ready & ~_writeIndexQueue_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_13_enq_bits),
    .empty        (_writeIndexQueue_fifo_13_empty),
    .almost_empty (writeIndexQueue_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_13_almostFull),
    .full         (_writeIndexQueue_fifo_13_full),
    .error        (_writeIndexQueue_fifo_13_error),
    .data_out     (writeIndexQueue_13_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_14_enq_ready & writeIndexQueue_14_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_14_deq_ready & ~_writeIndexQueue_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_14_enq_bits),
    .empty        (_writeIndexQueue_fifo_14_empty),
    .almost_empty (writeIndexQueue_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_14_almostFull),
    .full         (_writeIndexQueue_fifo_14_full),
    .error        (_writeIndexQueue_fifo_14_error),
    .data_out     (writeIndexQueue_14_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_15_enq_ready & writeIndexQueue_15_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_15_deq_ready & ~_writeIndexQueue_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_15_enq_bits),
    .empty        (_writeIndexQueue_fifo_15_empty),
    .almost_empty (writeIndexQueue_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_15_almostFull),
    .full         (_writeIndexQueue_fifo_15_full),
    .error        (_writeIndexQueue_fifo_15_error),
    .data_out     (writeIndexQueue_15_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(6)
  ) sourceQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sourceQueue_enq_ready & sourceQueue_enq_valid)),
    .pop_req_n    (~(sourceQueue_deq_ready & ~_sourceQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (sourceQueue_enq_bits),
    .empty        (_sourceQueue_fifo_empty),
    .almost_empty (sourceQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sourceQueue_almostFull),
    .full         (_sourceQueue_fifo_full),
    .error        (_sourceQueue_fifo_error),
    .data_out     (sourceQueue_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(2),
    .err_mode(2),
    .rst_mode(3),
    .width(614)
  ) dataQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(dataQueue_enq_ready & dataQueue_enq_valid)),
    .pop_req_n    (~(dataQueue_deq_ready & ~_dataQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (dataQueue_dataIn),
    .empty        (_dataQueue_fifo_empty),
    .almost_empty (dataQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (dataQueue_almostFull),
    .full         (_dataQueue_fifo_full),
    .error        (_dataQueue_fifo_error),
    .data_out     (_dataQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(9)
  ) simpleSourceQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(simpleSourceQueue_enq_ready & simpleSourceQueue_enq_valid)),
    .pop_req_n    (~(simpleSourceQueue_deq_ready & ~_simpleSourceQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (simpleSourceQueue_enq_bits),
    .empty        (_simpleSourceQueue_fifo_empty),
    .almost_empty (simpleSourceQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (simpleSourceQueue_almostFull),
    .full         (_simpleSourceQueue_fifo_full),
    .error        (_simpleSourceQueue_fifo_error),
    .data_out     (simpleSourceQueue_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(2),
    .err_mode(2),
    .rst_mode(3),
    .width(78)
  ) simpleDataQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(simpleDataQueue_enq_ready & simpleDataQueue_enq_valid)),
    .pop_req_n    (~(simpleDataQueue_deq_ready & ~_simpleDataQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (simpleDataQueue_dataIn),
    .empty        (_simpleDataQueue_fifo_empty),
    .almost_empty (simpleDataQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (simpleDataQueue_almostFull),
    .full         (_simpleDataQueue_fifo_full),
    .error        (_simpleDataQueue_fifo_error),
    .data_out     (_simpleDataQueue_fifo_data_out)
  );
  assign request_ready = request_ready_0;
  assign axi4Port_aw_valid = axi4Port_aw_valid_0;
  assign axi4Port_aw_bits_id = axi4Port_aw_bits_id_0;
  assign axi4Port_aw_bits_addr = axi4Port_aw_bits_addr_0;
  assign axi4Port_w_valid = axi4Port_w_valid_0;
  assign axi4Port_w_bits_data = axi4Port_w_bits_data_0;
  assign axi4Port_w_bits_strb = axi4Port_w_bits_strb_0;
  assign axi4Port_ar_valid = axi4Port_ar_valid_0;
  assign axi4Port_ar_bits_addr = axi4Port_ar_bits_addr_0;
  assign axi4Port_r_ready = axi4Port_r_ready_0;
  assign simpleAccessPorts_aw_valid = simpleAccessPorts_aw_valid_0;
  assign simpleAccessPorts_aw_bits_id = simpleAccessPorts_aw_bits_id_0;
  assign simpleAccessPorts_aw_bits_addr = simpleAccessPorts_aw_bits_addr_0;
  assign simpleAccessPorts_aw_bits_size = simpleAccessPorts_aw_bits_size_0;
  assign simpleAccessPorts_w_valid = simpleAccessPorts_w_valid_0;
  assign simpleAccessPorts_w_bits_data = simpleAccessPorts_w_bits_data_0;
  assign simpleAccessPorts_w_bits_strb = simpleAccessPorts_w_bits_strb_0;
  assign simpleAccessPorts_ar_valid = simpleAccessPorts_ar_valid_0;
  assign simpleAccessPorts_ar_bits_addr = simpleAccessPorts_ar_bits_addr_0;
  assign simpleAccessPorts_r_ready = simpleAccessPorts_r_ready_0;
  assign vrfReadDataPorts_0_valid = vrfReadDataPorts_0_valid_0;
  assign vrfReadDataPorts_0_bits_vs = vrfReadDataPorts_0_bits_vs_0;
  assign vrfReadDataPorts_0_bits_offset = vrfReadDataPorts_0_bits_offset_0;
  assign vrfReadDataPorts_0_bits_instructionIndex = vrfReadDataPorts_0_bits_instructionIndex_0;
  assign vrfReadDataPorts_1_valid = vrfReadDataPorts_1_valid_0;
  assign vrfReadDataPorts_1_bits_vs = vrfReadDataPorts_1_bits_vs_0;
  assign vrfReadDataPorts_1_bits_offset = vrfReadDataPorts_1_bits_offset_0;
  assign vrfReadDataPorts_1_bits_instructionIndex = vrfReadDataPorts_1_bits_instructionIndex_0;
  assign vrfReadDataPorts_2_valid = vrfReadDataPorts_2_valid_0;
  assign vrfReadDataPorts_2_bits_vs = vrfReadDataPorts_2_bits_vs_0;
  assign vrfReadDataPorts_2_bits_offset = vrfReadDataPorts_2_bits_offset_0;
  assign vrfReadDataPorts_2_bits_instructionIndex = vrfReadDataPorts_2_bits_instructionIndex_0;
  assign vrfReadDataPorts_3_valid = vrfReadDataPorts_3_valid_0;
  assign vrfReadDataPorts_3_bits_vs = vrfReadDataPorts_3_bits_vs_0;
  assign vrfReadDataPorts_3_bits_offset = vrfReadDataPorts_3_bits_offset_0;
  assign vrfReadDataPorts_3_bits_instructionIndex = vrfReadDataPorts_3_bits_instructionIndex_0;
  assign vrfReadDataPorts_4_valid = vrfReadDataPorts_4_valid_0;
  assign vrfReadDataPorts_4_bits_vs = vrfReadDataPorts_4_bits_vs_0;
  assign vrfReadDataPorts_4_bits_offset = vrfReadDataPorts_4_bits_offset_0;
  assign vrfReadDataPorts_4_bits_instructionIndex = vrfReadDataPorts_4_bits_instructionIndex_0;
  assign vrfReadDataPorts_5_valid = vrfReadDataPorts_5_valid_0;
  assign vrfReadDataPorts_5_bits_vs = vrfReadDataPorts_5_bits_vs_0;
  assign vrfReadDataPorts_5_bits_offset = vrfReadDataPorts_5_bits_offset_0;
  assign vrfReadDataPorts_5_bits_instructionIndex = vrfReadDataPorts_5_bits_instructionIndex_0;
  assign vrfReadDataPorts_6_valid = vrfReadDataPorts_6_valid_0;
  assign vrfReadDataPorts_6_bits_vs = vrfReadDataPorts_6_bits_vs_0;
  assign vrfReadDataPorts_6_bits_offset = vrfReadDataPorts_6_bits_offset_0;
  assign vrfReadDataPorts_6_bits_instructionIndex = vrfReadDataPorts_6_bits_instructionIndex_0;
  assign vrfReadDataPorts_7_valid = vrfReadDataPorts_7_valid_0;
  assign vrfReadDataPorts_7_bits_vs = vrfReadDataPorts_7_bits_vs_0;
  assign vrfReadDataPorts_7_bits_offset = vrfReadDataPorts_7_bits_offset_0;
  assign vrfReadDataPorts_7_bits_instructionIndex = vrfReadDataPorts_7_bits_instructionIndex_0;
  assign vrfReadDataPorts_8_valid = vrfReadDataPorts_8_valid_0;
  assign vrfReadDataPorts_8_bits_vs = vrfReadDataPorts_8_bits_vs_0;
  assign vrfReadDataPorts_8_bits_offset = vrfReadDataPorts_8_bits_offset_0;
  assign vrfReadDataPorts_8_bits_instructionIndex = vrfReadDataPorts_8_bits_instructionIndex_0;
  assign vrfReadDataPorts_9_valid = vrfReadDataPorts_9_valid_0;
  assign vrfReadDataPorts_9_bits_vs = vrfReadDataPorts_9_bits_vs_0;
  assign vrfReadDataPorts_9_bits_offset = vrfReadDataPorts_9_bits_offset_0;
  assign vrfReadDataPorts_9_bits_instructionIndex = vrfReadDataPorts_9_bits_instructionIndex_0;
  assign vrfReadDataPorts_10_valid = vrfReadDataPorts_10_valid_0;
  assign vrfReadDataPorts_10_bits_vs = vrfReadDataPorts_10_bits_vs_0;
  assign vrfReadDataPorts_10_bits_offset = vrfReadDataPorts_10_bits_offset_0;
  assign vrfReadDataPorts_10_bits_instructionIndex = vrfReadDataPorts_10_bits_instructionIndex_0;
  assign vrfReadDataPorts_11_valid = vrfReadDataPorts_11_valid_0;
  assign vrfReadDataPorts_11_bits_vs = vrfReadDataPorts_11_bits_vs_0;
  assign vrfReadDataPorts_11_bits_offset = vrfReadDataPorts_11_bits_offset_0;
  assign vrfReadDataPorts_11_bits_instructionIndex = vrfReadDataPorts_11_bits_instructionIndex_0;
  assign vrfReadDataPorts_12_valid = vrfReadDataPorts_12_valid_0;
  assign vrfReadDataPorts_12_bits_vs = vrfReadDataPorts_12_bits_vs_0;
  assign vrfReadDataPorts_12_bits_offset = vrfReadDataPorts_12_bits_offset_0;
  assign vrfReadDataPorts_12_bits_instructionIndex = vrfReadDataPorts_12_bits_instructionIndex_0;
  assign vrfReadDataPorts_13_valid = vrfReadDataPorts_13_valid_0;
  assign vrfReadDataPorts_13_bits_vs = vrfReadDataPorts_13_bits_vs_0;
  assign vrfReadDataPorts_13_bits_offset = vrfReadDataPorts_13_bits_offset_0;
  assign vrfReadDataPorts_13_bits_instructionIndex = vrfReadDataPorts_13_bits_instructionIndex_0;
  assign vrfReadDataPorts_14_valid = vrfReadDataPorts_14_valid_0;
  assign vrfReadDataPorts_14_bits_vs = vrfReadDataPorts_14_bits_vs_0;
  assign vrfReadDataPorts_14_bits_offset = vrfReadDataPorts_14_bits_offset_0;
  assign vrfReadDataPorts_14_bits_instructionIndex = vrfReadDataPorts_14_bits_instructionIndex_0;
  assign vrfReadDataPorts_15_valid = vrfReadDataPorts_15_valid_0;
  assign vrfReadDataPorts_15_bits_vs = vrfReadDataPorts_15_bits_vs_0;
  assign vrfReadDataPorts_15_bits_offset = vrfReadDataPorts_15_bits_offset_0;
  assign vrfReadDataPorts_15_bits_instructionIndex = vrfReadDataPorts_15_bits_instructionIndex_0;
  assign vrfWritePort_0_valid = vrfWritePort_0_valid_0;
  assign vrfWritePort_0_bits_vd = vrfWritePort_0_bits_vd_0;
  assign vrfWritePort_0_bits_offset = vrfWritePort_0_bits_offset_0;
  assign vrfWritePort_0_bits_mask = vrfWritePort_0_bits_mask_0;
  assign vrfWritePort_0_bits_data = vrfWritePort_0_bits_data_0;
  assign vrfWritePort_0_bits_last = vrfWritePort_0_bits_last_0;
  assign vrfWritePort_0_bits_instructionIndex = vrfWritePort_0_bits_instructionIndex_0;
  assign vrfWritePort_1_valid = vrfWritePort_1_valid_0;
  assign vrfWritePort_1_bits_vd = vrfWritePort_1_bits_vd_0;
  assign vrfWritePort_1_bits_offset = vrfWritePort_1_bits_offset_0;
  assign vrfWritePort_1_bits_mask = vrfWritePort_1_bits_mask_0;
  assign vrfWritePort_1_bits_data = vrfWritePort_1_bits_data_0;
  assign vrfWritePort_1_bits_last = vrfWritePort_1_bits_last_0;
  assign vrfWritePort_1_bits_instructionIndex = vrfWritePort_1_bits_instructionIndex_0;
  assign vrfWritePort_2_valid = vrfWritePort_2_valid_0;
  assign vrfWritePort_2_bits_vd = vrfWritePort_2_bits_vd_0;
  assign vrfWritePort_2_bits_offset = vrfWritePort_2_bits_offset_0;
  assign vrfWritePort_2_bits_mask = vrfWritePort_2_bits_mask_0;
  assign vrfWritePort_2_bits_data = vrfWritePort_2_bits_data_0;
  assign vrfWritePort_2_bits_last = vrfWritePort_2_bits_last_0;
  assign vrfWritePort_2_bits_instructionIndex = vrfWritePort_2_bits_instructionIndex_0;
  assign vrfWritePort_3_valid = vrfWritePort_3_valid_0;
  assign vrfWritePort_3_bits_vd = vrfWritePort_3_bits_vd_0;
  assign vrfWritePort_3_bits_offset = vrfWritePort_3_bits_offset_0;
  assign vrfWritePort_3_bits_mask = vrfWritePort_3_bits_mask_0;
  assign vrfWritePort_3_bits_data = vrfWritePort_3_bits_data_0;
  assign vrfWritePort_3_bits_last = vrfWritePort_3_bits_last_0;
  assign vrfWritePort_3_bits_instructionIndex = vrfWritePort_3_bits_instructionIndex_0;
  assign vrfWritePort_4_valid = vrfWritePort_4_valid_0;
  assign vrfWritePort_4_bits_vd = vrfWritePort_4_bits_vd_0;
  assign vrfWritePort_4_bits_offset = vrfWritePort_4_bits_offset_0;
  assign vrfWritePort_4_bits_mask = vrfWritePort_4_bits_mask_0;
  assign vrfWritePort_4_bits_data = vrfWritePort_4_bits_data_0;
  assign vrfWritePort_4_bits_last = vrfWritePort_4_bits_last_0;
  assign vrfWritePort_4_bits_instructionIndex = vrfWritePort_4_bits_instructionIndex_0;
  assign vrfWritePort_5_valid = vrfWritePort_5_valid_0;
  assign vrfWritePort_5_bits_vd = vrfWritePort_5_bits_vd_0;
  assign vrfWritePort_5_bits_offset = vrfWritePort_5_bits_offset_0;
  assign vrfWritePort_5_bits_mask = vrfWritePort_5_bits_mask_0;
  assign vrfWritePort_5_bits_data = vrfWritePort_5_bits_data_0;
  assign vrfWritePort_5_bits_last = vrfWritePort_5_bits_last_0;
  assign vrfWritePort_5_bits_instructionIndex = vrfWritePort_5_bits_instructionIndex_0;
  assign vrfWritePort_6_valid = vrfWritePort_6_valid_0;
  assign vrfWritePort_6_bits_vd = vrfWritePort_6_bits_vd_0;
  assign vrfWritePort_6_bits_offset = vrfWritePort_6_bits_offset_0;
  assign vrfWritePort_6_bits_mask = vrfWritePort_6_bits_mask_0;
  assign vrfWritePort_6_bits_data = vrfWritePort_6_bits_data_0;
  assign vrfWritePort_6_bits_last = vrfWritePort_6_bits_last_0;
  assign vrfWritePort_6_bits_instructionIndex = vrfWritePort_6_bits_instructionIndex_0;
  assign vrfWritePort_7_valid = vrfWritePort_7_valid_0;
  assign vrfWritePort_7_bits_vd = vrfWritePort_7_bits_vd_0;
  assign vrfWritePort_7_bits_offset = vrfWritePort_7_bits_offset_0;
  assign vrfWritePort_7_bits_mask = vrfWritePort_7_bits_mask_0;
  assign vrfWritePort_7_bits_data = vrfWritePort_7_bits_data_0;
  assign vrfWritePort_7_bits_last = vrfWritePort_7_bits_last_0;
  assign vrfWritePort_7_bits_instructionIndex = vrfWritePort_7_bits_instructionIndex_0;
  assign vrfWritePort_8_valid = vrfWritePort_8_valid_0;
  assign vrfWritePort_8_bits_vd = vrfWritePort_8_bits_vd_0;
  assign vrfWritePort_8_bits_offset = vrfWritePort_8_bits_offset_0;
  assign vrfWritePort_8_bits_mask = vrfWritePort_8_bits_mask_0;
  assign vrfWritePort_8_bits_data = vrfWritePort_8_bits_data_0;
  assign vrfWritePort_8_bits_last = vrfWritePort_8_bits_last_0;
  assign vrfWritePort_8_bits_instructionIndex = vrfWritePort_8_bits_instructionIndex_0;
  assign vrfWritePort_9_valid = vrfWritePort_9_valid_0;
  assign vrfWritePort_9_bits_vd = vrfWritePort_9_bits_vd_0;
  assign vrfWritePort_9_bits_offset = vrfWritePort_9_bits_offset_0;
  assign vrfWritePort_9_bits_mask = vrfWritePort_9_bits_mask_0;
  assign vrfWritePort_9_bits_data = vrfWritePort_9_bits_data_0;
  assign vrfWritePort_9_bits_last = vrfWritePort_9_bits_last_0;
  assign vrfWritePort_9_bits_instructionIndex = vrfWritePort_9_bits_instructionIndex_0;
  assign vrfWritePort_10_valid = vrfWritePort_10_valid_0;
  assign vrfWritePort_10_bits_vd = vrfWritePort_10_bits_vd_0;
  assign vrfWritePort_10_bits_offset = vrfWritePort_10_bits_offset_0;
  assign vrfWritePort_10_bits_mask = vrfWritePort_10_bits_mask_0;
  assign vrfWritePort_10_bits_data = vrfWritePort_10_bits_data_0;
  assign vrfWritePort_10_bits_last = vrfWritePort_10_bits_last_0;
  assign vrfWritePort_10_bits_instructionIndex = vrfWritePort_10_bits_instructionIndex_0;
  assign vrfWritePort_11_valid = vrfWritePort_11_valid_0;
  assign vrfWritePort_11_bits_vd = vrfWritePort_11_bits_vd_0;
  assign vrfWritePort_11_bits_offset = vrfWritePort_11_bits_offset_0;
  assign vrfWritePort_11_bits_mask = vrfWritePort_11_bits_mask_0;
  assign vrfWritePort_11_bits_data = vrfWritePort_11_bits_data_0;
  assign vrfWritePort_11_bits_last = vrfWritePort_11_bits_last_0;
  assign vrfWritePort_11_bits_instructionIndex = vrfWritePort_11_bits_instructionIndex_0;
  assign vrfWritePort_12_valid = vrfWritePort_12_valid_0;
  assign vrfWritePort_12_bits_vd = vrfWritePort_12_bits_vd_0;
  assign vrfWritePort_12_bits_offset = vrfWritePort_12_bits_offset_0;
  assign vrfWritePort_12_bits_mask = vrfWritePort_12_bits_mask_0;
  assign vrfWritePort_12_bits_data = vrfWritePort_12_bits_data_0;
  assign vrfWritePort_12_bits_last = vrfWritePort_12_bits_last_0;
  assign vrfWritePort_12_bits_instructionIndex = vrfWritePort_12_bits_instructionIndex_0;
  assign vrfWritePort_13_valid = vrfWritePort_13_valid_0;
  assign vrfWritePort_13_bits_vd = vrfWritePort_13_bits_vd_0;
  assign vrfWritePort_13_bits_offset = vrfWritePort_13_bits_offset_0;
  assign vrfWritePort_13_bits_mask = vrfWritePort_13_bits_mask_0;
  assign vrfWritePort_13_bits_data = vrfWritePort_13_bits_data_0;
  assign vrfWritePort_13_bits_last = vrfWritePort_13_bits_last_0;
  assign vrfWritePort_13_bits_instructionIndex = vrfWritePort_13_bits_instructionIndex_0;
  assign vrfWritePort_14_valid = vrfWritePort_14_valid_0;
  assign vrfWritePort_14_bits_vd = vrfWritePort_14_bits_vd_0;
  assign vrfWritePort_14_bits_offset = vrfWritePort_14_bits_offset_0;
  assign vrfWritePort_14_bits_mask = vrfWritePort_14_bits_mask_0;
  assign vrfWritePort_14_bits_data = vrfWritePort_14_bits_data_0;
  assign vrfWritePort_14_bits_last = vrfWritePort_14_bits_last_0;
  assign vrfWritePort_14_bits_instructionIndex = vrfWritePort_14_bits_instructionIndex_0;
  assign vrfWritePort_15_valid = vrfWritePort_15_valid_0;
  assign vrfWritePort_15_bits_vd = vrfWritePort_15_bits_vd_0;
  assign vrfWritePort_15_bits_offset = vrfWritePort_15_bits_offset_0;
  assign vrfWritePort_15_bits_mask = vrfWritePort_15_bits_mask_0;
  assign vrfWritePort_15_bits_data = vrfWritePort_15_bits_data_0;
  assign vrfWritePort_15_bits_last = vrfWritePort_15_bits_last_0;
  assign vrfWritePort_15_bits_instructionIndex = vrfWritePort_15_bits_instructionIndex_0;
  assign dataInWriteQueue_0 = {dataInWriteQueue_0_hi, dataInWriteQueue_0_lo} | dataInMSHR;
  assign dataInWriteQueue_1 = {dataInWriteQueue_1_hi, dataInWriteQueue_1_lo} | dataInMSHR;
  assign dataInWriteQueue_2 = {dataInWriteQueue_2_hi, dataInWriteQueue_2_lo} | dataInMSHR;
  assign dataInWriteQueue_3 = {dataInWriteQueue_3_hi, dataInWriteQueue_3_lo} | dataInMSHR;
  assign dataInWriteQueue_4 = {dataInWriteQueue_4_hi, dataInWriteQueue_4_lo} | dataInMSHR;
  assign dataInWriteQueue_5 = {dataInWriteQueue_5_hi, dataInWriteQueue_5_lo} | dataInMSHR;
  assign dataInWriteQueue_6 = {dataInWriteQueue_6_hi, dataInWriteQueue_6_lo} | dataInMSHR;
  assign dataInWriteQueue_7 = {dataInWriteQueue_7_hi, dataInWriteQueue_7_lo} | dataInMSHR;
  assign dataInWriteQueue_8 = {dataInWriteQueue_8_hi, dataInWriteQueue_8_lo} | dataInMSHR;
  assign dataInWriteQueue_9 = {dataInWriteQueue_9_hi, dataInWriteQueue_9_lo} | dataInMSHR;
  assign dataInWriteQueue_10 = {dataInWriteQueue_10_hi, dataInWriteQueue_10_lo} | dataInMSHR;
  assign dataInWriteQueue_11 = {dataInWriteQueue_11_hi, dataInWriteQueue_11_lo} | dataInMSHR;
  assign dataInWriteQueue_12 = {dataInWriteQueue_12_hi, dataInWriteQueue_12_lo} | dataInMSHR;
  assign dataInWriteQueue_13 = {dataInWriteQueue_13_hi, dataInWriteQueue_13_lo} | dataInMSHR;
  assign dataInWriteQueue_14 = {dataInWriteQueue_14_hi, dataInWriteQueue_14_lo} | dataInMSHR;
  assign dataInWriteQueue_15 = {dataInWriteQueue_15_hi, dataInWriteQueue_15_lo} | dataInMSHR;
  assign lastReport = (_loadUnit_status_last ? 8'h1 << _GEN_34 : 8'h0) | (_storeUnit_status_last ? 8'h1 << _storeUnit_status_instructionIndex : 8'h0) | (_otherUnit_status_last ? 8'h1 << _GEN_35 : 8'h0);
  assign tokenIO_offsetGroupRelease = {tokenIO_offsetGroupRelease_hi, tokenIO_offsetGroupRelease_lo};
endmodule

