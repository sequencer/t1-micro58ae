module Rsqrt7Fn(
  input  [31:0] in_data,
  input  [9:0]  in_classifyIn,
  output [31:0] out_data,
  output [4:0]  out_exceptionFlags
);

  wire         sign = in_data[31];
  wire [7:0]   expIn = in_data[30:23];
  wire [22:0]  fractIn = in_data[22:0];
  wire         inIsSub = expIn == 8'h0;
  wire         outNaN = |{in_classifyIn[2:0], in_classifyIn[9:8]};
  wire         outInf = in_classifyIn[3] | in_classifyIn[4];
  wire [7:0]   normDist =
    {3'h0,
     fractIn[22]
       ? 5'h0
       : fractIn[21]
           ? 5'h1
           : fractIn[20]
               ? 5'h2
               : fractIn[19]
                   ? 5'h3
                   : fractIn[18]
                       ? 5'h4
                       : fractIn[17]
                           ? 5'h5
                           : fractIn[16]
                               ? 5'h6
                               : fractIn[15]
                                   ? 5'h7
                                   : fractIn[14]
                                       ? 5'h8
                                       : fractIn[13]
                                           ? 5'h9
                                           : fractIn[12]
                                               ? 5'hA
                                               : fractIn[11]
                                                   ? 5'hB
                                                   : fractIn[10]
                                                       ? 5'hC
                                                       : fractIn[9]
                                                           ? 5'hD
                                                           : fractIn[8] ? 5'hE : fractIn[7] ? 5'hF : fractIn[6] ? 5'h10 : fractIn[5] ? 5'h11 : fractIn[4] ? 5'h12 : fractIn[3] ? 5'h13 : fractIn[2] ? 5'h14 : fractIn[1] ? 5'h15 : 5'h16};
  wire [7:0]   normExpIn = inIsSub ? 8'h0 - normDist : expIn;
  wire [278:0] _normSigIn_T_1 = {255'h0, fractIn, 1'h0} << normDist;
  wire [22:0]  normSigIn = inIsSub ? _normSigIn_T_1[22:0] : fractIn;
  wire [6:0]   sigOut_plaInput = {normExpIn[0], normSigIn[22:17]};
  wire [6:0]   sigOut_invInputs = ~sigOut_plaInput;
  wire [6:0]   sigOut_invMatrixOutputs;
  wire         sigOut_andMatrixOutputs_andMatrixInput_0 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_3 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_6 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_7 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_9 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_14 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_15 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_19 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_20 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_21 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_23 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_27 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_28 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_34 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_35 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_37 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_41 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_46 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_55 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_57 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_60 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_62 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_64 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_70 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_71 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_72 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_74 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_81 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_84 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_87 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_89 = sigOut_invInputs[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_1 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_3 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_5 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_8 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_9 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_10 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_14 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_16 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_17 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_19 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_23 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_27 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_30 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_31 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_32 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_37 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_41 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_42 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_44 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_49 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_50 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_51 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_52 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_55 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_57 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_59 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_60 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_64 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_65 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_67 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_68 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_70 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_73 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_74 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_75 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_77 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_81 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_83 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_87 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_90 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_91 = sigOut_invInputs[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_1 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_4 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_4 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_5 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_15 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_15 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_16 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_17 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_21 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_22 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_26 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_32 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_33 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_36 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_39 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_40 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_44 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_45 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_47 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_49 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_52 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_56 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_54 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_61 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_59 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_63 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_64 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_70 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_76 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_74 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_79 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_78 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_84 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_85 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_90 = sigOut_invInputs[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_1 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_2 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_4 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_4 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_5 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_6 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_7 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_8 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_11 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_12 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_20 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_21 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_22 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_24 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_24 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_31 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_31 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_32 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_33 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_35 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_43 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_44 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_48 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_48 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_51 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_52 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_56 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_58 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_59 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_57 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_61 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_60 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_61 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_69 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_78 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_76 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_80 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_83 = sigOut_invInputs[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_2 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_2 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_3 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_2 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_3 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_7 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_5 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_11 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_13 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_14 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_30 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_30 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_31 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_32 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_34 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_38 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_37 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_38 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_32 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_40 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_34 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_53 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_53 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_58 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_56 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_56 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_58 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_60 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_51 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_53 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_64 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_66 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_56 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_58 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_73 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_75 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_79 = sigOut_invInputs[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_79 = sigOut_invInputs[4];
  wire [1:0]   sigOut_andMatrixOutputs_lo = {sigOut_andMatrixOutputs_andMatrixInput_3, sigOut_andMatrixOutputs_andMatrixInput_4};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi = {sigOut_andMatrixOutputs_andMatrixInput_0, sigOut_andMatrixOutputs_andMatrixInput_1};
  wire [2:0]   sigOut_andMatrixOutputs_hi = {sigOut_andMatrixOutputs_hi_hi, sigOut_andMatrixOutputs_andMatrixInput_2};
  wire         sigOut_andMatrixOutputs_27_2 = &{sigOut_andMatrixOutputs_hi, sigOut_andMatrixOutputs_lo};
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_1 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_2 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_1 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_6 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_4 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_1 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_9 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_10 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_6 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_7 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_14 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_10 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_12 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_4 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_16 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_23 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_18 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_25 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_6 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_20 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_27 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_22 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_54 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_51 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_53 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_44 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_55 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_55 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_46 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_57 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_58 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_59 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_62 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_54 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_65 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_24 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_26 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_60 = sigOut_invInputs[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_62 = sigOut_invInputs[5];
  wire [1:0]   sigOut_andMatrixOutputs_lo_1 = {sigOut_andMatrixOutputs_andMatrixInput_2_1, sigOut_andMatrixOutputs_andMatrixInput_3_1};
  wire [1:0]   sigOut_andMatrixOutputs_hi_1 = {sigOut_andMatrixOutputs_andMatrixInput_0_1, sigOut_andMatrixOutputs_andMatrixInput_1_1};
  wire         sigOut_andMatrixOutputs_57_2 = &{sigOut_andMatrixOutputs_hi_1, sigOut_andMatrixOutputs_lo_1};
  wire         sigOut_andMatrixOutputs_92_2 = &{sigOut_andMatrixOutputs_andMatrixInput_0_2, sigOut_andMatrixOutputs_andMatrixInput_1_2};
  wire [1:0]   sigOut_andMatrixOutputs_lo_2 = {sigOut_andMatrixOutputs_andMatrixInput_3_2, sigOut_andMatrixOutputs_andMatrixInput_4_1};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_1 = {sigOut_andMatrixOutputs_andMatrixInput_0_3, sigOut_andMatrixOutputs_andMatrixInput_1_3};
  wire [2:0]   sigOut_andMatrixOutputs_hi_2 = {sigOut_andMatrixOutputs_hi_hi_1, sigOut_andMatrixOutputs_andMatrixInput_2_2};
  wire         sigOut_andMatrixOutputs_63_2 = &{sigOut_andMatrixOutputs_hi_2, sigOut_andMatrixOutputs_lo_2};
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_3 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_9 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_10 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_2 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_8 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_9 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_11 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_3 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_13 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_15 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_5 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_21 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_7 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_23 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_8 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_9 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_10 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_11 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_36 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_13 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_6 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_15 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_37 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_38 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_39 = sigOut_invInputs[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_16 = sigOut_invInputs[6];
  wire [1:0]   sigOut_andMatrixOutputs_lo_3 = {sigOut_andMatrixOutputs_andMatrixInput_2_3, sigOut_andMatrixOutputs_andMatrixInput_3_3};
  wire [1:0]   sigOut_andMatrixOutputs_hi_3 = {sigOut_andMatrixOutputs_andMatrixInput_0_4, sigOut_andMatrixOutputs_andMatrixInput_1_4};
  wire         sigOut_andMatrixOutputs_83_2 = &{sigOut_andMatrixOutputs_hi_3, sigOut_andMatrixOutputs_lo_3};
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_5 = sigOut_plaInput[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_12 = sigOut_plaInput[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_13 = sigOut_plaInput[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_16 = sigOut_plaInput[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_17 = sigOut_plaInput[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_18 = sigOut_plaInput[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_25 = sigOut_plaInput[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_33 = sigOut_plaInput[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_39 = sigOut_plaInput[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_43 = sigOut_plaInput[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_50 = sigOut_plaInput[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_51 = sigOut_plaInput[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_65 = sigOut_plaInput[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_66 = sigOut_plaInput[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_67 = sigOut_plaInput[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_68 = sigOut_plaInput[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_73 = sigOut_plaInput[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_75 = sigOut_plaInput[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_77 = sigOut_plaInput[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_78 = sigOut_plaInput[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_86 = sigOut_plaInput[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_88 = sigOut_plaInput[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_91 = sigOut_plaInput[0];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_92 = sigOut_plaInput[0];
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi = {sigOut_andMatrixOutputs_andMatrixInput_3_4, sigOut_andMatrixOutputs_andMatrixInput_4_2};
  wire [2:0]   sigOut_andMatrixOutputs_lo_4 = {sigOut_andMatrixOutputs_lo_hi, sigOut_andMatrixOutputs_andMatrixInput_5};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_2 = {sigOut_andMatrixOutputs_andMatrixInput_0_5, sigOut_andMatrixOutputs_andMatrixInput_1_5};
  wire [2:0]   sigOut_andMatrixOutputs_hi_4 = {sigOut_andMatrixOutputs_hi_hi_2, sigOut_andMatrixOutputs_andMatrixInput_2_4};
  wire         sigOut_andMatrixOutputs_90_2 = &{sigOut_andMatrixOutputs_hi_4, sigOut_andMatrixOutputs_lo_4};
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_6 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_12 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_13 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_18 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_20 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_22 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_34 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_35 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_36 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_40 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_43 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_45 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_46 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_47 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_48 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_62 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_63 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_66 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_69 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_71 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_72 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_76 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_79 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_82 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_85 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_86 = sigOut_plaInput[1];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_89 = sigOut_plaInput[1];
  wire [1:0]   sigOut_andMatrixOutputs_lo_5 = {sigOut_andMatrixOutputs_andMatrixInput_3_5, sigOut_andMatrixOutputs_andMatrixInput_4_3};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_3 = {sigOut_andMatrixOutputs_andMatrixInput_0_6, sigOut_andMatrixOutputs_andMatrixInput_1_6};
  wire [2:0]   sigOut_andMatrixOutputs_hi_5 = {sigOut_andMatrixOutputs_hi_hi_3, sigOut_andMatrixOutputs_andMatrixInput_2_5};
  wire         sigOut_andMatrixOutputs_2_2 = &{sigOut_andMatrixOutputs_hi_5, sigOut_andMatrixOutputs_lo_5};
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_7 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_8 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_8 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_10 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_11 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_11 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_12 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_18 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_19 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_22 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_24 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_25 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_28 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_29 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_30 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_33 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_34 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_36 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_40 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_42 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_42 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_49 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_50 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_61 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_62 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_63 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_67 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_68 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_69 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_71 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_72 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_80 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_83 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_84 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_88 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_86 = sigOut_plaInput[2];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_92 = sigOut_plaInput[2];
  wire [1:0]   sigOut_andMatrixOutputs_lo_6 = {sigOut_andMatrixOutputs_andMatrixInput_2_6, sigOut_andMatrixOutputs_andMatrixInput_3_6};
  wire [1:0]   sigOut_andMatrixOutputs_hi_6 = {sigOut_andMatrixOutputs_andMatrixInput_0_7, sigOut_andMatrixOutputs_andMatrixInput_1_7};
  wire         sigOut_andMatrixOutputs_16_2 = &{sigOut_andMatrixOutputs_hi_6, sigOut_andMatrixOutputs_lo_6};
  wire [1:0]   sigOut_andMatrixOutputs_lo_7 = {sigOut_andMatrixOutputs_andMatrixInput_3_7, sigOut_andMatrixOutputs_andMatrixInput_4_4};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_4 = {sigOut_andMatrixOutputs_andMatrixInput_0_8, sigOut_andMatrixOutputs_andMatrixInput_1_8};
  wire [2:0]   sigOut_andMatrixOutputs_hi_7 = {sigOut_andMatrixOutputs_hi_hi_4, sigOut_andMatrixOutputs_andMatrixInput_2_7};
  wire         sigOut_andMatrixOutputs_8_2 = &{sigOut_andMatrixOutputs_hi_7, sigOut_andMatrixOutputs_lo_7};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_1 = {sigOut_andMatrixOutputs_andMatrixInput_3_8, sigOut_andMatrixOutputs_andMatrixInput_4_5};
  wire [2:0]   sigOut_andMatrixOutputs_lo_8 = {sigOut_andMatrixOutputs_lo_hi_1, sigOut_andMatrixOutputs_andMatrixInput_5_1};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_5 = {sigOut_andMatrixOutputs_andMatrixInput_0_9, sigOut_andMatrixOutputs_andMatrixInput_1_9};
  wire [2:0]   sigOut_andMatrixOutputs_hi_8 = {sigOut_andMatrixOutputs_hi_hi_5, sigOut_andMatrixOutputs_andMatrixInput_2_8};
  wire         sigOut_andMatrixOutputs_78_2 = &{sigOut_andMatrixOutputs_hi_8, sigOut_andMatrixOutputs_lo_8};
  wire [1:0]   sigOut_andMatrixOutputs_lo_9 = {sigOut_andMatrixOutputs_andMatrixInput_2_9, sigOut_andMatrixOutputs_andMatrixInput_3_9};
  wire [1:0]   sigOut_andMatrixOutputs_hi_9 = {sigOut_andMatrixOutputs_andMatrixInput_0_10, sigOut_andMatrixOutputs_andMatrixInput_1_10};
  wire         sigOut_andMatrixOutputs_60_2 = &{sigOut_andMatrixOutputs_hi_9, sigOut_andMatrixOutputs_lo_9};
  wire [1:0]   sigOut_andMatrixOutputs_lo_10 = {sigOut_andMatrixOutputs_andMatrixInput_2_10, sigOut_andMatrixOutputs_andMatrixInput_3_10};
  wire [1:0]   sigOut_andMatrixOutputs_hi_10 = {sigOut_andMatrixOutputs_andMatrixInput_0_11, sigOut_andMatrixOutputs_andMatrixInput_1_11};
  wire         sigOut_andMatrixOutputs_49_2 = &{sigOut_andMatrixOutputs_hi_10, sigOut_andMatrixOutputs_lo_10};
  wire [1:0]   sigOut_andMatrixOutputs_lo_11 = {sigOut_andMatrixOutputs_andMatrixInput_3_11, sigOut_andMatrixOutputs_andMatrixInput_4_6};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_6 = {sigOut_andMatrixOutputs_andMatrixInput_0_12, sigOut_andMatrixOutputs_andMatrixInput_1_12};
  wire [2:0]   sigOut_andMatrixOutputs_hi_11 = {sigOut_andMatrixOutputs_hi_hi_6, sigOut_andMatrixOutputs_andMatrixInput_2_11};
  wire         sigOut_andMatrixOutputs_34_2 = &{sigOut_andMatrixOutputs_hi_11, sigOut_andMatrixOutputs_lo_11};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_2 = {sigOut_andMatrixOutputs_andMatrixInput_3_12, sigOut_andMatrixOutputs_andMatrixInput_4_7};
  wire [2:0]   sigOut_andMatrixOutputs_lo_12 = {sigOut_andMatrixOutputs_lo_hi_2, sigOut_andMatrixOutputs_andMatrixInput_5_2};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_7 = {sigOut_andMatrixOutputs_andMatrixInput_0_13, sigOut_andMatrixOutputs_andMatrixInput_1_13};
  wire [2:0]   sigOut_andMatrixOutputs_hi_12 = {sigOut_andMatrixOutputs_hi_hi_7, sigOut_andMatrixOutputs_andMatrixInput_2_12};
  wire         sigOut_andMatrixOutputs_19_2 = &{sigOut_andMatrixOutputs_hi_12, sigOut_andMatrixOutputs_lo_12};
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_13 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_14 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_15 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_16 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_17 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_18 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_19 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_26 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_25 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_27 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_29 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_29 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_35 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_0_38 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_38 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_39 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_39 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_41 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_41 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_48 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_49 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_63 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_65 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_69 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_66 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_67 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_68 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_73 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_77 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_82 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_80 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_87 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_88 = sigOut_plaInput[3];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_89 = sigOut_plaInput[3];
  wire [1:0]   sigOut_andMatrixOutputs_lo_13 = {sigOut_andMatrixOutputs_andMatrixInput_3_13, sigOut_andMatrixOutputs_andMatrixInput_4_8};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_8 = {sigOut_andMatrixOutputs_andMatrixInput_0_14, sigOut_andMatrixOutputs_andMatrixInput_1_14};
  wire [2:0]   sigOut_andMatrixOutputs_hi_13 = {sigOut_andMatrixOutputs_hi_hi_8, sigOut_andMatrixOutputs_andMatrixInput_2_13};
  wire         sigOut_andMatrixOutputs_80_2 = &{sigOut_andMatrixOutputs_hi_13, sigOut_andMatrixOutputs_lo_13};
  wire [1:0]   sigOut_andMatrixOutputs_lo_14 = {sigOut_andMatrixOutputs_andMatrixInput_3_14, sigOut_andMatrixOutputs_andMatrixInput_4_9};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_9 = {sigOut_andMatrixOutputs_andMatrixInput_0_15, sigOut_andMatrixOutputs_andMatrixInput_1_15};
  wire [2:0]   sigOut_andMatrixOutputs_hi_14 = {sigOut_andMatrixOutputs_hi_hi_9, sigOut_andMatrixOutputs_andMatrixInput_2_14};
  wire         sigOut_andMatrixOutputs_33_2 = &{sigOut_andMatrixOutputs_hi_14, sigOut_andMatrixOutputs_lo_14};
  wire [1:0]   sigOut_andMatrixOutputs_lo_15 = {sigOut_andMatrixOutputs_andMatrixInput_3_15, sigOut_andMatrixOutputs_andMatrixInput_4_10};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_10 = {sigOut_andMatrixOutputs_andMatrixInput_0_16, sigOut_andMatrixOutputs_andMatrixInput_1_16};
  wire [2:0]   sigOut_andMatrixOutputs_hi_15 = {sigOut_andMatrixOutputs_hi_hi_10, sigOut_andMatrixOutputs_andMatrixInput_2_15};
  wire         sigOut_andMatrixOutputs_77_2 = &{sigOut_andMatrixOutputs_hi_15, sigOut_andMatrixOutputs_lo_15};
  wire [1:0]   sigOut_andMatrixOutputs_lo_16 = {sigOut_andMatrixOutputs_andMatrixInput_3_16, sigOut_andMatrixOutputs_andMatrixInput_4_11};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_11 = {sigOut_andMatrixOutputs_andMatrixInput_0_17, sigOut_andMatrixOutputs_andMatrixInput_1_17};
  wire [2:0]   sigOut_andMatrixOutputs_hi_16 = {sigOut_andMatrixOutputs_hi_hi_11, sigOut_andMatrixOutputs_andMatrixInput_2_16};
  wire         sigOut_andMatrixOutputs_68_2 = &{sigOut_andMatrixOutputs_hi_16, sigOut_andMatrixOutputs_lo_16};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_3 = {sigOut_andMatrixOutputs_andMatrixInput_3_17, sigOut_andMatrixOutputs_andMatrixInput_4_12};
  wire [2:0]   sigOut_andMatrixOutputs_lo_17 = {sigOut_andMatrixOutputs_lo_hi_3, sigOut_andMatrixOutputs_andMatrixInput_5_3};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_12 = {sigOut_andMatrixOutputs_andMatrixInput_0_18, sigOut_andMatrixOutputs_andMatrixInput_1_18};
  wire [2:0]   sigOut_andMatrixOutputs_hi_17 = {sigOut_andMatrixOutputs_hi_hi_12, sigOut_andMatrixOutputs_andMatrixInput_2_17};
  wire         sigOut_andMatrixOutputs_4_2 = &{sigOut_andMatrixOutputs_hi_17, sigOut_andMatrixOutputs_lo_17};
  wire [1:0]   sigOut_andMatrixOutputs_lo_18 = {sigOut_andMatrixOutputs_andMatrixInput_3_18, sigOut_andMatrixOutputs_andMatrixInput_4_13};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_13 = {sigOut_andMatrixOutputs_andMatrixInput_0_19, sigOut_andMatrixOutputs_andMatrixInput_1_19};
  wire [2:0]   sigOut_andMatrixOutputs_hi_18 = {sigOut_andMatrixOutputs_hi_hi_13, sigOut_andMatrixOutputs_andMatrixInput_2_18};
  wire         sigOut_andMatrixOutputs_47_2 = &{sigOut_andMatrixOutputs_hi_18, sigOut_andMatrixOutputs_lo_18};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_4 = {sigOut_andMatrixOutputs_andMatrixInput_3_19, sigOut_andMatrixOutputs_andMatrixInput_4_14};
  wire [2:0]   sigOut_andMatrixOutputs_lo_19 = {sigOut_andMatrixOutputs_lo_hi_4, sigOut_andMatrixOutputs_andMatrixInput_5_4};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_14 = {sigOut_andMatrixOutputs_andMatrixInput_0_20, sigOut_andMatrixOutputs_andMatrixInput_1_20};
  wire [2:0]   sigOut_andMatrixOutputs_hi_19 = {sigOut_andMatrixOutputs_hi_hi_14, sigOut_andMatrixOutputs_andMatrixInput_2_19};
  wire         sigOut_andMatrixOutputs_45_2 = &{sigOut_andMatrixOutputs_hi_19, sigOut_andMatrixOutputs_lo_19};
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_20 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_21 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_17 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_23 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_24 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_26 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_19 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_26 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_28 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_28 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_42 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_43 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_45 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_46 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_47 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_47 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_41 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_42 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_59 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_70 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_71 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_72 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_81 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_82 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_82 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_83 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_85 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_85 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_86 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_87 = sigOut_plaInput[4];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_88 = sigOut_plaInput[4];
  wire [1:0]   sigOut_andMatrixOutputs_lo_20 = {sigOut_andMatrixOutputs_andMatrixInput_3_20, sigOut_andMatrixOutputs_andMatrixInput_4_15};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_15 = {sigOut_andMatrixOutputs_andMatrixInput_0_21, sigOut_andMatrixOutputs_andMatrixInput_1_21};
  wire [2:0]   sigOut_andMatrixOutputs_hi_20 = {sigOut_andMatrixOutputs_hi_hi_15, sigOut_andMatrixOutputs_andMatrixInput_2_20};
  wire         sigOut_andMatrixOutputs_69_2 = &{sigOut_andMatrixOutputs_hi_20, sigOut_andMatrixOutputs_lo_20};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_5 = {sigOut_andMatrixOutputs_andMatrixInput_3_21, sigOut_andMatrixOutputs_andMatrixInput_4_16};
  wire [2:0]   sigOut_andMatrixOutputs_lo_21 = {sigOut_andMatrixOutputs_lo_hi_5, sigOut_andMatrixOutputs_andMatrixInput_5_5};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_16 = {sigOut_andMatrixOutputs_andMatrixInput_0_22, sigOut_andMatrixOutputs_andMatrixInput_1_22};
  wire [2:0]   sigOut_andMatrixOutputs_hi_21 = {sigOut_andMatrixOutputs_hi_hi_16, sigOut_andMatrixOutputs_andMatrixInput_2_21};
  wire         sigOut_andMatrixOutputs_1_2 = &{sigOut_andMatrixOutputs_hi_21, sigOut_andMatrixOutputs_lo_21};
  wire [1:0]   sigOut_andMatrixOutputs_lo_22 = {sigOut_andMatrixOutputs_andMatrixInput_3_22, sigOut_andMatrixOutputs_andMatrixInput_4_17};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_17 = {sigOut_andMatrixOutputs_andMatrixInput_0_23, sigOut_andMatrixOutputs_andMatrixInput_1_23};
  wire [2:0]   sigOut_andMatrixOutputs_hi_22 = {sigOut_andMatrixOutputs_hi_hi_17, sigOut_andMatrixOutputs_andMatrixInput_2_22};
  wire         sigOut_andMatrixOutputs_44_2 = &{sigOut_andMatrixOutputs_hi_22, sigOut_andMatrixOutputs_lo_22};
  wire [1:0]   sigOut_andMatrixOutputs_lo_23 = {sigOut_andMatrixOutputs_andMatrixInput_2_23, sigOut_andMatrixOutputs_andMatrixInput_3_23};
  wire [1:0]   sigOut_andMatrixOutputs_hi_23 = {sigOut_andMatrixOutputs_andMatrixInput_0_24, sigOut_andMatrixOutputs_andMatrixInput_1_24};
  wire         sigOut_andMatrixOutputs_50_2 = &{sigOut_andMatrixOutputs_hi_23, sigOut_andMatrixOutputs_lo_23};
  wire [1:0]   sigOut_andMatrixOutputs_lo_24 = {sigOut_andMatrixOutputs_andMatrixInput_3_24, sigOut_andMatrixOutputs_andMatrixInput_4_18};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_18 = {sigOut_andMatrixOutputs_andMatrixInput_0_25, sigOut_andMatrixOutputs_andMatrixInput_1_25};
  wire [2:0]   sigOut_andMatrixOutputs_hi_24 = {sigOut_andMatrixOutputs_hi_hi_18, sigOut_andMatrixOutputs_andMatrixInput_2_24};
  wire         sigOut_andMatrixOutputs_24_2 = &{sigOut_andMatrixOutputs_hi_24, sigOut_andMatrixOutputs_lo_24};
  wire [1:0]   sigOut_andMatrixOutputs_hi_25 = {sigOut_andMatrixOutputs_andMatrixInput_0_26, sigOut_andMatrixOutputs_andMatrixInput_1_26};
  wire         sigOut_andMatrixOutputs_88_2 = &{sigOut_andMatrixOutputs_hi_25, sigOut_andMatrixOutputs_andMatrixInput_2_25};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_6 = {sigOut_andMatrixOutputs_andMatrixInput_3_25, sigOut_andMatrixOutputs_andMatrixInput_4_19};
  wire [2:0]   sigOut_andMatrixOutputs_lo_25 = {sigOut_andMatrixOutputs_lo_hi_6, sigOut_andMatrixOutputs_andMatrixInput_5_6};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_19 = {sigOut_andMatrixOutputs_andMatrixInput_0_27, sigOut_andMatrixOutputs_andMatrixInput_1_27};
  wire [2:0]   sigOut_andMatrixOutputs_hi_26 = {sigOut_andMatrixOutputs_hi_hi_19, sigOut_andMatrixOutputs_andMatrixInput_2_26};
  wire         sigOut_andMatrixOutputs_25_2 = &{sigOut_andMatrixOutputs_hi_26, sigOut_andMatrixOutputs_lo_25};
  wire [1:0]   sigOut_andMatrixOutputs_lo_26 = {sigOut_andMatrixOutputs_andMatrixInput_3_26, sigOut_andMatrixOutputs_andMatrixInput_4_20};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_20 = {sigOut_andMatrixOutputs_andMatrixInput_0_28, sigOut_andMatrixOutputs_andMatrixInput_1_28};
  wire [2:0]   sigOut_andMatrixOutputs_hi_27 = {sigOut_andMatrixOutputs_hi_hi_20, sigOut_andMatrixOutputs_andMatrixInput_2_27};
  wire         sigOut_andMatrixOutputs_30_2 = &{sigOut_andMatrixOutputs_hi_27, sigOut_andMatrixOutputs_lo_26};
  wire [1:0]   sigOut_andMatrixOutputs_lo_27 = {sigOut_andMatrixOutputs_andMatrixInput_3_27, sigOut_andMatrixOutputs_andMatrixInput_4_21};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_21 = {sigOut_andMatrixOutputs_andMatrixInput_0_29, sigOut_andMatrixOutputs_andMatrixInput_1_29};
  wire [2:0]   sigOut_andMatrixOutputs_hi_28 = {sigOut_andMatrixOutputs_hi_hi_21, sigOut_andMatrixOutputs_andMatrixInput_2_28};
  wire         sigOut_andMatrixOutputs_65_2 = &{sigOut_andMatrixOutputs_hi_28, sigOut_andMatrixOutputs_lo_27};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_7 = {sigOut_andMatrixOutputs_andMatrixInput_3_28, sigOut_andMatrixOutputs_andMatrixInput_4_22};
  wire [2:0]   sigOut_andMatrixOutputs_lo_28 = {sigOut_andMatrixOutputs_lo_hi_7, sigOut_andMatrixOutputs_andMatrixInput_5_7};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_22 = {sigOut_andMatrixOutputs_andMatrixInput_0_30, sigOut_andMatrixOutputs_andMatrixInput_1_30};
  wire [2:0]   sigOut_andMatrixOutputs_hi_29 = {sigOut_andMatrixOutputs_hi_hi_22, sigOut_andMatrixOutputs_andMatrixInput_2_29};
  wire         sigOut_andMatrixOutputs_12_2 = &{sigOut_andMatrixOutputs_hi_29, sigOut_andMatrixOutputs_lo_28};
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_29 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_24 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_25 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_26 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_27 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_28 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_29 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_37 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_30 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_31 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_12 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_33 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_14 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_35 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_36 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_44 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_45 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_46 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_40 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_17 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_18 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_63 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_74 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_75 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_2_77 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_66 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_78 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_68 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_80 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_81 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_71 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_72 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_84 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_74 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_75 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_76 = sigOut_plaInput[5];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_77 = sigOut_plaInput[5];
  wire [1:0]   sigOut_andMatrixOutputs_lo_29 = {sigOut_andMatrixOutputs_andMatrixInput_3_29, sigOut_andMatrixOutputs_andMatrixInput_4_23};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_23 = {sigOut_andMatrixOutputs_andMatrixInput_0_31, sigOut_andMatrixOutputs_andMatrixInput_1_31};
  wire [2:0]   sigOut_andMatrixOutputs_hi_30 = {sigOut_andMatrixOutputs_hi_hi_23, sigOut_andMatrixOutputs_andMatrixInput_2_30};
  wire         sigOut_andMatrixOutputs_15_2 = &{sigOut_andMatrixOutputs_hi_30, sigOut_andMatrixOutputs_lo_29};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_8 = {sigOut_andMatrixOutputs_andMatrixInput_3_30, sigOut_andMatrixOutputs_andMatrixInput_4_24};
  wire [2:0]   sigOut_andMatrixOutputs_lo_30 = {sigOut_andMatrixOutputs_lo_hi_8, sigOut_andMatrixOutputs_andMatrixInput_5_8};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_24 = {sigOut_andMatrixOutputs_andMatrixInput_0_32, sigOut_andMatrixOutputs_andMatrixInput_1_32};
  wire [2:0]   sigOut_andMatrixOutputs_hi_31 = {sigOut_andMatrixOutputs_hi_hi_24, sigOut_andMatrixOutputs_andMatrixInput_2_31};
  wire         sigOut_andMatrixOutputs_5_2 = &{sigOut_andMatrixOutputs_hi_31, sigOut_andMatrixOutputs_lo_30};
  wire [1:0]   sigOut_andMatrixOutputs_lo_31 = {sigOut_andMatrixOutputs_andMatrixInput_3_31, sigOut_andMatrixOutputs_andMatrixInput_4_25};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_25 = {sigOut_andMatrixOutputs_andMatrixInput_0_33, sigOut_andMatrixOutputs_andMatrixInput_1_33};
  wire [2:0]   sigOut_andMatrixOutputs_hi_32 = {sigOut_andMatrixOutputs_hi_hi_25, sigOut_andMatrixOutputs_andMatrixInput_2_32};
  wire         sigOut_andMatrixOutputs_59_2 = &{sigOut_andMatrixOutputs_hi_32, sigOut_andMatrixOutputs_lo_31};
  wire [1:0]   sigOut_andMatrixOutputs_lo_32 = {sigOut_andMatrixOutputs_andMatrixInput_3_32, sigOut_andMatrixOutputs_andMatrixInput_4_26};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_26 = {sigOut_andMatrixOutputs_andMatrixInput_0_34, sigOut_andMatrixOutputs_andMatrixInput_1_34};
  wire [2:0]   sigOut_andMatrixOutputs_hi_33 = {sigOut_andMatrixOutputs_hi_hi_26, sigOut_andMatrixOutputs_andMatrixInput_2_33};
  wire         sigOut_andMatrixOutputs_51_2 = &{sigOut_andMatrixOutputs_hi_33, sigOut_andMatrixOutputs_lo_32};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_9 = {sigOut_andMatrixOutputs_andMatrixInput_3_33, sigOut_andMatrixOutputs_andMatrixInput_4_27};
  wire [2:0]   sigOut_andMatrixOutputs_lo_33 = {sigOut_andMatrixOutputs_lo_hi_9, sigOut_andMatrixOutputs_andMatrixInput_5_9};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_27 = {sigOut_andMatrixOutputs_andMatrixInput_0_35, sigOut_andMatrixOutputs_andMatrixInput_1_35};
  wire [2:0]   sigOut_andMatrixOutputs_hi_34 = {sigOut_andMatrixOutputs_hi_hi_27, sigOut_andMatrixOutputs_andMatrixInput_2_34};
  wire         sigOut_andMatrixOutputs_29_2 = &{sigOut_andMatrixOutputs_hi_34, sigOut_andMatrixOutputs_lo_33};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_10 = {sigOut_andMatrixOutputs_andMatrixInput_3_34, sigOut_andMatrixOutputs_andMatrixInput_4_28};
  wire [2:0]   sigOut_andMatrixOutputs_lo_34 = {sigOut_andMatrixOutputs_lo_hi_10, sigOut_andMatrixOutputs_andMatrixInput_5_10};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_28 = {sigOut_andMatrixOutputs_andMatrixInput_0_36, sigOut_andMatrixOutputs_andMatrixInput_1_36};
  wire [2:0]   sigOut_andMatrixOutputs_hi_35 = {sigOut_andMatrixOutputs_hi_hi_28, sigOut_andMatrixOutputs_andMatrixInput_2_35};
  wire         sigOut_andMatrixOutputs_46_2 = &{sigOut_andMatrixOutputs_hi_35, sigOut_andMatrixOutputs_lo_34};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_11 = {sigOut_andMatrixOutputs_andMatrixInput_3_35, sigOut_andMatrixOutputs_andMatrixInput_4_29};
  wire [2:0]   sigOut_andMatrixOutputs_lo_35 = {sigOut_andMatrixOutputs_lo_hi_11, sigOut_andMatrixOutputs_andMatrixInput_5_11};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_29 = {sigOut_andMatrixOutputs_andMatrixInput_0_37, sigOut_andMatrixOutputs_andMatrixInput_1_37};
  wire [2:0]   sigOut_andMatrixOutputs_hi_36 = {sigOut_andMatrixOutputs_hi_hi_29, sigOut_andMatrixOutputs_andMatrixInput_2_36};
  wire         sigOut_andMatrixOutputs_73_2 = &{sigOut_andMatrixOutputs_hi_36, sigOut_andMatrixOutputs_lo_35};
  wire [1:0]   sigOut_andMatrixOutputs_lo_36 = {sigOut_andMatrixOutputs_andMatrixInput_2_37, sigOut_andMatrixOutputs_andMatrixInput_3_36};
  wire [1:0]   sigOut_andMatrixOutputs_hi_37 = {sigOut_andMatrixOutputs_andMatrixInput_0_38, sigOut_andMatrixOutputs_andMatrixInput_1_38};
  wire         sigOut_andMatrixOutputs_48_2 = &{sigOut_andMatrixOutputs_hi_37, sigOut_andMatrixOutputs_lo_36};
  wire [1:0]   sigOut_andMatrixOutputs_lo_37 = {sigOut_andMatrixOutputs_andMatrixInput_3_37, sigOut_andMatrixOutputs_andMatrixInput_4_30};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_30 = {sigOut_andMatrixOutputs_andMatrixInput_0_39, sigOut_andMatrixOutputs_andMatrixInput_1_39};
  wire [2:0]   sigOut_andMatrixOutputs_hi_38 = {sigOut_andMatrixOutputs_hi_hi_30, sigOut_andMatrixOutputs_andMatrixInput_2_38};
  wire         sigOut_andMatrixOutputs_81_2 = &{sigOut_andMatrixOutputs_hi_38, sigOut_andMatrixOutputs_lo_37};
  wire [1:0]   sigOut_andMatrixOutputs_lo_38 = {sigOut_andMatrixOutputs_andMatrixInput_3_38, sigOut_andMatrixOutputs_andMatrixInput_4_31};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_31 = {sigOut_andMatrixOutputs_andMatrixInput_0_40, sigOut_andMatrixOutputs_andMatrixInput_1_40};
  wire [2:0]   sigOut_andMatrixOutputs_hi_39 = {sigOut_andMatrixOutputs_hi_hi_31, sigOut_andMatrixOutputs_andMatrixInput_2_39};
  wire         sigOut_andMatrixOutputs_38_2 = &{sigOut_andMatrixOutputs_hi_39, sigOut_andMatrixOutputs_lo_38};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_12 = {sigOut_andMatrixOutputs_andMatrixInput_3_39, sigOut_andMatrixOutputs_andMatrixInput_4_32};
  wire [2:0]   sigOut_andMatrixOutputs_lo_39 = {sigOut_andMatrixOutputs_lo_hi_12, sigOut_andMatrixOutputs_andMatrixInput_5_12};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_32 = {sigOut_andMatrixOutputs_andMatrixInput_0_41, sigOut_andMatrixOutputs_andMatrixInput_1_41};
  wire [2:0]   sigOut_andMatrixOutputs_hi_40 = {sigOut_andMatrixOutputs_hi_hi_32, sigOut_andMatrixOutputs_andMatrixInput_2_40};
  wire         sigOut_andMatrixOutputs_53_2 = &{sigOut_andMatrixOutputs_hi_40, sigOut_andMatrixOutputs_lo_39};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_13 = {sigOut_andMatrixOutputs_andMatrixInput_3_40, sigOut_andMatrixOutputs_andMatrixInput_4_33};
  wire [2:0]   sigOut_andMatrixOutputs_lo_40 = {sigOut_andMatrixOutputs_lo_hi_13, sigOut_andMatrixOutputs_andMatrixInput_5_13};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_33 = {sigOut_andMatrixOutputs_andMatrixInput_0_42, sigOut_andMatrixOutputs_andMatrixInput_1_42};
  wire [2:0]   sigOut_andMatrixOutputs_hi_41 = {sigOut_andMatrixOutputs_hi_hi_33, sigOut_andMatrixOutputs_andMatrixInput_2_41};
  wire         sigOut_andMatrixOutputs_35_2 = &{sigOut_andMatrixOutputs_hi_41, sigOut_andMatrixOutputs_lo_40};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_14 = {sigOut_andMatrixOutputs_andMatrixInput_4_34, sigOut_andMatrixOutputs_andMatrixInput_5_14};
  wire [2:0]   sigOut_andMatrixOutputs_lo_41 = {sigOut_andMatrixOutputs_lo_hi_14, sigOut_andMatrixOutputs_andMatrixInput_6};
  wire [1:0]   sigOut_andMatrixOutputs_hi_lo = {sigOut_andMatrixOutputs_andMatrixInput_2_42, sigOut_andMatrixOutputs_andMatrixInput_3_41};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_34 = {sigOut_andMatrixOutputs_andMatrixInput_0_43, sigOut_andMatrixOutputs_andMatrixInput_1_43};
  wire [3:0]   sigOut_andMatrixOutputs_hi_42 = {sigOut_andMatrixOutputs_hi_hi_34, sigOut_andMatrixOutputs_hi_lo};
  wire         sigOut_andMatrixOutputs_17_2 = &{sigOut_andMatrixOutputs_hi_42, sigOut_andMatrixOutputs_lo_41};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_15 = {sigOut_andMatrixOutputs_andMatrixInput_3_42, sigOut_andMatrixOutputs_andMatrixInput_4_35};
  wire [2:0]   sigOut_andMatrixOutputs_lo_42 = {sigOut_andMatrixOutputs_lo_hi_15, sigOut_andMatrixOutputs_andMatrixInput_5_15};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_35 = {sigOut_andMatrixOutputs_andMatrixInput_0_44, sigOut_andMatrixOutputs_andMatrixInput_1_44};
  wire [2:0]   sigOut_andMatrixOutputs_hi_43 = {sigOut_andMatrixOutputs_hi_hi_35, sigOut_andMatrixOutputs_andMatrixInput_2_43};
  wire         sigOut_andMatrixOutputs_56_2 = &{sigOut_andMatrixOutputs_hi_43, sigOut_andMatrixOutputs_lo_42};
  wire [1:0]   sigOut_andMatrixOutputs_lo_43 = {sigOut_andMatrixOutputs_andMatrixInput_3_43, sigOut_andMatrixOutputs_andMatrixInput_4_36};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_36 = {sigOut_andMatrixOutputs_andMatrixInput_0_45, sigOut_andMatrixOutputs_andMatrixInput_1_45};
  wire [2:0]   sigOut_andMatrixOutputs_hi_44 = {sigOut_andMatrixOutputs_hi_hi_36, sigOut_andMatrixOutputs_andMatrixInput_2_44};
  wire         sigOut_andMatrixOutputs_13_2 = &{sigOut_andMatrixOutputs_hi_44, sigOut_andMatrixOutputs_lo_43};
  wire [1:0]   sigOut_andMatrixOutputs_lo_44 = {sigOut_andMatrixOutputs_andMatrixInput_3_44, sigOut_andMatrixOutputs_andMatrixInput_4_37};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_37 = {sigOut_andMatrixOutputs_andMatrixInput_0_46, sigOut_andMatrixOutputs_andMatrixInput_1_46};
  wire [2:0]   sigOut_andMatrixOutputs_hi_45 = {sigOut_andMatrixOutputs_hi_hi_37, sigOut_andMatrixOutputs_andMatrixInput_2_45};
  wire         sigOut_andMatrixOutputs_41_2 = &{sigOut_andMatrixOutputs_hi_45, sigOut_andMatrixOutputs_lo_44};
  wire [1:0]   sigOut_andMatrixOutputs_lo_45 = {sigOut_andMatrixOutputs_andMatrixInput_3_45, sigOut_andMatrixOutputs_andMatrixInput_4_38};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_38 = {sigOut_andMatrixOutputs_andMatrixInput_0_47, sigOut_andMatrixOutputs_andMatrixInput_1_47};
  wire [2:0]   sigOut_andMatrixOutputs_hi_46 = {sigOut_andMatrixOutputs_hi_hi_38, sigOut_andMatrixOutputs_andMatrixInput_2_46};
  wire         sigOut_andMatrixOutputs_62_2 = &{sigOut_andMatrixOutputs_hi_46, sigOut_andMatrixOutputs_lo_45};
  wire [1:0]   sigOut_andMatrixOutputs_lo_46 = {sigOut_andMatrixOutputs_andMatrixInput_3_46, sigOut_andMatrixOutputs_andMatrixInput_4_39};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_39 = {sigOut_andMatrixOutputs_andMatrixInput_0_48, sigOut_andMatrixOutputs_andMatrixInput_1_48};
  wire [2:0]   sigOut_andMatrixOutputs_hi_47 = {sigOut_andMatrixOutputs_hi_hi_39, sigOut_andMatrixOutputs_andMatrixInput_2_47};
  wire         sigOut_andMatrixOutputs_75_2 = &{sigOut_andMatrixOutputs_hi_47, sigOut_andMatrixOutputs_lo_46};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_16 = {sigOut_andMatrixOutputs_andMatrixInput_3_47, sigOut_andMatrixOutputs_andMatrixInput_4_40};
  wire [2:0]   sigOut_andMatrixOutputs_lo_47 = {sigOut_andMatrixOutputs_lo_hi_16, sigOut_andMatrixOutputs_andMatrixInput_5_16};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_40 = {sigOut_andMatrixOutputs_andMatrixInput_0_49, sigOut_andMatrixOutputs_andMatrixInput_1_49};
  wire [2:0]   sigOut_andMatrixOutputs_hi_48 = {sigOut_andMatrixOutputs_hi_hi_40, sigOut_andMatrixOutputs_andMatrixInput_2_48};
  wire         sigOut_andMatrixOutputs_86_2 = &{sigOut_andMatrixOutputs_hi_48, sigOut_andMatrixOutputs_lo_47};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_17 = {sigOut_andMatrixOutputs_andMatrixInput_3_48, sigOut_andMatrixOutputs_andMatrixInput_4_41};
  wire [2:0]   sigOut_andMatrixOutputs_lo_48 = {sigOut_andMatrixOutputs_lo_hi_17, sigOut_andMatrixOutputs_andMatrixInput_5_17};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_41 = {sigOut_andMatrixOutputs_andMatrixInput_0_50, sigOut_andMatrixOutputs_andMatrixInput_1_50};
  wire [2:0]   sigOut_andMatrixOutputs_hi_49 = {sigOut_andMatrixOutputs_hi_hi_41, sigOut_andMatrixOutputs_andMatrixInput_2_49};
  wire         sigOut_andMatrixOutputs_40_2 = &{sigOut_andMatrixOutputs_hi_49, sigOut_andMatrixOutputs_lo_48};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_18 = {sigOut_andMatrixOutputs_andMatrixInput_3_49, sigOut_andMatrixOutputs_andMatrixInput_4_42};
  wire [2:0]   sigOut_andMatrixOutputs_lo_49 = {sigOut_andMatrixOutputs_lo_hi_18, sigOut_andMatrixOutputs_andMatrixInput_5_18};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_42 = {sigOut_andMatrixOutputs_andMatrixInput_0_51, sigOut_andMatrixOutputs_andMatrixInput_1_51};
  wire [2:0]   sigOut_andMatrixOutputs_hi_50 = {sigOut_andMatrixOutputs_hi_hi_42, sigOut_andMatrixOutputs_andMatrixInput_2_50};
  wire         sigOut_andMatrixOutputs_18_2 = &{sigOut_andMatrixOutputs_hi_50, sigOut_andMatrixOutputs_lo_49};
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_50 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_53 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_1_54 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_43 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_52 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_19 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_54 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_45 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_20 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_47 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_48 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_49 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_50 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_21 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_52 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_22 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_23 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_55 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_6_1 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_57 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_25 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_6_2 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_27 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_61 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_28 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_29 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_64 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_65 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_3_76 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_30 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_67 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_31 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_69 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_70 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_32 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_33 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_4_73 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_34 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_35 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_36 = sigOut_plaInput[6];
  wire         sigOut_andMatrixOutputs_andMatrixInput_5_37 = sigOut_plaInput[6];
  wire [1:0]   sigOut_andMatrixOutputs_lo_50 = {sigOut_andMatrixOutputs_andMatrixInput_2_51, sigOut_andMatrixOutputs_andMatrixInput_3_50};
  wire [1:0]   sigOut_andMatrixOutputs_hi_51 = {sigOut_andMatrixOutputs_andMatrixInput_0_52, sigOut_andMatrixOutputs_andMatrixInput_1_52};
  wire         sigOut_andMatrixOutputs_66_2 = &{sigOut_andMatrixOutputs_hi_51, sigOut_andMatrixOutputs_lo_50};
  wire         sigOut_andMatrixOutputs_72_2 = &{sigOut_andMatrixOutputs_andMatrixInput_0_53, sigOut_andMatrixOutputs_andMatrixInput_1_53};
  wire         sigOut_andMatrixOutputs_55_2 = &{sigOut_andMatrixOutputs_andMatrixInput_0_54, sigOut_andMatrixOutputs_andMatrixInput_1_54};
  wire [1:0]   sigOut_andMatrixOutputs_lo_51 = {sigOut_andMatrixOutputs_andMatrixInput_3_51, sigOut_andMatrixOutputs_andMatrixInput_4_43};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_43 = {sigOut_andMatrixOutputs_andMatrixInput_0_55, sigOut_andMatrixOutputs_andMatrixInput_1_55};
  wire [2:0]   sigOut_andMatrixOutputs_hi_52 = {sigOut_andMatrixOutputs_hi_hi_43, sigOut_andMatrixOutputs_andMatrixInput_2_52};
  wire         sigOut_andMatrixOutputs_37_2 = &{sigOut_andMatrixOutputs_hi_52, sigOut_andMatrixOutputs_lo_51};
  wire [1:0]   sigOut_andMatrixOutputs_lo_52 = {sigOut_andMatrixOutputs_andMatrixInput_2_53, sigOut_andMatrixOutputs_andMatrixInput_3_52};
  wire [1:0]   sigOut_andMatrixOutputs_hi_53 = {sigOut_andMatrixOutputs_andMatrixInput_0_56, sigOut_andMatrixOutputs_andMatrixInput_1_56};
  wire         sigOut_andMatrixOutputs_32_2 = &{sigOut_andMatrixOutputs_hi_53, sigOut_andMatrixOutputs_lo_52};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_19 = {sigOut_andMatrixOutputs_andMatrixInput_3_53, sigOut_andMatrixOutputs_andMatrixInput_4_44};
  wire [2:0]   sigOut_andMatrixOutputs_lo_53 = {sigOut_andMatrixOutputs_lo_hi_19, sigOut_andMatrixOutputs_andMatrixInput_5_19};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_44 = {sigOut_andMatrixOutputs_andMatrixInput_0_57, sigOut_andMatrixOutputs_andMatrixInput_1_57};
  wire [2:0]   sigOut_andMatrixOutputs_hi_54 = {sigOut_andMatrixOutputs_hi_hi_44, sigOut_andMatrixOutputs_andMatrixInput_2_54};
  wire         sigOut_andMatrixOutputs_7_2 = &{sigOut_andMatrixOutputs_hi_54, sigOut_andMatrixOutputs_lo_53};
  wire [1:0]   sigOut_andMatrixOutputs_lo_54 = {sigOut_andMatrixOutputs_andMatrixInput_2_55, sigOut_andMatrixOutputs_andMatrixInput_3_54};
  wire [1:0]   sigOut_andMatrixOutputs_hi_55 = {sigOut_andMatrixOutputs_andMatrixInput_0_58, sigOut_andMatrixOutputs_andMatrixInput_1_58};
  wire         sigOut_andMatrixOutputs_84_2 = &{sigOut_andMatrixOutputs_hi_55, sigOut_andMatrixOutputs_lo_54};
  wire [1:0]   sigOut_andMatrixOutputs_lo_55 = {sigOut_andMatrixOutputs_andMatrixInput_3_55, sigOut_andMatrixOutputs_andMatrixInput_4_45};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_45 = {sigOut_andMatrixOutputs_andMatrixInput_0_59, sigOut_andMatrixOutputs_andMatrixInput_1_59};
  wire [2:0]   sigOut_andMatrixOutputs_hi_56 = {sigOut_andMatrixOutputs_hi_hi_45, sigOut_andMatrixOutputs_andMatrixInput_2_56};
  wire         sigOut_andMatrixOutputs_85_2 = &{sigOut_andMatrixOutputs_hi_56, sigOut_andMatrixOutputs_lo_55};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_20 = {sigOut_andMatrixOutputs_andMatrixInput_3_56, sigOut_andMatrixOutputs_andMatrixInput_4_46};
  wire [2:0]   sigOut_andMatrixOutputs_lo_56 = {sigOut_andMatrixOutputs_lo_hi_20, sigOut_andMatrixOutputs_andMatrixInput_5_20};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_46 = {sigOut_andMatrixOutputs_andMatrixInput_0_60, sigOut_andMatrixOutputs_andMatrixInput_1_60};
  wire [2:0]   sigOut_andMatrixOutputs_hi_57 = {sigOut_andMatrixOutputs_hi_hi_46, sigOut_andMatrixOutputs_andMatrixInput_2_57};
  wire         sigOut_andMatrixOutputs_71_2 = &{sigOut_andMatrixOutputs_hi_57, sigOut_andMatrixOutputs_lo_56};
  wire [1:0]   sigOut_andMatrixOutputs_lo_57 = {sigOut_andMatrixOutputs_andMatrixInput_3_57, sigOut_andMatrixOutputs_andMatrixInput_4_47};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_47 = {sigOut_andMatrixOutputs_andMatrixInput_0_61, sigOut_andMatrixOutputs_andMatrixInput_1_61};
  wire [2:0]   sigOut_andMatrixOutputs_hi_58 = {sigOut_andMatrixOutputs_hi_hi_47, sigOut_andMatrixOutputs_andMatrixInput_2_58};
  wire         sigOut_andMatrixOutputs_76_2 = &{sigOut_andMatrixOutputs_hi_58, sigOut_andMatrixOutputs_lo_57};
  wire [1:0]   sigOut_andMatrixOutputs_lo_58 = {sigOut_andMatrixOutputs_andMatrixInput_3_58, sigOut_andMatrixOutputs_andMatrixInput_4_48};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_48 = {sigOut_andMatrixOutputs_andMatrixInput_0_62, sigOut_andMatrixOutputs_andMatrixInput_1_62};
  wire [2:0]   sigOut_andMatrixOutputs_hi_59 = {sigOut_andMatrixOutputs_hi_hi_48, sigOut_andMatrixOutputs_andMatrixInput_2_59};
  wire         sigOut_andMatrixOutputs_0_2 = &{sigOut_andMatrixOutputs_hi_59, sigOut_andMatrixOutputs_lo_58};
  wire [1:0]   sigOut_andMatrixOutputs_lo_59 = {sigOut_andMatrixOutputs_andMatrixInput_3_59, sigOut_andMatrixOutputs_andMatrixInput_4_49};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_49 = {sigOut_andMatrixOutputs_andMatrixInput_0_63, sigOut_andMatrixOutputs_andMatrixInput_1_63};
  wire [2:0]   sigOut_andMatrixOutputs_hi_60 = {sigOut_andMatrixOutputs_hi_hi_49, sigOut_andMatrixOutputs_andMatrixInput_2_60};
  wire         sigOut_andMatrixOutputs_52_2 = &{sigOut_andMatrixOutputs_hi_60, sigOut_andMatrixOutputs_lo_59};
  wire [1:0]   sigOut_andMatrixOutputs_lo_60 = {sigOut_andMatrixOutputs_andMatrixInput_3_60, sigOut_andMatrixOutputs_andMatrixInput_4_50};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_50 = {sigOut_andMatrixOutputs_andMatrixInput_0_64, sigOut_andMatrixOutputs_andMatrixInput_1_64};
  wire [2:0]   sigOut_andMatrixOutputs_hi_61 = {sigOut_andMatrixOutputs_hi_hi_50, sigOut_andMatrixOutputs_andMatrixInput_2_61};
  wire         sigOut_andMatrixOutputs_26_2 = &{sigOut_andMatrixOutputs_hi_61, sigOut_andMatrixOutputs_lo_60};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_21 = {sigOut_andMatrixOutputs_andMatrixInput_3_61, sigOut_andMatrixOutputs_andMatrixInput_4_51};
  wire [2:0]   sigOut_andMatrixOutputs_lo_61 = {sigOut_andMatrixOutputs_lo_hi_21, sigOut_andMatrixOutputs_andMatrixInput_5_21};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_51 = {sigOut_andMatrixOutputs_andMatrixInput_0_65, sigOut_andMatrixOutputs_andMatrixInput_1_65};
  wire [2:0]   sigOut_andMatrixOutputs_hi_62 = {sigOut_andMatrixOutputs_hi_hi_51, sigOut_andMatrixOutputs_andMatrixInput_2_62};
  wire         sigOut_andMatrixOutputs_42_2 = &{sigOut_andMatrixOutputs_hi_62, sigOut_andMatrixOutputs_lo_61};
  wire [1:0]   sigOut_andMatrixOutputs_lo_62 = {sigOut_andMatrixOutputs_andMatrixInput_3_62, sigOut_andMatrixOutputs_andMatrixInput_4_52};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_52 = {sigOut_andMatrixOutputs_andMatrixInput_0_66, sigOut_andMatrixOutputs_andMatrixInput_1_66};
  wire [2:0]   sigOut_andMatrixOutputs_hi_63 = {sigOut_andMatrixOutputs_hi_hi_52, sigOut_andMatrixOutputs_andMatrixInput_2_63};
  wire         sigOut_andMatrixOutputs_70_2 = &{sigOut_andMatrixOutputs_hi_63, sigOut_andMatrixOutputs_lo_62};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_22 = {sigOut_andMatrixOutputs_andMatrixInput_3_63, sigOut_andMatrixOutputs_andMatrixInput_4_53};
  wire [2:0]   sigOut_andMatrixOutputs_lo_63 = {sigOut_andMatrixOutputs_lo_hi_22, sigOut_andMatrixOutputs_andMatrixInput_5_22};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_53 = {sigOut_andMatrixOutputs_andMatrixInput_0_67, sigOut_andMatrixOutputs_andMatrixInput_1_67};
  wire [2:0]   sigOut_andMatrixOutputs_hi_64 = {sigOut_andMatrixOutputs_hi_hi_53, sigOut_andMatrixOutputs_andMatrixInput_2_64};
  wire         sigOut_andMatrixOutputs_36_2 = &{sigOut_andMatrixOutputs_hi_64, sigOut_andMatrixOutputs_lo_63};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_23 = {sigOut_andMatrixOutputs_andMatrixInput_3_64, sigOut_andMatrixOutputs_andMatrixInput_4_54};
  wire [2:0]   sigOut_andMatrixOutputs_lo_64 = {sigOut_andMatrixOutputs_lo_hi_23, sigOut_andMatrixOutputs_andMatrixInput_5_23};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_54 = {sigOut_andMatrixOutputs_andMatrixInput_0_68, sigOut_andMatrixOutputs_andMatrixInput_1_68};
  wire [2:0]   sigOut_andMatrixOutputs_hi_65 = {sigOut_andMatrixOutputs_hi_hi_54, sigOut_andMatrixOutputs_andMatrixInput_2_65};
  wire         sigOut_andMatrixOutputs_39_2 = &{sigOut_andMatrixOutputs_hi_65, sigOut_andMatrixOutputs_lo_64};
  wire [1:0]   sigOut_andMatrixOutputs_lo_65 = {sigOut_andMatrixOutputs_andMatrixInput_3_65, sigOut_andMatrixOutputs_andMatrixInput_4_55};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_55 = {sigOut_andMatrixOutputs_andMatrixInput_0_69, sigOut_andMatrixOutputs_andMatrixInput_1_69};
  wire [2:0]   sigOut_andMatrixOutputs_hi_66 = {sigOut_andMatrixOutputs_hi_hi_55, sigOut_andMatrixOutputs_andMatrixInput_2_66};
  wire         sigOut_andMatrixOutputs_67_2 = &{sigOut_andMatrixOutputs_hi_66, sigOut_andMatrixOutputs_lo_65};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_24 = {sigOut_andMatrixOutputs_andMatrixInput_4_56, sigOut_andMatrixOutputs_andMatrixInput_5_24};
  wire [2:0]   sigOut_andMatrixOutputs_lo_66 = {sigOut_andMatrixOutputs_lo_hi_24, sigOut_andMatrixOutputs_andMatrixInput_6_1};
  wire [1:0]   sigOut_andMatrixOutputs_hi_lo_1 = {sigOut_andMatrixOutputs_andMatrixInput_2_67, sigOut_andMatrixOutputs_andMatrixInput_3_66};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_56 = {sigOut_andMatrixOutputs_andMatrixInput_0_70, sigOut_andMatrixOutputs_andMatrixInput_1_70};
  wire [3:0]   sigOut_andMatrixOutputs_hi_67 = {sigOut_andMatrixOutputs_hi_hi_56, sigOut_andMatrixOutputs_hi_lo_1};
  wire         sigOut_andMatrixOutputs_64_2 = &{sigOut_andMatrixOutputs_hi_67, sigOut_andMatrixOutputs_lo_66};
  wire [1:0]   sigOut_andMatrixOutputs_lo_67 = {sigOut_andMatrixOutputs_andMatrixInput_3_67, sigOut_andMatrixOutputs_andMatrixInput_4_57};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_57 = {sigOut_andMatrixOutputs_andMatrixInput_0_71, sigOut_andMatrixOutputs_andMatrixInput_1_71};
  wire [2:0]   sigOut_andMatrixOutputs_hi_68 = {sigOut_andMatrixOutputs_hi_hi_57, sigOut_andMatrixOutputs_andMatrixInput_2_68};
  wire         sigOut_andMatrixOutputs_10_2 = &{sigOut_andMatrixOutputs_hi_68, sigOut_andMatrixOutputs_lo_67};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_25 = {sigOut_andMatrixOutputs_andMatrixInput_3_68, sigOut_andMatrixOutputs_andMatrixInput_4_58};
  wire [2:0]   sigOut_andMatrixOutputs_lo_68 = {sigOut_andMatrixOutputs_lo_hi_25, sigOut_andMatrixOutputs_andMatrixInput_5_25};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_58 = {sigOut_andMatrixOutputs_andMatrixInput_0_72, sigOut_andMatrixOutputs_andMatrixInput_1_72};
  wire [2:0]   sigOut_andMatrixOutputs_hi_69 = {sigOut_andMatrixOutputs_hi_hi_58, sigOut_andMatrixOutputs_andMatrixInput_2_69};
  wire         sigOut_andMatrixOutputs_22_2 = &{sigOut_andMatrixOutputs_hi_69, sigOut_andMatrixOutputs_lo_68};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_26 = {sigOut_andMatrixOutputs_andMatrixInput_4_59, sigOut_andMatrixOutputs_andMatrixInput_5_26};
  wire [2:0]   sigOut_andMatrixOutputs_lo_69 = {sigOut_andMatrixOutputs_lo_hi_26, sigOut_andMatrixOutputs_andMatrixInput_6_2};
  wire [1:0]   sigOut_andMatrixOutputs_hi_lo_2 = {sigOut_andMatrixOutputs_andMatrixInput_2_70, sigOut_andMatrixOutputs_andMatrixInput_3_69};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_59 = {sigOut_andMatrixOutputs_andMatrixInput_0_73, sigOut_andMatrixOutputs_andMatrixInput_1_73};
  wire [3:0]   sigOut_andMatrixOutputs_hi_70 = {sigOut_andMatrixOutputs_hi_hi_59, sigOut_andMatrixOutputs_hi_lo_2};
  wire         sigOut_andMatrixOutputs_20_2 = &{sigOut_andMatrixOutputs_hi_70, sigOut_andMatrixOutputs_lo_69};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_27 = {sigOut_andMatrixOutputs_andMatrixInput_3_70, sigOut_andMatrixOutputs_andMatrixInput_4_60};
  wire [2:0]   sigOut_andMatrixOutputs_lo_70 = {sigOut_andMatrixOutputs_lo_hi_27, sigOut_andMatrixOutputs_andMatrixInput_5_27};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_60 = {sigOut_andMatrixOutputs_andMatrixInput_0_74, sigOut_andMatrixOutputs_andMatrixInput_1_74};
  wire [2:0]   sigOut_andMatrixOutputs_hi_71 = {sigOut_andMatrixOutputs_hi_hi_60, sigOut_andMatrixOutputs_andMatrixInput_2_71};
  wire         sigOut_andMatrixOutputs_31_2 = &{sigOut_andMatrixOutputs_hi_71, sigOut_andMatrixOutputs_lo_70};
  wire [1:0]   sigOut_andMatrixOutputs_lo_71 = {sigOut_andMatrixOutputs_andMatrixInput_3_71, sigOut_andMatrixOutputs_andMatrixInput_4_61};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_61 = {sigOut_andMatrixOutputs_andMatrixInput_0_75, sigOut_andMatrixOutputs_andMatrixInput_1_75};
  wire [2:0]   sigOut_andMatrixOutputs_hi_72 = {sigOut_andMatrixOutputs_hi_hi_61, sigOut_andMatrixOutputs_andMatrixInput_2_72};
  wire         sigOut_andMatrixOutputs_61_2 = &{sigOut_andMatrixOutputs_hi_72, sigOut_andMatrixOutputs_lo_71};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_28 = {sigOut_andMatrixOutputs_andMatrixInput_3_72, sigOut_andMatrixOutputs_andMatrixInput_4_62};
  wire [2:0]   sigOut_andMatrixOutputs_lo_72 = {sigOut_andMatrixOutputs_lo_hi_28, sigOut_andMatrixOutputs_andMatrixInput_5_28};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_62 = {sigOut_andMatrixOutputs_andMatrixInput_0_76, sigOut_andMatrixOutputs_andMatrixInput_1_76};
  wire [2:0]   sigOut_andMatrixOutputs_hi_73 = {sigOut_andMatrixOutputs_hi_hi_62, sigOut_andMatrixOutputs_andMatrixInput_2_73};
  wire         sigOut_andMatrixOutputs_87_2 = &{sigOut_andMatrixOutputs_hi_73, sigOut_andMatrixOutputs_lo_72};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_29 = {sigOut_andMatrixOutputs_andMatrixInput_3_73, sigOut_andMatrixOutputs_andMatrixInput_4_63};
  wire [2:0]   sigOut_andMatrixOutputs_lo_73 = {sigOut_andMatrixOutputs_lo_hi_29, sigOut_andMatrixOutputs_andMatrixInput_5_29};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_63 = {sigOut_andMatrixOutputs_andMatrixInput_0_77, sigOut_andMatrixOutputs_andMatrixInput_1_77};
  wire [2:0]   sigOut_andMatrixOutputs_hi_74 = {sigOut_andMatrixOutputs_hi_hi_63, sigOut_andMatrixOutputs_andMatrixInput_2_74};
  wire         sigOut_andMatrixOutputs_11_2 = &{sigOut_andMatrixOutputs_hi_74, sigOut_andMatrixOutputs_lo_73};
  wire [1:0]   sigOut_andMatrixOutputs_lo_74 = {sigOut_andMatrixOutputs_andMatrixInput_3_74, sigOut_andMatrixOutputs_andMatrixInput_4_64};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_64 = {sigOut_andMatrixOutputs_andMatrixInput_0_78, sigOut_andMatrixOutputs_andMatrixInput_1_78};
  wire [2:0]   sigOut_andMatrixOutputs_hi_75 = {sigOut_andMatrixOutputs_hi_hi_64, sigOut_andMatrixOutputs_andMatrixInput_2_75};
  wire         sigOut_andMatrixOutputs_91_2 = &{sigOut_andMatrixOutputs_hi_75, sigOut_andMatrixOutputs_lo_74};
  wire [1:0]   sigOut_andMatrixOutputs_lo_75 = {sigOut_andMatrixOutputs_andMatrixInput_3_75, sigOut_andMatrixOutputs_andMatrixInput_4_65};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_65 = {sigOut_andMatrixOutputs_andMatrixInput_0_79, sigOut_andMatrixOutputs_andMatrixInput_1_79};
  wire [2:0]   sigOut_andMatrixOutputs_hi_76 = {sigOut_andMatrixOutputs_hi_hi_65, sigOut_andMatrixOutputs_andMatrixInput_2_76};
  wire         sigOut_andMatrixOutputs_89_2 = &{sigOut_andMatrixOutputs_hi_76, sigOut_andMatrixOutputs_lo_75};
  wire [1:0]   sigOut_andMatrixOutputs_lo_76 = {sigOut_andMatrixOutputs_andMatrixInput_2_77, sigOut_andMatrixOutputs_andMatrixInput_3_76};
  wire [1:0]   sigOut_andMatrixOutputs_hi_77 = {sigOut_andMatrixOutputs_andMatrixInput_0_80, sigOut_andMatrixOutputs_andMatrixInput_1_80};
  wire         sigOut_andMatrixOutputs_58_2 = &{sigOut_andMatrixOutputs_hi_77, sigOut_andMatrixOutputs_lo_76};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_30 = {sigOut_andMatrixOutputs_andMatrixInput_3_77, sigOut_andMatrixOutputs_andMatrixInput_4_66};
  wire [2:0]   sigOut_andMatrixOutputs_lo_77 = {sigOut_andMatrixOutputs_lo_hi_30, sigOut_andMatrixOutputs_andMatrixInput_5_30};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_66 = {sigOut_andMatrixOutputs_andMatrixInput_0_81, sigOut_andMatrixOutputs_andMatrixInput_1_81};
  wire [2:0]   sigOut_andMatrixOutputs_hi_78 = {sigOut_andMatrixOutputs_hi_hi_66, sigOut_andMatrixOutputs_andMatrixInput_2_78};
  wire         sigOut_andMatrixOutputs_43_2 = &{sigOut_andMatrixOutputs_hi_78, sigOut_andMatrixOutputs_lo_77};
  wire [1:0]   sigOut_andMatrixOutputs_lo_78 = {sigOut_andMatrixOutputs_andMatrixInput_3_78, sigOut_andMatrixOutputs_andMatrixInput_4_67};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_67 = {sigOut_andMatrixOutputs_andMatrixInput_0_82, sigOut_andMatrixOutputs_andMatrixInput_1_82};
  wire [2:0]   sigOut_andMatrixOutputs_hi_79 = {sigOut_andMatrixOutputs_hi_hi_67, sigOut_andMatrixOutputs_andMatrixInput_2_79};
  wire         sigOut_andMatrixOutputs_3_2 = &{sigOut_andMatrixOutputs_hi_79, sigOut_andMatrixOutputs_lo_78};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_31 = {sigOut_andMatrixOutputs_andMatrixInput_3_79, sigOut_andMatrixOutputs_andMatrixInput_4_68};
  wire [2:0]   sigOut_andMatrixOutputs_lo_79 = {sigOut_andMatrixOutputs_lo_hi_31, sigOut_andMatrixOutputs_andMatrixInput_5_31};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_68 = {sigOut_andMatrixOutputs_andMatrixInput_0_83, sigOut_andMatrixOutputs_andMatrixInput_1_83};
  wire [2:0]   sigOut_andMatrixOutputs_hi_80 = {sigOut_andMatrixOutputs_hi_hi_68, sigOut_andMatrixOutputs_andMatrixInput_2_80};
  wire         sigOut_andMatrixOutputs_21_2 = &{sigOut_andMatrixOutputs_hi_80, sigOut_andMatrixOutputs_lo_79};
  wire [1:0]   sigOut_andMatrixOutputs_lo_80 = {sigOut_andMatrixOutputs_andMatrixInput_3_80, sigOut_andMatrixOutputs_andMatrixInput_4_69};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_69 = {sigOut_andMatrixOutputs_andMatrixInput_0_84, sigOut_andMatrixOutputs_andMatrixInput_1_84};
  wire [2:0]   sigOut_andMatrixOutputs_hi_81 = {sigOut_andMatrixOutputs_hi_hi_69, sigOut_andMatrixOutputs_andMatrixInput_2_81};
  wire         sigOut_andMatrixOutputs_79_2 = &{sigOut_andMatrixOutputs_hi_81, sigOut_andMatrixOutputs_lo_80};
  wire [1:0]   sigOut_andMatrixOutputs_lo_81 = {sigOut_andMatrixOutputs_andMatrixInput_3_81, sigOut_andMatrixOutputs_andMatrixInput_4_70};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_70 = {sigOut_andMatrixOutputs_andMatrixInput_0_85, sigOut_andMatrixOutputs_andMatrixInput_1_85};
  wire [2:0]   sigOut_andMatrixOutputs_hi_82 = {sigOut_andMatrixOutputs_hi_hi_70, sigOut_andMatrixOutputs_andMatrixInput_2_82};
  wire         sigOut_andMatrixOutputs_6_2 = &{sigOut_andMatrixOutputs_hi_82, sigOut_andMatrixOutputs_lo_81};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_32 = {sigOut_andMatrixOutputs_andMatrixInput_3_82, sigOut_andMatrixOutputs_andMatrixInput_4_71};
  wire [2:0]   sigOut_andMatrixOutputs_lo_82 = {sigOut_andMatrixOutputs_lo_hi_32, sigOut_andMatrixOutputs_andMatrixInput_5_32};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_71 = {sigOut_andMatrixOutputs_andMatrixInput_0_86, sigOut_andMatrixOutputs_andMatrixInput_1_86};
  wire [2:0]   sigOut_andMatrixOutputs_hi_83 = {sigOut_andMatrixOutputs_hi_hi_71, sigOut_andMatrixOutputs_andMatrixInput_2_83};
  wire         sigOut_andMatrixOutputs_54_2 = &{sigOut_andMatrixOutputs_hi_83, sigOut_andMatrixOutputs_lo_82};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_33 = {sigOut_andMatrixOutputs_andMatrixInput_3_83, sigOut_andMatrixOutputs_andMatrixInput_4_72};
  wire [2:0]   sigOut_andMatrixOutputs_lo_83 = {sigOut_andMatrixOutputs_lo_hi_33, sigOut_andMatrixOutputs_andMatrixInput_5_33};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_72 = {sigOut_andMatrixOutputs_andMatrixInput_0_87, sigOut_andMatrixOutputs_andMatrixInput_1_87};
  wire [2:0]   sigOut_andMatrixOutputs_hi_84 = {sigOut_andMatrixOutputs_hi_hi_72, sigOut_andMatrixOutputs_andMatrixInput_2_84};
  wire         sigOut_andMatrixOutputs_82_2 = &{sigOut_andMatrixOutputs_hi_84, sigOut_andMatrixOutputs_lo_83};
  wire [1:0]   sigOut_andMatrixOutputs_lo_84 = {sigOut_andMatrixOutputs_andMatrixInput_3_84, sigOut_andMatrixOutputs_andMatrixInput_4_73};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_73 = {sigOut_andMatrixOutputs_andMatrixInput_0_88, sigOut_andMatrixOutputs_andMatrixInput_1_88};
  wire [2:0]   sigOut_andMatrixOutputs_hi_85 = {sigOut_andMatrixOutputs_hi_hi_73, sigOut_andMatrixOutputs_andMatrixInput_2_85};
  wire         sigOut_andMatrixOutputs_14_2 = &{sigOut_andMatrixOutputs_hi_85, sigOut_andMatrixOutputs_lo_84};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_34 = {sigOut_andMatrixOutputs_andMatrixInput_3_85, sigOut_andMatrixOutputs_andMatrixInput_4_74};
  wire [2:0]   sigOut_andMatrixOutputs_lo_85 = {sigOut_andMatrixOutputs_lo_hi_34, sigOut_andMatrixOutputs_andMatrixInput_5_34};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_74 = {sigOut_andMatrixOutputs_andMatrixInput_0_89, sigOut_andMatrixOutputs_andMatrixInput_1_89};
  wire [2:0]   sigOut_andMatrixOutputs_hi_86 = {sigOut_andMatrixOutputs_hi_hi_74, sigOut_andMatrixOutputs_andMatrixInput_2_86};
  wire         sigOut_andMatrixOutputs_23_2 = &{sigOut_andMatrixOutputs_hi_86, sigOut_andMatrixOutputs_lo_85};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_35 = {sigOut_andMatrixOutputs_andMatrixInput_3_86, sigOut_andMatrixOutputs_andMatrixInput_4_75};
  wire [2:0]   sigOut_andMatrixOutputs_lo_86 = {sigOut_andMatrixOutputs_lo_hi_35, sigOut_andMatrixOutputs_andMatrixInput_5_35};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_75 = {sigOut_andMatrixOutputs_andMatrixInput_0_90, sigOut_andMatrixOutputs_andMatrixInput_1_90};
  wire [2:0]   sigOut_andMatrixOutputs_hi_87 = {sigOut_andMatrixOutputs_hi_hi_75, sigOut_andMatrixOutputs_andMatrixInput_2_87};
  wire         sigOut_andMatrixOutputs_74_2 = &{sigOut_andMatrixOutputs_hi_87, sigOut_andMatrixOutputs_lo_86};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_36 = {sigOut_andMatrixOutputs_andMatrixInput_3_87, sigOut_andMatrixOutputs_andMatrixInput_4_76};
  wire [2:0]   sigOut_andMatrixOutputs_lo_87 = {sigOut_andMatrixOutputs_lo_hi_36, sigOut_andMatrixOutputs_andMatrixInput_5_36};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_76 = {sigOut_andMatrixOutputs_andMatrixInput_0_91, sigOut_andMatrixOutputs_andMatrixInput_1_91};
  wire [2:0]   sigOut_andMatrixOutputs_hi_88 = {sigOut_andMatrixOutputs_hi_hi_76, sigOut_andMatrixOutputs_andMatrixInput_2_88};
  wire         sigOut_andMatrixOutputs_9_2 = &{sigOut_andMatrixOutputs_hi_88, sigOut_andMatrixOutputs_lo_87};
  wire [1:0]   sigOut_andMatrixOutputs_lo_hi_37 = {sigOut_andMatrixOutputs_andMatrixInput_3_88, sigOut_andMatrixOutputs_andMatrixInput_4_77};
  wire [2:0]   sigOut_andMatrixOutputs_lo_88 = {sigOut_andMatrixOutputs_lo_hi_37, sigOut_andMatrixOutputs_andMatrixInput_5_37};
  wire [1:0]   sigOut_andMatrixOutputs_hi_hi_77 = {sigOut_andMatrixOutputs_andMatrixInput_0_92, sigOut_andMatrixOutputs_andMatrixInput_1_92};
  wire [2:0]   sigOut_andMatrixOutputs_hi_89 = {sigOut_andMatrixOutputs_hi_hi_77, sigOut_andMatrixOutputs_andMatrixInput_2_89};
  wire         sigOut_andMatrixOutputs_28_2 = &{sigOut_andMatrixOutputs_hi_89, sigOut_andMatrixOutputs_lo_88};
  wire [1:0]   sigOut_orMatrixOutputs_lo_lo_lo_hi = {sigOut_andMatrixOutputs_91_2, sigOut_andMatrixOutputs_79_2};
  wire [2:0]   sigOut_orMatrixOutputs_lo_lo_lo = {sigOut_orMatrixOutputs_lo_lo_lo_hi, sigOut_andMatrixOutputs_14_2};
  wire [1:0]   sigOut_orMatrixOutputs_lo_lo_hi_lo = {sigOut_andMatrixOutputs_31_2, sigOut_andMatrixOutputs_11_2};
  wire [1:0]   sigOut_orMatrixOutputs_lo_lo_hi_hi = {sigOut_andMatrixOutputs_22_2, sigOut_andMatrixOutputs_20_2};
  wire [3:0]   sigOut_orMatrixOutputs_lo_lo_hi = {sigOut_orMatrixOutputs_lo_lo_hi_hi, sigOut_orMatrixOutputs_lo_lo_hi_lo};
  wire [6:0]   sigOut_orMatrixOutputs_lo_lo = {sigOut_orMatrixOutputs_lo_lo_hi, sigOut_orMatrixOutputs_lo_lo_lo};
  wire [1:0]   sigOut_orMatrixOutputs_lo_hi_lo_hi = {sigOut_andMatrixOutputs_76_2, sigOut_andMatrixOutputs_0_2};
  wire [2:0]   sigOut_orMatrixOutputs_lo_hi_lo = {sigOut_orMatrixOutputs_lo_hi_lo_hi, sigOut_andMatrixOutputs_39_2};
  wire [1:0]   sigOut_orMatrixOutputs_lo_hi_hi_lo = {sigOut_andMatrixOutputs_18_2, sigOut_andMatrixOutputs_7_2};
  wire [1:0]   sigOut_orMatrixOutputs_lo_hi_hi_hi = {sigOut_andMatrixOutputs_13_2, sigOut_andMatrixOutputs_41_2};
  wire [3:0]   sigOut_orMatrixOutputs_lo_hi_hi = {sigOut_orMatrixOutputs_lo_hi_hi_hi, sigOut_orMatrixOutputs_lo_hi_hi_lo};
  wire [6:0]   sigOut_orMatrixOutputs_lo_hi = {sigOut_orMatrixOutputs_lo_hi_hi, sigOut_orMatrixOutputs_lo_hi_lo};
  wire [13:0]  sigOut_orMatrixOutputs_lo = {sigOut_orMatrixOutputs_lo_hi, sigOut_orMatrixOutputs_lo_lo};
  wire [1:0]   sigOut_orMatrixOutputs_hi_lo_lo_hi = {sigOut_andMatrixOutputs_29_2, sigOut_andMatrixOutputs_53_2};
  wire [2:0]   sigOut_orMatrixOutputs_hi_lo_lo = {sigOut_orMatrixOutputs_hi_lo_lo_hi, sigOut_andMatrixOutputs_17_2};
  wire [1:0]   sigOut_orMatrixOutputs_hi_lo_hi_lo = {sigOut_andMatrixOutputs_5_2, sigOut_andMatrixOutputs_59_2};
  wire [1:0]   sigOut_orMatrixOutputs_hi_lo_hi_hi = {sigOut_andMatrixOutputs_24_2, sigOut_andMatrixOutputs_30_2};
  wire [3:0]   sigOut_orMatrixOutputs_hi_lo_hi = {sigOut_orMatrixOutputs_hi_lo_hi_hi, sigOut_orMatrixOutputs_hi_lo_hi_lo};
  wire [6:0]   sigOut_orMatrixOutputs_hi_lo = {sigOut_orMatrixOutputs_hi_lo_hi, sigOut_orMatrixOutputs_hi_lo_lo};
  wire [1:0]   sigOut_orMatrixOutputs_hi_hi_lo_hi = {sigOut_andMatrixOutputs_4_2, sigOut_andMatrixOutputs_45_2};
  wire [2:0]   sigOut_orMatrixOutputs_hi_hi_lo = {sigOut_orMatrixOutputs_hi_hi_lo_hi, sigOut_andMatrixOutputs_69_2};
  wire [1:0]   sigOut_orMatrixOutputs_hi_hi_hi_lo = {sigOut_andMatrixOutputs_19_2, sigOut_andMatrixOutputs_68_2};
  wire [1:0]   sigOut_orMatrixOutputs_hi_hi_hi_hi = {sigOut_andMatrixOutputs_90_2, sigOut_andMatrixOutputs_78_2};
  wire [3:0]   sigOut_orMatrixOutputs_hi_hi_hi = {sigOut_orMatrixOutputs_hi_hi_hi_hi, sigOut_orMatrixOutputs_hi_hi_hi_lo};
  wire [6:0]   sigOut_orMatrixOutputs_hi_hi = {sigOut_orMatrixOutputs_hi_hi_hi, sigOut_orMatrixOutputs_hi_hi_lo};
  wire [13:0]  sigOut_orMatrixOutputs_hi = {sigOut_orMatrixOutputs_hi_hi, sigOut_orMatrixOutputs_hi_lo};
  wire [1:0]   sigOut_orMatrixOutputs_lo_lo_lo_lo = {sigOut_andMatrixOutputs_74_2, sigOut_andMatrixOutputs_9_2};
  wire [1:0]   sigOut_orMatrixOutputs_lo_lo_lo_hi_1 = {sigOut_andMatrixOutputs_3_2, sigOut_andMatrixOutputs_54_2};
  wire [3:0]   sigOut_orMatrixOutputs_lo_lo_lo_1 = {sigOut_orMatrixOutputs_lo_lo_lo_hi_1, sigOut_orMatrixOutputs_lo_lo_lo_lo};
  wire [1:0]   _GEN = {sigOut_andMatrixOutputs_87_2, sigOut_andMatrixOutputs_11_2};
  wire [1:0]   sigOut_orMatrixOutputs_lo_lo_hi_lo_1;
  assign sigOut_orMatrixOutputs_lo_lo_hi_lo_1 = _GEN;
  wire [1:0]   sigOut_orMatrixOutputs_lo_lo_hi_hi_2;
  assign sigOut_orMatrixOutputs_lo_lo_hi_hi_2 = _GEN;
  wire [1:0]   sigOut_orMatrixOutputs_lo_lo_hi_hi_1 = {sigOut_andMatrixOutputs_10_2, sigOut_andMatrixOutputs_20_2};
  wire [3:0]   sigOut_orMatrixOutputs_lo_lo_hi_1 = {sigOut_orMatrixOutputs_lo_lo_hi_hi_1, sigOut_orMatrixOutputs_lo_lo_hi_lo_1};
  wire [7:0]   sigOut_orMatrixOutputs_lo_lo_1 = {sigOut_orMatrixOutputs_lo_lo_hi_1, sigOut_orMatrixOutputs_lo_lo_lo_1};
  wire [1:0]   sigOut_orMatrixOutputs_lo_hi_lo_lo = {sigOut_andMatrixOutputs_36_2, sigOut_andMatrixOutputs_64_2};
  wire [1:0]   sigOut_orMatrixOutputs_lo_hi_lo_hi_1 = {sigOut_andMatrixOutputs_42_2, sigOut_andMatrixOutputs_70_2};
  wire [3:0]   sigOut_orMatrixOutputs_lo_hi_lo_1 = {sigOut_orMatrixOutputs_lo_hi_lo_hi_1, sigOut_orMatrixOutputs_lo_hi_lo_lo};
  wire [1:0]   sigOut_orMatrixOutputs_lo_hi_hi_lo_1 = {sigOut_andMatrixOutputs_40_2, sigOut_andMatrixOutputs_71_2};
  wire [1:0]   sigOut_orMatrixOutputs_lo_hi_hi_hi_hi = {sigOut_andMatrixOutputs_13_2, sigOut_andMatrixOutputs_62_2};
  wire [2:0]   sigOut_orMatrixOutputs_lo_hi_hi_hi_1 = {sigOut_orMatrixOutputs_lo_hi_hi_hi_hi, sigOut_andMatrixOutputs_86_2};
  wire [4:0]   sigOut_orMatrixOutputs_lo_hi_hi_1 = {sigOut_orMatrixOutputs_lo_hi_hi_hi_1, sigOut_orMatrixOutputs_lo_hi_hi_lo_1};
  wire [8:0]   sigOut_orMatrixOutputs_lo_hi_1 = {sigOut_orMatrixOutputs_lo_hi_hi_1, sigOut_orMatrixOutputs_lo_hi_lo_1};
  wire [16:0]  sigOut_orMatrixOutputs_lo_1 = {sigOut_orMatrixOutputs_lo_hi_1, sigOut_orMatrixOutputs_lo_lo_1};
  wire [1:0]   sigOut_orMatrixOutputs_hi_lo_lo_lo = {sigOut_andMatrixOutputs_46_2, sigOut_andMatrixOutputs_35_2};
  wire [1:0]   sigOut_orMatrixOutputs_hi_lo_lo_hi_1 = {sigOut_andMatrixOutputs_5_2, sigOut_andMatrixOutputs_51_2};
  wire [3:0]   sigOut_orMatrixOutputs_hi_lo_lo_1 = {sigOut_orMatrixOutputs_hi_lo_lo_hi_1, sigOut_orMatrixOutputs_hi_lo_lo_lo};
  wire [1:0]   sigOut_orMatrixOutputs_hi_lo_hi_lo_1 = {sigOut_andMatrixOutputs_25_2, sigOut_andMatrixOutputs_12_2};
  wire [1:0]   sigOut_orMatrixOutputs_hi_lo_hi_hi_1 = {sigOut_andMatrixOutputs_1_2, sigOut_andMatrixOutputs_44_2};
  wire [3:0]   sigOut_orMatrixOutputs_hi_lo_hi_1 = {sigOut_orMatrixOutputs_hi_lo_hi_hi_1, sigOut_orMatrixOutputs_hi_lo_hi_lo_1};
  wire [7:0]   sigOut_orMatrixOutputs_hi_lo_1 = {sigOut_orMatrixOutputs_hi_lo_hi_1, sigOut_orMatrixOutputs_hi_lo_lo_1};
  wire [1:0]   sigOut_orMatrixOutputs_hi_hi_lo_lo = {sigOut_andMatrixOutputs_47_2, sigOut_andMatrixOutputs_45_2};
  wire [1:0]   sigOut_orMatrixOutputs_hi_hi_lo_hi_1 = {sigOut_andMatrixOutputs_80_2, sigOut_andMatrixOutputs_4_2};
  wire [3:0]   sigOut_orMatrixOutputs_hi_hi_lo_1 = {sigOut_orMatrixOutputs_hi_hi_lo_hi_1, sigOut_orMatrixOutputs_hi_hi_lo_lo};
  wire [1:0]   sigOut_orMatrixOutputs_hi_hi_hi_lo_1 = {sigOut_andMatrixOutputs_34_2, sigOut_andMatrixOutputs_19_2};
  wire [1:0]   sigOut_orMatrixOutputs_hi_hi_hi_hi_hi = {sigOut_andMatrixOutputs_90_2, sigOut_andMatrixOutputs_2_2};
  wire [2:0]   sigOut_orMatrixOutputs_hi_hi_hi_hi_1 = {sigOut_orMatrixOutputs_hi_hi_hi_hi_hi, sigOut_andMatrixOutputs_8_2};
  wire [4:0]   sigOut_orMatrixOutputs_hi_hi_hi_1 = {sigOut_orMatrixOutputs_hi_hi_hi_hi_1, sigOut_orMatrixOutputs_hi_hi_hi_lo_1};
  wire [8:0]   sigOut_orMatrixOutputs_hi_hi_1 = {sigOut_orMatrixOutputs_hi_hi_hi_1, sigOut_orMatrixOutputs_hi_hi_lo_1};
  wire [16:0]  sigOut_orMatrixOutputs_hi_1 = {sigOut_orMatrixOutputs_hi_hi_1, sigOut_orMatrixOutputs_hi_lo_1};
  wire [1:0]   sigOut_orMatrixOutputs_lo_lo_lo_hi_2 = {sigOut_andMatrixOutputs_21_2, sigOut_andMatrixOutputs_23_2};
  wire [2:0]   sigOut_orMatrixOutputs_lo_lo_lo_2 = {sigOut_orMatrixOutputs_lo_lo_lo_hi_2, sigOut_andMatrixOutputs_28_2};
  wire [2:0]   sigOut_orMatrixOutputs_lo_lo_hi_2 = {sigOut_orMatrixOutputs_lo_lo_hi_hi_2, sigOut_andMatrixOutputs_89_2};
  wire [5:0]   sigOut_orMatrixOutputs_lo_lo_2 = {sigOut_orMatrixOutputs_lo_lo_hi_2, sigOut_orMatrixOutputs_lo_lo_lo_2};
  wire [1:0]   sigOut_orMatrixOutputs_lo_hi_lo_hi_2 = {sigOut_andMatrixOutputs_67_2, sigOut_andMatrixOutputs_31_2};
  wire [2:0]   sigOut_orMatrixOutputs_lo_hi_lo_2 = {sigOut_orMatrixOutputs_lo_hi_lo_hi_2, sigOut_andMatrixOutputs_61_2};
  wire [1:0]   sigOut_orMatrixOutputs_lo_hi_hi_hi_2 = {sigOut_andMatrixOutputs_85_2, sigOut_andMatrixOutputs_26_2};
  wire [2:0]   sigOut_orMatrixOutputs_lo_hi_hi_2 = {sigOut_orMatrixOutputs_lo_hi_hi_hi_2, sigOut_andMatrixOutputs_36_2};
  wire [5:0]   sigOut_orMatrixOutputs_lo_hi_2 = {sigOut_orMatrixOutputs_lo_hi_hi_2, sigOut_orMatrixOutputs_lo_hi_lo_2};
  wire [11:0]  sigOut_orMatrixOutputs_lo_2 = {sigOut_orMatrixOutputs_lo_hi_2, sigOut_orMatrixOutputs_lo_lo_2};
  wire [1:0]   sigOut_orMatrixOutputs_hi_lo_lo_hi_2 = {sigOut_andMatrixOutputs_75_2, sigOut_andMatrixOutputs_86_2};
  wire [2:0]   sigOut_orMatrixOutputs_hi_lo_lo_2 = {sigOut_orMatrixOutputs_hi_lo_lo_hi_2, sigOut_andMatrixOutputs_37_2};
  wire [1:0]   sigOut_orMatrixOutputs_hi_lo_hi_hi_2 = {sigOut_andMatrixOutputs_73_2, sigOut_andMatrixOutputs_81_2};
  wire [2:0]   sigOut_orMatrixOutputs_hi_lo_hi_2 = {sigOut_orMatrixOutputs_hi_lo_hi_hi_2, sigOut_andMatrixOutputs_38_2};
  wire [5:0]   sigOut_orMatrixOutputs_hi_lo_2 = {sigOut_orMatrixOutputs_hi_lo_hi_2, sigOut_orMatrixOutputs_hi_lo_lo_2};
  wire [1:0]   sigOut_orMatrixOutputs_hi_hi_lo_hi_2 = {sigOut_andMatrixOutputs_1_2, sigOut_andMatrixOutputs_65_2};
  wire [2:0]   sigOut_orMatrixOutputs_hi_hi_lo_2 = {sigOut_orMatrixOutputs_hi_hi_lo_hi_2, sigOut_andMatrixOutputs_46_2};
  wire [1:0]   sigOut_orMatrixOutputs_hi_hi_hi_lo_2 = {sigOut_andMatrixOutputs_60_2, sigOut_andMatrixOutputs_4_2};
  wire [1:0]   sigOut_orMatrixOutputs_hi_hi_hi_hi_2 = {sigOut_andMatrixOutputs_63_2, sigOut_andMatrixOutputs_16_2};
  wire [3:0]   sigOut_orMatrixOutputs_hi_hi_hi_2 = {sigOut_orMatrixOutputs_hi_hi_hi_hi_2, sigOut_orMatrixOutputs_hi_hi_hi_lo_2};
  wire [6:0]   sigOut_orMatrixOutputs_hi_hi_2 = {sigOut_orMatrixOutputs_hi_hi_hi_2, sigOut_orMatrixOutputs_hi_hi_lo_2};
  wire [12:0]  sigOut_orMatrixOutputs_hi_2 = {sigOut_orMatrixOutputs_hi_hi_2, sigOut_orMatrixOutputs_hi_lo_2};
  wire [1:0]   sigOut_orMatrixOutputs_lo_lo_lo_3 = {sigOut_andMatrixOutputs_82_2, sigOut_andMatrixOutputs_74_2};
  wire [1:0]   sigOut_orMatrixOutputs_lo_lo_hi_hi_3 = {sigOut_andMatrixOutputs_58_2, sigOut_andMatrixOutputs_43_2};
  wire [2:0]   sigOut_orMatrixOutputs_lo_lo_hi_3 = {sigOut_orMatrixOutputs_lo_lo_hi_hi_3, sigOut_andMatrixOutputs_6_2};
  wire [4:0]   sigOut_orMatrixOutputs_lo_lo_3 = {sigOut_orMatrixOutputs_lo_lo_hi_3, sigOut_orMatrixOutputs_lo_lo_lo_3};
  wire [1:0]   sigOut_orMatrixOutputs_lo_hi_lo_3 = {sigOut_andMatrixOutputs_91_2, sigOut_andMatrixOutputs_89_2};
  wire [1:0]   sigOut_orMatrixOutputs_lo_hi_hi_hi_3 = {sigOut_andMatrixOutputs_52_2, sigOut_andMatrixOutputs_39_2};
  wire [2:0]   sigOut_orMatrixOutputs_lo_hi_hi_3 = {sigOut_orMatrixOutputs_lo_hi_hi_hi_3, sigOut_andMatrixOutputs_64_2};
  wire [4:0]   sigOut_orMatrixOutputs_lo_hi_3 = {sigOut_orMatrixOutputs_lo_hi_hi_3, sigOut_orMatrixOutputs_lo_hi_lo_3};
  wire [9:0]   sigOut_orMatrixOutputs_lo_3 = {sigOut_orMatrixOutputs_lo_hi_3, sigOut_orMatrixOutputs_lo_lo_3};
  wire [1:0]   sigOut_orMatrixOutputs_hi_lo_lo_3 = {sigOut_andMatrixOutputs_56_2, sigOut_andMatrixOutputs_76_2};
  wire [1:0]   sigOut_orMatrixOutputs_hi_lo_hi_hi_3 = {sigOut_andMatrixOutputs_25_2, sigOut_andMatrixOutputs_46_2};
  wire [2:0]   sigOut_orMatrixOutputs_hi_lo_hi_3 = {sigOut_orMatrixOutputs_hi_lo_hi_hi_3, sigOut_andMatrixOutputs_48_2};
  wire [4:0]   sigOut_orMatrixOutputs_hi_lo_3 = {sigOut_orMatrixOutputs_hi_lo_hi_3, sigOut_orMatrixOutputs_hi_lo_lo_3};
  wire [1:0]   _GEN_0 = {sigOut_andMatrixOutputs_1_2, sigOut_andMatrixOutputs_50_2};
  wire [1:0]   sigOut_orMatrixOutputs_hi_hi_lo_3;
  assign sigOut_orMatrixOutputs_hi_hi_lo_3 = _GEN_0;
  wire [1:0]   sigOut_orMatrixOutputs_hi_hi_lo_4;
  assign sigOut_orMatrixOutputs_hi_hi_lo_4 = _GEN_0;
  wire [1:0]   sigOut_orMatrixOutputs_hi_hi_hi_hi_3 = {sigOut_andMatrixOutputs_49_2, sigOut_andMatrixOutputs_33_2};
  wire [2:0]   sigOut_orMatrixOutputs_hi_hi_hi_3 = {sigOut_orMatrixOutputs_hi_hi_hi_hi_3, sigOut_andMatrixOutputs_77_2};
  wire [4:0]   sigOut_orMatrixOutputs_hi_hi_3 = {sigOut_orMatrixOutputs_hi_hi_hi_3, sigOut_orMatrixOutputs_hi_hi_lo_3};
  wire [9:0]   sigOut_orMatrixOutputs_hi_3 = {sigOut_orMatrixOutputs_hi_hi_3, sigOut_orMatrixOutputs_hi_lo_3};
  wire [1:0]   sigOut_orMatrixOutputs_lo_lo_hi_4 = {sigOut_andMatrixOutputs_14_2, sigOut_andMatrixOutputs_23_2};
  wire [2:0]   sigOut_orMatrixOutputs_lo_lo_4 = {sigOut_orMatrixOutputs_lo_lo_hi_4, sigOut_andMatrixOutputs_74_2};
  wire [1:0]   sigOut_orMatrixOutputs_lo_hi_hi_4 = {sigOut_andMatrixOutputs_84_2, sigOut_andMatrixOutputs_6_2};
  wire [2:0]   sigOut_orMatrixOutputs_lo_hi_4 = {sigOut_orMatrixOutputs_lo_hi_hi_4, sigOut_andMatrixOutputs_82_2};
  wire [5:0]   sigOut_orMatrixOutputs_lo_4 = {sigOut_orMatrixOutputs_lo_hi_4, sigOut_orMatrixOutputs_lo_lo_4};
  wire [1:0]   sigOut_orMatrixOutputs_hi_lo_hi_4 = {sigOut_andMatrixOutputs_88_2, sigOut_andMatrixOutputs_15_2};
  wire [2:0]   sigOut_orMatrixOutputs_hi_lo_4 = {sigOut_orMatrixOutputs_hi_lo_hi_4, sigOut_andMatrixOutputs_7_2};
  wire [1:0]   sigOut_orMatrixOutputs_hi_hi_hi_4 = {sigOut_andMatrixOutputs_27_2, sigOut_andMatrixOutputs_83_2};
  wire [3:0]   sigOut_orMatrixOutputs_hi_hi_4 = {sigOut_orMatrixOutputs_hi_hi_hi_4, sigOut_orMatrixOutputs_hi_hi_lo_4};
  wire [6:0]   sigOut_orMatrixOutputs_hi_4 = {sigOut_orMatrixOutputs_hi_hi_4, sigOut_orMatrixOutputs_hi_lo_4};
  wire [1:0]   sigOut_orMatrixOutputs_lo_lo_5 = {sigOut_andMatrixOutputs_23_2, sigOut_andMatrixOutputs_74_2};
  wire [1:0]   sigOut_orMatrixOutputs_lo_hi_5 = {sigOut_andMatrixOutputs_82_2, sigOut_andMatrixOutputs_14_2};
  wire [3:0]   sigOut_orMatrixOutputs_lo_5 = {sigOut_orMatrixOutputs_lo_hi_5, sigOut_orMatrixOutputs_lo_lo_5};
  wire [1:0]   sigOut_orMatrixOutputs_hi_lo_5 = {sigOut_andMatrixOutputs_32_2, sigOut_andMatrixOutputs_6_2};
  wire [1:0]   sigOut_orMatrixOutputs_hi_hi_5 = {sigOut_andMatrixOutputs_57_2, sigOut_andMatrixOutputs_92_2};
  wire [3:0]   sigOut_orMatrixOutputs_hi_5 = {sigOut_orMatrixOutputs_hi_hi_5, sigOut_orMatrixOutputs_hi_lo_5};
  wire [1:0]   sigOut_orMatrixOutputs_hi_6 = {sigOut_andMatrixOutputs_66_2, sigOut_andMatrixOutputs_72_2};
  wire [1:0]   sigOut_orMatrixOutputs_lo_hi_6 = {|{sigOut_orMatrixOutputs_hi_2, sigOut_orMatrixOutputs_lo_2}, |{sigOut_orMatrixOutputs_hi_1, sigOut_orMatrixOutputs_lo_1}};
  wire [2:0]   sigOut_orMatrixOutputs_lo_6 = {sigOut_orMatrixOutputs_lo_hi_6, |{sigOut_orMatrixOutputs_hi, sigOut_orMatrixOutputs_lo}};
  wire [1:0]   sigOut_orMatrixOutputs_hi_lo_6 = {|{sigOut_orMatrixOutputs_hi_4, sigOut_orMatrixOutputs_lo_4}, |{sigOut_orMatrixOutputs_hi_3, sigOut_orMatrixOutputs_lo_3}};
  wire [1:0]   sigOut_orMatrixOutputs_hi_hi_6 = {|{sigOut_orMatrixOutputs_hi_6, sigOut_andMatrixOutputs_55_2}, |{sigOut_orMatrixOutputs_hi_5, sigOut_orMatrixOutputs_lo_5}};
  wire [3:0]   sigOut_orMatrixOutputs_hi_7 = {sigOut_orMatrixOutputs_hi_hi_6, sigOut_orMatrixOutputs_hi_lo_6};
  wire [6:0]   sigOut_orMatrixOutputs = {sigOut_orMatrixOutputs_hi_7, sigOut_orMatrixOutputs_lo_6};
  wire [1:0]   sigOut_invMatrixOutputs_lo_hi = sigOut_orMatrixOutputs[2:1];
  wire [2:0]   sigOut_invMatrixOutputs_lo = {sigOut_invMatrixOutputs_lo_hi, sigOut_orMatrixOutputs[0]};
  wire [1:0]   sigOut_invMatrixOutputs_hi_lo = sigOut_orMatrixOutputs[4:3];
  wire [1:0]   sigOut_invMatrixOutputs_hi_hi = sigOut_orMatrixOutputs[6:5];
  wire [3:0]   sigOut_invMatrixOutputs_hi = {sigOut_invMatrixOutputs_hi_hi, sigOut_invMatrixOutputs_hi_lo};
  assign sigOut_invMatrixOutputs = {sigOut_invMatrixOutputs_hi, sigOut_invMatrixOutputs_lo};
  wire [6:0]   sigOut_plaOutput = sigOut_invMatrixOutputs;
  wire [22:0]  sigOut = {sigOut_plaOutput, 16'h0};
  wire [8:0]   _expOut_T = {1'h0, normDist} - 9'h84;
  wire [8:0]   _expOut_T_2 = 9'h17C - {1'h0, expIn};
  wire [7:0]   expOut = inIsSub ? _expOut_T[8:1] : _expOut_T_2[8:1];
  wire [8:0]   view__out_data_hi = {sign, expOut};
  assign out_data = outNaN ? 32'h7FC00000 : outInf ? {sign, 31'h7F800000} : {view__out_data_hi, sigOut};
  assign out_exceptionFlags = outNaN ? 5'h10 : {1'h0, outInf, 3'h0};
endmodule

