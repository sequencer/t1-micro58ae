
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module SimpleAccessUnit(
  input          clock,
                 reset,
                 lsuRequest_valid,
  input  [2:0]   lsuRequest_bits_instructionInformation_nf,
  input          lsuRequest_bits_instructionInformation_mew,
  input  [1:0]   lsuRequest_bits_instructionInformation_mop,
  input  [4:0]   lsuRequest_bits_instructionInformation_lumop,
  input  [1:0]   lsuRequest_bits_instructionInformation_eew,
  input  [4:0]   lsuRequest_bits_instructionInformation_vs3,
  input          lsuRequest_bits_instructionInformation_isStore,
                 lsuRequest_bits_instructionInformation_maskedLoadStore,
  input  [31:0]  lsuRequest_bits_rs1Data,
                 lsuRequest_bits_rs2Data,
  input  [2:0]   lsuRequest_bits_instructionIndex,
  input          vrfReadDataPorts_ready,
  output         vrfReadDataPorts_valid,
  output [4:0]   vrfReadDataPorts_bits_vs,
  output         vrfReadDataPorts_bits_offset,
  output [2:0]   vrfReadDataPorts_bits_instructionIndex,
  input          vrfReadResults_valid,
  input  [31:0]  vrfReadResults_bits,
  input          offsetReadResult_0_valid,
  input  [31:0]  offsetReadResult_0_bits,
  input          offsetReadResult_1_valid,
  input  [31:0]  offsetReadResult_1_bits,
  input          offsetReadResult_2_valid,
  input  [31:0]  offsetReadResult_2_bits,
  input          offsetReadResult_3_valid,
  input  [31:0]  offsetReadResult_3_bits,
  input          offsetReadResult_4_valid,
  input  [31:0]  offsetReadResult_4_bits,
  input          offsetReadResult_5_valid,
  input  [31:0]  offsetReadResult_5_bits,
  input          offsetReadResult_6_valid,
  input  [31:0]  offsetReadResult_6_bits,
  input          offsetReadResult_7_valid,
  input  [31:0]  offsetReadResult_7_bits,
  input          offsetReadResult_8_valid,
  input  [31:0]  offsetReadResult_8_bits,
  input          offsetReadResult_9_valid,
  input  [31:0]  offsetReadResult_9_bits,
  input          offsetReadResult_10_valid,
  input  [31:0]  offsetReadResult_10_bits,
  input          offsetReadResult_11_valid,
  input  [31:0]  offsetReadResult_11_bits,
  input          offsetReadResult_12_valid,
  input  [31:0]  offsetReadResult_12_bits,
  input          offsetReadResult_13_valid,
  input  [31:0]  offsetReadResult_13_bits,
  input          offsetReadResult_14_valid,
  input  [31:0]  offsetReadResult_14_bits,
  input          offsetReadResult_15_valid,
  input  [31:0]  offsetReadResult_15_bits,
  input          offsetReadResult_16_valid,
  input  [31:0]  offsetReadResult_16_bits,
  input          offsetReadResult_17_valid,
  input  [31:0]  offsetReadResult_17_bits,
  input          offsetReadResult_18_valid,
  input  [31:0]  offsetReadResult_18_bits,
  input          offsetReadResult_19_valid,
  input  [31:0]  offsetReadResult_19_bits,
  input          offsetReadResult_20_valid,
  input  [31:0]  offsetReadResult_20_bits,
  input          offsetReadResult_21_valid,
  input  [31:0]  offsetReadResult_21_bits,
  input          offsetReadResult_22_valid,
  input  [31:0]  offsetReadResult_22_bits,
  input          offsetReadResult_23_valid,
  input  [31:0]  offsetReadResult_23_bits,
  input          offsetReadResult_24_valid,
  input  [31:0]  offsetReadResult_24_bits,
  input          offsetReadResult_25_valid,
  input  [31:0]  offsetReadResult_25_bits,
  input          offsetReadResult_26_valid,
  input  [31:0]  offsetReadResult_26_bits,
  input          offsetReadResult_27_valid,
  input  [31:0]  offsetReadResult_27_bits,
  input          offsetReadResult_28_valid,
  input  [31:0]  offsetReadResult_28_bits,
  input          offsetReadResult_29_valid,
  input  [31:0]  offsetReadResult_29_bits,
  input          offsetReadResult_30_valid,
  input  [31:0]  offsetReadResult_30_bits,
  input          offsetReadResult_31_valid,
  input  [31:0]  offsetReadResult_31_bits,
  input  [127:0] maskInput,
  output         maskSelect_valid,
  output [3:0]   maskSelect_bits,
  input          memReadRequest_ready,
  output         memReadRequest_valid,
  output [31:0]  memReadRequest_bits_address,
  output [9:0]   memReadRequest_bits_source,
  output         memReadResponse_ready,
  input          memReadResponse_valid,
  input  [31:0]  memReadResponse_bits_data,
  input  [9:0]   memReadResponse_bits_source,
  input          memWriteRequest_ready,
  output         memWriteRequest_valid,
  output [31:0]  memWriteRequest_bits_data,
  output [3:0]   memWriteRequest_bits_mask,
  output [7:0]   memWriteRequest_bits_source,
  output [31:0]  memWriteRequest_bits_address,
  output [1:0]   memWriteRequest_bits_size,
  input          vrfWritePort_ready,
  output         vrfWritePort_valid,
  output [4:0]   vrfWritePort_bits_vd,
  output         vrfWritePort_bits_offset,
  output [3:0]   vrfWritePort_bits_mask,
  output [31:0]  vrfWritePort_bits_data,
  output         vrfWritePort_bits_last,
  output [2:0]   vrfWritePort_bits_instructionIndex,
  input  [11:0]  csrInterface_vl,
                 csrInterface_vStart,
  input  [2:0]   csrInterface_vlmul,
  input  [1:0]   csrInterface_vSew,
                 csrInterface_vxrm,
  input          csrInterface_vta,
                 csrInterface_vma,
  output         status_idle,
                 status_last,
  output [2:0]   status_instructionIndex,
  output [31:0]  status_targetLane,
  output         status_isStore,
                 offsetRelease_0,
                 offsetRelease_1,
                 offsetRelease_2,
                 offsetRelease_3,
                 offsetRelease_4,
                 offsetRelease_5,
                 offsetRelease_6,
                 offsetRelease_7,
                 offsetRelease_8,
                 offsetRelease_9,
                 offsetRelease_10,
                 offsetRelease_11,
                 offsetRelease_12,
                 offsetRelease_13,
                 offsetRelease_14,
                 offsetRelease_15,
                 offsetRelease_16,
                 offsetRelease_17,
                 offsetRelease_18,
                 offsetRelease_19,
                 offsetRelease_20,
                 offsetRelease_21,
                 offsetRelease_22,
                 offsetRelease_23,
                 offsetRelease_24,
                 offsetRelease_25,
                 offsetRelease_26,
                 offsetRelease_27,
                 offsetRelease_28,
                 offsetRelease_29,
                 offsetRelease_30,
                 offsetRelease_31
);

  wire              _s1EnqDataQueue_fifo_empty;
  wire              _s1EnqDataQueue_fifo_full;
  wire              _s1EnqDataQueue_fifo_error;
  wire              _s1EnqQueue_fifo_empty;
  wire              _s1EnqQueue_fifo_full;
  wire              _s1EnqQueue_fifo_error;
  wire [73:0]       _s1EnqQueue_fifo_data_out;
  wire              _offsetQueueVec_queue_fifo_31_empty;
  wire              _offsetQueueVec_queue_fifo_31_full;
  wire              _offsetQueueVec_queue_fifo_31_error;
  wire              _offsetQueueVec_queue_fifo_30_empty;
  wire              _offsetQueueVec_queue_fifo_30_full;
  wire              _offsetQueueVec_queue_fifo_30_error;
  wire              _offsetQueueVec_queue_fifo_29_empty;
  wire              _offsetQueueVec_queue_fifo_29_full;
  wire              _offsetQueueVec_queue_fifo_29_error;
  wire              _offsetQueueVec_queue_fifo_28_empty;
  wire              _offsetQueueVec_queue_fifo_28_full;
  wire              _offsetQueueVec_queue_fifo_28_error;
  wire              _offsetQueueVec_queue_fifo_27_empty;
  wire              _offsetQueueVec_queue_fifo_27_full;
  wire              _offsetQueueVec_queue_fifo_27_error;
  wire              _offsetQueueVec_queue_fifo_26_empty;
  wire              _offsetQueueVec_queue_fifo_26_full;
  wire              _offsetQueueVec_queue_fifo_26_error;
  wire              _offsetQueueVec_queue_fifo_25_empty;
  wire              _offsetQueueVec_queue_fifo_25_full;
  wire              _offsetQueueVec_queue_fifo_25_error;
  wire              _offsetQueueVec_queue_fifo_24_empty;
  wire              _offsetQueueVec_queue_fifo_24_full;
  wire              _offsetQueueVec_queue_fifo_24_error;
  wire              _offsetQueueVec_queue_fifo_23_empty;
  wire              _offsetQueueVec_queue_fifo_23_full;
  wire              _offsetQueueVec_queue_fifo_23_error;
  wire              _offsetQueueVec_queue_fifo_22_empty;
  wire              _offsetQueueVec_queue_fifo_22_full;
  wire              _offsetQueueVec_queue_fifo_22_error;
  wire              _offsetQueueVec_queue_fifo_21_empty;
  wire              _offsetQueueVec_queue_fifo_21_full;
  wire              _offsetQueueVec_queue_fifo_21_error;
  wire              _offsetQueueVec_queue_fifo_20_empty;
  wire              _offsetQueueVec_queue_fifo_20_full;
  wire              _offsetQueueVec_queue_fifo_20_error;
  wire              _offsetQueueVec_queue_fifo_19_empty;
  wire              _offsetQueueVec_queue_fifo_19_full;
  wire              _offsetQueueVec_queue_fifo_19_error;
  wire              _offsetQueueVec_queue_fifo_18_empty;
  wire              _offsetQueueVec_queue_fifo_18_full;
  wire              _offsetQueueVec_queue_fifo_18_error;
  wire              _offsetQueueVec_queue_fifo_17_empty;
  wire              _offsetQueueVec_queue_fifo_17_full;
  wire              _offsetQueueVec_queue_fifo_17_error;
  wire              _offsetQueueVec_queue_fifo_16_empty;
  wire              _offsetQueueVec_queue_fifo_16_full;
  wire              _offsetQueueVec_queue_fifo_16_error;
  wire              _offsetQueueVec_queue_fifo_15_empty;
  wire              _offsetQueueVec_queue_fifo_15_full;
  wire              _offsetQueueVec_queue_fifo_15_error;
  wire              _offsetQueueVec_queue_fifo_14_empty;
  wire              _offsetQueueVec_queue_fifo_14_full;
  wire              _offsetQueueVec_queue_fifo_14_error;
  wire              _offsetQueueVec_queue_fifo_13_empty;
  wire              _offsetQueueVec_queue_fifo_13_full;
  wire              _offsetQueueVec_queue_fifo_13_error;
  wire              _offsetQueueVec_queue_fifo_12_empty;
  wire              _offsetQueueVec_queue_fifo_12_full;
  wire              _offsetQueueVec_queue_fifo_12_error;
  wire              _offsetQueueVec_queue_fifo_11_empty;
  wire              _offsetQueueVec_queue_fifo_11_full;
  wire              _offsetQueueVec_queue_fifo_11_error;
  wire              _offsetQueueVec_queue_fifo_10_empty;
  wire              _offsetQueueVec_queue_fifo_10_full;
  wire              _offsetQueueVec_queue_fifo_10_error;
  wire              _offsetQueueVec_queue_fifo_9_empty;
  wire              _offsetQueueVec_queue_fifo_9_full;
  wire              _offsetQueueVec_queue_fifo_9_error;
  wire              _offsetQueueVec_queue_fifo_8_empty;
  wire              _offsetQueueVec_queue_fifo_8_full;
  wire              _offsetQueueVec_queue_fifo_8_error;
  wire              _offsetQueueVec_queue_fifo_7_empty;
  wire              _offsetQueueVec_queue_fifo_7_full;
  wire              _offsetQueueVec_queue_fifo_7_error;
  wire              _offsetQueueVec_queue_fifo_6_empty;
  wire              _offsetQueueVec_queue_fifo_6_full;
  wire              _offsetQueueVec_queue_fifo_6_error;
  wire              _offsetQueueVec_queue_fifo_5_empty;
  wire              _offsetQueueVec_queue_fifo_5_full;
  wire              _offsetQueueVec_queue_fifo_5_error;
  wire              _offsetQueueVec_queue_fifo_4_empty;
  wire              _offsetQueueVec_queue_fifo_4_full;
  wire              _offsetQueueVec_queue_fifo_4_error;
  wire              _offsetQueueVec_queue_fifo_3_empty;
  wire              _offsetQueueVec_queue_fifo_3_full;
  wire              _offsetQueueVec_queue_fifo_3_error;
  wire              _offsetQueueVec_queue_fifo_2_empty;
  wire              _offsetQueueVec_queue_fifo_2_full;
  wire              _offsetQueueVec_queue_fifo_2_error;
  wire              _offsetQueueVec_queue_fifo_1_empty;
  wire              _offsetQueueVec_queue_fifo_1_full;
  wire              _offsetQueueVec_queue_fifo_1_error;
  wire              _offsetQueueVec_queue_fifo_empty;
  wire              _offsetQueueVec_queue_fifo_full;
  wire              _offsetQueueVec_queue_fifo_error;
  wire              s1EnqDataQueue_almostFull;
  wire              s1EnqDataQueue_almostEmpty;
  wire              s1EnqQueue_almostFull;
  wire              s1EnqQueue_almostEmpty;
  wire              offsetQueueVec_31_almostFull;
  wire              offsetQueueVec_31_almostEmpty;
  wire              offsetQueueVec_30_almostFull;
  wire              offsetQueueVec_30_almostEmpty;
  wire              offsetQueueVec_29_almostFull;
  wire              offsetQueueVec_29_almostEmpty;
  wire              offsetQueueVec_28_almostFull;
  wire              offsetQueueVec_28_almostEmpty;
  wire              offsetQueueVec_27_almostFull;
  wire              offsetQueueVec_27_almostEmpty;
  wire              offsetQueueVec_26_almostFull;
  wire              offsetQueueVec_26_almostEmpty;
  wire              offsetQueueVec_25_almostFull;
  wire              offsetQueueVec_25_almostEmpty;
  wire              offsetQueueVec_24_almostFull;
  wire              offsetQueueVec_24_almostEmpty;
  wire              offsetQueueVec_23_almostFull;
  wire              offsetQueueVec_23_almostEmpty;
  wire              offsetQueueVec_22_almostFull;
  wire              offsetQueueVec_22_almostEmpty;
  wire              offsetQueueVec_21_almostFull;
  wire              offsetQueueVec_21_almostEmpty;
  wire              offsetQueueVec_20_almostFull;
  wire              offsetQueueVec_20_almostEmpty;
  wire              offsetQueueVec_19_almostFull;
  wire              offsetQueueVec_19_almostEmpty;
  wire              offsetQueueVec_18_almostFull;
  wire              offsetQueueVec_18_almostEmpty;
  wire              offsetQueueVec_17_almostFull;
  wire              offsetQueueVec_17_almostEmpty;
  wire              offsetQueueVec_16_almostFull;
  wire              offsetQueueVec_16_almostEmpty;
  wire              offsetQueueVec_15_almostFull;
  wire              offsetQueueVec_15_almostEmpty;
  wire              offsetQueueVec_14_almostFull;
  wire              offsetQueueVec_14_almostEmpty;
  wire              offsetQueueVec_13_almostFull;
  wire              offsetQueueVec_13_almostEmpty;
  wire              offsetQueueVec_12_almostFull;
  wire              offsetQueueVec_12_almostEmpty;
  wire              offsetQueueVec_11_almostFull;
  wire              offsetQueueVec_11_almostEmpty;
  wire              offsetQueueVec_10_almostFull;
  wire              offsetQueueVec_10_almostEmpty;
  wire              offsetQueueVec_9_almostFull;
  wire              offsetQueueVec_9_almostEmpty;
  wire              offsetQueueVec_8_almostFull;
  wire              offsetQueueVec_8_almostEmpty;
  wire              offsetQueueVec_7_almostFull;
  wire              offsetQueueVec_7_almostEmpty;
  wire              offsetQueueVec_6_almostFull;
  wire              offsetQueueVec_6_almostEmpty;
  wire              offsetQueueVec_5_almostFull;
  wire              offsetQueueVec_5_almostEmpty;
  wire              offsetQueueVec_4_almostFull;
  wire              offsetQueueVec_4_almostEmpty;
  wire              offsetQueueVec_3_almostFull;
  wire              offsetQueueVec_3_almostEmpty;
  wire              offsetQueueVec_2_almostFull;
  wire              offsetQueueVec_2_almostEmpty;
  wire              offsetQueueVec_1_almostFull;
  wire              offsetQueueVec_1_almostEmpty;
  wire              offsetQueueVec_0_almostFull;
  wire              offsetQueueVec_0_almostEmpty;
  wire [31:0]       s1EnqDataQueue_deq_bits;
  wire              s1EnqueueReady;
  wire [31:0]       s1EnqQueue_deq_bits_address;
  wire [2:0]        s1EnqQueue_deq_bits_segmentIndex;
  wire [6:0]        s1EnqQueue_deq_bits_indexInMaskGroup;
  wire              vrfReadDataPorts_ready_0 = vrfReadDataPorts_ready;
  wire              memReadRequest_ready_0 = memReadRequest_ready;
  wire              memReadResponse_valid_0 = memReadResponse_valid;
  wire [31:0]       memReadResponse_bits_data_0 = memReadResponse_bits_data;
  wire [9:0]        memReadResponse_bits_source_0 = memReadResponse_bits_source;
  wire              memWriteRequest_ready_0 = memWriteRequest_ready;
  wire              vrfWritePort_ready_0 = vrfWritePort_ready;
  wire              offsetQueueVec_0_enq_valid = offsetReadResult_0_valid;
  wire [31:0]       offsetQueueVec_0_enq_bits = offsetReadResult_0_bits;
  wire              offsetQueueVec_1_enq_valid = offsetReadResult_1_valid;
  wire [31:0]       offsetQueueVec_1_enq_bits = offsetReadResult_1_bits;
  wire              offsetQueueVec_2_enq_valid = offsetReadResult_2_valid;
  wire [31:0]       offsetQueueVec_2_enq_bits = offsetReadResult_2_bits;
  wire              offsetQueueVec_3_enq_valid = offsetReadResult_3_valid;
  wire [31:0]       offsetQueueVec_3_enq_bits = offsetReadResult_3_bits;
  wire              offsetQueueVec_4_enq_valid = offsetReadResult_4_valid;
  wire [31:0]       offsetQueueVec_4_enq_bits = offsetReadResult_4_bits;
  wire              offsetQueueVec_5_enq_valid = offsetReadResult_5_valid;
  wire [31:0]       offsetQueueVec_5_enq_bits = offsetReadResult_5_bits;
  wire              offsetQueueVec_6_enq_valid = offsetReadResult_6_valid;
  wire [31:0]       offsetQueueVec_6_enq_bits = offsetReadResult_6_bits;
  wire              offsetQueueVec_7_enq_valid = offsetReadResult_7_valid;
  wire [31:0]       offsetQueueVec_7_enq_bits = offsetReadResult_7_bits;
  wire              offsetQueueVec_8_enq_valid = offsetReadResult_8_valid;
  wire [31:0]       offsetQueueVec_8_enq_bits = offsetReadResult_8_bits;
  wire              offsetQueueVec_9_enq_valid = offsetReadResult_9_valid;
  wire [31:0]       offsetQueueVec_9_enq_bits = offsetReadResult_9_bits;
  wire              offsetQueueVec_10_enq_valid = offsetReadResult_10_valid;
  wire [31:0]       offsetQueueVec_10_enq_bits = offsetReadResult_10_bits;
  wire              offsetQueueVec_11_enq_valid = offsetReadResult_11_valid;
  wire [31:0]       offsetQueueVec_11_enq_bits = offsetReadResult_11_bits;
  wire              offsetQueueVec_12_enq_valid = offsetReadResult_12_valid;
  wire [31:0]       offsetQueueVec_12_enq_bits = offsetReadResult_12_bits;
  wire              offsetQueueVec_13_enq_valid = offsetReadResult_13_valid;
  wire [31:0]       offsetQueueVec_13_enq_bits = offsetReadResult_13_bits;
  wire              offsetQueueVec_14_enq_valid = offsetReadResult_14_valid;
  wire [31:0]       offsetQueueVec_14_enq_bits = offsetReadResult_14_bits;
  wire              offsetQueueVec_15_enq_valid = offsetReadResult_15_valid;
  wire [31:0]       offsetQueueVec_15_enq_bits = offsetReadResult_15_bits;
  wire              offsetQueueVec_16_enq_valid = offsetReadResult_16_valid;
  wire [31:0]       offsetQueueVec_16_enq_bits = offsetReadResult_16_bits;
  wire              offsetQueueVec_17_enq_valid = offsetReadResult_17_valid;
  wire [31:0]       offsetQueueVec_17_enq_bits = offsetReadResult_17_bits;
  wire              offsetQueueVec_18_enq_valid = offsetReadResult_18_valid;
  wire [31:0]       offsetQueueVec_18_enq_bits = offsetReadResult_18_bits;
  wire              offsetQueueVec_19_enq_valid = offsetReadResult_19_valid;
  wire [31:0]       offsetQueueVec_19_enq_bits = offsetReadResult_19_bits;
  wire              offsetQueueVec_20_enq_valid = offsetReadResult_20_valid;
  wire [31:0]       offsetQueueVec_20_enq_bits = offsetReadResult_20_bits;
  wire              offsetQueueVec_21_enq_valid = offsetReadResult_21_valid;
  wire [31:0]       offsetQueueVec_21_enq_bits = offsetReadResult_21_bits;
  wire              offsetQueueVec_22_enq_valid = offsetReadResult_22_valid;
  wire [31:0]       offsetQueueVec_22_enq_bits = offsetReadResult_22_bits;
  wire              offsetQueueVec_23_enq_valid = offsetReadResult_23_valid;
  wire [31:0]       offsetQueueVec_23_enq_bits = offsetReadResult_23_bits;
  wire              offsetQueueVec_24_enq_valid = offsetReadResult_24_valid;
  wire [31:0]       offsetQueueVec_24_enq_bits = offsetReadResult_24_bits;
  wire              offsetQueueVec_25_enq_valid = offsetReadResult_25_valid;
  wire [31:0]       offsetQueueVec_25_enq_bits = offsetReadResult_25_bits;
  wire              offsetQueueVec_26_enq_valid = offsetReadResult_26_valid;
  wire [31:0]       offsetQueueVec_26_enq_bits = offsetReadResult_26_bits;
  wire              offsetQueueVec_27_enq_valid = offsetReadResult_27_valid;
  wire [31:0]       offsetQueueVec_27_enq_bits = offsetReadResult_27_bits;
  wire              offsetQueueVec_28_enq_valid = offsetReadResult_28_valid;
  wire [31:0]       offsetQueueVec_28_enq_bits = offsetReadResult_28_bits;
  wire              offsetQueueVec_29_enq_valid = offsetReadResult_29_valid;
  wire [31:0]       offsetQueueVec_29_enq_bits = offsetReadResult_29_bits;
  wire              offsetQueueVec_30_enq_valid = offsetReadResult_30_valid;
  wire [31:0]       offsetQueueVec_30_enq_bits = offsetReadResult_30_bits;
  wire              offsetQueueVec_31_enq_valid = offsetReadResult_31_valid;
  wire [31:0]       offsetQueueVec_31_enq_bits = offsetReadResult_31_bits;
  wire              s1EnqDataQueue_enq_valid = vrfReadResults_valid;
  wire [31:0]       s1EnqDataQueue_enq_bits = vrfReadResults_bits;
  wire [1:0]        vrfReadDataPorts_bits_readSource = 2'h2;
  wire [1:0]        memReadRequest_bits_size = 2'h2;
  wire [31:0]       s1EnqQueue_enq_bits_readData = 32'h0;
  wire [9:0]        memoryRequestSource;
  wire              vrfWritePort_valid_0 = memReadResponse_valid_0;
  wire [3:0]        storeMask;
  wire [1:0]        dataEEW;
  wire              memReadResponse_ready_0 = vrfWritePort_ready_0;
  wire              writeOffset;
  wire              last;
  wire              offsetQueueVec_0_deq_valid;
  assign offsetQueueVec_0_deq_valid = ~_offsetQueueVec_queue_fifo_empty;
  wire              offsetQueueVec_0_enq_ready = ~_offsetQueueVec_queue_fifo_full;
  wire              offsetQueueVec_0_deq_ready;
  reg               offsetQueueVec_deqLock;
  wire              waitQueueDeq_0 = offsetQueueVec_deqLock;
  wire              _allElementsMasked_T_1 = offsetQueueVec_0_deq_ready & offsetQueueVec_0_deq_valid;
  wire              stateIdle;
  assign offsetQueueVec_0_deq_ready = ~offsetQueueVec_deqLock | stateIdle;
  wire              offsetQueueVec_1_deq_valid;
  assign offsetQueueVec_1_deq_valid = ~_offsetQueueVec_queue_fifo_1_empty;
  wire              offsetQueueVec_1_enq_ready = ~_offsetQueueVec_queue_fifo_1_full;
  wire              offsetQueueVec_1_deq_ready;
  reg               offsetQueueVec_deqLock_1;
  wire              waitQueueDeq_1 = offsetQueueVec_deqLock_1;
  wire              _allElementsMasked_T_2 = offsetQueueVec_1_deq_ready & offsetQueueVec_1_deq_valid;
  assign offsetQueueVec_1_deq_ready = ~offsetQueueVec_deqLock_1 | stateIdle;
  wire              offsetQueueVec_2_deq_valid;
  assign offsetQueueVec_2_deq_valid = ~_offsetQueueVec_queue_fifo_2_empty;
  wire              offsetQueueVec_2_enq_ready = ~_offsetQueueVec_queue_fifo_2_full;
  wire              offsetQueueVec_2_deq_ready;
  reg               offsetQueueVec_deqLock_2;
  wire              waitQueueDeq_2 = offsetQueueVec_deqLock_2;
  wire              _allElementsMasked_T_3 = offsetQueueVec_2_deq_ready & offsetQueueVec_2_deq_valid;
  assign offsetQueueVec_2_deq_ready = ~offsetQueueVec_deqLock_2 | stateIdle;
  wire              offsetQueueVec_3_deq_valid;
  assign offsetQueueVec_3_deq_valid = ~_offsetQueueVec_queue_fifo_3_empty;
  wire              offsetQueueVec_3_enq_ready = ~_offsetQueueVec_queue_fifo_3_full;
  wire              offsetQueueVec_3_deq_ready;
  reg               offsetQueueVec_deqLock_3;
  wire              waitQueueDeq_3 = offsetQueueVec_deqLock_3;
  wire              _allElementsMasked_T_4 = offsetQueueVec_3_deq_ready & offsetQueueVec_3_deq_valid;
  assign offsetQueueVec_3_deq_ready = ~offsetQueueVec_deqLock_3 | stateIdle;
  wire              offsetQueueVec_4_deq_valid;
  assign offsetQueueVec_4_deq_valid = ~_offsetQueueVec_queue_fifo_4_empty;
  wire              offsetQueueVec_4_enq_ready = ~_offsetQueueVec_queue_fifo_4_full;
  wire              offsetQueueVec_4_deq_ready;
  reg               offsetQueueVec_deqLock_4;
  wire              waitQueueDeq_4 = offsetQueueVec_deqLock_4;
  wire              _allElementsMasked_T_5 = offsetQueueVec_4_deq_ready & offsetQueueVec_4_deq_valid;
  assign offsetQueueVec_4_deq_ready = ~offsetQueueVec_deqLock_4 | stateIdle;
  wire              offsetQueueVec_5_deq_valid;
  assign offsetQueueVec_5_deq_valid = ~_offsetQueueVec_queue_fifo_5_empty;
  wire              offsetQueueVec_5_enq_ready = ~_offsetQueueVec_queue_fifo_5_full;
  wire              offsetQueueVec_5_deq_ready;
  reg               offsetQueueVec_deqLock_5;
  wire              waitQueueDeq_5 = offsetQueueVec_deqLock_5;
  wire              _allElementsMasked_T_6 = offsetQueueVec_5_deq_ready & offsetQueueVec_5_deq_valid;
  assign offsetQueueVec_5_deq_ready = ~offsetQueueVec_deqLock_5 | stateIdle;
  wire              offsetQueueVec_6_deq_valid;
  assign offsetQueueVec_6_deq_valid = ~_offsetQueueVec_queue_fifo_6_empty;
  wire              offsetQueueVec_6_enq_ready = ~_offsetQueueVec_queue_fifo_6_full;
  wire              offsetQueueVec_6_deq_ready;
  reg               offsetQueueVec_deqLock_6;
  wire              waitQueueDeq_6 = offsetQueueVec_deqLock_6;
  wire              _allElementsMasked_T_7 = offsetQueueVec_6_deq_ready & offsetQueueVec_6_deq_valid;
  assign offsetQueueVec_6_deq_ready = ~offsetQueueVec_deqLock_6 | stateIdle;
  wire              offsetQueueVec_7_deq_valid;
  assign offsetQueueVec_7_deq_valid = ~_offsetQueueVec_queue_fifo_7_empty;
  wire              offsetQueueVec_7_enq_ready = ~_offsetQueueVec_queue_fifo_7_full;
  wire              offsetQueueVec_7_deq_ready;
  reg               offsetQueueVec_deqLock_7;
  wire              waitQueueDeq_7 = offsetQueueVec_deqLock_7;
  wire              _allElementsMasked_T_8 = offsetQueueVec_7_deq_ready & offsetQueueVec_7_deq_valid;
  assign offsetQueueVec_7_deq_ready = ~offsetQueueVec_deqLock_7 | stateIdle;
  wire              offsetQueueVec_8_deq_valid;
  assign offsetQueueVec_8_deq_valid = ~_offsetQueueVec_queue_fifo_8_empty;
  wire              offsetQueueVec_8_enq_ready = ~_offsetQueueVec_queue_fifo_8_full;
  wire              offsetQueueVec_8_deq_ready;
  reg               offsetQueueVec_deqLock_8;
  wire              waitQueueDeq_8 = offsetQueueVec_deqLock_8;
  wire              _allElementsMasked_T_9 = offsetQueueVec_8_deq_ready & offsetQueueVec_8_deq_valid;
  assign offsetQueueVec_8_deq_ready = ~offsetQueueVec_deqLock_8 | stateIdle;
  wire              offsetQueueVec_9_deq_valid;
  assign offsetQueueVec_9_deq_valid = ~_offsetQueueVec_queue_fifo_9_empty;
  wire              offsetQueueVec_9_enq_ready = ~_offsetQueueVec_queue_fifo_9_full;
  wire              offsetQueueVec_9_deq_ready;
  reg               offsetQueueVec_deqLock_9;
  wire              waitQueueDeq_9 = offsetQueueVec_deqLock_9;
  wire              _allElementsMasked_T_10 = offsetQueueVec_9_deq_ready & offsetQueueVec_9_deq_valid;
  assign offsetQueueVec_9_deq_ready = ~offsetQueueVec_deqLock_9 | stateIdle;
  wire              offsetQueueVec_10_deq_valid;
  assign offsetQueueVec_10_deq_valid = ~_offsetQueueVec_queue_fifo_10_empty;
  wire              offsetQueueVec_10_enq_ready = ~_offsetQueueVec_queue_fifo_10_full;
  wire              offsetQueueVec_10_deq_ready;
  reg               offsetQueueVec_deqLock_10;
  wire              waitQueueDeq_10 = offsetQueueVec_deqLock_10;
  wire              _allElementsMasked_T_11 = offsetQueueVec_10_deq_ready & offsetQueueVec_10_deq_valid;
  assign offsetQueueVec_10_deq_ready = ~offsetQueueVec_deqLock_10 | stateIdle;
  wire              offsetQueueVec_11_deq_valid;
  assign offsetQueueVec_11_deq_valid = ~_offsetQueueVec_queue_fifo_11_empty;
  wire              offsetQueueVec_11_enq_ready = ~_offsetQueueVec_queue_fifo_11_full;
  wire              offsetQueueVec_11_deq_ready;
  reg               offsetQueueVec_deqLock_11;
  wire              waitQueueDeq_11 = offsetQueueVec_deqLock_11;
  wire              _allElementsMasked_T_12 = offsetQueueVec_11_deq_ready & offsetQueueVec_11_deq_valid;
  assign offsetQueueVec_11_deq_ready = ~offsetQueueVec_deqLock_11 | stateIdle;
  wire              offsetQueueVec_12_deq_valid;
  assign offsetQueueVec_12_deq_valid = ~_offsetQueueVec_queue_fifo_12_empty;
  wire              offsetQueueVec_12_enq_ready = ~_offsetQueueVec_queue_fifo_12_full;
  wire              offsetQueueVec_12_deq_ready;
  reg               offsetQueueVec_deqLock_12;
  wire              waitQueueDeq_12 = offsetQueueVec_deqLock_12;
  wire              _allElementsMasked_T_13 = offsetQueueVec_12_deq_ready & offsetQueueVec_12_deq_valid;
  assign offsetQueueVec_12_deq_ready = ~offsetQueueVec_deqLock_12 | stateIdle;
  wire              offsetQueueVec_13_deq_valid;
  assign offsetQueueVec_13_deq_valid = ~_offsetQueueVec_queue_fifo_13_empty;
  wire              offsetQueueVec_13_enq_ready = ~_offsetQueueVec_queue_fifo_13_full;
  wire              offsetQueueVec_13_deq_ready;
  reg               offsetQueueVec_deqLock_13;
  wire              waitQueueDeq_13 = offsetQueueVec_deqLock_13;
  wire              _allElementsMasked_T_14 = offsetQueueVec_13_deq_ready & offsetQueueVec_13_deq_valid;
  assign offsetQueueVec_13_deq_ready = ~offsetQueueVec_deqLock_13 | stateIdle;
  wire              offsetQueueVec_14_deq_valid;
  assign offsetQueueVec_14_deq_valid = ~_offsetQueueVec_queue_fifo_14_empty;
  wire              offsetQueueVec_14_enq_ready = ~_offsetQueueVec_queue_fifo_14_full;
  wire              offsetQueueVec_14_deq_ready;
  reg               offsetQueueVec_deqLock_14;
  wire              waitQueueDeq_14 = offsetQueueVec_deqLock_14;
  wire              _allElementsMasked_T_15 = offsetQueueVec_14_deq_ready & offsetQueueVec_14_deq_valid;
  assign offsetQueueVec_14_deq_ready = ~offsetQueueVec_deqLock_14 | stateIdle;
  wire              offsetQueueVec_15_deq_valid;
  assign offsetQueueVec_15_deq_valid = ~_offsetQueueVec_queue_fifo_15_empty;
  wire              offsetQueueVec_15_enq_ready = ~_offsetQueueVec_queue_fifo_15_full;
  wire              offsetQueueVec_15_deq_ready;
  reg               offsetQueueVec_deqLock_15;
  wire              waitQueueDeq_15 = offsetQueueVec_deqLock_15;
  wire              _allElementsMasked_T_16 = offsetQueueVec_15_deq_ready & offsetQueueVec_15_deq_valid;
  assign offsetQueueVec_15_deq_ready = ~offsetQueueVec_deqLock_15 | stateIdle;
  wire              offsetQueueVec_16_deq_valid;
  assign offsetQueueVec_16_deq_valid = ~_offsetQueueVec_queue_fifo_16_empty;
  wire              offsetQueueVec_16_enq_ready = ~_offsetQueueVec_queue_fifo_16_full;
  wire              offsetQueueVec_16_deq_ready;
  reg               offsetQueueVec_deqLock_16;
  wire              waitQueueDeq_16 = offsetQueueVec_deqLock_16;
  wire              _allElementsMasked_T_17 = offsetQueueVec_16_deq_ready & offsetQueueVec_16_deq_valid;
  assign offsetQueueVec_16_deq_ready = ~offsetQueueVec_deqLock_16 | stateIdle;
  wire              offsetQueueVec_17_deq_valid;
  assign offsetQueueVec_17_deq_valid = ~_offsetQueueVec_queue_fifo_17_empty;
  wire              offsetQueueVec_17_enq_ready = ~_offsetQueueVec_queue_fifo_17_full;
  wire              offsetQueueVec_17_deq_ready;
  reg               offsetQueueVec_deqLock_17;
  wire              waitQueueDeq_17 = offsetQueueVec_deqLock_17;
  wire              _allElementsMasked_T_18 = offsetQueueVec_17_deq_ready & offsetQueueVec_17_deq_valid;
  assign offsetQueueVec_17_deq_ready = ~offsetQueueVec_deqLock_17 | stateIdle;
  wire              offsetQueueVec_18_deq_valid;
  assign offsetQueueVec_18_deq_valid = ~_offsetQueueVec_queue_fifo_18_empty;
  wire              offsetQueueVec_18_enq_ready = ~_offsetQueueVec_queue_fifo_18_full;
  wire              offsetQueueVec_18_deq_ready;
  reg               offsetQueueVec_deqLock_18;
  wire              waitQueueDeq_18 = offsetQueueVec_deqLock_18;
  wire              _allElementsMasked_T_19 = offsetQueueVec_18_deq_ready & offsetQueueVec_18_deq_valid;
  assign offsetQueueVec_18_deq_ready = ~offsetQueueVec_deqLock_18 | stateIdle;
  wire              offsetQueueVec_19_deq_valid;
  assign offsetQueueVec_19_deq_valid = ~_offsetQueueVec_queue_fifo_19_empty;
  wire              offsetQueueVec_19_enq_ready = ~_offsetQueueVec_queue_fifo_19_full;
  wire              offsetQueueVec_19_deq_ready;
  reg               offsetQueueVec_deqLock_19;
  wire              waitQueueDeq_19 = offsetQueueVec_deqLock_19;
  wire              _allElementsMasked_T_20 = offsetQueueVec_19_deq_ready & offsetQueueVec_19_deq_valid;
  assign offsetQueueVec_19_deq_ready = ~offsetQueueVec_deqLock_19 | stateIdle;
  wire              offsetQueueVec_20_deq_valid;
  assign offsetQueueVec_20_deq_valid = ~_offsetQueueVec_queue_fifo_20_empty;
  wire              offsetQueueVec_20_enq_ready = ~_offsetQueueVec_queue_fifo_20_full;
  wire              offsetQueueVec_20_deq_ready;
  reg               offsetQueueVec_deqLock_20;
  wire              waitQueueDeq_20 = offsetQueueVec_deqLock_20;
  wire              _allElementsMasked_T_21 = offsetQueueVec_20_deq_ready & offsetQueueVec_20_deq_valid;
  assign offsetQueueVec_20_deq_ready = ~offsetQueueVec_deqLock_20 | stateIdle;
  wire              offsetQueueVec_21_deq_valid;
  assign offsetQueueVec_21_deq_valid = ~_offsetQueueVec_queue_fifo_21_empty;
  wire              offsetQueueVec_21_enq_ready = ~_offsetQueueVec_queue_fifo_21_full;
  wire              offsetQueueVec_21_deq_ready;
  reg               offsetQueueVec_deqLock_21;
  wire              waitQueueDeq_21 = offsetQueueVec_deqLock_21;
  wire              _allElementsMasked_T_22 = offsetQueueVec_21_deq_ready & offsetQueueVec_21_deq_valid;
  assign offsetQueueVec_21_deq_ready = ~offsetQueueVec_deqLock_21 | stateIdle;
  wire              offsetQueueVec_22_deq_valid;
  assign offsetQueueVec_22_deq_valid = ~_offsetQueueVec_queue_fifo_22_empty;
  wire              offsetQueueVec_22_enq_ready = ~_offsetQueueVec_queue_fifo_22_full;
  wire              offsetQueueVec_22_deq_ready;
  reg               offsetQueueVec_deqLock_22;
  wire              waitQueueDeq_22 = offsetQueueVec_deqLock_22;
  wire              _allElementsMasked_T_23 = offsetQueueVec_22_deq_ready & offsetQueueVec_22_deq_valid;
  assign offsetQueueVec_22_deq_ready = ~offsetQueueVec_deqLock_22 | stateIdle;
  wire              offsetQueueVec_23_deq_valid;
  assign offsetQueueVec_23_deq_valid = ~_offsetQueueVec_queue_fifo_23_empty;
  wire              offsetQueueVec_23_enq_ready = ~_offsetQueueVec_queue_fifo_23_full;
  wire              offsetQueueVec_23_deq_ready;
  reg               offsetQueueVec_deqLock_23;
  wire              waitQueueDeq_23 = offsetQueueVec_deqLock_23;
  wire              _allElementsMasked_T_24 = offsetQueueVec_23_deq_ready & offsetQueueVec_23_deq_valid;
  assign offsetQueueVec_23_deq_ready = ~offsetQueueVec_deqLock_23 | stateIdle;
  wire              offsetQueueVec_24_deq_valid;
  assign offsetQueueVec_24_deq_valid = ~_offsetQueueVec_queue_fifo_24_empty;
  wire              offsetQueueVec_24_enq_ready = ~_offsetQueueVec_queue_fifo_24_full;
  wire              offsetQueueVec_24_deq_ready;
  reg               offsetQueueVec_deqLock_24;
  wire              waitQueueDeq_24 = offsetQueueVec_deqLock_24;
  wire              _allElementsMasked_T_25 = offsetQueueVec_24_deq_ready & offsetQueueVec_24_deq_valid;
  assign offsetQueueVec_24_deq_ready = ~offsetQueueVec_deqLock_24 | stateIdle;
  wire              offsetQueueVec_25_deq_valid;
  assign offsetQueueVec_25_deq_valid = ~_offsetQueueVec_queue_fifo_25_empty;
  wire              offsetQueueVec_25_enq_ready = ~_offsetQueueVec_queue_fifo_25_full;
  wire              offsetQueueVec_25_deq_ready;
  reg               offsetQueueVec_deqLock_25;
  wire              waitQueueDeq_25 = offsetQueueVec_deqLock_25;
  wire              _allElementsMasked_T_26 = offsetQueueVec_25_deq_ready & offsetQueueVec_25_deq_valid;
  assign offsetQueueVec_25_deq_ready = ~offsetQueueVec_deqLock_25 | stateIdle;
  wire              offsetQueueVec_26_deq_valid;
  assign offsetQueueVec_26_deq_valid = ~_offsetQueueVec_queue_fifo_26_empty;
  wire              offsetQueueVec_26_enq_ready = ~_offsetQueueVec_queue_fifo_26_full;
  wire              offsetQueueVec_26_deq_ready;
  reg               offsetQueueVec_deqLock_26;
  wire              waitQueueDeq_26 = offsetQueueVec_deqLock_26;
  wire              _allElementsMasked_T_27 = offsetQueueVec_26_deq_ready & offsetQueueVec_26_deq_valid;
  assign offsetQueueVec_26_deq_ready = ~offsetQueueVec_deqLock_26 | stateIdle;
  wire              offsetQueueVec_27_deq_valid;
  assign offsetQueueVec_27_deq_valid = ~_offsetQueueVec_queue_fifo_27_empty;
  wire              offsetQueueVec_27_enq_ready = ~_offsetQueueVec_queue_fifo_27_full;
  wire              offsetQueueVec_27_deq_ready;
  reg               offsetQueueVec_deqLock_27;
  wire              waitQueueDeq_27 = offsetQueueVec_deqLock_27;
  wire              _allElementsMasked_T_28 = offsetQueueVec_27_deq_ready & offsetQueueVec_27_deq_valid;
  assign offsetQueueVec_27_deq_ready = ~offsetQueueVec_deqLock_27 | stateIdle;
  wire              offsetQueueVec_28_deq_valid;
  assign offsetQueueVec_28_deq_valid = ~_offsetQueueVec_queue_fifo_28_empty;
  wire              offsetQueueVec_28_enq_ready = ~_offsetQueueVec_queue_fifo_28_full;
  wire              offsetQueueVec_28_deq_ready;
  reg               offsetQueueVec_deqLock_28;
  wire              waitQueueDeq_28 = offsetQueueVec_deqLock_28;
  wire              _allElementsMasked_T_29 = offsetQueueVec_28_deq_ready & offsetQueueVec_28_deq_valid;
  assign offsetQueueVec_28_deq_ready = ~offsetQueueVec_deqLock_28 | stateIdle;
  wire              offsetQueueVec_29_deq_valid;
  assign offsetQueueVec_29_deq_valid = ~_offsetQueueVec_queue_fifo_29_empty;
  wire              offsetQueueVec_29_enq_ready = ~_offsetQueueVec_queue_fifo_29_full;
  wire              offsetQueueVec_29_deq_ready;
  reg               offsetQueueVec_deqLock_29;
  wire              waitQueueDeq_29 = offsetQueueVec_deqLock_29;
  wire              _allElementsMasked_T_30 = offsetQueueVec_29_deq_ready & offsetQueueVec_29_deq_valid;
  assign offsetQueueVec_29_deq_ready = ~offsetQueueVec_deqLock_29 | stateIdle;
  wire              offsetQueueVec_30_deq_valid;
  assign offsetQueueVec_30_deq_valid = ~_offsetQueueVec_queue_fifo_30_empty;
  wire              offsetQueueVec_30_enq_ready = ~_offsetQueueVec_queue_fifo_30_full;
  wire              offsetQueueVec_30_deq_ready;
  reg               offsetQueueVec_deqLock_30;
  wire              waitQueueDeq_30 = offsetQueueVec_deqLock_30;
  wire              _allElementsMasked_T_31 = offsetQueueVec_30_deq_ready & offsetQueueVec_30_deq_valid;
  assign offsetQueueVec_30_deq_ready = ~offsetQueueVec_deqLock_30 | stateIdle;
  wire              offsetQueueVec_31_deq_valid;
  assign offsetQueueVec_31_deq_valid = ~_offsetQueueVec_queue_fifo_31_empty;
  wire              offsetQueueVec_31_enq_ready = ~_offsetQueueVec_queue_fifo_31_full;
  wire              offsetQueueVec_31_deq_ready;
  reg               offsetQueueVec_deqLock_31;
  wire              waitQueueDeq_31 = offsetQueueVec_deqLock_31;
  wire              _allElementsMasked_T_32 = offsetQueueVec_31_deq_ready & offsetQueueVec_31_deq_valid;
  assign offsetQueueVec_31_deq_ready = ~offsetQueueVec_deqLock_31 | stateIdle;
  wire              memReadRequest_valid_0;
  wire              _outstandingTLDMessages_T_4 = memReadRequest_ready_0 & memReadRequest_valid_0;
  wire              memWriteRequest_valid_0;
  wire              _probeWire_valid_T = memWriteRequest_ready_0 & memWriteRequest_valid_0;
  wire              memRequestFire = _outstandingTLDMessages_T_4 | _probeWire_valid_T;
  reg  [2:0]        lsuRequestReg_instructionInformation_nf;
  reg               lsuRequestReg_instructionInformation_mew;
  reg  [1:0]        lsuRequestReg_instructionInformation_mop;
  reg  [4:0]        lsuRequestReg_instructionInformation_lumop;
  reg  [1:0]        lsuRequestReg_instructionInformation_eew;
  reg  [4:0]        lsuRequestReg_instructionInformation_vs3;
  reg               lsuRequestReg_instructionInformation_isStore;
  reg               lsuRequestReg_instructionInformation_maskedLoadStore;
  reg  [31:0]       lsuRequestReg_rs1Data;
  reg  [31:0]       lsuRequestReg_rs2Data;
  reg  [2:0]        lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfWritePort_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  reg  [11:0]       csrInterfaceReg_vl;
  reg  [11:0]       csrInterfaceReg_vStart;
  reg  [2:0]        csrInterfaceReg_vlmul;
  reg  [1:0]        csrInterfaceReg_vSew;
  reg  [1:0]        csrInterfaceReg_vxrm;
  reg               csrInterfaceReg_vta;
  reg               csrInterfaceReg_vma;
  wire              _isMaskLoadStore_T = lsuRequestReg_instructionInformation_mop == 2'h0;
  wire              isWholeRegisterLoadStore = _isMaskLoadStore_T & lsuRequestReg_instructionInformation_lumop == 5'h8;
  wire              isSegmentLoadStore = (|lsuRequestReg_instructionInformation_nf) & ~isWholeRegisterLoadStore;
  wire              isMaskLoadStore = _isMaskLoadStore_T & lsuRequestReg_instructionInformation_lumop[0];
  wire              isIndexedLoadStore = lsuRequestReg_instructionInformation_mop[0];
  wire              _waitFirstMemoryResponseForFaultOnlyFirst_T = lsuRequest_bits_instructionInformation_mop == 2'h0;
  wire              requestIsWholeRegisterLoadStore = _waitFirstMemoryResponseForFaultOnlyFirst_T & lsuRequest_bits_instructionInformation_lumop == 5'h8;
  wire              requestIsMaskLoadStore = _waitFirstMemoryResponseForFaultOnlyFirst_T & lsuRequest_bits_instructionInformation_lumop[0];
  wire [1:0]        requestEEW = lsuRequest_bits_instructionInformation_mop[0] ? csrInterface_vSew : requestIsMaskLoadStore ? 2'h0 : requestIsWholeRegisterLoadStore ? 2'h2 : lsuRequest_bits_instructionInformation_eew;
  wire [2:0]        requestNF = requestIsWholeRegisterLoadStore ? 3'h0 : lsuRequest_bits_instructionInformation_nf;
  reg  [6:0]        dataWidthForSegmentLoadStore;
  reg  [2:0]        elementByteWidth;
  reg  [3:0]        segmentInstructionIndexInterval;
  reg  [127:0]      outstandingTLDMessages;
  wire              noOutstandingMessages = outstandingTLDMessages == 128'h0;
  reg               indexedInstructionOffsets_0_valid;
  reg  [31:0]       indexedInstructionOffsets_0_bits;
  reg               indexedInstructionOffsets_1_valid;
  reg  [31:0]       indexedInstructionOffsets_1_bits;
  reg               indexedInstructionOffsets_2_valid;
  reg  [31:0]       indexedInstructionOffsets_2_bits;
  reg               indexedInstructionOffsets_3_valid;
  reg  [31:0]       indexedInstructionOffsets_3_bits;
  reg               indexedInstructionOffsets_4_valid;
  reg  [31:0]       indexedInstructionOffsets_4_bits;
  reg               indexedInstructionOffsets_5_valid;
  reg  [31:0]       indexedInstructionOffsets_5_bits;
  reg               indexedInstructionOffsets_6_valid;
  reg  [31:0]       indexedInstructionOffsets_6_bits;
  reg               indexedInstructionOffsets_7_valid;
  reg  [31:0]       indexedInstructionOffsets_7_bits;
  reg               indexedInstructionOffsets_8_valid;
  reg  [31:0]       indexedInstructionOffsets_8_bits;
  reg               indexedInstructionOffsets_9_valid;
  reg  [31:0]       indexedInstructionOffsets_9_bits;
  reg               indexedInstructionOffsets_10_valid;
  reg  [31:0]       indexedInstructionOffsets_10_bits;
  reg               indexedInstructionOffsets_11_valid;
  reg  [31:0]       indexedInstructionOffsets_11_bits;
  reg               indexedInstructionOffsets_12_valid;
  reg  [31:0]       indexedInstructionOffsets_12_bits;
  reg               indexedInstructionOffsets_13_valid;
  reg  [31:0]       indexedInstructionOffsets_13_bits;
  reg               indexedInstructionOffsets_14_valid;
  reg  [31:0]       indexedInstructionOffsets_14_bits;
  reg               indexedInstructionOffsets_15_valid;
  reg  [31:0]       indexedInstructionOffsets_15_bits;
  reg               indexedInstructionOffsets_16_valid;
  reg  [31:0]       indexedInstructionOffsets_16_bits;
  reg               indexedInstructionOffsets_17_valid;
  reg  [31:0]       indexedInstructionOffsets_17_bits;
  reg               indexedInstructionOffsets_18_valid;
  reg  [31:0]       indexedInstructionOffsets_18_bits;
  reg               indexedInstructionOffsets_19_valid;
  reg  [31:0]       indexedInstructionOffsets_19_bits;
  reg               indexedInstructionOffsets_20_valid;
  reg  [31:0]       indexedInstructionOffsets_20_bits;
  reg               indexedInstructionOffsets_21_valid;
  reg  [31:0]       indexedInstructionOffsets_21_bits;
  reg               indexedInstructionOffsets_22_valid;
  reg  [31:0]       indexedInstructionOffsets_22_bits;
  reg               indexedInstructionOffsets_23_valid;
  reg  [31:0]       indexedInstructionOffsets_23_bits;
  reg               indexedInstructionOffsets_24_valid;
  reg  [31:0]       indexedInstructionOffsets_24_bits;
  reg               indexedInstructionOffsets_25_valid;
  reg  [31:0]       indexedInstructionOffsets_25_bits;
  reg               indexedInstructionOffsets_26_valid;
  reg  [31:0]       indexedInstructionOffsets_26_bits;
  reg               indexedInstructionOffsets_27_valid;
  reg  [31:0]       indexedInstructionOffsets_27_bits;
  reg               indexedInstructionOffsets_28_valid;
  reg  [31:0]       indexedInstructionOffsets_28_bits;
  reg               indexedInstructionOffsets_29_valid;
  reg  [31:0]       indexedInstructionOffsets_29_bits;
  reg               indexedInstructionOffsets_30_valid;
  reg  [31:0]       indexedInstructionOffsets_30_bits;
  reg               indexedInstructionOffsets_31_valid;
  reg  [31:0]       indexedInstructionOffsets_31_bits;
  reg  [4:0]        groupIndex;
  wire [4:0]        nextGroupIndex = lsuRequest_valid ? 5'h0 : groupIndex + 5'h1;
  reg  [1:0]        indexOfIndexedInstructionOffsets;
  wire [1:0]        indexOfIndexedInstructionOffsetsNext = lsuRequest_valid ? 2'h3 : indexOfIndexedInstructionOffsets + 2'h1;
  reg  [127:0]      maskReg;
  reg  [2:0]        segmentIndex;
  wire [2:0]        s0Wire_segmentIndex = segmentIndex;
  wire [2:0]        segmentIndexNext = segmentIndex + 3'h1;
  wire              segmentEnd = segmentIndex == lsuRequestReg_instructionInformation_nf;
  wire              lastElementForSegment = ~isSegmentLoadStore | segmentEnd;
  wire              s0Fire;
  wire              segmentEndWithHandshake = s0Fire & lastElementForSegment;
  reg  [1:0]        state;
  reg  [127:0]      sentMemoryRequests;
  wire [127:0]      unsentMemoryRequests = ~sentMemoryRequests;
  wire [127:0]      maskedUnsentMemoryRequests = maskReg & unsentMemoryRequests;
  wire [126:0]      _findFirstMaskedUnsentMemoryRequests_T_2 = maskedUnsentMemoryRequests[126:0] | {maskedUnsentMemoryRequests[125:0], 1'h0};
  wire [126:0]      _findFirstMaskedUnsentMemoryRequests_T_5 = _findFirstMaskedUnsentMemoryRequests_T_2 | {_findFirstMaskedUnsentMemoryRequests_T_2[124:0], 2'h0};
  wire [126:0]      _findFirstMaskedUnsentMemoryRequests_T_8 = _findFirstMaskedUnsentMemoryRequests_T_5 | {_findFirstMaskedUnsentMemoryRequests_T_5[122:0], 4'h0};
  wire [126:0]      _findFirstMaskedUnsentMemoryRequests_T_11 = _findFirstMaskedUnsentMemoryRequests_T_8 | {_findFirstMaskedUnsentMemoryRequests_T_8[118:0], 8'h0};
  wire [126:0]      _findFirstMaskedUnsentMemoryRequests_T_14 = _findFirstMaskedUnsentMemoryRequests_T_11 | {_findFirstMaskedUnsentMemoryRequests_T_11[110:0], 16'h0};
  wire [126:0]      _findFirstMaskedUnsentMemoryRequests_T_17 = _findFirstMaskedUnsentMemoryRequests_T_14 | {_findFirstMaskedUnsentMemoryRequests_T_14[94:0], 32'h0};
  wire [127:0]      findFirstMaskedUnsentMemoryRequests = {~(_findFirstMaskedUnsentMemoryRequests_T_17 | {_findFirstMaskedUnsentMemoryRequests_T_17[62:0], 64'h0}), 1'h1} & maskedUnsentMemoryRequests;
  wire [128:0]      findFirstUnsentMemoryRequestsNext = {1'h0, {sentMemoryRequests[126:0], 1'h1} & unsentMemoryRequests};
  wire [127:0]      nextElementForMemoryRequest = lsuRequestReg_instructionInformation_maskedLoadStore ? findFirstMaskedUnsentMemoryRequests : findFirstUnsentMemoryRequestsNext[127:0];
  wire [63:0]       nextElementForMemoryRequestIndex_hi = nextElementForMemoryRequest[127:64];
  wire [63:0]       nextElementForMemoryRequestIndex_lo = nextElementForMemoryRequest[63:0];
  wire [63:0]       _nextElementForMemoryRequestIndex_T_1 = nextElementForMemoryRequestIndex_hi | nextElementForMemoryRequestIndex_lo;
  wire [31:0]       nextElementForMemoryRequestIndex_hi_1 = _nextElementForMemoryRequestIndex_T_1[63:32];
  wire [31:0]       nextElementForMemoryRequestIndex_lo_1 = _nextElementForMemoryRequestIndex_T_1[31:0];
  wire [31:0]       _nextElementForMemoryRequestIndex_T_3 = nextElementForMemoryRequestIndex_hi_1 | nextElementForMemoryRequestIndex_lo_1;
  wire [15:0]       nextElementForMemoryRequestIndex_hi_2 = _nextElementForMemoryRequestIndex_T_3[31:16];
  wire [15:0]       nextElementForMemoryRequestIndex_lo_2 = _nextElementForMemoryRequestIndex_T_3[15:0];
  wire [15:0]       _nextElementForMemoryRequestIndex_T_5 = nextElementForMemoryRequestIndex_hi_2 | nextElementForMemoryRequestIndex_lo_2;
  wire [7:0]        nextElementForMemoryRequestIndex_hi_3 = _nextElementForMemoryRequestIndex_T_5[15:8];
  wire [7:0]        nextElementForMemoryRequestIndex_lo_3 = _nextElementForMemoryRequestIndex_T_5[7:0];
  wire [7:0]        _nextElementForMemoryRequestIndex_T_7 = nextElementForMemoryRequestIndex_hi_3 | nextElementForMemoryRequestIndex_lo_3;
  wire [3:0]        nextElementForMemoryRequestIndex_hi_4 = _nextElementForMemoryRequestIndex_T_7[7:4];
  wire [3:0]        nextElementForMemoryRequestIndex_lo_4 = _nextElementForMemoryRequestIndex_T_7[3:0];
  wire [3:0]        _nextElementForMemoryRequestIndex_T_9 = nextElementForMemoryRequestIndex_hi_4 | nextElementForMemoryRequestIndex_lo_4;
  wire [1:0]        nextElementForMemoryRequestIndex_hi_5 = _nextElementForMemoryRequestIndex_T_9[3:2];
  wire [1:0]        nextElementForMemoryRequestIndex_lo_5 = _nextElementForMemoryRequestIndex_T_9[1:0];
  wire [6:0]        nextElementForMemoryRequestIndex =
    {|nextElementForMemoryRequestIndex_hi,
     |nextElementForMemoryRequestIndex_hi_1,
     |nextElementForMemoryRequestIndex_hi_2,
     |nextElementForMemoryRequestIndex_hi_3,
     |nextElementForMemoryRequestIndex_hi_4,
     |nextElementForMemoryRequestIndex_hi_5,
     nextElementForMemoryRequestIndex_hi_5[1] | nextElementForMemoryRequestIndex_lo_5[1]};
  wire [6:0]        s0Wire_indexInGroup = nextElementForMemoryRequestIndex;
  assign dataEEW = isIndexedLoadStore ? csrInterfaceReg_vSew : isMaskLoadStore ? 2'h0 : isWholeRegisterLoadStore ? 2'h2 : lsuRequestReg_instructionInformation_eew;
  wire [1:0]        memWriteRequest_bits_size_0 = dataEEW;
  wire [3:0]        dataEEWOH = 4'h1 << dataEEW;
  wire              noMoreMaskedUnsentMemoryRequests = maskedUnsentMemoryRequests == 128'h0;
  wire              maskGroupEndAndRequestNewMask = (noMoreMaskedUnsentMemoryRequests | nextElementForMemoryRequest[127] & segmentEndWithHandshake) & lsuRequestReg_instructionInformation_maskedLoadStore;
  wire              maskGroupEnd = maskGroupEndAndRequestNewMask | nextElementForMemoryRequest[127] & segmentEndWithHandshake;
  wire [3:0]        _offsetEEWOH_T = 4'h1 << lsuRequestReg_instructionInformation_eew;
  wire [2:0]        offsetEEWOH = _offsetEEWOH_T[2:0];
  wire [11:0]       _offsetForStride_T = {groupIndex, nextElementForMemoryRequestIndex};
  wire [11:0]       offsetForUnitStride;
  assign offsetForUnitStride = _offsetForStride_T;
  wire [11:0]       s0ElementIndex;
  assign s0ElementIndex = _offsetForStride_T;
  wire [14:0]       _globalOffsetOfIndexedInstructionOffsets_T_1 = {3'h0, groupIndex, nextElementForMemoryRequestIndex} << lsuRequestReg_instructionInformation_eew;
  wire [8:0]        globalOffsetOfIndexedInstructionOffsets = _globalOffsetOfIndexedInstructionOffsets_T_1[8:0];
  wire [1:0]        offsetGroupIndexOfMemoryRequest = globalOffsetOfIndexedInstructionOffsets[8:7];
  wire [6:0]        offsetOfOffsetGroup = globalOffsetOfIndexedInstructionOffsets[6:0];
  wire [63:0]       offsetOfCurrentMemoryRequest_lo_lo_lo_lo = {indexedInstructionOffsets_1_bits, indexedInstructionOffsets_0_bits};
  wire [63:0]       offsetOfCurrentMemoryRequest_lo_lo_lo_hi = {indexedInstructionOffsets_3_bits, indexedInstructionOffsets_2_bits};
  wire [127:0]      offsetOfCurrentMemoryRequest_lo_lo_lo = {offsetOfCurrentMemoryRequest_lo_lo_lo_hi, offsetOfCurrentMemoryRequest_lo_lo_lo_lo};
  wire [63:0]       offsetOfCurrentMemoryRequest_lo_lo_hi_lo = {indexedInstructionOffsets_5_bits, indexedInstructionOffsets_4_bits};
  wire [63:0]       offsetOfCurrentMemoryRequest_lo_lo_hi_hi = {indexedInstructionOffsets_7_bits, indexedInstructionOffsets_6_bits};
  wire [127:0]      offsetOfCurrentMemoryRequest_lo_lo_hi = {offsetOfCurrentMemoryRequest_lo_lo_hi_hi, offsetOfCurrentMemoryRequest_lo_lo_hi_lo};
  wire [255:0]      offsetOfCurrentMemoryRequest_lo_lo = {offsetOfCurrentMemoryRequest_lo_lo_hi, offsetOfCurrentMemoryRequest_lo_lo_lo};
  wire [63:0]       offsetOfCurrentMemoryRequest_lo_hi_lo_lo = {indexedInstructionOffsets_9_bits, indexedInstructionOffsets_8_bits};
  wire [63:0]       offsetOfCurrentMemoryRequest_lo_hi_lo_hi = {indexedInstructionOffsets_11_bits, indexedInstructionOffsets_10_bits};
  wire [127:0]      offsetOfCurrentMemoryRequest_lo_hi_lo = {offsetOfCurrentMemoryRequest_lo_hi_lo_hi, offsetOfCurrentMemoryRequest_lo_hi_lo_lo};
  wire [63:0]       offsetOfCurrentMemoryRequest_lo_hi_hi_lo = {indexedInstructionOffsets_13_bits, indexedInstructionOffsets_12_bits};
  wire [63:0]       offsetOfCurrentMemoryRequest_lo_hi_hi_hi = {indexedInstructionOffsets_15_bits, indexedInstructionOffsets_14_bits};
  wire [127:0]      offsetOfCurrentMemoryRequest_lo_hi_hi = {offsetOfCurrentMemoryRequest_lo_hi_hi_hi, offsetOfCurrentMemoryRequest_lo_hi_hi_lo};
  wire [255:0]      offsetOfCurrentMemoryRequest_lo_hi = {offsetOfCurrentMemoryRequest_lo_hi_hi, offsetOfCurrentMemoryRequest_lo_hi_lo};
  wire [511:0]      offsetOfCurrentMemoryRequest_lo = {offsetOfCurrentMemoryRequest_lo_hi, offsetOfCurrentMemoryRequest_lo_lo};
  wire [63:0]       offsetOfCurrentMemoryRequest_hi_lo_lo_lo = {indexedInstructionOffsets_17_bits, indexedInstructionOffsets_16_bits};
  wire [63:0]       offsetOfCurrentMemoryRequest_hi_lo_lo_hi = {indexedInstructionOffsets_19_bits, indexedInstructionOffsets_18_bits};
  wire [127:0]      offsetOfCurrentMemoryRequest_hi_lo_lo = {offsetOfCurrentMemoryRequest_hi_lo_lo_hi, offsetOfCurrentMemoryRequest_hi_lo_lo_lo};
  wire [63:0]       offsetOfCurrentMemoryRequest_hi_lo_hi_lo = {indexedInstructionOffsets_21_bits, indexedInstructionOffsets_20_bits};
  wire [63:0]       offsetOfCurrentMemoryRequest_hi_lo_hi_hi = {indexedInstructionOffsets_23_bits, indexedInstructionOffsets_22_bits};
  wire [127:0]      offsetOfCurrentMemoryRequest_hi_lo_hi = {offsetOfCurrentMemoryRequest_hi_lo_hi_hi, offsetOfCurrentMemoryRequest_hi_lo_hi_lo};
  wire [255:0]      offsetOfCurrentMemoryRequest_hi_lo = {offsetOfCurrentMemoryRequest_hi_lo_hi, offsetOfCurrentMemoryRequest_hi_lo_lo};
  wire [63:0]       offsetOfCurrentMemoryRequest_hi_hi_lo_lo = {indexedInstructionOffsets_25_bits, indexedInstructionOffsets_24_bits};
  wire [63:0]       offsetOfCurrentMemoryRequest_hi_hi_lo_hi = {indexedInstructionOffsets_27_bits, indexedInstructionOffsets_26_bits};
  wire [127:0]      offsetOfCurrentMemoryRequest_hi_hi_lo = {offsetOfCurrentMemoryRequest_hi_hi_lo_hi, offsetOfCurrentMemoryRequest_hi_hi_lo_lo};
  wire [63:0]       offsetOfCurrentMemoryRequest_hi_hi_hi_lo = {indexedInstructionOffsets_29_bits, indexedInstructionOffsets_28_bits};
  wire [63:0]       offsetOfCurrentMemoryRequest_hi_hi_hi_hi = {indexedInstructionOffsets_31_bits, indexedInstructionOffsets_30_bits};
  wire [127:0]      offsetOfCurrentMemoryRequest_hi_hi_hi = {offsetOfCurrentMemoryRequest_hi_hi_hi_hi, offsetOfCurrentMemoryRequest_hi_hi_hi_lo};
  wire [255:0]      offsetOfCurrentMemoryRequest_hi_hi = {offsetOfCurrentMemoryRequest_hi_hi_hi, offsetOfCurrentMemoryRequest_hi_hi_lo};
  wire [511:0]      offsetOfCurrentMemoryRequest_hi = {offsetOfCurrentMemoryRequest_hi_hi, offsetOfCurrentMemoryRequest_hi_lo};
  wire [1023:0]     _offsetOfCurrentMemoryRequest_T_2 = {offsetOfCurrentMemoryRequest_hi, offsetOfCurrentMemoryRequest_lo} >> {1014'h0, offsetOfOffsetGroup, 3'h0};
  wire [15:0]       offsetOfCurrentMemoryRequest_lo_1 = {{8{~(offsetEEWOH[0])}}, 8'hFF};
  wire [15:0]       offsetOfCurrentMemoryRequest_hi_1 = {16{offsetEEWOH[2]}};
  wire [31:0]       offsetOfCurrentMemoryRequest = _offsetOfCurrentMemoryRequest_T_2[31:0] & {offsetOfCurrentMemoryRequest_hi_1, offsetOfCurrentMemoryRequest_lo_1};
  wire [1:0]        offsetValidCheck_lo_lo_lo_lo = {indexedInstructionOffsets_1_valid, indexedInstructionOffsets_0_valid};
  wire [1:0]        offsetValidCheck_lo_lo_lo_hi = {indexedInstructionOffsets_3_valid, indexedInstructionOffsets_2_valid};
  wire [3:0]        offsetValidCheck_lo_lo_lo = {offsetValidCheck_lo_lo_lo_hi, offsetValidCheck_lo_lo_lo_lo};
  wire [1:0]        offsetValidCheck_lo_lo_hi_lo = {indexedInstructionOffsets_5_valid, indexedInstructionOffsets_4_valid};
  wire [1:0]        offsetValidCheck_lo_lo_hi_hi = {indexedInstructionOffsets_7_valid, indexedInstructionOffsets_6_valid};
  wire [3:0]        offsetValidCheck_lo_lo_hi = {offsetValidCheck_lo_lo_hi_hi, offsetValidCheck_lo_lo_hi_lo};
  wire [7:0]        offsetValidCheck_lo_lo = {offsetValidCheck_lo_lo_hi, offsetValidCheck_lo_lo_lo};
  wire [1:0]        offsetValidCheck_lo_hi_lo_lo = {indexedInstructionOffsets_9_valid, indexedInstructionOffsets_8_valid};
  wire [1:0]        offsetValidCheck_lo_hi_lo_hi = {indexedInstructionOffsets_11_valid, indexedInstructionOffsets_10_valid};
  wire [3:0]        offsetValidCheck_lo_hi_lo = {offsetValidCheck_lo_hi_lo_hi, offsetValidCheck_lo_hi_lo_lo};
  wire [1:0]        offsetValidCheck_lo_hi_hi_lo = {indexedInstructionOffsets_13_valid, indexedInstructionOffsets_12_valid};
  wire [1:0]        offsetValidCheck_lo_hi_hi_hi = {indexedInstructionOffsets_15_valid, indexedInstructionOffsets_14_valid};
  wire [3:0]        offsetValidCheck_lo_hi_hi = {offsetValidCheck_lo_hi_hi_hi, offsetValidCheck_lo_hi_hi_lo};
  wire [7:0]        offsetValidCheck_lo_hi = {offsetValidCheck_lo_hi_hi, offsetValidCheck_lo_hi_lo};
  wire [15:0]       offsetValidCheck_lo = {offsetValidCheck_lo_hi, offsetValidCheck_lo_lo};
  wire [1:0]        offsetValidCheck_hi_lo_lo_lo = {indexedInstructionOffsets_17_valid, indexedInstructionOffsets_16_valid};
  wire [1:0]        offsetValidCheck_hi_lo_lo_hi = {indexedInstructionOffsets_19_valid, indexedInstructionOffsets_18_valid};
  wire [3:0]        offsetValidCheck_hi_lo_lo = {offsetValidCheck_hi_lo_lo_hi, offsetValidCheck_hi_lo_lo_lo};
  wire [1:0]        offsetValidCheck_hi_lo_hi_lo = {indexedInstructionOffsets_21_valid, indexedInstructionOffsets_20_valid};
  wire [1:0]        offsetValidCheck_hi_lo_hi_hi = {indexedInstructionOffsets_23_valid, indexedInstructionOffsets_22_valid};
  wire [3:0]        offsetValidCheck_hi_lo_hi = {offsetValidCheck_hi_lo_hi_hi, offsetValidCheck_hi_lo_hi_lo};
  wire [7:0]        offsetValidCheck_hi_lo = {offsetValidCheck_hi_lo_hi, offsetValidCheck_hi_lo_lo};
  wire [1:0]        offsetValidCheck_hi_hi_lo_lo = {indexedInstructionOffsets_25_valid, indexedInstructionOffsets_24_valid};
  wire [1:0]        offsetValidCheck_hi_hi_lo_hi = {indexedInstructionOffsets_27_valid, indexedInstructionOffsets_26_valid};
  wire [3:0]        offsetValidCheck_hi_hi_lo = {offsetValidCheck_hi_hi_lo_hi, offsetValidCheck_hi_hi_lo_lo};
  wire [1:0]        offsetValidCheck_hi_hi_hi_lo = {indexedInstructionOffsets_29_valid, indexedInstructionOffsets_28_valid};
  wire [1:0]        offsetValidCheck_hi_hi_hi_hi = {indexedInstructionOffsets_31_valid, indexedInstructionOffsets_30_valid};
  wire [3:0]        offsetValidCheck_hi_hi_hi = {offsetValidCheck_hi_hi_hi_hi, offsetValidCheck_hi_hi_hi_lo};
  wire [7:0]        offsetValidCheck_hi_hi = {offsetValidCheck_hi_hi_hi, offsetValidCheck_hi_hi_lo};
  wire [15:0]       offsetValidCheck_hi = {offsetValidCheck_hi_hi, offsetValidCheck_hi_lo};
  wire [31:0]       _offsetValidCheck_T_2 = {offsetValidCheck_hi, offsetValidCheck_lo} >> offsetOfOffsetGroup[6:2];
  wire              offsetValidCheck = _offsetValidCheck_T_2[0];
  wire [1:0]        offsetGroupMatch = offsetGroupIndexOfMemoryRequest ^ indexOfIndexedInstructionOffsets;
  wire              offsetGroupCheck = (~(lsuRequestReg_instructionInformation_eew[0]) | ~(offsetGroupMatch[0])) & (~(lsuRequestReg_instructionInformation_eew[1]) | offsetGroupMatch == 2'h0);
  wire [43:0]       offsetForStride = {32'h0, groupIndex, nextElementForMemoryRequestIndex} * {12'h0, lsuRequestReg_rs2Data};
  wire [43:0]       baseOffsetForElement =
    isIndexedLoadStore ? {12'h0, offsetOfCurrentMemoryRequest} : lsuRequestReg_instructionInformation_mop[1] ? offsetForStride : {25'h0, {7'h0, offsetForUnitStride} * {12'h0, dataWidthForSegmentLoadStore}};
  wire [31:0]       laneOfOffsetOfOffsetGroup = 32'h1 << offsetOfOffsetGroup[6:2];
  wire              indexedInstructionOffsetExhausted = offsetEEWOH[0] & (&(offsetOfOffsetGroup[1:0])) | offsetEEWOH[1] & offsetOfOffsetGroup[1] | offsetEEWOH[2];
  wire              _GEN = segmentEndWithHandshake & indexedInstructionOffsetExhausted;
  wire [1:0]        _GEN_0 = {waitQueueDeq_1, waitQueueDeq_0};
  wire [1:0]        usedIndexedInstructionOffsets_0_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_0_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_1_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_1_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_2_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_2_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_3_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_3_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_4_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_4_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_5_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_5_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_6_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_6_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_7_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_7_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_8_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_8_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_9_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_9_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_10_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_10_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_11_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_11_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_12_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_12_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_13_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_13_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_14_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_14_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_15_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_15_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_16_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_16_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_17_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_17_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_18_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_18_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_19_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_19_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_20_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_20_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_21_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_21_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_22_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_22_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_23_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_23_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_24_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_24_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_25_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_25_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_26_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_26_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_27_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_27_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_28_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_28_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_29_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_29_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_30_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_30_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        usedIndexedInstructionOffsets_31_lo_lo_lo_lo;
  assign usedIndexedInstructionOffsets_31_lo_lo_lo_lo = _GEN_0;
  wire [1:0]        _GEN_1 = {waitQueueDeq_3, waitQueueDeq_2};
  wire [1:0]        usedIndexedInstructionOffsets_0_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_0_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_1_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_1_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_2_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_2_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_3_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_3_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_4_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_4_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_5_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_5_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_6_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_6_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_7_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_7_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_8_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_8_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_9_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_9_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_10_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_10_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_11_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_11_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_12_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_12_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_13_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_13_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_14_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_14_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_15_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_15_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_16_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_16_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_17_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_17_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_18_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_18_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_19_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_19_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_20_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_20_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_21_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_21_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_22_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_22_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_23_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_23_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_24_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_24_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_25_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_25_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_26_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_26_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_27_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_27_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_28_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_28_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_29_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_29_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_30_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_30_lo_lo_lo_hi = _GEN_1;
  wire [1:0]        usedIndexedInstructionOffsets_31_lo_lo_lo_hi;
  assign usedIndexedInstructionOffsets_31_lo_lo_lo_hi = _GEN_1;
  wire [3:0]        usedIndexedInstructionOffsets_0_lo_lo_lo = {usedIndexedInstructionOffsets_0_lo_lo_lo_hi, usedIndexedInstructionOffsets_0_lo_lo_lo_lo};
  wire [1:0]        _GEN_2 = {waitQueueDeq_5, waitQueueDeq_4};
  wire [1:0]        usedIndexedInstructionOffsets_0_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_0_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_1_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_1_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_2_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_2_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_3_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_3_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_4_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_4_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_5_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_5_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_6_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_6_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_7_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_7_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_8_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_8_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_9_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_9_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_10_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_10_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_11_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_11_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_12_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_12_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_13_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_13_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_14_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_14_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_15_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_15_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_16_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_16_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_17_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_17_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_18_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_18_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_19_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_19_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_20_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_20_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_21_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_21_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_22_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_22_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_23_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_23_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_24_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_24_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_25_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_25_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_26_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_26_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_27_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_27_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_28_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_28_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_29_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_29_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_30_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_30_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        usedIndexedInstructionOffsets_31_lo_lo_hi_lo;
  assign usedIndexedInstructionOffsets_31_lo_lo_hi_lo = _GEN_2;
  wire [1:0]        _GEN_3 = {waitQueueDeq_7, waitQueueDeq_6};
  wire [1:0]        usedIndexedInstructionOffsets_0_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_0_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_1_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_1_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_2_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_2_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_3_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_3_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_4_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_4_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_5_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_5_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_6_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_6_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_7_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_7_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_8_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_8_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_9_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_9_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_10_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_10_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_11_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_11_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_12_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_12_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_13_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_13_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_14_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_14_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_15_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_15_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_16_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_16_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_17_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_17_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_18_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_18_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_19_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_19_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_20_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_20_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_21_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_21_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_22_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_22_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_23_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_23_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_24_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_24_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_25_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_25_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_26_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_26_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_27_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_27_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_28_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_28_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_29_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_29_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_30_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_30_lo_lo_hi_hi = _GEN_3;
  wire [1:0]        usedIndexedInstructionOffsets_31_lo_lo_hi_hi;
  assign usedIndexedInstructionOffsets_31_lo_lo_hi_hi = _GEN_3;
  wire [3:0]        usedIndexedInstructionOffsets_0_lo_lo_hi = {usedIndexedInstructionOffsets_0_lo_lo_hi_hi, usedIndexedInstructionOffsets_0_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_0_lo_lo = {usedIndexedInstructionOffsets_0_lo_lo_hi, usedIndexedInstructionOffsets_0_lo_lo_lo};
  wire [1:0]        _GEN_4 = {waitQueueDeq_9, waitQueueDeq_8};
  wire [1:0]        usedIndexedInstructionOffsets_0_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_0_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_1_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_1_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_2_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_2_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_3_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_3_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_4_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_4_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_5_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_5_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_6_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_6_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_7_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_7_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_8_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_8_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_9_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_9_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_10_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_10_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_11_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_11_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_12_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_12_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_13_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_13_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_14_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_14_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_15_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_15_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_16_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_16_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_17_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_17_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_18_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_18_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_19_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_19_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_20_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_20_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_21_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_21_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_22_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_22_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_23_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_23_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_24_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_24_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_25_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_25_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_26_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_26_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_27_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_27_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_28_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_28_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_29_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_29_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_30_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_30_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        usedIndexedInstructionOffsets_31_lo_hi_lo_lo;
  assign usedIndexedInstructionOffsets_31_lo_hi_lo_lo = _GEN_4;
  wire [1:0]        _GEN_5 = {waitQueueDeq_11, waitQueueDeq_10};
  wire [1:0]        usedIndexedInstructionOffsets_0_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_0_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_1_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_1_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_2_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_2_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_3_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_3_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_4_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_4_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_5_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_5_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_6_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_6_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_7_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_7_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_8_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_8_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_9_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_9_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_10_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_10_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_11_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_11_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_12_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_12_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_13_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_13_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_14_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_14_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_15_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_15_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_16_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_16_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_17_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_17_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_18_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_18_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_19_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_19_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_20_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_20_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_21_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_21_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_22_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_22_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_23_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_23_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_24_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_24_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_25_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_25_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_26_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_26_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_27_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_27_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_28_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_28_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_29_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_29_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_30_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_30_lo_hi_lo_hi = _GEN_5;
  wire [1:0]        usedIndexedInstructionOffsets_31_lo_hi_lo_hi;
  assign usedIndexedInstructionOffsets_31_lo_hi_lo_hi = _GEN_5;
  wire [3:0]        usedIndexedInstructionOffsets_0_lo_hi_lo = {usedIndexedInstructionOffsets_0_lo_hi_lo_hi, usedIndexedInstructionOffsets_0_lo_hi_lo_lo};
  wire [1:0]        _GEN_6 = {waitQueueDeq_13, waitQueueDeq_12};
  wire [1:0]        usedIndexedInstructionOffsets_0_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_0_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_1_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_1_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_2_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_2_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_3_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_3_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_4_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_4_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_5_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_5_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_6_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_6_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_7_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_7_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_8_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_8_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_9_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_9_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_10_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_10_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_11_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_11_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_12_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_12_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_13_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_13_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_14_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_14_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_15_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_15_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_16_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_16_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_17_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_17_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_18_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_18_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_19_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_19_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_20_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_20_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_21_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_21_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_22_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_22_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_23_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_23_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_24_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_24_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_25_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_25_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_26_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_26_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_27_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_27_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_28_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_28_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_29_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_29_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_30_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_30_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        usedIndexedInstructionOffsets_31_lo_hi_hi_lo;
  assign usedIndexedInstructionOffsets_31_lo_hi_hi_lo = _GEN_6;
  wire [1:0]        _GEN_7 = {waitQueueDeq_15, waitQueueDeq_14};
  wire [1:0]        usedIndexedInstructionOffsets_0_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_0_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_1_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_1_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_2_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_2_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_3_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_3_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_4_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_4_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_5_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_5_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_6_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_6_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_7_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_7_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_8_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_8_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_9_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_9_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_10_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_10_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_11_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_11_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_12_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_12_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_13_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_13_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_14_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_14_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_15_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_15_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_16_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_16_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_17_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_17_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_18_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_18_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_19_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_19_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_20_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_20_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_21_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_21_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_22_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_22_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_23_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_23_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_24_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_24_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_25_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_25_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_26_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_26_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_27_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_27_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_28_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_28_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_29_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_29_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_30_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_30_lo_hi_hi_hi = _GEN_7;
  wire [1:0]        usedIndexedInstructionOffsets_31_lo_hi_hi_hi;
  assign usedIndexedInstructionOffsets_31_lo_hi_hi_hi = _GEN_7;
  wire [3:0]        usedIndexedInstructionOffsets_0_lo_hi_hi = {usedIndexedInstructionOffsets_0_lo_hi_hi_hi, usedIndexedInstructionOffsets_0_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_0_lo_hi = {usedIndexedInstructionOffsets_0_lo_hi_hi, usedIndexedInstructionOffsets_0_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_0_lo = {usedIndexedInstructionOffsets_0_lo_hi, usedIndexedInstructionOffsets_0_lo_lo};
  wire [1:0]        _GEN_8 = {waitQueueDeq_17, waitQueueDeq_16};
  wire [1:0]        usedIndexedInstructionOffsets_0_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_0_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_1_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_1_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_2_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_2_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_3_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_3_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_4_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_4_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_5_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_5_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_6_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_6_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_7_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_7_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_8_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_8_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_9_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_9_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_10_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_10_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_11_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_11_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_12_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_12_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_13_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_13_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_14_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_14_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_15_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_15_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_16_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_16_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_17_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_17_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_18_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_18_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_19_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_19_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_20_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_20_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_21_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_21_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_22_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_22_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_23_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_23_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_24_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_24_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_25_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_25_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_26_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_26_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_27_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_27_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_28_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_28_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_29_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_29_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_30_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_30_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        usedIndexedInstructionOffsets_31_hi_lo_lo_lo;
  assign usedIndexedInstructionOffsets_31_hi_lo_lo_lo = _GEN_8;
  wire [1:0]        _GEN_9 = {waitQueueDeq_19, waitQueueDeq_18};
  wire [1:0]        usedIndexedInstructionOffsets_0_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_0_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_1_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_1_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_2_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_2_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_3_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_3_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_4_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_4_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_5_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_5_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_6_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_6_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_7_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_7_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_8_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_8_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_9_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_9_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_10_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_10_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_11_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_11_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_12_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_12_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_13_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_13_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_14_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_14_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_15_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_15_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_16_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_16_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_17_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_17_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_18_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_18_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_19_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_19_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_20_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_20_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_21_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_21_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_22_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_22_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_23_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_23_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_24_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_24_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_25_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_25_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_26_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_26_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_27_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_27_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_28_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_28_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_29_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_29_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_30_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_30_hi_lo_lo_hi = _GEN_9;
  wire [1:0]        usedIndexedInstructionOffsets_31_hi_lo_lo_hi;
  assign usedIndexedInstructionOffsets_31_hi_lo_lo_hi = _GEN_9;
  wire [3:0]        usedIndexedInstructionOffsets_0_hi_lo_lo = {usedIndexedInstructionOffsets_0_hi_lo_lo_hi, usedIndexedInstructionOffsets_0_hi_lo_lo_lo};
  wire [1:0]        _GEN_10 = {waitQueueDeq_21, waitQueueDeq_20};
  wire [1:0]        usedIndexedInstructionOffsets_0_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_0_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_1_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_1_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_2_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_2_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_3_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_3_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_4_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_4_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_5_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_5_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_6_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_6_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_7_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_7_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_8_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_8_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_9_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_9_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_10_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_10_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_11_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_11_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_12_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_12_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_13_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_13_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_14_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_14_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_15_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_15_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_16_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_16_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_17_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_17_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_18_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_18_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_19_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_19_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_20_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_20_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_21_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_21_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_22_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_22_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_23_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_23_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_24_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_24_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_25_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_25_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_26_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_26_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_27_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_27_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_28_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_28_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_29_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_29_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_30_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_30_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        usedIndexedInstructionOffsets_31_hi_lo_hi_lo;
  assign usedIndexedInstructionOffsets_31_hi_lo_hi_lo = _GEN_10;
  wire [1:0]        _GEN_11 = {waitQueueDeq_23, waitQueueDeq_22};
  wire [1:0]        usedIndexedInstructionOffsets_0_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_0_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_1_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_1_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_2_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_2_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_3_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_3_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_4_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_4_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_5_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_5_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_6_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_6_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_7_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_7_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_8_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_8_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_9_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_9_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_10_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_10_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_11_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_11_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_12_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_12_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_13_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_13_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_14_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_14_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_15_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_15_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_16_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_16_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_17_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_17_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_18_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_18_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_19_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_19_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_20_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_20_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_21_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_21_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_22_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_22_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_23_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_23_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_24_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_24_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_25_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_25_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_26_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_26_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_27_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_27_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_28_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_28_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_29_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_29_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_30_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_30_hi_lo_hi_hi = _GEN_11;
  wire [1:0]        usedIndexedInstructionOffsets_31_hi_lo_hi_hi;
  assign usedIndexedInstructionOffsets_31_hi_lo_hi_hi = _GEN_11;
  wire [3:0]        usedIndexedInstructionOffsets_0_hi_lo_hi = {usedIndexedInstructionOffsets_0_hi_lo_hi_hi, usedIndexedInstructionOffsets_0_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_0_hi_lo = {usedIndexedInstructionOffsets_0_hi_lo_hi, usedIndexedInstructionOffsets_0_hi_lo_lo};
  wire [1:0]        _GEN_12 = {waitQueueDeq_25, waitQueueDeq_24};
  wire [1:0]        usedIndexedInstructionOffsets_0_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_0_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_1_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_1_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_2_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_2_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_3_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_3_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_4_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_4_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_5_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_5_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_6_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_6_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_7_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_7_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_8_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_8_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_9_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_9_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_10_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_10_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_11_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_11_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_12_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_12_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_13_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_13_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_14_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_14_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_15_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_15_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_16_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_16_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_17_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_17_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_18_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_18_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_19_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_19_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_20_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_20_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_21_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_21_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_22_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_22_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_23_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_23_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_24_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_24_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_25_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_25_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_26_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_26_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_27_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_27_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_28_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_28_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_29_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_29_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_30_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_30_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        usedIndexedInstructionOffsets_31_hi_hi_lo_lo;
  assign usedIndexedInstructionOffsets_31_hi_hi_lo_lo = _GEN_12;
  wire [1:0]        _GEN_13 = {waitQueueDeq_27, waitQueueDeq_26};
  wire [1:0]        usedIndexedInstructionOffsets_0_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_0_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_1_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_1_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_2_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_2_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_3_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_3_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_4_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_4_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_5_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_5_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_6_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_6_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_7_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_7_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_8_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_8_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_9_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_9_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_10_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_10_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_11_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_11_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_12_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_12_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_13_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_13_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_14_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_14_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_15_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_15_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_16_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_16_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_17_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_17_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_18_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_18_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_19_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_19_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_20_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_20_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_21_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_21_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_22_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_22_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_23_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_23_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_24_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_24_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_25_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_25_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_26_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_26_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_27_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_27_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_28_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_28_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_29_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_29_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_30_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_30_hi_hi_lo_hi = _GEN_13;
  wire [1:0]        usedIndexedInstructionOffsets_31_hi_hi_lo_hi;
  assign usedIndexedInstructionOffsets_31_hi_hi_lo_hi = _GEN_13;
  wire [3:0]        usedIndexedInstructionOffsets_0_hi_hi_lo = {usedIndexedInstructionOffsets_0_hi_hi_lo_hi, usedIndexedInstructionOffsets_0_hi_hi_lo_lo};
  wire [1:0]        _GEN_14 = {waitQueueDeq_29, waitQueueDeq_28};
  wire [1:0]        usedIndexedInstructionOffsets_0_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_0_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_1_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_1_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_2_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_2_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_3_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_3_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_4_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_4_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_5_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_5_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_6_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_6_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_7_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_7_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_8_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_8_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_9_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_9_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_10_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_10_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_11_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_11_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_12_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_12_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_13_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_13_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_14_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_14_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_15_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_15_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_16_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_16_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_17_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_17_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_18_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_18_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_19_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_19_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_20_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_20_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_21_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_21_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_22_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_22_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_23_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_23_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_24_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_24_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_25_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_25_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_26_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_26_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_27_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_27_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_28_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_28_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_29_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_29_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_30_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_30_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        usedIndexedInstructionOffsets_31_hi_hi_hi_lo;
  assign usedIndexedInstructionOffsets_31_hi_hi_hi_lo = _GEN_14;
  wire [1:0]        _GEN_15 = {waitQueueDeq_31, waitQueueDeq_30};
  wire [1:0]        usedIndexedInstructionOffsets_0_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_0_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_1_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_1_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_2_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_2_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_3_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_3_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_4_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_4_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_5_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_5_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_6_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_6_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_7_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_7_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_8_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_8_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_9_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_9_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_10_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_10_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_11_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_11_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_12_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_12_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_13_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_13_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_14_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_14_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_15_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_15_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_16_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_16_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_17_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_17_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_18_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_18_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_19_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_19_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_20_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_20_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_21_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_21_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_22_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_22_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_23_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_23_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_24_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_24_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_25_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_25_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_26_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_26_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_27_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_27_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_28_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_28_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_29_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_29_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_30_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_30_hi_hi_hi_hi = _GEN_15;
  wire [1:0]        usedIndexedInstructionOffsets_31_hi_hi_hi_hi;
  assign usedIndexedInstructionOffsets_31_hi_hi_hi_hi = _GEN_15;
  wire [3:0]        usedIndexedInstructionOffsets_0_hi_hi_hi = {usedIndexedInstructionOffsets_0_hi_hi_hi_hi, usedIndexedInstructionOffsets_0_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_0_hi_hi = {usedIndexedInstructionOffsets_0_hi_hi_hi, usedIndexedInstructionOffsets_0_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_0_hi = {usedIndexedInstructionOffsets_0_hi_hi, usedIndexedInstructionOffsets_0_hi_lo};
  wire              requestOffset;
  wire              usedIndexedInstructionOffsets_0 = laneOfOffsetOfOffsetGroup[0] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_0_hi, usedIndexedInstructionOffsets_0_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_1_lo_lo_lo = {usedIndexedInstructionOffsets_1_lo_lo_lo_hi, usedIndexedInstructionOffsets_1_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_1_lo_lo_hi = {usedIndexedInstructionOffsets_1_lo_lo_hi_hi, usedIndexedInstructionOffsets_1_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_1_lo_lo = {usedIndexedInstructionOffsets_1_lo_lo_hi, usedIndexedInstructionOffsets_1_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_1_lo_hi_lo = {usedIndexedInstructionOffsets_1_lo_hi_lo_hi, usedIndexedInstructionOffsets_1_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_1_lo_hi_hi = {usedIndexedInstructionOffsets_1_lo_hi_hi_hi, usedIndexedInstructionOffsets_1_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_1_lo_hi = {usedIndexedInstructionOffsets_1_lo_hi_hi, usedIndexedInstructionOffsets_1_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_1_lo = {usedIndexedInstructionOffsets_1_lo_hi, usedIndexedInstructionOffsets_1_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_1_hi_lo_lo = {usedIndexedInstructionOffsets_1_hi_lo_lo_hi, usedIndexedInstructionOffsets_1_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_1_hi_lo_hi = {usedIndexedInstructionOffsets_1_hi_lo_hi_hi, usedIndexedInstructionOffsets_1_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_1_hi_lo = {usedIndexedInstructionOffsets_1_hi_lo_hi, usedIndexedInstructionOffsets_1_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_1_hi_hi_lo = {usedIndexedInstructionOffsets_1_hi_hi_lo_hi, usedIndexedInstructionOffsets_1_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_1_hi_hi_hi = {usedIndexedInstructionOffsets_1_hi_hi_hi_hi, usedIndexedInstructionOffsets_1_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_1_hi_hi = {usedIndexedInstructionOffsets_1_hi_hi_hi, usedIndexedInstructionOffsets_1_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_1_hi = {usedIndexedInstructionOffsets_1_hi_hi, usedIndexedInstructionOffsets_1_hi_lo};
  wire              usedIndexedInstructionOffsets_1 = laneOfOffsetOfOffsetGroup[1] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_1_hi, usedIndexedInstructionOffsets_1_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_2_lo_lo_lo = {usedIndexedInstructionOffsets_2_lo_lo_lo_hi, usedIndexedInstructionOffsets_2_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_2_lo_lo_hi = {usedIndexedInstructionOffsets_2_lo_lo_hi_hi, usedIndexedInstructionOffsets_2_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_2_lo_lo = {usedIndexedInstructionOffsets_2_lo_lo_hi, usedIndexedInstructionOffsets_2_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_2_lo_hi_lo = {usedIndexedInstructionOffsets_2_lo_hi_lo_hi, usedIndexedInstructionOffsets_2_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_2_lo_hi_hi = {usedIndexedInstructionOffsets_2_lo_hi_hi_hi, usedIndexedInstructionOffsets_2_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_2_lo_hi = {usedIndexedInstructionOffsets_2_lo_hi_hi, usedIndexedInstructionOffsets_2_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_2_lo = {usedIndexedInstructionOffsets_2_lo_hi, usedIndexedInstructionOffsets_2_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_2_hi_lo_lo = {usedIndexedInstructionOffsets_2_hi_lo_lo_hi, usedIndexedInstructionOffsets_2_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_2_hi_lo_hi = {usedIndexedInstructionOffsets_2_hi_lo_hi_hi, usedIndexedInstructionOffsets_2_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_2_hi_lo = {usedIndexedInstructionOffsets_2_hi_lo_hi, usedIndexedInstructionOffsets_2_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_2_hi_hi_lo = {usedIndexedInstructionOffsets_2_hi_hi_lo_hi, usedIndexedInstructionOffsets_2_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_2_hi_hi_hi = {usedIndexedInstructionOffsets_2_hi_hi_hi_hi, usedIndexedInstructionOffsets_2_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_2_hi_hi = {usedIndexedInstructionOffsets_2_hi_hi_hi, usedIndexedInstructionOffsets_2_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_2_hi = {usedIndexedInstructionOffsets_2_hi_hi, usedIndexedInstructionOffsets_2_hi_lo};
  wire              usedIndexedInstructionOffsets_2 = laneOfOffsetOfOffsetGroup[2] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_2_hi, usedIndexedInstructionOffsets_2_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_3_lo_lo_lo = {usedIndexedInstructionOffsets_3_lo_lo_lo_hi, usedIndexedInstructionOffsets_3_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_3_lo_lo_hi = {usedIndexedInstructionOffsets_3_lo_lo_hi_hi, usedIndexedInstructionOffsets_3_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_3_lo_lo = {usedIndexedInstructionOffsets_3_lo_lo_hi, usedIndexedInstructionOffsets_3_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_3_lo_hi_lo = {usedIndexedInstructionOffsets_3_lo_hi_lo_hi, usedIndexedInstructionOffsets_3_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_3_lo_hi_hi = {usedIndexedInstructionOffsets_3_lo_hi_hi_hi, usedIndexedInstructionOffsets_3_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_3_lo_hi = {usedIndexedInstructionOffsets_3_lo_hi_hi, usedIndexedInstructionOffsets_3_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_3_lo = {usedIndexedInstructionOffsets_3_lo_hi, usedIndexedInstructionOffsets_3_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_3_hi_lo_lo = {usedIndexedInstructionOffsets_3_hi_lo_lo_hi, usedIndexedInstructionOffsets_3_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_3_hi_lo_hi = {usedIndexedInstructionOffsets_3_hi_lo_hi_hi, usedIndexedInstructionOffsets_3_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_3_hi_lo = {usedIndexedInstructionOffsets_3_hi_lo_hi, usedIndexedInstructionOffsets_3_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_3_hi_hi_lo = {usedIndexedInstructionOffsets_3_hi_hi_lo_hi, usedIndexedInstructionOffsets_3_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_3_hi_hi_hi = {usedIndexedInstructionOffsets_3_hi_hi_hi_hi, usedIndexedInstructionOffsets_3_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_3_hi_hi = {usedIndexedInstructionOffsets_3_hi_hi_hi, usedIndexedInstructionOffsets_3_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_3_hi = {usedIndexedInstructionOffsets_3_hi_hi, usedIndexedInstructionOffsets_3_hi_lo};
  wire              usedIndexedInstructionOffsets_3 = laneOfOffsetOfOffsetGroup[3] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_3_hi, usedIndexedInstructionOffsets_3_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_4_lo_lo_lo = {usedIndexedInstructionOffsets_4_lo_lo_lo_hi, usedIndexedInstructionOffsets_4_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_4_lo_lo_hi = {usedIndexedInstructionOffsets_4_lo_lo_hi_hi, usedIndexedInstructionOffsets_4_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_4_lo_lo = {usedIndexedInstructionOffsets_4_lo_lo_hi, usedIndexedInstructionOffsets_4_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_4_lo_hi_lo = {usedIndexedInstructionOffsets_4_lo_hi_lo_hi, usedIndexedInstructionOffsets_4_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_4_lo_hi_hi = {usedIndexedInstructionOffsets_4_lo_hi_hi_hi, usedIndexedInstructionOffsets_4_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_4_lo_hi = {usedIndexedInstructionOffsets_4_lo_hi_hi, usedIndexedInstructionOffsets_4_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_4_lo = {usedIndexedInstructionOffsets_4_lo_hi, usedIndexedInstructionOffsets_4_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_4_hi_lo_lo = {usedIndexedInstructionOffsets_4_hi_lo_lo_hi, usedIndexedInstructionOffsets_4_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_4_hi_lo_hi = {usedIndexedInstructionOffsets_4_hi_lo_hi_hi, usedIndexedInstructionOffsets_4_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_4_hi_lo = {usedIndexedInstructionOffsets_4_hi_lo_hi, usedIndexedInstructionOffsets_4_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_4_hi_hi_lo = {usedIndexedInstructionOffsets_4_hi_hi_lo_hi, usedIndexedInstructionOffsets_4_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_4_hi_hi_hi = {usedIndexedInstructionOffsets_4_hi_hi_hi_hi, usedIndexedInstructionOffsets_4_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_4_hi_hi = {usedIndexedInstructionOffsets_4_hi_hi_hi, usedIndexedInstructionOffsets_4_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_4_hi = {usedIndexedInstructionOffsets_4_hi_hi, usedIndexedInstructionOffsets_4_hi_lo};
  wire              usedIndexedInstructionOffsets_4 = laneOfOffsetOfOffsetGroup[4] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_4_hi, usedIndexedInstructionOffsets_4_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_5_lo_lo_lo = {usedIndexedInstructionOffsets_5_lo_lo_lo_hi, usedIndexedInstructionOffsets_5_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_5_lo_lo_hi = {usedIndexedInstructionOffsets_5_lo_lo_hi_hi, usedIndexedInstructionOffsets_5_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_5_lo_lo = {usedIndexedInstructionOffsets_5_lo_lo_hi, usedIndexedInstructionOffsets_5_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_5_lo_hi_lo = {usedIndexedInstructionOffsets_5_lo_hi_lo_hi, usedIndexedInstructionOffsets_5_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_5_lo_hi_hi = {usedIndexedInstructionOffsets_5_lo_hi_hi_hi, usedIndexedInstructionOffsets_5_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_5_lo_hi = {usedIndexedInstructionOffsets_5_lo_hi_hi, usedIndexedInstructionOffsets_5_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_5_lo = {usedIndexedInstructionOffsets_5_lo_hi, usedIndexedInstructionOffsets_5_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_5_hi_lo_lo = {usedIndexedInstructionOffsets_5_hi_lo_lo_hi, usedIndexedInstructionOffsets_5_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_5_hi_lo_hi = {usedIndexedInstructionOffsets_5_hi_lo_hi_hi, usedIndexedInstructionOffsets_5_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_5_hi_lo = {usedIndexedInstructionOffsets_5_hi_lo_hi, usedIndexedInstructionOffsets_5_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_5_hi_hi_lo = {usedIndexedInstructionOffsets_5_hi_hi_lo_hi, usedIndexedInstructionOffsets_5_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_5_hi_hi_hi = {usedIndexedInstructionOffsets_5_hi_hi_hi_hi, usedIndexedInstructionOffsets_5_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_5_hi_hi = {usedIndexedInstructionOffsets_5_hi_hi_hi, usedIndexedInstructionOffsets_5_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_5_hi = {usedIndexedInstructionOffsets_5_hi_hi, usedIndexedInstructionOffsets_5_hi_lo};
  wire              usedIndexedInstructionOffsets_5 = laneOfOffsetOfOffsetGroup[5] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_5_hi, usedIndexedInstructionOffsets_5_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_6_lo_lo_lo = {usedIndexedInstructionOffsets_6_lo_lo_lo_hi, usedIndexedInstructionOffsets_6_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_6_lo_lo_hi = {usedIndexedInstructionOffsets_6_lo_lo_hi_hi, usedIndexedInstructionOffsets_6_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_6_lo_lo = {usedIndexedInstructionOffsets_6_lo_lo_hi, usedIndexedInstructionOffsets_6_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_6_lo_hi_lo = {usedIndexedInstructionOffsets_6_lo_hi_lo_hi, usedIndexedInstructionOffsets_6_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_6_lo_hi_hi = {usedIndexedInstructionOffsets_6_lo_hi_hi_hi, usedIndexedInstructionOffsets_6_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_6_lo_hi = {usedIndexedInstructionOffsets_6_lo_hi_hi, usedIndexedInstructionOffsets_6_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_6_lo = {usedIndexedInstructionOffsets_6_lo_hi, usedIndexedInstructionOffsets_6_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_6_hi_lo_lo = {usedIndexedInstructionOffsets_6_hi_lo_lo_hi, usedIndexedInstructionOffsets_6_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_6_hi_lo_hi = {usedIndexedInstructionOffsets_6_hi_lo_hi_hi, usedIndexedInstructionOffsets_6_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_6_hi_lo = {usedIndexedInstructionOffsets_6_hi_lo_hi, usedIndexedInstructionOffsets_6_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_6_hi_hi_lo = {usedIndexedInstructionOffsets_6_hi_hi_lo_hi, usedIndexedInstructionOffsets_6_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_6_hi_hi_hi = {usedIndexedInstructionOffsets_6_hi_hi_hi_hi, usedIndexedInstructionOffsets_6_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_6_hi_hi = {usedIndexedInstructionOffsets_6_hi_hi_hi, usedIndexedInstructionOffsets_6_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_6_hi = {usedIndexedInstructionOffsets_6_hi_hi, usedIndexedInstructionOffsets_6_hi_lo};
  wire              usedIndexedInstructionOffsets_6 = laneOfOffsetOfOffsetGroup[6] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_6_hi, usedIndexedInstructionOffsets_6_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_7_lo_lo_lo = {usedIndexedInstructionOffsets_7_lo_lo_lo_hi, usedIndexedInstructionOffsets_7_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_7_lo_lo_hi = {usedIndexedInstructionOffsets_7_lo_lo_hi_hi, usedIndexedInstructionOffsets_7_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_7_lo_lo = {usedIndexedInstructionOffsets_7_lo_lo_hi, usedIndexedInstructionOffsets_7_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_7_lo_hi_lo = {usedIndexedInstructionOffsets_7_lo_hi_lo_hi, usedIndexedInstructionOffsets_7_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_7_lo_hi_hi = {usedIndexedInstructionOffsets_7_lo_hi_hi_hi, usedIndexedInstructionOffsets_7_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_7_lo_hi = {usedIndexedInstructionOffsets_7_lo_hi_hi, usedIndexedInstructionOffsets_7_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_7_lo = {usedIndexedInstructionOffsets_7_lo_hi, usedIndexedInstructionOffsets_7_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_7_hi_lo_lo = {usedIndexedInstructionOffsets_7_hi_lo_lo_hi, usedIndexedInstructionOffsets_7_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_7_hi_lo_hi = {usedIndexedInstructionOffsets_7_hi_lo_hi_hi, usedIndexedInstructionOffsets_7_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_7_hi_lo = {usedIndexedInstructionOffsets_7_hi_lo_hi, usedIndexedInstructionOffsets_7_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_7_hi_hi_lo = {usedIndexedInstructionOffsets_7_hi_hi_lo_hi, usedIndexedInstructionOffsets_7_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_7_hi_hi_hi = {usedIndexedInstructionOffsets_7_hi_hi_hi_hi, usedIndexedInstructionOffsets_7_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_7_hi_hi = {usedIndexedInstructionOffsets_7_hi_hi_hi, usedIndexedInstructionOffsets_7_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_7_hi = {usedIndexedInstructionOffsets_7_hi_hi, usedIndexedInstructionOffsets_7_hi_lo};
  wire              usedIndexedInstructionOffsets_7 = laneOfOffsetOfOffsetGroup[7] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_7_hi, usedIndexedInstructionOffsets_7_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_8_lo_lo_lo = {usedIndexedInstructionOffsets_8_lo_lo_lo_hi, usedIndexedInstructionOffsets_8_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_8_lo_lo_hi = {usedIndexedInstructionOffsets_8_lo_lo_hi_hi, usedIndexedInstructionOffsets_8_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_8_lo_lo = {usedIndexedInstructionOffsets_8_lo_lo_hi, usedIndexedInstructionOffsets_8_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_8_lo_hi_lo = {usedIndexedInstructionOffsets_8_lo_hi_lo_hi, usedIndexedInstructionOffsets_8_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_8_lo_hi_hi = {usedIndexedInstructionOffsets_8_lo_hi_hi_hi, usedIndexedInstructionOffsets_8_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_8_lo_hi = {usedIndexedInstructionOffsets_8_lo_hi_hi, usedIndexedInstructionOffsets_8_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_8_lo = {usedIndexedInstructionOffsets_8_lo_hi, usedIndexedInstructionOffsets_8_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_8_hi_lo_lo = {usedIndexedInstructionOffsets_8_hi_lo_lo_hi, usedIndexedInstructionOffsets_8_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_8_hi_lo_hi = {usedIndexedInstructionOffsets_8_hi_lo_hi_hi, usedIndexedInstructionOffsets_8_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_8_hi_lo = {usedIndexedInstructionOffsets_8_hi_lo_hi, usedIndexedInstructionOffsets_8_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_8_hi_hi_lo = {usedIndexedInstructionOffsets_8_hi_hi_lo_hi, usedIndexedInstructionOffsets_8_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_8_hi_hi_hi = {usedIndexedInstructionOffsets_8_hi_hi_hi_hi, usedIndexedInstructionOffsets_8_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_8_hi_hi = {usedIndexedInstructionOffsets_8_hi_hi_hi, usedIndexedInstructionOffsets_8_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_8_hi = {usedIndexedInstructionOffsets_8_hi_hi, usedIndexedInstructionOffsets_8_hi_lo};
  wire              usedIndexedInstructionOffsets_8 = laneOfOffsetOfOffsetGroup[8] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_8_hi, usedIndexedInstructionOffsets_8_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_9_lo_lo_lo = {usedIndexedInstructionOffsets_9_lo_lo_lo_hi, usedIndexedInstructionOffsets_9_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_9_lo_lo_hi = {usedIndexedInstructionOffsets_9_lo_lo_hi_hi, usedIndexedInstructionOffsets_9_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_9_lo_lo = {usedIndexedInstructionOffsets_9_lo_lo_hi, usedIndexedInstructionOffsets_9_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_9_lo_hi_lo = {usedIndexedInstructionOffsets_9_lo_hi_lo_hi, usedIndexedInstructionOffsets_9_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_9_lo_hi_hi = {usedIndexedInstructionOffsets_9_lo_hi_hi_hi, usedIndexedInstructionOffsets_9_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_9_lo_hi = {usedIndexedInstructionOffsets_9_lo_hi_hi, usedIndexedInstructionOffsets_9_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_9_lo = {usedIndexedInstructionOffsets_9_lo_hi, usedIndexedInstructionOffsets_9_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_9_hi_lo_lo = {usedIndexedInstructionOffsets_9_hi_lo_lo_hi, usedIndexedInstructionOffsets_9_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_9_hi_lo_hi = {usedIndexedInstructionOffsets_9_hi_lo_hi_hi, usedIndexedInstructionOffsets_9_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_9_hi_lo = {usedIndexedInstructionOffsets_9_hi_lo_hi, usedIndexedInstructionOffsets_9_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_9_hi_hi_lo = {usedIndexedInstructionOffsets_9_hi_hi_lo_hi, usedIndexedInstructionOffsets_9_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_9_hi_hi_hi = {usedIndexedInstructionOffsets_9_hi_hi_hi_hi, usedIndexedInstructionOffsets_9_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_9_hi_hi = {usedIndexedInstructionOffsets_9_hi_hi_hi, usedIndexedInstructionOffsets_9_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_9_hi = {usedIndexedInstructionOffsets_9_hi_hi, usedIndexedInstructionOffsets_9_hi_lo};
  wire              usedIndexedInstructionOffsets_9 = laneOfOffsetOfOffsetGroup[9] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_9_hi, usedIndexedInstructionOffsets_9_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_10_lo_lo_lo = {usedIndexedInstructionOffsets_10_lo_lo_lo_hi, usedIndexedInstructionOffsets_10_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_10_lo_lo_hi = {usedIndexedInstructionOffsets_10_lo_lo_hi_hi, usedIndexedInstructionOffsets_10_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_10_lo_lo = {usedIndexedInstructionOffsets_10_lo_lo_hi, usedIndexedInstructionOffsets_10_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_10_lo_hi_lo = {usedIndexedInstructionOffsets_10_lo_hi_lo_hi, usedIndexedInstructionOffsets_10_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_10_lo_hi_hi = {usedIndexedInstructionOffsets_10_lo_hi_hi_hi, usedIndexedInstructionOffsets_10_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_10_lo_hi = {usedIndexedInstructionOffsets_10_lo_hi_hi, usedIndexedInstructionOffsets_10_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_10_lo = {usedIndexedInstructionOffsets_10_lo_hi, usedIndexedInstructionOffsets_10_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_10_hi_lo_lo = {usedIndexedInstructionOffsets_10_hi_lo_lo_hi, usedIndexedInstructionOffsets_10_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_10_hi_lo_hi = {usedIndexedInstructionOffsets_10_hi_lo_hi_hi, usedIndexedInstructionOffsets_10_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_10_hi_lo = {usedIndexedInstructionOffsets_10_hi_lo_hi, usedIndexedInstructionOffsets_10_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_10_hi_hi_lo = {usedIndexedInstructionOffsets_10_hi_hi_lo_hi, usedIndexedInstructionOffsets_10_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_10_hi_hi_hi = {usedIndexedInstructionOffsets_10_hi_hi_hi_hi, usedIndexedInstructionOffsets_10_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_10_hi_hi = {usedIndexedInstructionOffsets_10_hi_hi_hi, usedIndexedInstructionOffsets_10_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_10_hi = {usedIndexedInstructionOffsets_10_hi_hi, usedIndexedInstructionOffsets_10_hi_lo};
  wire              usedIndexedInstructionOffsets_10 = laneOfOffsetOfOffsetGroup[10] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_10_hi, usedIndexedInstructionOffsets_10_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_11_lo_lo_lo = {usedIndexedInstructionOffsets_11_lo_lo_lo_hi, usedIndexedInstructionOffsets_11_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_11_lo_lo_hi = {usedIndexedInstructionOffsets_11_lo_lo_hi_hi, usedIndexedInstructionOffsets_11_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_11_lo_lo = {usedIndexedInstructionOffsets_11_lo_lo_hi, usedIndexedInstructionOffsets_11_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_11_lo_hi_lo = {usedIndexedInstructionOffsets_11_lo_hi_lo_hi, usedIndexedInstructionOffsets_11_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_11_lo_hi_hi = {usedIndexedInstructionOffsets_11_lo_hi_hi_hi, usedIndexedInstructionOffsets_11_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_11_lo_hi = {usedIndexedInstructionOffsets_11_lo_hi_hi, usedIndexedInstructionOffsets_11_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_11_lo = {usedIndexedInstructionOffsets_11_lo_hi, usedIndexedInstructionOffsets_11_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_11_hi_lo_lo = {usedIndexedInstructionOffsets_11_hi_lo_lo_hi, usedIndexedInstructionOffsets_11_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_11_hi_lo_hi = {usedIndexedInstructionOffsets_11_hi_lo_hi_hi, usedIndexedInstructionOffsets_11_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_11_hi_lo = {usedIndexedInstructionOffsets_11_hi_lo_hi, usedIndexedInstructionOffsets_11_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_11_hi_hi_lo = {usedIndexedInstructionOffsets_11_hi_hi_lo_hi, usedIndexedInstructionOffsets_11_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_11_hi_hi_hi = {usedIndexedInstructionOffsets_11_hi_hi_hi_hi, usedIndexedInstructionOffsets_11_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_11_hi_hi = {usedIndexedInstructionOffsets_11_hi_hi_hi, usedIndexedInstructionOffsets_11_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_11_hi = {usedIndexedInstructionOffsets_11_hi_hi, usedIndexedInstructionOffsets_11_hi_lo};
  wire              usedIndexedInstructionOffsets_11 = laneOfOffsetOfOffsetGroup[11] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_11_hi, usedIndexedInstructionOffsets_11_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_12_lo_lo_lo = {usedIndexedInstructionOffsets_12_lo_lo_lo_hi, usedIndexedInstructionOffsets_12_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_12_lo_lo_hi = {usedIndexedInstructionOffsets_12_lo_lo_hi_hi, usedIndexedInstructionOffsets_12_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_12_lo_lo = {usedIndexedInstructionOffsets_12_lo_lo_hi, usedIndexedInstructionOffsets_12_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_12_lo_hi_lo = {usedIndexedInstructionOffsets_12_lo_hi_lo_hi, usedIndexedInstructionOffsets_12_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_12_lo_hi_hi = {usedIndexedInstructionOffsets_12_lo_hi_hi_hi, usedIndexedInstructionOffsets_12_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_12_lo_hi = {usedIndexedInstructionOffsets_12_lo_hi_hi, usedIndexedInstructionOffsets_12_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_12_lo = {usedIndexedInstructionOffsets_12_lo_hi, usedIndexedInstructionOffsets_12_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_12_hi_lo_lo = {usedIndexedInstructionOffsets_12_hi_lo_lo_hi, usedIndexedInstructionOffsets_12_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_12_hi_lo_hi = {usedIndexedInstructionOffsets_12_hi_lo_hi_hi, usedIndexedInstructionOffsets_12_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_12_hi_lo = {usedIndexedInstructionOffsets_12_hi_lo_hi, usedIndexedInstructionOffsets_12_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_12_hi_hi_lo = {usedIndexedInstructionOffsets_12_hi_hi_lo_hi, usedIndexedInstructionOffsets_12_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_12_hi_hi_hi = {usedIndexedInstructionOffsets_12_hi_hi_hi_hi, usedIndexedInstructionOffsets_12_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_12_hi_hi = {usedIndexedInstructionOffsets_12_hi_hi_hi, usedIndexedInstructionOffsets_12_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_12_hi = {usedIndexedInstructionOffsets_12_hi_hi, usedIndexedInstructionOffsets_12_hi_lo};
  wire              usedIndexedInstructionOffsets_12 = laneOfOffsetOfOffsetGroup[12] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_12_hi, usedIndexedInstructionOffsets_12_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_13_lo_lo_lo = {usedIndexedInstructionOffsets_13_lo_lo_lo_hi, usedIndexedInstructionOffsets_13_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_13_lo_lo_hi = {usedIndexedInstructionOffsets_13_lo_lo_hi_hi, usedIndexedInstructionOffsets_13_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_13_lo_lo = {usedIndexedInstructionOffsets_13_lo_lo_hi, usedIndexedInstructionOffsets_13_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_13_lo_hi_lo = {usedIndexedInstructionOffsets_13_lo_hi_lo_hi, usedIndexedInstructionOffsets_13_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_13_lo_hi_hi = {usedIndexedInstructionOffsets_13_lo_hi_hi_hi, usedIndexedInstructionOffsets_13_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_13_lo_hi = {usedIndexedInstructionOffsets_13_lo_hi_hi, usedIndexedInstructionOffsets_13_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_13_lo = {usedIndexedInstructionOffsets_13_lo_hi, usedIndexedInstructionOffsets_13_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_13_hi_lo_lo = {usedIndexedInstructionOffsets_13_hi_lo_lo_hi, usedIndexedInstructionOffsets_13_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_13_hi_lo_hi = {usedIndexedInstructionOffsets_13_hi_lo_hi_hi, usedIndexedInstructionOffsets_13_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_13_hi_lo = {usedIndexedInstructionOffsets_13_hi_lo_hi, usedIndexedInstructionOffsets_13_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_13_hi_hi_lo = {usedIndexedInstructionOffsets_13_hi_hi_lo_hi, usedIndexedInstructionOffsets_13_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_13_hi_hi_hi = {usedIndexedInstructionOffsets_13_hi_hi_hi_hi, usedIndexedInstructionOffsets_13_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_13_hi_hi = {usedIndexedInstructionOffsets_13_hi_hi_hi, usedIndexedInstructionOffsets_13_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_13_hi = {usedIndexedInstructionOffsets_13_hi_hi, usedIndexedInstructionOffsets_13_hi_lo};
  wire              usedIndexedInstructionOffsets_13 = laneOfOffsetOfOffsetGroup[13] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_13_hi, usedIndexedInstructionOffsets_13_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_14_lo_lo_lo = {usedIndexedInstructionOffsets_14_lo_lo_lo_hi, usedIndexedInstructionOffsets_14_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_14_lo_lo_hi = {usedIndexedInstructionOffsets_14_lo_lo_hi_hi, usedIndexedInstructionOffsets_14_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_14_lo_lo = {usedIndexedInstructionOffsets_14_lo_lo_hi, usedIndexedInstructionOffsets_14_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_14_lo_hi_lo = {usedIndexedInstructionOffsets_14_lo_hi_lo_hi, usedIndexedInstructionOffsets_14_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_14_lo_hi_hi = {usedIndexedInstructionOffsets_14_lo_hi_hi_hi, usedIndexedInstructionOffsets_14_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_14_lo_hi = {usedIndexedInstructionOffsets_14_lo_hi_hi, usedIndexedInstructionOffsets_14_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_14_lo = {usedIndexedInstructionOffsets_14_lo_hi, usedIndexedInstructionOffsets_14_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_14_hi_lo_lo = {usedIndexedInstructionOffsets_14_hi_lo_lo_hi, usedIndexedInstructionOffsets_14_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_14_hi_lo_hi = {usedIndexedInstructionOffsets_14_hi_lo_hi_hi, usedIndexedInstructionOffsets_14_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_14_hi_lo = {usedIndexedInstructionOffsets_14_hi_lo_hi, usedIndexedInstructionOffsets_14_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_14_hi_hi_lo = {usedIndexedInstructionOffsets_14_hi_hi_lo_hi, usedIndexedInstructionOffsets_14_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_14_hi_hi_hi = {usedIndexedInstructionOffsets_14_hi_hi_hi_hi, usedIndexedInstructionOffsets_14_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_14_hi_hi = {usedIndexedInstructionOffsets_14_hi_hi_hi, usedIndexedInstructionOffsets_14_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_14_hi = {usedIndexedInstructionOffsets_14_hi_hi, usedIndexedInstructionOffsets_14_hi_lo};
  wire              usedIndexedInstructionOffsets_14 = laneOfOffsetOfOffsetGroup[14] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_14_hi, usedIndexedInstructionOffsets_14_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_15_lo_lo_lo = {usedIndexedInstructionOffsets_15_lo_lo_lo_hi, usedIndexedInstructionOffsets_15_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_15_lo_lo_hi = {usedIndexedInstructionOffsets_15_lo_lo_hi_hi, usedIndexedInstructionOffsets_15_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_15_lo_lo = {usedIndexedInstructionOffsets_15_lo_lo_hi, usedIndexedInstructionOffsets_15_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_15_lo_hi_lo = {usedIndexedInstructionOffsets_15_lo_hi_lo_hi, usedIndexedInstructionOffsets_15_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_15_lo_hi_hi = {usedIndexedInstructionOffsets_15_lo_hi_hi_hi, usedIndexedInstructionOffsets_15_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_15_lo_hi = {usedIndexedInstructionOffsets_15_lo_hi_hi, usedIndexedInstructionOffsets_15_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_15_lo = {usedIndexedInstructionOffsets_15_lo_hi, usedIndexedInstructionOffsets_15_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_15_hi_lo_lo = {usedIndexedInstructionOffsets_15_hi_lo_lo_hi, usedIndexedInstructionOffsets_15_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_15_hi_lo_hi = {usedIndexedInstructionOffsets_15_hi_lo_hi_hi, usedIndexedInstructionOffsets_15_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_15_hi_lo = {usedIndexedInstructionOffsets_15_hi_lo_hi, usedIndexedInstructionOffsets_15_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_15_hi_hi_lo = {usedIndexedInstructionOffsets_15_hi_hi_lo_hi, usedIndexedInstructionOffsets_15_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_15_hi_hi_hi = {usedIndexedInstructionOffsets_15_hi_hi_hi_hi, usedIndexedInstructionOffsets_15_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_15_hi_hi = {usedIndexedInstructionOffsets_15_hi_hi_hi, usedIndexedInstructionOffsets_15_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_15_hi = {usedIndexedInstructionOffsets_15_hi_hi, usedIndexedInstructionOffsets_15_hi_lo};
  wire              usedIndexedInstructionOffsets_15 = laneOfOffsetOfOffsetGroup[15] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_15_hi, usedIndexedInstructionOffsets_15_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_16_lo_lo_lo = {usedIndexedInstructionOffsets_16_lo_lo_lo_hi, usedIndexedInstructionOffsets_16_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_16_lo_lo_hi = {usedIndexedInstructionOffsets_16_lo_lo_hi_hi, usedIndexedInstructionOffsets_16_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_16_lo_lo = {usedIndexedInstructionOffsets_16_lo_lo_hi, usedIndexedInstructionOffsets_16_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_16_lo_hi_lo = {usedIndexedInstructionOffsets_16_lo_hi_lo_hi, usedIndexedInstructionOffsets_16_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_16_lo_hi_hi = {usedIndexedInstructionOffsets_16_lo_hi_hi_hi, usedIndexedInstructionOffsets_16_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_16_lo_hi = {usedIndexedInstructionOffsets_16_lo_hi_hi, usedIndexedInstructionOffsets_16_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_16_lo = {usedIndexedInstructionOffsets_16_lo_hi, usedIndexedInstructionOffsets_16_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_16_hi_lo_lo = {usedIndexedInstructionOffsets_16_hi_lo_lo_hi, usedIndexedInstructionOffsets_16_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_16_hi_lo_hi = {usedIndexedInstructionOffsets_16_hi_lo_hi_hi, usedIndexedInstructionOffsets_16_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_16_hi_lo = {usedIndexedInstructionOffsets_16_hi_lo_hi, usedIndexedInstructionOffsets_16_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_16_hi_hi_lo = {usedIndexedInstructionOffsets_16_hi_hi_lo_hi, usedIndexedInstructionOffsets_16_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_16_hi_hi_hi = {usedIndexedInstructionOffsets_16_hi_hi_hi_hi, usedIndexedInstructionOffsets_16_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_16_hi_hi = {usedIndexedInstructionOffsets_16_hi_hi_hi, usedIndexedInstructionOffsets_16_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_16_hi = {usedIndexedInstructionOffsets_16_hi_hi, usedIndexedInstructionOffsets_16_hi_lo};
  wire              usedIndexedInstructionOffsets_16 = laneOfOffsetOfOffsetGroup[16] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_16_hi, usedIndexedInstructionOffsets_16_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_17_lo_lo_lo = {usedIndexedInstructionOffsets_17_lo_lo_lo_hi, usedIndexedInstructionOffsets_17_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_17_lo_lo_hi = {usedIndexedInstructionOffsets_17_lo_lo_hi_hi, usedIndexedInstructionOffsets_17_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_17_lo_lo = {usedIndexedInstructionOffsets_17_lo_lo_hi, usedIndexedInstructionOffsets_17_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_17_lo_hi_lo = {usedIndexedInstructionOffsets_17_lo_hi_lo_hi, usedIndexedInstructionOffsets_17_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_17_lo_hi_hi = {usedIndexedInstructionOffsets_17_lo_hi_hi_hi, usedIndexedInstructionOffsets_17_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_17_lo_hi = {usedIndexedInstructionOffsets_17_lo_hi_hi, usedIndexedInstructionOffsets_17_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_17_lo = {usedIndexedInstructionOffsets_17_lo_hi, usedIndexedInstructionOffsets_17_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_17_hi_lo_lo = {usedIndexedInstructionOffsets_17_hi_lo_lo_hi, usedIndexedInstructionOffsets_17_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_17_hi_lo_hi = {usedIndexedInstructionOffsets_17_hi_lo_hi_hi, usedIndexedInstructionOffsets_17_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_17_hi_lo = {usedIndexedInstructionOffsets_17_hi_lo_hi, usedIndexedInstructionOffsets_17_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_17_hi_hi_lo = {usedIndexedInstructionOffsets_17_hi_hi_lo_hi, usedIndexedInstructionOffsets_17_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_17_hi_hi_hi = {usedIndexedInstructionOffsets_17_hi_hi_hi_hi, usedIndexedInstructionOffsets_17_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_17_hi_hi = {usedIndexedInstructionOffsets_17_hi_hi_hi, usedIndexedInstructionOffsets_17_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_17_hi = {usedIndexedInstructionOffsets_17_hi_hi, usedIndexedInstructionOffsets_17_hi_lo};
  wire              usedIndexedInstructionOffsets_17 = laneOfOffsetOfOffsetGroup[17] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_17_hi, usedIndexedInstructionOffsets_17_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_18_lo_lo_lo = {usedIndexedInstructionOffsets_18_lo_lo_lo_hi, usedIndexedInstructionOffsets_18_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_18_lo_lo_hi = {usedIndexedInstructionOffsets_18_lo_lo_hi_hi, usedIndexedInstructionOffsets_18_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_18_lo_lo = {usedIndexedInstructionOffsets_18_lo_lo_hi, usedIndexedInstructionOffsets_18_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_18_lo_hi_lo = {usedIndexedInstructionOffsets_18_lo_hi_lo_hi, usedIndexedInstructionOffsets_18_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_18_lo_hi_hi = {usedIndexedInstructionOffsets_18_lo_hi_hi_hi, usedIndexedInstructionOffsets_18_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_18_lo_hi = {usedIndexedInstructionOffsets_18_lo_hi_hi, usedIndexedInstructionOffsets_18_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_18_lo = {usedIndexedInstructionOffsets_18_lo_hi, usedIndexedInstructionOffsets_18_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_18_hi_lo_lo = {usedIndexedInstructionOffsets_18_hi_lo_lo_hi, usedIndexedInstructionOffsets_18_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_18_hi_lo_hi = {usedIndexedInstructionOffsets_18_hi_lo_hi_hi, usedIndexedInstructionOffsets_18_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_18_hi_lo = {usedIndexedInstructionOffsets_18_hi_lo_hi, usedIndexedInstructionOffsets_18_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_18_hi_hi_lo = {usedIndexedInstructionOffsets_18_hi_hi_lo_hi, usedIndexedInstructionOffsets_18_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_18_hi_hi_hi = {usedIndexedInstructionOffsets_18_hi_hi_hi_hi, usedIndexedInstructionOffsets_18_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_18_hi_hi = {usedIndexedInstructionOffsets_18_hi_hi_hi, usedIndexedInstructionOffsets_18_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_18_hi = {usedIndexedInstructionOffsets_18_hi_hi, usedIndexedInstructionOffsets_18_hi_lo};
  wire              usedIndexedInstructionOffsets_18 = laneOfOffsetOfOffsetGroup[18] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_18_hi, usedIndexedInstructionOffsets_18_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_19_lo_lo_lo = {usedIndexedInstructionOffsets_19_lo_lo_lo_hi, usedIndexedInstructionOffsets_19_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_19_lo_lo_hi = {usedIndexedInstructionOffsets_19_lo_lo_hi_hi, usedIndexedInstructionOffsets_19_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_19_lo_lo = {usedIndexedInstructionOffsets_19_lo_lo_hi, usedIndexedInstructionOffsets_19_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_19_lo_hi_lo = {usedIndexedInstructionOffsets_19_lo_hi_lo_hi, usedIndexedInstructionOffsets_19_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_19_lo_hi_hi = {usedIndexedInstructionOffsets_19_lo_hi_hi_hi, usedIndexedInstructionOffsets_19_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_19_lo_hi = {usedIndexedInstructionOffsets_19_lo_hi_hi, usedIndexedInstructionOffsets_19_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_19_lo = {usedIndexedInstructionOffsets_19_lo_hi, usedIndexedInstructionOffsets_19_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_19_hi_lo_lo = {usedIndexedInstructionOffsets_19_hi_lo_lo_hi, usedIndexedInstructionOffsets_19_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_19_hi_lo_hi = {usedIndexedInstructionOffsets_19_hi_lo_hi_hi, usedIndexedInstructionOffsets_19_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_19_hi_lo = {usedIndexedInstructionOffsets_19_hi_lo_hi, usedIndexedInstructionOffsets_19_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_19_hi_hi_lo = {usedIndexedInstructionOffsets_19_hi_hi_lo_hi, usedIndexedInstructionOffsets_19_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_19_hi_hi_hi = {usedIndexedInstructionOffsets_19_hi_hi_hi_hi, usedIndexedInstructionOffsets_19_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_19_hi_hi = {usedIndexedInstructionOffsets_19_hi_hi_hi, usedIndexedInstructionOffsets_19_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_19_hi = {usedIndexedInstructionOffsets_19_hi_hi, usedIndexedInstructionOffsets_19_hi_lo};
  wire              usedIndexedInstructionOffsets_19 = laneOfOffsetOfOffsetGroup[19] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_19_hi, usedIndexedInstructionOffsets_19_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_20_lo_lo_lo = {usedIndexedInstructionOffsets_20_lo_lo_lo_hi, usedIndexedInstructionOffsets_20_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_20_lo_lo_hi = {usedIndexedInstructionOffsets_20_lo_lo_hi_hi, usedIndexedInstructionOffsets_20_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_20_lo_lo = {usedIndexedInstructionOffsets_20_lo_lo_hi, usedIndexedInstructionOffsets_20_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_20_lo_hi_lo = {usedIndexedInstructionOffsets_20_lo_hi_lo_hi, usedIndexedInstructionOffsets_20_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_20_lo_hi_hi = {usedIndexedInstructionOffsets_20_lo_hi_hi_hi, usedIndexedInstructionOffsets_20_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_20_lo_hi = {usedIndexedInstructionOffsets_20_lo_hi_hi, usedIndexedInstructionOffsets_20_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_20_lo = {usedIndexedInstructionOffsets_20_lo_hi, usedIndexedInstructionOffsets_20_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_20_hi_lo_lo = {usedIndexedInstructionOffsets_20_hi_lo_lo_hi, usedIndexedInstructionOffsets_20_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_20_hi_lo_hi = {usedIndexedInstructionOffsets_20_hi_lo_hi_hi, usedIndexedInstructionOffsets_20_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_20_hi_lo = {usedIndexedInstructionOffsets_20_hi_lo_hi, usedIndexedInstructionOffsets_20_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_20_hi_hi_lo = {usedIndexedInstructionOffsets_20_hi_hi_lo_hi, usedIndexedInstructionOffsets_20_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_20_hi_hi_hi = {usedIndexedInstructionOffsets_20_hi_hi_hi_hi, usedIndexedInstructionOffsets_20_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_20_hi_hi = {usedIndexedInstructionOffsets_20_hi_hi_hi, usedIndexedInstructionOffsets_20_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_20_hi = {usedIndexedInstructionOffsets_20_hi_hi, usedIndexedInstructionOffsets_20_hi_lo};
  wire              usedIndexedInstructionOffsets_20 = laneOfOffsetOfOffsetGroup[20] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_20_hi, usedIndexedInstructionOffsets_20_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_21_lo_lo_lo = {usedIndexedInstructionOffsets_21_lo_lo_lo_hi, usedIndexedInstructionOffsets_21_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_21_lo_lo_hi = {usedIndexedInstructionOffsets_21_lo_lo_hi_hi, usedIndexedInstructionOffsets_21_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_21_lo_lo = {usedIndexedInstructionOffsets_21_lo_lo_hi, usedIndexedInstructionOffsets_21_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_21_lo_hi_lo = {usedIndexedInstructionOffsets_21_lo_hi_lo_hi, usedIndexedInstructionOffsets_21_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_21_lo_hi_hi = {usedIndexedInstructionOffsets_21_lo_hi_hi_hi, usedIndexedInstructionOffsets_21_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_21_lo_hi = {usedIndexedInstructionOffsets_21_lo_hi_hi, usedIndexedInstructionOffsets_21_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_21_lo = {usedIndexedInstructionOffsets_21_lo_hi, usedIndexedInstructionOffsets_21_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_21_hi_lo_lo = {usedIndexedInstructionOffsets_21_hi_lo_lo_hi, usedIndexedInstructionOffsets_21_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_21_hi_lo_hi = {usedIndexedInstructionOffsets_21_hi_lo_hi_hi, usedIndexedInstructionOffsets_21_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_21_hi_lo = {usedIndexedInstructionOffsets_21_hi_lo_hi, usedIndexedInstructionOffsets_21_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_21_hi_hi_lo = {usedIndexedInstructionOffsets_21_hi_hi_lo_hi, usedIndexedInstructionOffsets_21_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_21_hi_hi_hi = {usedIndexedInstructionOffsets_21_hi_hi_hi_hi, usedIndexedInstructionOffsets_21_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_21_hi_hi = {usedIndexedInstructionOffsets_21_hi_hi_hi, usedIndexedInstructionOffsets_21_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_21_hi = {usedIndexedInstructionOffsets_21_hi_hi, usedIndexedInstructionOffsets_21_hi_lo};
  wire              usedIndexedInstructionOffsets_21 = laneOfOffsetOfOffsetGroup[21] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_21_hi, usedIndexedInstructionOffsets_21_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_22_lo_lo_lo = {usedIndexedInstructionOffsets_22_lo_lo_lo_hi, usedIndexedInstructionOffsets_22_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_22_lo_lo_hi = {usedIndexedInstructionOffsets_22_lo_lo_hi_hi, usedIndexedInstructionOffsets_22_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_22_lo_lo = {usedIndexedInstructionOffsets_22_lo_lo_hi, usedIndexedInstructionOffsets_22_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_22_lo_hi_lo = {usedIndexedInstructionOffsets_22_lo_hi_lo_hi, usedIndexedInstructionOffsets_22_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_22_lo_hi_hi = {usedIndexedInstructionOffsets_22_lo_hi_hi_hi, usedIndexedInstructionOffsets_22_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_22_lo_hi = {usedIndexedInstructionOffsets_22_lo_hi_hi, usedIndexedInstructionOffsets_22_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_22_lo = {usedIndexedInstructionOffsets_22_lo_hi, usedIndexedInstructionOffsets_22_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_22_hi_lo_lo = {usedIndexedInstructionOffsets_22_hi_lo_lo_hi, usedIndexedInstructionOffsets_22_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_22_hi_lo_hi = {usedIndexedInstructionOffsets_22_hi_lo_hi_hi, usedIndexedInstructionOffsets_22_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_22_hi_lo = {usedIndexedInstructionOffsets_22_hi_lo_hi, usedIndexedInstructionOffsets_22_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_22_hi_hi_lo = {usedIndexedInstructionOffsets_22_hi_hi_lo_hi, usedIndexedInstructionOffsets_22_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_22_hi_hi_hi = {usedIndexedInstructionOffsets_22_hi_hi_hi_hi, usedIndexedInstructionOffsets_22_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_22_hi_hi = {usedIndexedInstructionOffsets_22_hi_hi_hi, usedIndexedInstructionOffsets_22_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_22_hi = {usedIndexedInstructionOffsets_22_hi_hi, usedIndexedInstructionOffsets_22_hi_lo};
  wire              usedIndexedInstructionOffsets_22 = laneOfOffsetOfOffsetGroup[22] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_22_hi, usedIndexedInstructionOffsets_22_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_23_lo_lo_lo = {usedIndexedInstructionOffsets_23_lo_lo_lo_hi, usedIndexedInstructionOffsets_23_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_23_lo_lo_hi = {usedIndexedInstructionOffsets_23_lo_lo_hi_hi, usedIndexedInstructionOffsets_23_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_23_lo_lo = {usedIndexedInstructionOffsets_23_lo_lo_hi, usedIndexedInstructionOffsets_23_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_23_lo_hi_lo = {usedIndexedInstructionOffsets_23_lo_hi_lo_hi, usedIndexedInstructionOffsets_23_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_23_lo_hi_hi = {usedIndexedInstructionOffsets_23_lo_hi_hi_hi, usedIndexedInstructionOffsets_23_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_23_lo_hi = {usedIndexedInstructionOffsets_23_lo_hi_hi, usedIndexedInstructionOffsets_23_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_23_lo = {usedIndexedInstructionOffsets_23_lo_hi, usedIndexedInstructionOffsets_23_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_23_hi_lo_lo = {usedIndexedInstructionOffsets_23_hi_lo_lo_hi, usedIndexedInstructionOffsets_23_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_23_hi_lo_hi = {usedIndexedInstructionOffsets_23_hi_lo_hi_hi, usedIndexedInstructionOffsets_23_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_23_hi_lo = {usedIndexedInstructionOffsets_23_hi_lo_hi, usedIndexedInstructionOffsets_23_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_23_hi_hi_lo = {usedIndexedInstructionOffsets_23_hi_hi_lo_hi, usedIndexedInstructionOffsets_23_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_23_hi_hi_hi = {usedIndexedInstructionOffsets_23_hi_hi_hi_hi, usedIndexedInstructionOffsets_23_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_23_hi_hi = {usedIndexedInstructionOffsets_23_hi_hi_hi, usedIndexedInstructionOffsets_23_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_23_hi = {usedIndexedInstructionOffsets_23_hi_hi, usedIndexedInstructionOffsets_23_hi_lo};
  wire              usedIndexedInstructionOffsets_23 = laneOfOffsetOfOffsetGroup[23] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_23_hi, usedIndexedInstructionOffsets_23_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_24_lo_lo_lo = {usedIndexedInstructionOffsets_24_lo_lo_lo_hi, usedIndexedInstructionOffsets_24_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_24_lo_lo_hi = {usedIndexedInstructionOffsets_24_lo_lo_hi_hi, usedIndexedInstructionOffsets_24_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_24_lo_lo = {usedIndexedInstructionOffsets_24_lo_lo_hi, usedIndexedInstructionOffsets_24_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_24_lo_hi_lo = {usedIndexedInstructionOffsets_24_lo_hi_lo_hi, usedIndexedInstructionOffsets_24_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_24_lo_hi_hi = {usedIndexedInstructionOffsets_24_lo_hi_hi_hi, usedIndexedInstructionOffsets_24_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_24_lo_hi = {usedIndexedInstructionOffsets_24_lo_hi_hi, usedIndexedInstructionOffsets_24_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_24_lo = {usedIndexedInstructionOffsets_24_lo_hi, usedIndexedInstructionOffsets_24_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_24_hi_lo_lo = {usedIndexedInstructionOffsets_24_hi_lo_lo_hi, usedIndexedInstructionOffsets_24_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_24_hi_lo_hi = {usedIndexedInstructionOffsets_24_hi_lo_hi_hi, usedIndexedInstructionOffsets_24_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_24_hi_lo = {usedIndexedInstructionOffsets_24_hi_lo_hi, usedIndexedInstructionOffsets_24_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_24_hi_hi_lo = {usedIndexedInstructionOffsets_24_hi_hi_lo_hi, usedIndexedInstructionOffsets_24_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_24_hi_hi_hi = {usedIndexedInstructionOffsets_24_hi_hi_hi_hi, usedIndexedInstructionOffsets_24_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_24_hi_hi = {usedIndexedInstructionOffsets_24_hi_hi_hi, usedIndexedInstructionOffsets_24_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_24_hi = {usedIndexedInstructionOffsets_24_hi_hi, usedIndexedInstructionOffsets_24_hi_lo};
  wire              usedIndexedInstructionOffsets_24 = laneOfOffsetOfOffsetGroup[24] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_24_hi, usedIndexedInstructionOffsets_24_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_25_lo_lo_lo = {usedIndexedInstructionOffsets_25_lo_lo_lo_hi, usedIndexedInstructionOffsets_25_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_25_lo_lo_hi = {usedIndexedInstructionOffsets_25_lo_lo_hi_hi, usedIndexedInstructionOffsets_25_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_25_lo_lo = {usedIndexedInstructionOffsets_25_lo_lo_hi, usedIndexedInstructionOffsets_25_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_25_lo_hi_lo = {usedIndexedInstructionOffsets_25_lo_hi_lo_hi, usedIndexedInstructionOffsets_25_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_25_lo_hi_hi = {usedIndexedInstructionOffsets_25_lo_hi_hi_hi, usedIndexedInstructionOffsets_25_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_25_lo_hi = {usedIndexedInstructionOffsets_25_lo_hi_hi, usedIndexedInstructionOffsets_25_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_25_lo = {usedIndexedInstructionOffsets_25_lo_hi, usedIndexedInstructionOffsets_25_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_25_hi_lo_lo = {usedIndexedInstructionOffsets_25_hi_lo_lo_hi, usedIndexedInstructionOffsets_25_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_25_hi_lo_hi = {usedIndexedInstructionOffsets_25_hi_lo_hi_hi, usedIndexedInstructionOffsets_25_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_25_hi_lo = {usedIndexedInstructionOffsets_25_hi_lo_hi, usedIndexedInstructionOffsets_25_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_25_hi_hi_lo = {usedIndexedInstructionOffsets_25_hi_hi_lo_hi, usedIndexedInstructionOffsets_25_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_25_hi_hi_hi = {usedIndexedInstructionOffsets_25_hi_hi_hi_hi, usedIndexedInstructionOffsets_25_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_25_hi_hi = {usedIndexedInstructionOffsets_25_hi_hi_hi, usedIndexedInstructionOffsets_25_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_25_hi = {usedIndexedInstructionOffsets_25_hi_hi, usedIndexedInstructionOffsets_25_hi_lo};
  wire              usedIndexedInstructionOffsets_25 = laneOfOffsetOfOffsetGroup[25] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_25_hi, usedIndexedInstructionOffsets_25_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_26_lo_lo_lo = {usedIndexedInstructionOffsets_26_lo_lo_lo_hi, usedIndexedInstructionOffsets_26_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_26_lo_lo_hi = {usedIndexedInstructionOffsets_26_lo_lo_hi_hi, usedIndexedInstructionOffsets_26_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_26_lo_lo = {usedIndexedInstructionOffsets_26_lo_lo_hi, usedIndexedInstructionOffsets_26_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_26_lo_hi_lo = {usedIndexedInstructionOffsets_26_lo_hi_lo_hi, usedIndexedInstructionOffsets_26_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_26_lo_hi_hi = {usedIndexedInstructionOffsets_26_lo_hi_hi_hi, usedIndexedInstructionOffsets_26_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_26_lo_hi = {usedIndexedInstructionOffsets_26_lo_hi_hi, usedIndexedInstructionOffsets_26_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_26_lo = {usedIndexedInstructionOffsets_26_lo_hi, usedIndexedInstructionOffsets_26_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_26_hi_lo_lo = {usedIndexedInstructionOffsets_26_hi_lo_lo_hi, usedIndexedInstructionOffsets_26_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_26_hi_lo_hi = {usedIndexedInstructionOffsets_26_hi_lo_hi_hi, usedIndexedInstructionOffsets_26_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_26_hi_lo = {usedIndexedInstructionOffsets_26_hi_lo_hi, usedIndexedInstructionOffsets_26_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_26_hi_hi_lo = {usedIndexedInstructionOffsets_26_hi_hi_lo_hi, usedIndexedInstructionOffsets_26_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_26_hi_hi_hi = {usedIndexedInstructionOffsets_26_hi_hi_hi_hi, usedIndexedInstructionOffsets_26_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_26_hi_hi = {usedIndexedInstructionOffsets_26_hi_hi_hi, usedIndexedInstructionOffsets_26_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_26_hi = {usedIndexedInstructionOffsets_26_hi_hi, usedIndexedInstructionOffsets_26_hi_lo};
  wire              usedIndexedInstructionOffsets_26 = laneOfOffsetOfOffsetGroup[26] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_26_hi, usedIndexedInstructionOffsets_26_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_27_lo_lo_lo = {usedIndexedInstructionOffsets_27_lo_lo_lo_hi, usedIndexedInstructionOffsets_27_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_27_lo_lo_hi = {usedIndexedInstructionOffsets_27_lo_lo_hi_hi, usedIndexedInstructionOffsets_27_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_27_lo_lo = {usedIndexedInstructionOffsets_27_lo_lo_hi, usedIndexedInstructionOffsets_27_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_27_lo_hi_lo = {usedIndexedInstructionOffsets_27_lo_hi_lo_hi, usedIndexedInstructionOffsets_27_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_27_lo_hi_hi = {usedIndexedInstructionOffsets_27_lo_hi_hi_hi, usedIndexedInstructionOffsets_27_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_27_lo_hi = {usedIndexedInstructionOffsets_27_lo_hi_hi, usedIndexedInstructionOffsets_27_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_27_lo = {usedIndexedInstructionOffsets_27_lo_hi, usedIndexedInstructionOffsets_27_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_27_hi_lo_lo = {usedIndexedInstructionOffsets_27_hi_lo_lo_hi, usedIndexedInstructionOffsets_27_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_27_hi_lo_hi = {usedIndexedInstructionOffsets_27_hi_lo_hi_hi, usedIndexedInstructionOffsets_27_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_27_hi_lo = {usedIndexedInstructionOffsets_27_hi_lo_hi, usedIndexedInstructionOffsets_27_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_27_hi_hi_lo = {usedIndexedInstructionOffsets_27_hi_hi_lo_hi, usedIndexedInstructionOffsets_27_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_27_hi_hi_hi = {usedIndexedInstructionOffsets_27_hi_hi_hi_hi, usedIndexedInstructionOffsets_27_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_27_hi_hi = {usedIndexedInstructionOffsets_27_hi_hi_hi, usedIndexedInstructionOffsets_27_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_27_hi = {usedIndexedInstructionOffsets_27_hi_hi, usedIndexedInstructionOffsets_27_hi_lo};
  wire              usedIndexedInstructionOffsets_27 = laneOfOffsetOfOffsetGroup[27] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_27_hi, usedIndexedInstructionOffsets_27_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_28_lo_lo_lo = {usedIndexedInstructionOffsets_28_lo_lo_lo_hi, usedIndexedInstructionOffsets_28_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_28_lo_lo_hi = {usedIndexedInstructionOffsets_28_lo_lo_hi_hi, usedIndexedInstructionOffsets_28_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_28_lo_lo = {usedIndexedInstructionOffsets_28_lo_lo_hi, usedIndexedInstructionOffsets_28_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_28_lo_hi_lo = {usedIndexedInstructionOffsets_28_lo_hi_lo_hi, usedIndexedInstructionOffsets_28_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_28_lo_hi_hi = {usedIndexedInstructionOffsets_28_lo_hi_hi_hi, usedIndexedInstructionOffsets_28_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_28_lo_hi = {usedIndexedInstructionOffsets_28_lo_hi_hi, usedIndexedInstructionOffsets_28_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_28_lo = {usedIndexedInstructionOffsets_28_lo_hi, usedIndexedInstructionOffsets_28_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_28_hi_lo_lo = {usedIndexedInstructionOffsets_28_hi_lo_lo_hi, usedIndexedInstructionOffsets_28_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_28_hi_lo_hi = {usedIndexedInstructionOffsets_28_hi_lo_hi_hi, usedIndexedInstructionOffsets_28_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_28_hi_lo = {usedIndexedInstructionOffsets_28_hi_lo_hi, usedIndexedInstructionOffsets_28_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_28_hi_hi_lo = {usedIndexedInstructionOffsets_28_hi_hi_lo_hi, usedIndexedInstructionOffsets_28_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_28_hi_hi_hi = {usedIndexedInstructionOffsets_28_hi_hi_hi_hi, usedIndexedInstructionOffsets_28_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_28_hi_hi = {usedIndexedInstructionOffsets_28_hi_hi_hi, usedIndexedInstructionOffsets_28_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_28_hi = {usedIndexedInstructionOffsets_28_hi_hi, usedIndexedInstructionOffsets_28_hi_lo};
  wire              usedIndexedInstructionOffsets_28 = laneOfOffsetOfOffsetGroup[28] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_28_hi, usedIndexedInstructionOffsets_28_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_29_lo_lo_lo = {usedIndexedInstructionOffsets_29_lo_lo_lo_hi, usedIndexedInstructionOffsets_29_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_29_lo_lo_hi = {usedIndexedInstructionOffsets_29_lo_lo_hi_hi, usedIndexedInstructionOffsets_29_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_29_lo_lo = {usedIndexedInstructionOffsets_29_lo_lo_hi, usedIndexedInstructionOffsets_29_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_29_lo_hi_lo = {usedIndexedInstructionOffsets_29_lo_hi_lo_hi, usedIndexedInstructionOffsets_29_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_29_lo_hi_hi = {usedIndexedInstructionOffsets_29_lo_hi_hi_hi, usedIndexedInstructionOffsets_29_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_29_lo_hi = {usedIndexedInstructionOffsets_29_lo_hi_hi, usedIndexedInstructionOffsets_29_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_29_lo = {usedIndexedInstructionOffsets_29_lo_hi, usedIndexedInstructionOffsets_29_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_29_hi_lo_lo = {usedIndexedInstructionOffsets_29_hi_lo_lo_hi, usedIndexedInstructionOffsets_29_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_29_hi_lo_hi = {usedIndexedInstructionOffsets_29_hi_lo_hi_hi, usedIndexedInstructionOffsets_29_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_29_hi_lo = {usedIndexedInstructionOffsets_29_hi_lo_hi, usedIndexedInstructionOffsets_29_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_29_hi_hi_lo = {usedIndexedInstructionOffsets_29_hi_hi_lo_hi, usedIndexedInstructionOffsets_29_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_29_hi_hi_hi = {usedIndexedInstructionOffsets_29_hi_hi_hi_hi, usedIndexedInstructionOffsets_29_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_29_hi_hi = {usedIndexedInstructionOffsets_29_hi_hi_hi, usedIndexedInstructionOffsets_29_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_29_hi = {usedIndexedInstructionOffsets_29_hi_hi, usedIndexedInstructionOffsets_29_hi_lo};
  wire              usedIndexedInstructionOffsets_29 = laneOfOffsetOfOffsetGroup[29] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_29_hi, usedIndexedInstructionOffsets_29_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_30_lo_lo_lo = {usedIndexedInstructionOffsets_30_lo_lo_lo_hi, usedIndexedInstructionOffsets_30_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_30_lo_lo_hi = {usedIndexedInstructionOffsets_30_lo_lo_hi_hi, usedIndexedInstructionOffsets_30_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_30_lo_lo = {usedIndexedInstructionOffsets_30_lo_lo_hi, usedIndexedInstructionOffsets_30_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_30_lo_hi_lo = {usedIndexedInstructionOffsets_30_lo_hi_lo_hi, usedIndexedInstructionOffsets_30_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_30_lo_hi_hi = {usedIndexedInstructionOffsets_30_lo_hi_hi_hi, usedIndexedInstructionOffsets_30_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_30_lo_hi = {usedIndexedInstructionOffsets_30_lo_hi_hi, usedIndexedInstructionOffsets_30_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_30_lo = {usedIndexedInstructionOffsets_30_lo_hi, usedIndexedInstructionOffsets_30_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_30_hi_lo_lo = {usedIndexedInstructionOffsets_30_hi_lo_lo_hi, usedIndexedInstructionOffsets_30_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_30_hi_lo_hi = {usedIndexedInstructionOffsets_30_hi_lo_hi_hi, usedIndexedInstructionOffsets_30_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_30_hi_lo = {usedIndexedInstructionOffsets_30_hi_lo_hi, usedIndexedInstructionOffsets_30_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_30_hi_hi_lo = {usedIndexedInstructionOffsets_30_hi_hi_lo_hi, usedIndexedInstructionOffsets_30_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_30_hi_hi_hi = {usedIndexedInstructionOffsets_30_hi_hi_hi_hi, usedIndexedInstructionOffsets_30_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_30_hi_hi = {usedIndexedInstructionOffsets_30_hi_hi_hi, usedIndexedInstructionOffsets_30_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_30_hi = {usedIndexedInstructionOffsets_30_hi_hi, usedIndexedInstructionOffsets_30_hi_lo};
  wire              usedIndexedInstructionOffsets_30 = laneOfOffsetOfOffsetGroup[30] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_30_hi, usedIndexedInstructionOffsets_30_lo}) | maskGroupEndAndRequestNewMask;
  wire [3:0]        usedIndexedInstructionOffsets_31_lo_lo_lo = {usedIndexedInstructionOffsets_31_lo_lo_lo_hi, usedIndexedInstructionOffsets_31_lo_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_31_lo_lo_hi = {usedIndexedInstructionOffsets_31_lo_lo_hi_hi, usedIndexedInstructionOffsets_31_lo_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_31_lo_lo = {usedIndexedInstructionOffsets_31_lo_lo_hi, usedIndexedInstructionOffsets_31_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_31_lo_hi_lo = {usedIndexedInstructionOffsets_31_lo_hi_lo_hi, usedIndexedInstructionOffsets_31_lo_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_31_lo_hi_hi = {usedIndexedInstructionOffsets_31_lo_hi_hi_hi, usedIndexedInstructionOffsets_31_lo_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_31_lo_hi = {usedIndexedInstructionOffsets_31_lo_hi_hi, usedIndexedInstructionOffsets_31_lo_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_31_lo = {usedIndexedInstructionOffsets_31_lo_hi, usedIndexedInstructionOffsets_31_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_31_hi_lo_lo = {usedIndexedInstructionOffsets_31_hi_lo_lo_hi, usedIndexedInstructionOffsets_31_hi_lo_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_31_hi_lo_hi = {usedIndexedInstructionOffsets_31_hi_lo_hi_hi, usedIndexedInstructionOffsets_31_hi_lo_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_31_hi_lo = {usedIndexedInstructionOffsets_31_hi_lo_hi, usedIndexedInstructionOffsets_31_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_31_hi_hi_lo = {usedIndexedInstructionOffsets_31_hi_hi_lo_hi, usedIndexedInstructionOffsets_31_hi_hi_lo_lo};
  wire [3:0]        usedIndexedInstructionOffsets_31_hi_hi_hi = {usedIndexedInstructionOffsets_31_hi_hi_hi_hi, usedIndexedInstructionOffsets_31_hi_hi_hi_lo};
  wire [7:0]        usedIndexedInstructionOffsets_31_hi_hi = {usedIndexedInstructionOffsets_31_hi_hi_hi, usedIndexedInstructionOffsets_31_hi_hi_lo};
  wire [15:0]       usedIndexedInstructionOffsets_31_hi = {usedIndexedInstructionOffsets_31_hi_hi, usedIndexedInstructionOffsets_31_hi_lo};
  wire              usedIndexedInstructionOffsets_31 = laneOfOffsetOfOffsetGroup[31] & _GEN | requestOffset & (&{usedIndexedInstructionOffsets_31_hi, usedIndexedInstructionOffsets_31_lo}) | maskGroupEndAndRequestNewMask;
  wire [127:0]      memoryRequestSourceOH;
  wire              sourceFree = (memoryRequestSourceOH & outstandingTLDMessages) == 128'h0;
  wire              stateIsRequest = state == 2'h1;
  wire [11:0]       nextElementIndex = {stateIsRequest ? groupIndex : nextGroupIndex, stateIsRequest ? nextElementForMemoryRequestIndex : 7'h0};
  wire [9:0]        wholeEvl = {{1'h0, lsuRequestReg_instructionInformation_nf} + 4'h1, 6'h0};
  wire [11:0]       evl = isWholeRegisterLoadStore ? {2'h0, wholeEvl} : isMaskLoadStore ? {3'h0, csrInterfaceReg_vl[11:3] + {8'h0, |(csrInterfaceReg_vl[2:0])}} : csrInterfaceReg_vl;
  assign last = nextElementIndex >= evl;
  wire              vrfWritePort_bits_last_0 = last;
  wire              maskCheck = ~lsuRequestReg_instructionInformation_maskedLoadStore | ~noMoreMaskedUnsentMemoryRequests;
  wire              indexCheck = ~isIndexedLoadStore | offsetValidCheck & offsetGroupCheck;
  reg               firstMemoryRequestOfInstruction;
  reg               waitFirstMemoryResponseForFaultOnlyFirst;
  wire              fofCheck = firstMemoryRequestOfInstruction | ~waitFirstMemoryResponseForFaultOnlyFirst;
  wire              _requestOffset_T = stateIsRequest & maskCheck;
  wire              stateReady = _requestOffset_T & indexCheck & fofCheck;
  assign requestOffset = _requestOffset_T & ~indexCheck & fofCheck;
  wire              s0EnqueueValid = stateReady & ~last;
  reg               s0Valid;
  reg  [4:0]        s0Reg_readVS;
  wire [4:0]        vrfReadDataPorts_bits_vs_0 = s0Reg_readVS;
  reg               s0Reg_offsetForVSInLane;
  wire              vrfReadDataPorts_bits_offset_0 = s0Reg_offsetForVSInLane;
  reg  [31:0]       s0Reg_addressOffset;
  reg  [2:0]        s0Reg_segmentIndex;
  wire [2:0]        s1EnqQueue_enq_bits_segmentIndex = s0Reg_segmentIndex;
  reg  [4:0]        s0Reg_offsetForLane;
  reg  [6:0]        s0Reg_indexInGroup;
  wire [6:0]        s1EnqQueue_enq_bits_indexInMaskGroup = s0Reg_indexInGroup;
  wire              s1EnqDataQueue_deq_ready = s1EnqueueReady;
  wire              s1EnqQueue_deq_valid;
  assign s1EnqQueue_deq_valid = ~_s1EnqQueue_fifo_empty;
  wire [6:0]        s1EnqQueue_dataOut_indexInMaskGroup;
  wire [2:0]        s1EnqQueue_dataOut_segmentIndex;
  wire [6:0]        s1Wire_indexInMaskGroup = s1EnqQueue_deq_bits_indexInMaskGroup;
  wire [31:0]       s1EnqQueue_dataOut_address;
  wire [2:0]        s1Wire_segmentIndex = s1EnqQueue_deq_bits_segmentIndex;
  wire [31:0]       s1EnqQueue_dataOut_readData;
  wire [31:0]       s1Wire_address = s1EnqQueue_deq_bits_address;
  wire [31:0]       s1EnqQueue_enq_bits_address;
  wire [63:0]       s1EnqQueue_dataIn_lo = {s1EnqQueue_enq_bits_address, 32'h0};
  wire [9:0]        s1EnqQueue_dataIn_hi = {s1EnqQueue_enq_bits_indexInMaskGroup, s1EnqQueue_enq_bits_segmentIndex};
  wire [73:0]       s1EnqQueue_dataIn = {s1EnqQueue_dataIn_hi, s1EnqQueue_dataIn_lo};
  assign s1EnqQueue_dataOut_readData = _s1EnqQueue_fifo_data_out[31:0];
  assign s1EnqQueue_dataOut_address = _s1EnqQueue_fifo_data_out[63:32];
  assign s1EnqQueue_dataOut_segmentIndex = _s1EnqQueue_fifo_data_out[66:64];
  assign s1EnqQueue_dataOut_indexInMaskGroup = _s1EnqQueue_fifo_data_out[73:67];
  assign s1EnqQueue_deq_bits_indexInMaskGroup = s1EnqQueue_dataOut_indexInMaskGroup;
  assign s1EnqQueue_deq_bits_segmentIndex = s1EnqQueue_dataOut_segmentIndex;
  assign s1EnqQueue_deq_bits_address = s1EnqQueue_dataOut_address;
  wire [31:0]       s1EnqQueue_deq_bits_readData = s1EnqQueue_dataOut_readData;
  wire              s1EnqQueue_enq_ready = ~_s1EnqQueue_fifo_full;
  wire              s1EnqQueue_enq_valid;
  wire              s0DequeueFire = s1EnqQueue_enq_ready & s1EnqQueue_enq_valid;
  wire              s1EnqQueue_deq_ready;
  wire              s1EnqDataQueue_deq_valid;
  assign s1EnqDataQueue_deq_valid = ~_s1EnqDataQueue_fifo_empty;
  wire [31:0]       s1Wire_readData = s1EnqDataQueue_deq_bits;
  wire              s1EnqDataQueue_enq_ready = ~_s1EnqDataQueue_fifo_full;
  wire [14:0]       _GEN_16 = {13'h0, dataEEW};
  wire [14:0]       _storeBaseByteOffset_T = {3'h0, s0ElementIndex} << _GEN_16;
  wire [10:0]       storeBaseByteOffset = _storeBaseByteOffset_T[10:0];
  wire [4:0]        _GEN_17 = {1'h0, segmentInstructionIndexInterval};
  wire [4:0]        s0Wire_readVS = lsuRequestReg_instructionInformation_vs3 + (isSegmentLoadStore ? {2'h0, segmentIndex} * _GEN_17 : 5'h0) + {2'h0, storeBaseByteOffset[10:8]};
  wire              s0Wire_offsetForVSInLane = storeBaseByteOffset[7];
  wire [31:0]       s0Wire_addressOffset = baseOffsetForElement[31:0] + {26'h0, {3'h0, elementByteWidth} * {3'h0, segmentIndex}};
  wire [4:0]        s0Wire_offsetForLane = storeBaseByteOffset[6:2];
  wire              vrfReadDataPorts_valid_0 = s0Valid & lsuRequestReg_instructionInformation_isStore & s1EnqQueue_enq_ready;
  wire              readReady = ~lsuRequestReg_instructionInformation_isStore | vrfReadDataPorts_ready_0;
  reg               s1Valid;
  reg  [6:0]        s1Reg_indexInMaskGroup;
  reg  [2:0]        s1Reg_segmentIndex;
  reg  [31:0]       s1Reg_address;
  wire [31:0]       memWriteRequest_bits_address_0 = s1Reg_address;
  reg  [31:0]       s1Reg_readData;
  wire              memRequestReady = lsuRequestReg_instructionInformation_isStore ? memWriteRequest_ready_0 : memReadRequest_ready_0;
  wire              s2EnqueueReady = memRequestReady & sourceFree;
  assign s1EnqueueReady = s2EnqueueReady | ~s1Valid;
  wire              s0EnqueueReady = s1EnqQueue_enq_ready & readReady | ~s0Valid;
  assign s0Fire = s0EnqueueReady & s0EnqueueValid;
  wire              pipelineClear = ~s0Valid & ~s1Valid & ~s1EnqQueue_deq_valid;
  assign s1EnqQueue_enq_valid = s0Valid & readReady;
  assign s1EnqQueue_enq_bits_address = lsuRequestReg_rs1Data + s0Reg_addressOffset;
  wire              s1DataEnqValid = s1EnqDataQueue_deq_valid | ~lsuRequestReg_instructionInformation_isStore;
  wire              s1EnqValid = s1DataEnqValid & s1EnqQueue_deq_valid;
  wire              s1Fire = s1EnqValid & s1EnqueueReady;
  assign s1EnqQueue_deq_ready = s1EnqueueReady & s1DataEnqValid;
  wire [1:0]        addressInBeatByte = s1Reg_address[1:0];
  wire [3:0]        baseMask = {{2{dataEEWOH[2]}}, ~(dataEEWOH[0]), 1'h1};
  wire [6:0]        _storeMask_T = {3'h0, baseMask} << addressInBeatByte;
  assign storeMask = _storeMask_T[3:0];
  wire [3:0]        memWriteRequest_bits_mask_0 = storeMask;
  wire [4:0]        _storeOffsetByIndex_T_1 = {3'h0, s1Reg_indexInMaskGroup[1:0]} << dataEEW;
  wire [1:0]        storeOffsetByIndex = _storeOffsetByIndex_T_1[1:0];
  wire [62:0]       storeData = {31'h0, s1Reg_readData} << {58'h0, addressInBeatByte, 3'h0} >> {58'h0, storeOffsetByIndex, 3'h0};
  assign memoryRequestSource = isSegmentLoadStore ? {s1Reg_indexInMaskGroup, s1Reg_segmentIndex} : {3'h0, s1Reg_indexInMaskGroup};
  wire [9:0]        memReadRequest_bits_source_0 = memoryRequestSource;
  assign memoryRequestSourceOH = 128'h1 << memoryRequestSource[6:0];
  wire [31:0]       memReadRequest_bits_address_0 = {s1Reg_address[31:2], 2'h0};
  wire              _memWriteRequest_valid_T = s1Valid & sourceFree;
  assign memReadRequest_valid_0 = _memWriteRequest_valid_T & ~lsuRequestReg_instructionInformation_isStore;
  assign memWriteRequest_valid_0 = _memWriteRequest_valid_T & lsuRequestReg_instructionInformation_isStore;
  wire [31:0]       memWriteRequest_bits_data_0 = storeData[31:0];
  wire [7:0]        memWriteRequest_bits_source_0 = memoryRequestSource[7:0];
  reg  [1:0]        offsetRecord_0;
  reg  [1:0]        offsetRecord_1;
  reg  [1:0]        offsetRecord_2;
  reg  [1:0]        offsetRecord_3;
  reg  [1:0]        offsetRecord_4;
  reg  [1:0]        offsetRecord_5;
  reg  [1:0]        offsetRecord_6;
  reg  [1:0]        offsetRecord_7;
  reg  [1:0]        offsetRecord_8;
  reg  [1:0]        offsetRecord_9;
  reg  [1:0]        offsetRecord_10;
  reg  [1:0]        offsetRecord_11;
  reg  [1:0]        offsetRecord_12;
  reg  [1:0]        offsetRecord_13;
  reg  [1:0]        offsetRecord_14;
  reg  [1:0]        offsetRecord_15;
  reg  [1:0]        offsetRecord_16;
  reg  [1:0]        offsetRecord_17;
  reg  [1:0]        offsetRecord_18;
  reg  [1:0]        offsetRecord_19;
  reg  [1:0]        offsetRecord_20;
  reg  [1:0]        offsetRecord_21;
  reg  [1:0]        offsetRecord_22;
  reg  [1:0]        offsetRecord_23;
  reg  [1:0]        offsetRecord_24;
  reg  [1:0]        offsetRecord_25;
  reg  [1:0]        offsetRecord_26;
  reg  [1:0]        offsetRecord_27;
  reg  [1:0]        offsetRecord_28;
  reg  [1:0]        offsetRecord_29;
  reg  [1:0]        offsetRecord_30;
  reg  [1:0]        offsetRecord_31;
  reg  [1:0]        offsetRecord_32;
  reg  [1:0]        offsetRecord_33;
  reg  [1:0]        offsetRecord_34;
  reg  [1:0]        offsetRecord_35;
  reg  [1:0]        offsetRecord_36;
  reg  [1:0]        offsetRecord_37;
  reg  [1:0]        offsetRecord_38;
  reg  [1:0]        offsetRecord_39;
  reg  [1:0]        offsetRecord_40;
  reg  [1:0]        offsetRecord_41;
  reg  [1:0]        offsetRecord_42;
  reg  [1:0]        offsetRecord_43;
  reg  [1:0]        offsetRecord_44;
  reg  [1:0]        offsetRecord_45;
  reg  [1:0]        offsetRecord_46;
  reg  [1:0]        offsetRecord_47;
  reg  [1:0]        offsetRecord_48;
  reg  [1:0]        offsetRecord_49;
  reg  [1:0]        offsetRecord_50;
  reg  [1:0]        offsetRecord_51;
  reg  [1:0]        offsetRecord_52;
  reg  [1:0]        offsetRecord_53;
  reg  [1:0]        offsetRecord_54;
  reg  [1:0]        offsetRecord_55;
  reg  [1:0]        offsetRecord_56;
  reg  [1:0]        offsetRecord_57;
  reg  [1:0]        offsetRecord_58;
  reg  [1:0]        offsetRecord_59;
  reg  [1:0]        offsetRecord_60;
  reg  [1:0]        offsetRecord_61;
  reg  [1:0]        offsetRecord_62;
  reg  [1:0]        offsetRecord_63;
  reg  [1:0]        offsetRecord_64;
  reg  [1:0]        offsetRecord_65;
  reg  [1:0]        offsetRecord_66;
  reg  [1:0]        offsetRecord_67;
  reg  [1:0]        offsetRecord_68;
  reg  [1:0]        offsetRecord_69;
  reg  [1:0]        offsetRecord_70;
  reg  [1:0]        offsetRecord_71;
  reg  [1:0]        offsetRecord_72;
  reg  [1:0]        offsetRecord_73;
  reg  [1:0]        offsetRecord_74;
  reg  [1:0]        offsetRecord_75;
  reg  [1:0]        offsetRecord_76;
  reg  [1:0]        offsetRecord_77;
  reg  [1:0]        offsetRecord_78;
  reg  [1:0]        offsetRecord_79;
  reg  [1:0]        offsetRecord_80;
  reg  [1:0]        offsetRecord_81;
  reg  [1:0]        offsetRecord_82;
  reg  [1:0]        offsetRecord_83;
  reg  [1:0]        offsetRecord_84;
  reg  [1:0]        offsetRecord_85;
  reg  [1:0]        offsetRecord_86;
  reg  [1:0]        offsetRecord_87;
  reg  [1:0]        offsetRecord_88;
  reg  [1:0]        offsetRecord_89;
  reg  [1:0]        offsetRecord_90;
  reg  [1:0]        offsetRecord_91;
  reg  [1:0]        offsetRecord_92;
  reg  [1:0]        offsetRecord_93;
  reg  [1:0]        offsetRecord_94;
  reg  [1:0]        offsetRecord_95;
  reg  [1:0]        offsetRecord_96;
  reg  [1:0]        offsetRecord_97;
  reg  [1:0]        offsetRecord_98;
  reg  [1:0]        offsetRecord_99;
  reg  [1:0]        offsetRecord_100;
  reg  [1:0]        offsetRecord_101;
  reg  [1:0]        offsetRecord_102;
  reg  [1:0]        offsetRecord_103;
  reg  [1:0]        offsetRecord_104;
  reg  [1:0]        offsetRecord_105;
  reg  [1:0]        offsetRecord_106;
  reg  [1:0]        offsetRecord_107;
  reg  [1:0]        offsetRecord_108;
  reg  [1:0]        offsetRecord_109;
  reg  [1:0]        offsetRecord_110;
  reg  [1:0]        offsetRecord_111;
  reg  [1:0]        offsetRecord_112;
  reg  [1:0]        offsetRecord_113;
  reg  [1:0]        offsetRecord_114;
  reg  [1:0]        offsetRecord_115;
  reg  [1:0]        offsetRecord_116;
  reg  [1:0]        offsetRecord_117;
  reg  [1:0]        offsetRecord_118;
  reg  [1:0]        offsetRecord_119;
  reg  [1:0]        offsetRecord_120;
  reg  [1:0]        offsetRecord_121;
  reg  [1:0]        offsetRecord_122;
  reg  [1:0]        offsetRecord_123;
  reg  [1:0]        offsetRecord_124;
  reg  [1:0]        offsetRecord_125;
  reg  [1:0]        offsetRecord_126;
  reg  [1:0]        offsetRecord_127;
  wire [6:0]        indexInMaskGroupResponse = isSegmentLoadStore ? memReadResponse_bits_source_0[9:3] : memReadResponse_bits_source_0[6:0];
  wire [127:0]      responseSourceLSBOH = 128'h1 << memReadResponse_bits_source_0[6:0];
  wire [14:0]       loadBaseByteOffset = {3'h0, groupIndex, indexInMaskGroupResponse} << _GEN_16;
  wire [127:0][1:0] _GEN_18 =
    {{offsetRecord_127},
     {offsetRecord_126},
     {offsetRecord_125},
     {offsetRecord_124},
     {offsetRecord_123},
     {offsetRecord_122},
     {offsetRecord_121},
     {offsetRecord_120},
     {offsetRecord_119},
     {offsetRecord_118},
     {offsetRecord_117},
     {offsetRecord_116},
     {offsetRecord_115},
     {offsetRecord_114},
     {offsetRecord_113},
     {offsetRecord_112},
     {offsetRecord_111},
     {offsetRecord_110},
     {offsetRecord_109},
     {offsetRecord_108},
     {offsetRecord_107},
     {offsetRecord_106},
     {offsetRecord_105},
     {offsetRecord_104},
     {offsetRecord_103},
     {offsetRecord_102},
     {offsetRecord_101},
     {offsetRecord_100},
     {offsetRecord_99},
     {offsetRecord_98},
     {offsetRecord_97},
     {offsetRecord_96},
     {offsetRecord_95},
     {offsetRecord_94},
     {offsetRecord_93},
     {offsetRecord_92},
     {offsetRecord_91},
     {offsetRecord_90},
     {offsetRecord_89},
     {offsetRecord_88},
     {offsetRecord_87},
     {offsetRecord_86},
     {offsetRecord_85},
     {offsetRecord_84},
     {offsetRecord_83},
     {offsetRecord_82},
     {offsetRecord_81},
     {offsetRecord_80},
     {offsetRecord_79},
     {offsetRecord_78},
     {offsetRecord_77},
     {offsetRecord_76},
     {offsetRecord_75},
     {offsetRecord_74},
     {offsetRecord_73},
     {offsetRecord_72},
     {offsetRecord_71},
     {offsetRecord_70},
     {offsetRecord_69},
     {offsetRecord_68},
     {offsetRecord_67},
     {offsetRecord_66},
     {offsetRecord_65},
     {offsetRecord_64},
     {offsetRecord_63},
     {offsetRecord_62},
     {offsetRecord_61},
     {offsetRecord_60},
     {offsetRecord_59},
     {offsetRecord_58},
     {offsetRecord_57},
     {offsetRecord_56},
     {offsetRecord_55},
     {offsetRecord_54},
     {offsetRecord_53},
     {offsetRecord_52},
     {offsetRecord_51},
     {offsetRecord_50},
     {offsetRecord_49},
     {offsetRecord_48},
     {offsetRecord_47},
     {offsetRecord_46},
     {offsetRecord_45},
     {offsetRecord_44},
     {offsetRecord_43},
     {offsetRecord_42},
     {offsetRecord_41},
     {offsetRecord_40},
     {offsetRecord_39},
     {offsetRecord_38},
     {offsetRecord_37},
     {offsetRecord_36},
     {offsetRecord_35},
     {offsetRecord_34},
     {offsetRecord_33},
     {offsetRecord_32},
     {offsetRecord_31},
     {offsetRecord_30},
     {offsetRecord_29},
     {offsetRecord_28},
     {offsetRecord_27},
     {offsetRecord_26},
     {offsetRecord_25},
     {offsetRecord_24},
     {offsetRecord_23},
     {offsetRecord_22},
     {offsetRecord_21},
     {offsetRecord_20},
     {offsetRecord_19},
     {offsetRecord_18},
     {offsetRecord_17},
     {offsetRecord_16},
     {offsetRecord_15},
     {offsetRecord_14},
     {offsetRecord_13},
     {offsetRecord_12},
     {offsetRecord_11},
     {offsetRecord_10},
     {offsetRecord_9},
     {offsetRecord_8},
     {offsetRecord_7},
     {offsetRecord_6},
     {offsetRecord_5},
     {offsetRecord_4},
     {offsetRecord_3},
     {offsetRecord_2},
     {offsetRecord_1},
     {offsetRecord_0}};
  wire [4:0]        addressOffset = {_GEN_18[memReadResponse_bits_source_0[6:0]], 3'h0};
  wire [62:0]       _vrfWritePort_bits_data_T_3 = {31'h0, memReadResponse_bits_data_0 >> addressOffset} << {58'h0, loadBaseByteOffset[1:0], 3'h0};
  wire [31:0]       vrfWritePort_bits_data_0 = _vrfWritePort_bits_data_T_3[31:0];
  wire [3:0]        vrfWritePort_bits_mask_0 = (dataEEWOH[0] ? 4'h1 << loadBaseByteOffset[1:0] : 4'h0) | (dataEEWOH[1] ? {{2{loadBaseByteOffset[1]}}, ~(loadBaseByteOffset[1]), ~(loadBaseByteOffset[1])} : 4'h0) | {4{dataEEWOH[2]}};
  wire [4:0]        vrfWritePort_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + (isSegmentLoadStore ? {2'h0, memReadResponse_bits_source_0[2:0]} * _GEN_17 : 5'h0) + {2'h0, loadBaseByteOffset[10:8]};
  assign writeOffset = loadBaseByteOffset[7];
  wire              vrfWritePort_bits_offset_0 = writeOffset;
  wire              _GEN_19 = state == 2'h2 & noOutstandingMessages & pipelineClear & ~memReadResponse_valid_0;
  wire              invalidInstruction = csrInterface_vl == 12'h0 & ~requestIsWholeRegisterLoadStore & lsuRequest_valid;
  reg               invalidInstructionNext;
  assign stateIdle = state == 2'h0;
  wire              allElementsMasked =
    stateIdle
    & (_allElementsMasked_T_1 | _allElementsMasked_T_2 | _allElementsMasked_T_3 | _allElementsMasked_T_4 | _allElementsMasked_T_5 | _allElementsMasked_T_6 | _allElementsMasked_T_7 | _allElementsMasked_T_8 | _allElementsMasked_T_9
       | _allElementsMasked_T_10 | _allElementsMasked_T_11 | _allElementsMasked_T_12 | _allElementsMasked_T_13 | _allElementsMasked_T_14 | _allElementsMasked_T_15 | _allElementsMasked_T_16 | _allElementsMasked_T_17 | _allElementsMasked_T_18
       | _allElementsMasked_T_19 | _allElementsMasked_T_20 | _allElementsMasked_T_21 | _allElementsMasked_T_22 | _allElementsMasked_T_23 | _allElementsMasked_T_24 | _allElementsMasked_T_25 | _allElementsMasked_T_26 | _allElementsMasked_T_27
       | _allElementsMasked_T_28 | _allElementsMasked_T_29 | _allElementsMasked_T_30 | _allElementsMasked_T_31 | _allElementsMasked_T_32);
  wire              _GEN_26 = lsuRequest_valid & ~invalidInstruction;
  wire              updateOffsetGroupEnable = _GEN_26 | _GEN_19 & ~last;
  reg               status_last_REG;
  wire              _status_last_output = ~status_last_REG & stateIdle | invalidInstructionNext | allElementsMasked;
  wire [9:0]        _dataOffset_T = {3'h0, s1EnqQueue_deq_bits_indexInMaskGroup} << dataEEW;
  wire [4:0]        dataOffset = {_dataOffset_T[1:0], 3'h0};
  wire [31:0]       offsetQueueVec_0_deq_bits;
  wire [31:0]       offsetQueueVec_1_deq_bits;
  wire [31:0]       offsetQueueVec_2_deq_bits;
  wire [31:0]       offsetQueueVec_3_deq_bits;
  wire [31:0]       offsetQueueVec_4_deq_bits;
  wire [31:0]       offsetQueueVec_5_deq_bits;
  wire [31:0]       offsetQueueVec_6_deq_bits;
  wire [31:0]       offsetQueueVec_7_deq_bits;
  wire [31:0]       offsetQueueVec_8_deq_bits;
  wire [31:0]       offsetQueueVec_9_deq_bits;
  wire [31:0]       offsetQueueVec_10_deq_bits;
  wire [31:0]       offsetQueueVec_11_deq_bits;
  wire [31:0]       offsetQueueVec_12_deq_bits;
  wire [31:0]       offsetQueueVec_13_deq_bits;
  wire [31:0]       offsetQueueVec_14_deq_bits;
  wire [31:0]       offsetQueueVec_15_deq_bits;
  wire [31:0]       offsetQueueVec_16_deq_bits;
  wire [31:0]       offsetQueueVec_17_deq_bits;
  wire [31:0]       offsetQueueVec_18_deq_bits;
  wire [31:0]       offsetQueueVec_19_deq_bits;
  wire [31:0]       offsetQueueVec_20_deq_bits;
  wire [31:0]       offsetQueueVec_21_deq_bits;
  wire [31:0]       offsetQueueVec_22_deq_bits;
  wire [31:0]       offsetQueueVec_23_deq_bits;
  wire [31:0]       offsetQueueVec_24_deq_bits;
  wire [31:0]       offsetQueueVec_25_deq_bits;
  wire [31:0]       offsetQueueVec_26_deq_bits;
  wire [31:0]       offsetQueueVec_27_deq_bits;
  wire [31:0]       offsetQueueVec_28_deq_bits;
  wire [31:0]       offsetQueueVec_29_deq_bits;
  wire [31:0]       offsetQueueVec_30_deq_bits;
  wire [31:0]       offsetQueueVec_31_deq_bits;
  always @(posedge clock) begin
    if (reset) begin
      offsetQueueVec_deqLock <= 1'h0;
      offsetQueueVec_deqLock_1 <= 1'h0;
      offsetQueueVec_deqLock_2 <= 1'h0;
      offsetQueueVec_deqLock_3 <= 1'h0;
      offsetQueueVec_deqLock_4 <= 1'h0;
      offsetQueueVec_deqLock_5 <= 1'h0;
      offsetQueueVec_deqLock_6 <= 1'h0;
      offsetQueueVec_deqLock_7 <= 1'h0;
      offsetQueueVec_deqLock_8 <= 1'h0;
      offsetQueueVec_deqLock_9 <= 1'h0;
      offsetQueueVec_deqLock_10 <= 1'h0;
      offsetQueueVec_deqLock_11 <= 1'h0;
      offsetQueueVec_deqLock_12 <= 1'h0;
      offsetQueueVec_deqLock_13 <= 1'h0;
      offsetQueueVec_deqLock_14 <= 1'h0;
      offsetQueueVec_deqLock_15 <= 1'h0;
      offsetQueueVec_deqLock_16 <= 1'h0;
      offsetQueueVec_deqLock_17 <= 1'h0;
      offsetQueueVec_deqLock_18 <= 1'h0;
      offsetQueueVec_deqLock_19 <= 1'h0;
      offsetQueueVec_deqLock_20 <= 1'h0;
      offsetQueueVec_deqLock_21 <= 1'h0;
      offsetQueueVec_deqLock_22 <= 1'h0;
      offsetQueueVec_deqLock_23 <= 1'h0;
      offsetQueueVec_deqLock_24 <= 1'h0;
      offsetQueueVec_deqLock_25 <= 1'h0;
      offsetQueueVec_deqLock_26 <= 1'h0;
      offsetQueueVec_deqLock_27 <= 1'h0;
      offsetQueueVec_deqLock_28 <= 1'h0;
      offsetQueueVec_deqLock_29 <= 1'h0;
      offsetQueueVec_deqLock_30 <= 1'h0;
      offsetQueueVec_deqLock_31 <= 1'h0;
      lsuRequestReg_instructionInformation_nf <= 3'h0;
      lsuRequestReg_instructionInformation_mew <= 1'h0;
      lsuRequestReg_instructionInformation_mop <= 2'h0;
      lsuRequestReg_instructionInformation_lumop <= 5'h0;
      lsuRequestReg_instructionInformation_eew <= 2'h0;
      lsuRequestReg_instructionInformation_vs3 <= 5'h0;
      lsuRequestReg_instructionInformation_isStore <= 1'h0;
      lsuRequestReg_instructionInformation_maskedLoadStore <= 1'h0;
      lsuRequestReg_rs1Data <= 32'h0;
      lsuRequestReg_rs2Data <= 32'h0;
      lsuRequestReg_instructionIndex <= 3'h0;
      csrInterfaceReg_vl <= 12'h0;
      csrInterfaceReg_vStart <= 12'h0;
      csrInterfaceReg_vlmul <= 3'h0;
      csrInterfaceReg_vSew <= 2'h0;
      csrInterfaceReg_vxrm <= 2'h0;
      csrInterfaceReg_vta <= 1'h0;
      csrInterfaceReg_vma <= 1'h0;
      dataWidthForSegmentLoadStore <= 7'h0;
      elementByteWidth <= 3'h0;
      segmentInstructionIndexInterval <= 4'h0;
      outstandingTLDMessages <= 128'h0;
      indexedInstructionOffsets_0_valid <= 1'h0;
      indexedInstructionOffsets_0_bits <= 32'h0;
      indexedInstructionOffsets_1_valid <= 1'h0;
      indexedInstructionOffsets_1_bits <= 32'h0;
      indexedInstructionOffsets_2_valid <= 1'h0;
      indexedInstructionOffsets_2_bits <= 32'h0;
      indexedInstructionOffsets_3_valid <= 1'h0;
      indexedInstructionOffsets_3_bits <= 32'h0;
      indexedInstructionOffsets_4_valid <= 1'h0;
      indexedInstructionOffsets_4_bits <= 32'h0;
      indexedInstructionOffsets_5_valid <= 1'h0;
      indexedInstructionOffsets_5_bits <= 32'h0;
      indexedInstructionOffsets_6_valid <= 1'h0;
      indexedInstructionOffsets_6_bits <= 32'h0;
      indexedInstructionOffsets_7_valid <= 1'h0;
      indexedInstructionOffsets_7_bits <= 32'h0;
      indexedInstructionOffsets_8_valid <= 1'h0;
      indexedInstructionOffsets_8_bits <= 32'h0;
      indexedInstructionOffsets_9_valid <= 1'h0;
      indexedInstructionOffsets_9_bits <= 32'h0;
      indexedInstructionOffsets_10_valid <= 1'h0;
      indexedInstructionOffsets_10_bits <= 32'h0;
      indexedInstructionOffsets_11_valid <= 1'h0;
      indexedInstructionOffsets_11_bits <= 32'h0;
      indexedInstructionOffsets_12_valid <= 1'h0;
      indexedInstructionOffsets_12_bits <= 32'h0;
      indexedInstructionOffsets_13_valid <= 1'h0;
      indexedInstructionOffsets_13_bits <= 32'h0;
      indexedInstructionOffsets_14_valid <= 1'h0;
      indexedInstructionOffsets_14_bits <= 32'h0;
      indexedInstructionOffsets_15_valid <= 1'h0;
      indexedInstructionOffsets_15_bits <= 32'h0;
      indexedInstructionOffsets_16_valid <= 1'h0;
      indexedInstructionOffsets_16_bits <= 32'h0;
      indexedInstructionOffsets_17_valid <= 1'h0;
      indexedInstructionOffsets_17_bits <= 32'h0;
      indexedInstructionOffsets_18_valid <= 1'h0;
      indexedInstructionOffsets_18_bits <= 32'h0;
      indexedInstructionOffsets_19_valid <= 1'h0;
      indexedInstructionOffsets_19_bits <= 32'h0;
      indexedInstructionOffsets_20_valid <= 1'h0;
      indexedInstructionOffsets_20_bits <= 32'h0;
      indexedInstructionOffsets_21_valid <= 1'h0;
      indexedInstructionOffsets_21_bits <= 32'h0;
      indexedInstructionOffsets_22_valid <= 1'h0;
      indexedInstructionOffsets_22_bits <= 32'h0;
      indexedInstructionOffsets_23_valid <= 1'h0;
      indexedInstructionOffsets_23_bits <= 32'h0;
      indexedInstructionOffsets_24_valid <= 1'h0;
      indexedInstructionOffsets_24_bits <= 32'h0;
      indexedInstructionOffsets_25_valid <= 1'h0;
      indexedInstructionOffsets_25_bits <= 32'h0;
      indexedInstructionOffsets_26_valid <= 1'h0;
      indexedInstructionOffsets_26_bits <= 32'h0;
      indexedInstructionOffsets_27_valid <= 1'h0;
      indexedInstructionOffsets_27_bits <= 32'h0;
      indexedInstructionOffsets_28_valid <= 1'h0;
      indexedInstructionOffsets_28_bits <= 32'h0;
      indexedInstructionOffsets_29_valid <= 1'h0;
      indexedInstructionOffsets_29_bits <= 32'h0;
      indexedInstructionOffsets_30_valid <= 1'h0;
      indexedInstructionOffsets_30_bits <= 32'h0;
      indexedInstructionOffsets_31_valid <= 1'h0;
      indexedInstructionOffsets_31_bits <= 32'h0;
      groupIndex <= 5'h0;
      maskReg <= 128'h0;
      segmentIndex <= 3'h0;
      state <= 2'h0;
      sentMemoryRequests <= 128'h0;
      firstMemoryRequestOfInstruction <= 1'h0;
      waitFirstMemoryResponseForFaultOnlyFirst <= 1'h0;
      s0Valid <= 1'h0;
      s0Reg_readVS <= 5'h0;
      s0Reg_offsetForVSInLane <= 1'h0;
      s0Reg_addressOffset <= 32'h0;
      s0Reg_segmentIndex <= 3'h0;
      s0Reg_offsetForLane <= 5'h0;
      s0Reg_indexInGroup <= 7'h0;
      s1Valid <= 1'h0;
      s1Reg_indexInMaskGroup <= 7'h0;
      s1Reg_segmentIndex <= 3'h0;
      s1Reg_address <= 32'h0;
      s1Reg_readData <= 32'h0;
      offsetRecord_0 <= 2'h0;
      offsetRecord_1 <= 2'h0;
      offsetRecord_2 <= 2'h0;
      offsetRecord_3 <= 2'h0;
      offsetRecord_4 <= 2'h0;
      offsetRecord_5 <= 2'h0;
      offsetRecord_6 <= 2'h0;
      offsetRecord_7 <= 2'h0;
      offsetRecord_8 <= 2'h0;
      offsetRecord_9 <= 2'h0;
      offsetRecord_10 <= 2'h0;
      offsetRecord_11 <= 2'h0;
      offsetRecord_12 <= 2'h0;
      offsetRecord_13 <= 2'h0;
      offsetRecord_14 <= 2'h0;
      offsetRecord_15 <= 2'h0;
      offsetRecord_16 <= 2'h0;
      offsetRecord_17 <= 2'h0;
      offsetRecord_18 <= 2'h0;
      offsetRecord_19 <= 2'h0;
      offsetRecord_20 <= 2'h0;
      offsetRecord_21 <= 2'h0;
      offsetRecord_22 <= 2'h0;
      offsetRecord_23 <= 2'h0;
      offsetRecord_24 <= 2'h0;
      offsetRecord_25 <= 2'h0;
      offsetRecord_26 <= 2'h0;
      offsetRecord_27 <= 2'h0;
      offsetRecord_28 <= 2'h0;
      offsetRecord_29 <= 2'h0;
      offsetRecord_30 <= 2'h0;
      offsetRecord_31 <= 2'h0;
      offsetRecord_32 <= 2'h0;
      offsetRecord_33 <= 2'h0;
      offsetRecord_34 <= 2'h0;
      offsetRecord_35 <= 2'h0;
      offsetRecord_36 <= 2'h0;
      offsetRecord_37 <= 2'h0;
      offsetRecord_38 <= 2'h0;
      offsetRecord_39 <= 2'h0;
      offsetRecord_40 <= 2'h0;
      offsetRecord_41 <= 2'h0;
      offsetRecord_42 <= 2'h0;
      offsetRecord_43 <= 2'h0;
      offsetRecord_44 <= 2'h0;
      offsetRecord_45 <= 2'h0;
      offsetRecord_46 <= 2'h0;
      offsetRecord_47 <= 2'h0;
      offsetRecord_48 <= 2'h0;
      offsetRecord_49 <= 2'h0;
      offsetRecord_50 <= 2'h0;
      offsetRecord_51 <= 2'h0;
      offsetRecord_52 <= 2'h0;
      offsetRecord_53 <= 2'h0;
      offsetRecord_54 <= 2'h0;
      offsetRecord_55 <= 2'h0;
      offsetRecord_56 <= 2'h0;
      offsetRecord_57 <= 2'h0;
      offsetRecord_58 <= 2'h0;
      offsetRecord_59 <= 2'h0;
      offsetRecord_60 <= 2'h0;
      offsetRecord_61 <= 2'h0;
      offsetRecord_62 <= 2'h0;
      offsetRecord_63 <= 2'h0;
      offsetRecord_64 <= 2'h0;
      offsetRecord_65 <= 2'h0;
      offsetRecord_66 <= 2'h0;
      offsetRecord_67 <= 2'h0;
      offsetRecord_68 <= 2'h0;
      offsetRecord_69 <= 2'h0;
      offsetRecord_70 <= 2'h0;
      offsetRecord_71 <= 2'h0;
      offsetRecord_72 <= 2'h0;
      offsetRecord_73 <= 2'h0;
      offsetRecord_74 <= 2'h0;
      offsetRecord_75 <= 2'h0;
      offsetRecord_76 <= 2'h0;
      offsetRecord_77 <= 2'h0;
      offsetRecord_78 <= 2'h0;
      offsetRecord_79 <= 2'h0;
      offsetRecord_80 <= 2'h0;
      offsetRecord_81 <= 2'h0;
      offsetRecord_82 <= 2'h0;
      offsetRecord_83 <= 2'h0;
      offsetRecord_84 <= 2'h0;
      offsetRecord_85 <= 2'h0;
      offsetRecord_86 <= 2'h0;
      offsetRecord_87 <= 2'h0;
      offsetRecord_88 <= 2'h0;
      offsetRecord_89 <= 2'h0;
      offsetRecord_90 <= 2'h0;
      offsetRecord_91 <= 2'h0;
      offsetRecord_92 <= 2'h0;
      offsetRecord_93 <= 2'h0;
      offsetRecord_94 <= 2'h0;
      offsetRecord_95 <= 2'h0;
      offsetRecord_96 <= 2'h0;
      offsetRecord_97 <= 2'h0;
      offsetRecord_98 <= 2'h0;
      offsetRecord_99 <= 2'h0;
      offsetRecord_100 <= 2'h0;
      offsetRecord_101 <= 2'h0;
      offsetRecord_102 <= 2'h0;
      offsetRecord_103 <= 2'h0;
      offsetRecord_104 <= 2'h0;
      offsetRecord_105 <= 2'h0;
      offsetRecord_106 <= 2'h0;
      offsetRecord_107 <= 2'h0;
      offsetRecord_108 <= 2'h0;
      offsetRecord_109 <= 2'h0;
      offsetRecord_110 <= 2'h0;
      offsetRecord_111 <= 2'h0;
      offsetRecord_112 <= 2'h0;
      offsetRecord_113 <= 2'h0;
      offsetRecord_114 <= 2'h0;
      offsetRecord_115 <= 2'h0;
      offsetRecord_116 <= 2'h0;
      offsetRecord_117 <= 2'h0;
      offsetRecord_118 <= 2'h0;
      offsetRecord_119 <= 2'h0;
      offsetRecord_120 <= 2'h0;
      offsetRecord_121 <= 2'h0;
      offsetRecord_122 <= 2'h0;
      offsetRecord_123 <= 2'h0;
      offsetRecord_124 <= 2'h0;
      offsetRecord_125 <= 2'h0;
      offsetRecord_126 <= 2'h0;
      offsetRecord_127 <= 2'h0;
    end
    else begin
      automatic logic _offsetQueueVec_T_93 = lsuRequest_valid | requestOffset;
      automatic logic _outstandingTLDMessages_T;
      _outstandingTLDMessages_T = memReadResponse_ready_0 & memReadResponse_valid_0;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_1)
        offsetQueueVec_deqLock <= _allElementsMasked_T_1;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_2)
        offsetQueueVec_deqLock_1 <= _allElementsMasked_T_2;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_3)
        offsetQueueVec_deqLock_2 <= _allElementsMasked_T_3;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_4)
        offsetQueueVec_deqLock_3 <= _allElementsMasked_T_4;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_5)
        offsetQueueVec_deqLock_4 <= _allElementsMasked_T_5;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_6)
        offsetQueueVec_deqLock_5 <= _allElementsMasked_T_6;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_7)
        offsetQueueVec_deqLock_6 <= _allElementsMasked_T_7;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_8)
        offsetQueueVec_deqLock_7 <= _allElementsMasked_T_8;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_9)
        offsetQueueVec_deqLock_8 <= _allElementsMasked_T_9;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_10)
        offsetQueueVec_deqLock_9 <= _allElementsMasked_T_10;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_11)
        offsetQueueVec_deqLock_10 <= _allElementsMasked_T_11;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_12)
        offsetQueueVec_deqLock_11 <= _allElementsMasked_T_12;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_13)
        offsetQueueVec_deqLock_12 <= _allElementsMasked_T_13;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_14)
        offsetQueueVec_deqLock_13 <= _allElementsMasked_T_14;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_15)
        offsetQueueVec_deqLock_14 <= _allElementsMasked_T_15;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_16)
        offsetQueueVec_deqLock_15 <= _allElementsMasked_T_16;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_17)
        offsetQueueVec_deqLock_16 <= _allElementsMasked_T_17;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_18)
        offsetQueueVec_deqLock_17 <= _allElementsMasked_T_18;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_19)
        offsetQueueVec_deqLock_18 <= _allElementsMasked_T_19;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_20)
        offsetQueueVec_deqLock_19 <= _allElementsMasked_T_20;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_21)
        offsetQueueVec_deqLock_20 <= _allElementsMasked_T_21;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_22)
        offsetQueueVec_deqLock_21 <= _allElementsMasked_T_22;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_23)
        offsetQueueVec_deqLock_22 <= _allElementsMasked_T_23;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_24)
        offsetQueueVec_deqLock_23 <= _allElementsMasked_T_24;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_25)
        offsetQueueVec_deqLock_24 <= _allElementsMasked_T_25;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_26)
        offsetQueueVec_deqLock_25 <= _allElementsMasked_T_26;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_27)
        offsetQueueVec_deqLock_26 <= _allElementsMasked_T_27;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_28)
        offsetQueueVec_deqLock_27 <= _allElementsMasked_T_28;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_29)
        offsetQueueVec_deqLock_28 <= _allElementsMasked_T_29;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_30)
        offsetQueueVec_deqLock_29 <= _allElementsMasked_T_30;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_31)
        offsetQueueVec_deqLock_30 <= _allElementsMasked_T_31;
      if (_offsetQueueVec_T_93 | _allElementsMasked_T_32)
        offsetQueueVec_deqLock_31 <= _allElementsMasked_T_32;
      if (lsuRequest_valid) begin
        automatic logic [3:0] _elementByteWidth_T = 4'h1 << requestEEW;
        lsuRequestReg_instructionInformation_nf <= lsuRequest_bits_instructionInformation_nf;
        lsuRequestReg_instructionInformation_mew <= lsuRequest_bits_instructionInformation_mew;
        lsuRequestReg_instructionInformation_mop <= lsuRequest_bits_instructionInformation_mop;
        lsuRequestReg_instructionInformation_lumop <= lsuRequest_bits_instructionInformation_lumop;
        lsuRequestReg_instructionInformation_eew <= lsuRequest_bits_instructionInformation_eew;
        lsuRequestReg_instructionInformation_vs3 <= lsuRequest_bits_instructionInformation_vs3;
        lsuRequestReg_instructionInformation_isStore <= lsuRequest_bits_instructionInformation_isStore;
        lsuRequestReg_instructionInformation_maskedLoadStore <= lsuRequest_bits_instructionInformation_maskedLoadStore;
        lsuRequestReg_rs1Data <= lsuRequest_bits_rs1Data;
        lsuRequestReg_rs2Data <= lsuRequest_bits_rs2Data;
        lsuRequestReg_instructionIndex <= lsuRequest_bits_instructionIndex;
        csrInterfaceReg_vl <= csrInterface_vl;
        csrInterfaceReg_vStart <= csrInterface_vStart;
        csrInterfaceReg_vlmul <= csrInterface_vlmul;
        csrInterfaceReg_vSew <= csrInterface_vSew;
        csrInterfaceReg_vxrm <= csrInterface_vxrm;
        csrInterfaceReg_vta <= csrInterface_vta;
        csrInterfaceReg_vma <= csrInterface_vma;
        dataWidthForSegmentLoadStore <= {3'h0, {1'h0, requestNF} + 4'h1} * {4'h0, _elementByteWidth_T[2:0]};
        elementByteWidth <= _elementByteWidth_T[2:0];
        segmentInstructionIndexInterval <= csrInterface_vlmul[2] ? 4'h1 : 4'h1 << csrInterface_vlmul[1:0];
      end
      if ((_outstandingTLDMessages_T | _outstandingTLDMessages_T_4) & ~lsuRequestReg_instructionInformation_isStore)
        outstandingTLDMessages <= outstandingTLDMessages & ~(_outstandingTLDMessages_T ? responseSourceLSBOH : 128'h0) | (_outstandingTLDMessages_T_4 ? memoryRequestSourceOH : 128'h0);
      indexedInstructionOffsets_0_valid <= _allElementsMasked_T_1 | indexedInstructionOffsets_0_valid & ~usedIndexedInstructionOffsets_0 & ~_status_last_output;
      if (_allElementsMasked_T_1)
        indexedInstructionOffsets_0_bits <= offsetQueueVec_0_deq_bits;
      indexedInstructionOffsets_1_valid <= _allElementsMasked_T_2 | indexedInstructionOffsets_1_valid & ~usedIndexedInstructionOffsets_1 & ~_status_last_output;
      if (_allElementsMasked_T_2)
        indexedInstructionOffsets_1_bits <= offsetQueueVec_1_deq_bits;
      indexedInstructionOffsets_2_valid <= _allElementsMasked_T_3 | indexedInstructionOffsets_2_valid & ~usedIndexedInstructionOffsets_2 & ~_status_last_output;
      if (_allElementsMasked_T_3)
        indexedInstructionOffsets_2_bits <= offsetQueueVec_2_deq_bits;
      indexedInstructionOffsets_3_valid <= _allElementsMasked_T_4 | indexedInstructionOffsets_3_valid & ~usedIndexedInstructionOffsets_3 & ~_status_last_output;
      if (_allElementsMasked_T_4)
        indexedInstructionOffsets_3_bits <= offsetQueueVec_3_deq_bits;
      indexedInstructionOffsets_4_valid <= _allElementsMasked_T_5 | indexedInstructionOffsets_4_valid & ~usedIndexedInstructionOffsets_4 & ~_status_last_output;
      if (_allElementsMasked_T_5)
        indexedInstructionOffsets_4_bits <= offsetQueueVec_4_deq_bits;
      indexedInstructionOffsets_5_valid <= _allElementsMasked_T_6 | indexedInstructionOffsets_5_valid & ~usedIndexedInstructionOffsets_5 & ~_status_last_output;
      if (_allElementsMasked_T_6)
        indexedInstructionOffsets_5_bits <= offsetQueueVec_5_deq_bits;
      indexedInstructionOffsets_6_valid <= _allElementsMasked_T_7 | indexedInstructionOffsets_6_valid & ~usedIndexedInstructionOffsets_6 & ~_status_last_output;
      if (_allElementsMasked_T_7)
        indexedInstructionOffsets_6_bits <= offsetQueueVec_6_deq_bits;
      indexedInstructionOffsets_7_valid <= _allElementsMasked_T_8 | indexedInstructionOffsets_7_valid & ~usedIndexedInstructionOffsets_7 & ~_status_last_output;
      if (_allElementsMasked_T_8)
        indexedInstructionOffsets_7_bits <= offsetQueueVec_7_deq_bits;
      indexedInstructionOffsets_8_valid <= _allElementsMasked_T_9 | indexedInstructionOffsets_8_valid & ~usedIndexedInstructionOffsets_8 & ~_status_last_output;
      if (_allElementsMasked_T_9)
        indexedInstructionOffsets_8_bits <= offsetQueueVec_8_deq_bits;
      indexedInstructionOffsets_9_valid <= _allElementsMasked_T_10 | indexedInstructionOffsets_9_valid & ~usedIndexedInstructionOffsets_9 & ~_status_last_output;
      if (_allElementsMasked_T_10)
        indexedInstructionOffsets_9_bits <= offsetQueueVec_9_deq_bits;
      indexedInstructionOffsets_10_valid <= _allElementsMasked_T_11 | indexedInstructionOffsets_10_valid & ~usedIndexedInstructionOffsets_10 & ~_status_last_output;
      if (_allElementsMasked_T_11)
        indexedInstructionOffsets_10_bits <= offsetQueueVec_10_deq_bits;
      indexedInstructionOffsets_11_valid <= _allElementsMasked_T_12 | indexedInstructionOffsets_11_valid & ~usedIndexedInstructionOffsets_11 & ~_status_last_output;
      if (_allElementsMasked_T_12)
        indexedInstructionOffsets_11_bits <= offsetQueueVec_11_deq_bits;
      indexedInstructionOffsets_12_valid <= _allElementsMasked_T_13 | indexedInstructionOffsets_12_valid & ~usedIndexedInstructionOffsets_12 & ~_status_last_output;
      if (_allElementsMasked_T_13)
        indexedInstructionOffsets_12_bits <= offsetQueueVec_12_deq_bits;
      indexedInstructionOffsets_13_valid <= _allElementsMasked_T_14 | indexedInstructionOffsets_13_valid & ~usedIndexedInstructionOffsets_13 & ~_status_last_output;
      if (_allElementsMasked_T_14)
        indexedInstructionOffsets_13_bits <= offsetQueueVec_13_deq_bits;
      indexedInstructionOffsets_14_valid <= _allElementsMasked_T_15 | indexedInstructionOffsets_14_valid & ~usedIndexedInstructionOffsets_14 & ~_status_last_output;
      if (_allElementsMasked_T_15)
        indexedInstructionOffsets_14_bits <= offsetQueueVec_14_deq_bits;
      indexedInstructionOffsets_15_valid <= _allElementsMasked_T_16 | indexedInstructionOffsets_15_valid & ~usedIndexedInstructionOffsets_15 & ~_status_last_output;
      if (_allElementsMasked_T_16)
        indexedInstructionOffsets_15_bits <= offsetQueueVec_15_deq_bits;
      indexedInstructionOffsets_16_valid <= _allElementsMasked_T_17 | indexedInstructionOffsets_16_valid & ~usedIndexedInstructionOffsets_16 & ~_status_last_output;
      if (_allElementsMasked_T_17)
        indexedInstructionOffsets_16_bits <= offsetQueueVec_16_deq_bits;
      indexedInstructionOffsets_17_valid <= _allElementsMasked_T_18 | indexedInstructionOffsets_17_valid & ~usedIndexedInstructionOffsets_17 & ~_status_last_output;
      if (_allElementsMasked_T_18)
        indexedInstructionOffsets_17_bits <= offsetQueueVec_17_deq_bits;
      indexedInstructionOffsets_18_valid <= _allElementsMasked_T_19 | indexedInstructionOffsets_18_valid & ~usedIndexedInstructionOffsets_18 & ~_status_last_output;
      if (_allElementsMasked_T_19)
        indexedInstructionOffsets_18_bits <= offsetQueueVec_18_deq_bits;
      indexedInstructionOffsets_19_valid <= _allElementsMasked_T_20 | indexedInstructionOffsets_19_valid & ~usedIndexedInstructionOffsets_19 & ~_status_last_output;
      if (_allElementsMasked_T_20)
        indexedInstructionOffsets_19_bits <= offsetQueueVec_19_deq_bits;
      indexedInstructionOffsets_20_valid <= _allElementsMasked_T_21 | indexedInstructionOffsets_20_valid & ~usedIndexedInstructionOffsets_20 & ~_status_last_output;
      if (_allElementsMasked_T_21)
        indexedInstructionOffsets_20_bits <= offsetQueueVec_20_deq_bits;
      indexedInstructionOffsets_21_valid <= _allElementsMasked_T_22 | indexedInstructionOffsets_21_valid & ~usedIndexedInstructionOffsets_21 & ~_status_last_output;
      if (_allElementsMasked_T_22)
        indexedInstructionOffsets_21_bits <= offsetQueueVec_21_deq_bits;
      indexedInstructionOffsets_22_valid <= _allElementsMasked_T_23 | indexedInstructionOffsets_22_valid & ~usedIndexedInstructionOffsets_22 & ~_status_last_output;
      if (_allElementsMasked_T_23)
        indexedInstructionOffsets_22_bits <= offsetQueueVec_22_deq_bits;
      indexedInstructionOffsets_23_valid <= _allElementsMasked_T_24 | indexedInstructionOffsets_23_valid & ~usedIndexedInstructionOffsets_23 & ~_status_last_output;
      if (_allElementsMasked_T_24)
        indexedInstructionOffsets_23_bits <= offsetQueueVec_23_deq_bits;
      indexedInstructionOffsets_24_valid <= _allElementsMasked_T_25 | indexedInstructionOffsets_24_valid & ~usedIndexedInstructionOffsets_24 & ~_status_last_output;
      if (_allElementsMasked_T_25)
        indexedInstructionOffsets_24_bits <= offsetQueueVec_24_deq_bits;
      indexedInstructionOffsets_25_valid <= _allElementsMasked_T_26 | indexedInstructionOffsets_25_valid & ~usedIndexedInstructionOffsets_25 & ~_status_last_output;
      if (_allElementsMasked_T_26)
        indexedInstructionOffsets_25_bits <= offsetQueueVec_25_deq_bits;
      indexedInstructionOffsets_26_valid <= _allElementsMasked_T_27 | indexedInstructionOffsets_26_valid & ~usedIndexedInstructionOffsets_26 & ~_status_last_output;
      if (_allElementsMasked_T_27)
        indexedInstructionOffsets_26_bits <= offsetQueueVec_26_deq_bits;
      indexedInstructionOffsets_27_valid <= _allElementsMasked_T_28 | indexedInstructionOffsets_27_valid & ~usedIndexedInstructionOffsets_27 & ~_status_last_output;
      if (_allElementsMasked_T_28)
        indexedInstructionOffsets_27_bits <= offsetQueueVec_27_deq_bits;
      indexedInstructionOffsets_28_valid <= _allElementsMasked_T_29 | indexedInstructionOffsets_28_valid & ~usedIndexedInstructionOffsets_28 & ~_status_last_output;
      if (_allElementsMasked_T_29)
        indexedInstructionOffsets_28_bits <= offsetQueueVec_28_deq_bits;
      indexedInstructionOffsets_29_valid <= _allElementsMasked_T_30 | indexedInstructionOffsets_29_valid & ~usedIndexedInstructionOffsets_29 & ~_status_last_output;
      if (_allElementsMasked_T_30)
        indexedInstructionOffsets_29_bits <= offsetQueueVec_29_deq_bits;
      indexedInstructionOffsets_30_valid <= _allElementsMasked_T_31 | indexedInstructionOffsets_30_valid & ~usedIndexedInstructionOffsets_30 & ~_status_last_output;
      if (_allElementsMasked_T_31)
        indexedInstructionOffsets_30_bits <= offsetQueueVec_30_deq_bits;
      indexedInstructionOffsets_31_valid <= _allElementsMasked_T_32 | indexedInstructionOffsets_31_valid & ~usedIndexedInstructionOffsets_31 & ~_status_last_output;
      if (_allElementsMasked_T_32)
        indexedInstructionOffsets_31_bits <= offsetQueueVec_31_deq_bits;
      if (updateOffsetGroupEnable)
        groupIndex <= nextGroupIndex;
      if (maskGroupEndAndRequestNewMask | lsuRequest_valid)
        maskReg <= maskInput;
      if (isSegmentLoadStore & s0Fire | lsuRequest_valid)
        segmentIndex <= segmentEnd | lsuRequest_valid ? 3'h0 : segmentIndexNext;
      if (_GEN_26)
        state <= 2'h1;
      else if (_GEN_19)
        state <= {1'h0, ~last};
      else if (stateIsRequest & (last | maskGroupEnd))
        state <= 2'h2;
      if (segmentEndWithHandshake | updateOffsetGroupEnable) begin
        automatic logic [126:0] _GEN_20 = nextElementForMemoryRequest[126:0] | nextElementForMemoryRequest[127:1];
        automatic logic [125:0] _GEN_21 = _GEN_20[125:0] | {nextElementForMemoryRequest[127], _GEN_20[126:2]};
        automatic logic [123:0] _GEN_22 = _GEN_21[123:0] | {nextElementForMemoryRequest[127], _GEN_20[126], _GEN_21[125:4]};
        automatic logic [119:0] _GEN_23 = _GEN_22[119:0] | {nextElementForMemoryRequest[127], _GEN_20[126], _GEN_21[125:124], _GEN_22[123:8]};
        automatic logic [111:0] _GEN_24 = _GEN_23[111:0] | {nextElementForMemoryRequest[127], _GEN_20[126], _GEN_21[125:124], _GEN_22[123:120], _GEN_23[119:16]};
        automatic logic [95:0]  _GEN_25 = _GEN_24[95:0] | {nextElementForMemoryRequest[127], _GEN_20[126], _GEN_21[125:124], _GEN_22[123:120], _GEN_23[119:112], _GEN_24[111:32]};
        sentMemoryRequests <=
          updateOffsetGroupEnable
            ? 128'h0
            : {nextElementForMemoryRequest[127],
               _GEN_20[126],
               _GEN_21[125:124],
               _GEN_22[123:120],
               _GEN_23[119:112],
               _GEN_24[111:96],
               _GEN_25[95:64],
               _GEN_25[63:0] | {nextElementForMemoryRequest[127], _GEN_20[126], _GEN_21[125:124], _GEN_22[123:120], _GEN_23[119:112], _GEN_24[111:96], _GEN_25[95:64]}};
      end
      if (lsuRequest_valid | _outstandingTLDMessages_T_4)
        firstMemoryRequestOfInstruction <= lsuRequest_valid;
      if (lsuRequest_valid | _outstandingTLDMessages_T)
        waitFirstMemoryResponseForFaultOnlyFirst <= lsuRequest_valid & _waitFirstMemoryResponseForFaultOnlyFirst_T & lsuRequest_bits_instructionInformation_lumop[4] & ~lsuRequest_bits_instructionInformation_isStore;
      if (s0Fire ^ s0DequeueFire)
        s0Valid <= s0Fire;
      if (s0Fire) begin
        s0Reg_readVS <= s0Wire_readVS;
        s0Reg_offsetForVSInLane <= s0Wire_offsetForVSInLane;
        s0Reg_addressOffset <= s0Wire_addressOffset;
        s0Reg_segmentIndex <= s0Wire_segmentIndex;
        s0Reg_offsetForLane <= s0Wire_offsetForLane;
        s0Reg_indexInGroup <= s0Wire_indexInGroup;
      end
      if (s1Fire ^ memRequestFire)
        s1Valid <= s1Fire;
      if (s1Fire) begin
        s1Reg_indexInMaskGroup <= s1Wire_indexInMaskGroup;
        s1Reg_segmentIndex <= s1Wire_segmentIndex;
        s1Reg_address <= s1Wire_address;
        s1Reg_readData <= s1Wire_readData;
      end
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[0])
        offsetRecord_0 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[1])
        offsetRecord_1 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[2])
        offsetRecord_2 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[3])
        offsetRecord_3 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[4])
        offsetRecord_4 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[5])
        offsetRecord_5 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[6])
        offsetRecord_6 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[7])
        offsetRecord_7 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[8])
        offsetRecord_8 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[9])
        offsetRecord_9 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[10])
        offsetRecord_10 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[11])
        offsetRecord_11 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[12])
        offsetRecord_12 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[13])
        offsetRecord_13 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[14])
        offsetRecord_14 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[15])
        offsetRecord_15 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[16])
        offsetRecord_16 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[17])
        offsetRecord_17 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[18])
        offsetRecord_18 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[19])
        offsetRecord_19 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[20])
        offsetRecord_20 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[21])
        offsetRecord_21 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[22])
        offsetRecord_22 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[23])
        offsetRecord_23 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[24])
        offsetRecord_24 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[25])
        offsetRecord_25 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[26])
        offsetRecord_26 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[27])
        offsetRecord_27 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[28])
        offsetRecord_28 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[29])
        offsetRecord_29 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[30])
        offsetRecord_30 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[31])
        offsetRecord_31 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[32])
        offsetRecord_32 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[33])
        offsetRecord_33 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[34])
        offsetRecord_34 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[35])
        offsetRecord_35 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[36])
        offsetRecord_36 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[37])
        offsetRecord_37 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[38])
        offsetRecord_38 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[39])
        offsetRecord_39 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[40])
        offsetRecord_40 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[41])
        offsetRecord_41 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[42])
        offsetRecord_42 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[43])
        offsetRecord_43 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[44])
        offsetRecord_44 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[45])
        offsetRecord_45 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[46])
        offsetRecord_46 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[47])
        offsetRecord_47 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[48])
        offsetRecord_48 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[49])
        offsetRecord_49 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[50])
        offsetRecord_50 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[51])
        offsetRecord_51 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[52])
        offsetRecord_52 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[53])
        offsetRecord_53 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[54])
        offsetRecord_54 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[55])
        offsetRecord_55 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[56])
        offsetRecord_56 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[57])
        offsetRecord_57 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[58])
        offsetRecord_58 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[59])
        offsetRecord_59 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[60])
        offsetRecord_60 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[61])
        offsetRecord_61 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[62])
        offsetRecord_62 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[63])
        offsetRecord_63 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[64])
        offsetRecord_64 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[65])
        offsetRecord_65 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[66])
        offsetRecord_66 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[67])
        offsetRecord_67 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[68])
        offsetRecord_68 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[69])
        offsetRecord_69 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[70])
        offsetRecord_70 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[71])
        offsetRecord_71 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[72])
        offsetRecord_72 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[73])
        offsetRecord_73 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[74])
        offsetRecord_74 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[75])
        offsetRecord_75 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[76])
        offsetRecord_76 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[77])
        offsetRecord_77 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[78])
        offsetRecord_78 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[79])
        offsetRecord_79 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[80])
        offsetRecord_80 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[81])
        offsetRecord_81 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[82])
        offsetRecord_82 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[83])
        offsetRecord_83 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[84])
        offsetRecord_84 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[85])
        offsetRecord_85 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[86])
        offsetRecord_86 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[87])
        offsetRecord_87 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[88])
        offsetRecord_88 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[89])
        offsetRecord_89 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[90])
        offsetRecord_90 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[91])
        offsetRecord_91 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[92])
        offsetRecord_92 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[93])
        offsetRecord_93 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[94])
        offsetRecord_94 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[95])
        offsetRecord_95 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[96])
        offsetRecord_96 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[97])
        offsetRecord_97 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[98])
        offsetRecord_98 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[99])
        offsetRecord_99 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[100])
        offsetRecord_100 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[101])
        offsetRecord_101 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[102])
        offsetRecord_102 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[103])
        offsetRecord_103 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[104])
        offsetRecord_104 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[105])
        offsetRecord_105 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[106])
        offsetRecord_106 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[107])
        offsetRecord_107 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[108])
        offsetRecord_108 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[109])
        offsetRecord_109 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[110])
        offsetRecord_110 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[111])
        offsetRecord_111 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[112])
        offsetRecord_112 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[113])
        offsetRecord_113 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[114])
        offsetRecord_114 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[115])
        offsetRecord_115 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[116])
        offsetRecord_116 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[117])
        offsetRecord_117 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[118])
        offsetRecord_118 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[119])
        offsetRecord_119 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[120])
        offsetRecord_120 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[121])
        offsetRecord_121 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[122])
        offsetRecord_122 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[123])
        offsetRecord_123 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[124])
        offsetRecord_124 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[125])
        offsetRecord_125 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[126])
        offsetRecord_126 <= addressInBeatByte;
      if (_outstandingTLDMessages_T_4 & memoryRequestSourceOH[127])
        offsetRecord_127 <= addressInBeatByte;
    end
    if (lsuRequest_valid | _allElementsMasked_T_1)
      indexOfIndexedInstructionOffsets <= indexOfIndexedInstructionOffsetsNext;
    invalidInstructionNext <= invalidInstruction;
    status_last_REG <= stateIdle;
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:62];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [5:0] i = 6'h0; i < 6'h3F; i += 6'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        offsetQueueVec_deqLock = _RANDOM[6'h0][0];
        offsetQueueVec_deqLock_1 = _RANDOM[6'h0][1];
        offsetQueueVec_deqLock_2 = _RANDOM[6'h0][2];
        offsetQueueVec_deqLock_3 = _RANDOM[6'h0][3];
        offsetQueueVec_deqLock_4 = _RANDOM[6'h0][4];
        offsetQueueVec_deqLock_5 = _RANDOM[6'h0][5];
        offsetQueueVec_deqLock_6 = _RANDOM[6'h0][6];
        offsetQueueVec_deqLock_7 = _RANDOM[6'h0][7];
        offsetQueueVec_deqLock_8 = _RANDOM[6'h0][8];
        offsetQueueVec_deqLock_9 = _RANDOM[6'h0][9];
        offsetQueueVec_deqLock_10 = _RANDOM[6'h0][10];
        offsetQueueVec_deqLock_11 = _RANDOM[6'h0][11];
        offsetQueueVec_deqLock_12 = _RANDOM[6'h0][12];
        offsetQueueVec_deqLock_13 = _RANDOM[6'h0][13];
        offsetQueueVec_deqLock_14 = _RANDOM[6'h0][14];
        offsetQueueVec_deqLock_15 = _RANDOM[6'h0][15];
        offsetQueueVec_deqLock_16 = _RANDOM[6'h0][16];
        offsetQueueVec_deqLock_17 = _RANDOM[6'h0][17];
        offsetQueueVec_deqLock_18 = _RANDOM[6'h0][18];
        offsetQueueVec_deqLock_19 = _RANDOM[6'h0][19];
        offsetQueueVec_deqLock_20 = _RANDOM[6'h0][20];
        offsetQueueVec_deqLock_21 = _RANDOM[6'h0][21];
        offsetQueueVec_deqLock_22 = _RANDOM[6'h0][22];
        offsetQueueVec_deqLock_23 = _RANDOM[6'h0][23];
        offsetQueueVec_deqLock_24 = _RANDOM[6'h0][24];
        offsetQueueVec_deqLock_25 = _RANDOM[6'h0][25];
        offsetQueueVec_deqLock_26 = _RANDOM[6'h0][26];
        offsetQueueVec_deqLock_27 = _RANDOM[6'h0][27];
        offsetQueueVec_deqLock_28 = _RANDOM[6'h0][28];
        offsetQueueVec_deqLock_29 = _RANDOM[6'h0][29];
        offsetQueueVec_deqLock_30 = _RANDOM[6'h0][30];
        offsetQueueVec_deqLock_31 = _RANDOM[6'h0][31];
        lsuRequestReg_instructionInformation_nf = _RANDOM[6'h1][2:0];
        lsuRequestReg_instructionInformation_mew = _RANDOM[6'h1][3];
        lsuRequestReg_instructionInformation_mop = _RANDOM[6'h1][5:4];
        lsuRequestReg_instructionInformation_lumop = _RANDOM[6'h1][10:6];
        lsuRequestReg_instructionInformation_eew = _RANDOM[6'h1][12:11];
        lsuRequestReg_instructionInformation_vs3 = _RANDOM[6'h1][17:13];
        lsuRequestReg_instructionInformation_isStore = _RANDOM[6'h1][18];
        lsuRequestReg_instructionInformation_maskedLoadStore = _RANDOM[6'h1][19];
        lsuRequestReg_rs1Data = {_RANDOM[6'h1][31:20], _RANDOM[6'h2][19:0]};
        lsuRequestReg_rs2Data = {_RANDOM[6'h2][31:20], _RANDOM[6'h3][19:0]};
        lsuRequestReg_instructionIndex = _RANDOM[6'h3][22:20];
        csrInterfaceReg_vl = {_RANDOM[6'h3][31:23], _RANDOM[6'h4][2:0]};
        csrInterfaceReg_vStart = _RANDOM[6'h4][14:3];
        csrInterfaceReg_vlmul = _RANDOM[6'h4][17:15];
        csrInterfaceReg_vSew = _RANDOM[6'h4][19:18];
        csrInterfaceReg_vxrm = _RANDOM[6'h4][21:20];
        csrInterfaceReg_vta = _RANDOM[6'h4][22];
        csrInterfaceReg_vma = _RANDOM[6'h4][23];
        dataWidthForSegmentLoadStore = _RANDOM[6'h4][30:24];
        elementByteWidth = {_RANDOM[6'h4][31], _RANDOM[6'h5][1:0]};
        segmentInstructionIndexInterval = _RANDOM[6'h5][5:2];
        outstandingTLDMessages = {_RANDOM[6'h5][31:6], _RANDOM[6'h6], _RANDOM[6'h7], _RANDOM[6'h8], _RANDOM[6'h9][5:0]};
        indexedInstructionOffsets_0_valid = _RANDOM[6'h9][6];
        indexedInstructionOffsets_0_bits = {_RANDOM[6'h9][31:7], _RANDOM[6'hA][6:0]};
        indexedInstructionOffsets_1_valid = _RANDOM[6'hA][7];
        indexedInstructionOffsets_1_bits = {_RANDOM[6'hA][31:8], _RANDOM[6'hB][7:0]};
        indexedInstructionOffsets_2_valid = _RANDOM[6'hB][8];
        indexedInstructionOffsets_2_bits = {_RANDOM[6'hB][31:9], _RANDOM[6'hC][8:0]};
        indexedInstructionOffsets_3_valid = _RANDOM[6'hC][9];
        indexedInstructionOffsets_3_bits = {_RANDOM[6'hC][31:10], _RANDOM[6'hD][9:0]};
        indexedInstructionOffsets_4_valid = _RANDOM[6'hD][10];
        indexedInstructionOffsets_4_bits = {_RANDOM[6'hD][31:11], _RANDOM[6'hE][10:0]};
        indexedInstructionOffsets_5_valid = _RANDOM[6'hE][11];
        indexedInstructionOffsets_5_bits = {_RANDOM[6'hE][31:12], _RANDOM[6'hF][11:0]};
        indexedInstructionOffsets_6_valid = _RANDOM[6'hF][12];
        indexedInstructionOffsets_6_bits = {_RANDOM[6'hF][31:13], _RANDOM[6'h10][12:0]};
        indexedInstructionOffsets_7_valid = _RANDOM[6'h10][13];
        indexedInstructionOffsets_7_bits = {_RANDOM[6'h10][31:14], _RANDOM[6'h11][13:0]};
        indexedInstructionOffsets_8_valid = _RANDOM[6'h11][14];
        indexedInstructionOffsets_8_bits = {_RANDOM[6'h11][31:15], _RANDOM[6'h12][14:0]};
        indexedInstructionOffsets_9_valid = _RANDOM[6'h12][15];
        indexedInstructionOffsets_9_bits = {_RANDOM[6'h12][31:16], _RANDOM[6'h13][15:0]};
        indexedInstructionOffsets_10_valid = _RANDOM[6'h13][16];
        indexedInstructionOffsets_10_bits = {_RANDOM[6'h13][31:17], _RANDOM[6'h14][16:0]};
        indexedInstructionOffsets_11_valid = _RANDOM[6'h14][17];
        indexedInstructionOffsets_11_bits = {_RANDOM[6'h14][31:18], _RANDOM[6'h15][17:0]};
        indexedInstructionOffsets_12_valid = _RANDOM[6'h15][18];
        indexedInstructionOffsets_12_bits = {_RANDOM[6'h15][31:19], _RANDOM[6'h16][18:0]};
        indexedInstructionOffsets_13_valid = _RANDOM[6'h16][19];
        indexedInstructionOffsets_13_bits = {_RANDOM[6'h16][31:20], _RANDOM[6'h17][19:0]};
        indexedInstructionOffsets_14_valid = _RANDOM[6'h17][20];
        indexedInstructionOffsets_14_bits = {_RANDOM[6'h17][31:21], _RANDOM[6'h18][20:0]};
        indexedInstructionOffsets_15_valid = _RANDOM[6'h18][21];
        indexedInstructionOffsets_15_bits = {_RANDOM[6'h18][31:22], _RANDOM[6'h19][21:0]};
        indexedInstructionOffsets_16_valid = _RANDOM[6'h19][22];
        indexedInstructionOffsets_16_bits = {_RANDOM[6'h19][31:23], _RANDOM[6'h1A][22:0]};
        indexedInstructionOffsets_17_valid = _RANDOM[6'h1A][23];
        indexedInstructionOffsets_17_bits = {_RANDOM[6'h1A][31:24], _RANDOM[6'h1B][23:0]};
        indexedInstructionOffsets_18_valid = _RANDOM[6'h1B][24];
        indexedInstructionOffsets_18_bits = {_RANDOM[6'h1B][31:25], _RANDOM[6'h1C][24:0]};
        indexedInstructionOffsets_19_valid = _RANDOM[6'h1C][25];
        indexedInstructionOffsets_19_bits = {_RANDOM[6'h1C][31:26], _RANDOM[6'h1D][25:0]};
        indexedInstructionOffsets_20_valid = _RANDOM[6'h1D][26];
        indexedInstructionOffsets_20_bits = {_RANDOM[6'h1D][31:27], _RANDOM[6'h1E][26:0]};
        indexedInstructionOffsets_21_valid = _RANDOM[6'h1E][27];
        indexedInstructionOffsets_21_bits = {_RANDOM[6'h1E][31:28], _RANDOM[6'h1F][27:0]};
        indexedInstructionOffsets_22_valid = _RANDOM[6'h1F][28];
        indexedInstructionOffsets_22_bits = {_RANDOM[6'h1F][31:29], _RANDOM[6'h20][28:0]};
        indexedInstructionOffsets_23_valid = _RANDOM[6'h20][29];
        indexedInstructionOffsets_23_bits = {_RANDOM[6'h20][31:30], _RANDOM[6'h21][29:0]};
        indexedInstructionOffsets_24_valid = _RANDOM[6'h21][30];
        indexedInstructionOffsets_24_bits = {_RANDOM[6'h21][31], _RANDOM[6'h22][30:0]};
        indexedInstructionOffsets_25_valid = _RANDOM[6'h22][31];
        indexedInstructionOffsets_25_bits = _RANDOM[6'h23];
        indexedInstructionOffsets_26_valid = _RANDOM[6'h24][0];
        indexedInstructionOffsets_26_bits = {_RANDOM[6'h24][31:1], _RANDOM[6'h25][0]};
        indexedInstructionOffsets_27_valid = _RANDOM[6'h25][1];
        indexedInstructionOffsets_27_bits = {_RANDOM[6'h25][31:2], _RANDOM[6'h26][1:0]};
        indexedInstructionOffsets_28_valid = _RANDOM[6'h26][2];
        indexedInstructionOffsets_28_bits = {_RANDOM[6'h26][31:3], _RANDOM[6'h27][2:0]};
        indexedInstructionOffsets_29_valid = _RANDOM[6'h27][3];
        indexedInstructionOffsets_29_bits = {_RANDOM[6'h27][31:4], _RANDOM[6'h28][3:0]};
        indexedInstructionOffsets_30_valid = _RANDOM[6'h28][4];
        indexedInstructionOffsets_30_bits = {_RANDOM[6'h28][31:5], _RANDOM[6'h29][4:0]};
        indexedInstructionOffsets_31_valid = _RANDOM[6'h29][5];
        indexedInstructionOffsets_31_bits = {_RANDOM[6'h29][31:6], _RANDOM[6'h2A][5:0]};
        groupIndex = _RANDOM[6'h2A][10:6];
        indexOfIndexedInstructionOffsets = _RANDOM[6'h2A][12:11];
        maskReg = {_RANDOM[6'h2A][31:13], _RANDOM[6'h2B], _RANDOM[6'h2C], _RANDOM[6'h2D], _RANDOM[6'h2E][12:0]};
        segmentIndex = _RANDOM[6'h2E][15:13];
        state = _RANDOM[6'h2E][17:16];
        sentMemoryRequests = {_RANDOM[6'h2E][31:18], _RANDOM[6'h2F], _RANDOM[6'h30], _RANDOM[6'h31], _RANDOM[6'h32][17:0]};
        firstMemoryRequestOfInstruction = _RANDOM[6'h32][18];
        waitFirstMemoryResponseForFaultOnlyFirst = _RANDOM[6'h32][19];
        s0Valid = _RANDOM[6'h32][20];
        s0Reg_readVS = _RANDOM[6'h32][25:21];
        s0Reg_offsetForVSInLane = _RANDOM[6'h32][26];
        s0Reg_addressOffset = {_RANDOM[6'h32][31:27], _RANDOM[6'h33][26:0]};
        s0Reg_segmentIndex = _RANDOM[6'h33][29:27];
        s0Reg_offsetForLane = {_RANDOM[6'h33][31:30], _RANDOM[6'h34][2:0]};
        s0Reg_indexInGroup = _RANDOM[6'h34][9:3];
        s1Valid = _RANDOM[6'h34][10];
        s1Reg_indexInMaskGroup = _RANDOM[6'h34][17:11];
        s1Reg_segmentIndex = _RANDOM[6'h34][20:18];
        s1Reg_address = {_RANDOM[6'h34][31:21], _RANDOM[6'h35][20:0]};
        s1Reg_readData = {_RANDOM[6'h35][31:21], _RANDOM[6'h36][20:0]};
        offsetRecord_0 = _RANDOM[6'h36][22:21];
        offsetRecord_1 = _RANDOM[6'h36][24:23];
        offsetRecord_2 = _RANDOM[6'h36][26:25];
        offsetRecord_3 = _RANDOM[6'h36][28:27];
        offsetRecord_4 = _RANDOM[6'h36][30:29];
        offsetRecord_5 = {_RANDOM[6'h36][31], _RANDOM[6'h37][0]};
        offsetRecord_6 = _RANDOM[6'h37][2:1];
        offsetRecord_7 = _RANDOM[6'h37][4:3];
        offsetRecord_8 = _RANDOM[6'h37][6:5];
        offsetRecord_9 = _RANDOM[6'h37][8:7];
        offsetRecord_10 = _RANDOM[6'h37][10:9];
        offsetRecord_11 = _RANDOM[6'h37][12:11];
        offsetRecord_12 = _RANDOM[6'h37][14:13];
        offsetRecord_13 = _RANDOM[6'h37][16:15];
        offsetRecord_14 = _RANDOM[6'h37][18:17];
        offsetRecord_15 = _RANDOM[6'h37][20:19];
        offsetRecord_16 = _RANDOM[6'h37][22:21];
        offsetRecord_17 = _RANDOM[6'h37][24:23];
        offsetRecord_18 = _RANDOM[6'h37][26:25];
        offsetRecord_19 = _RANDOM[6'h37][28:27];
        offsetRecord_20 = _RANDOM[6'h37][30:29];
        offsetRecord_21 = {_RANDOM[6'h37][31], _RANDOM[6'h38][0]};
        offsetRecord_22 = _RANDOM[6'h38][2:1];
        offsetRecord_23 = _RANDOM[6'h38][4:3];
        offsetRecord_24 = _RANDOM[6'h38][6:5];
        offsetRecord_25 = _RANDOM[6'h38][8:7];
        offsetRecord_26 = _RANDOM[6'h38][10:9];
        offsetRecord_27 = _RANDOM[6'h38][12:11];
        offsetRecord_28 = _RANDOM[6'h38][14:13];
        offsetRecord_29 = _RANDOM[6'h38][16:15];
        offsetRecord_30 = _RANDOM[6'h38][18:17];
        offsetRecord_31 = _RANDOM[6'h38][20:19];
        offsetRecord_32 = _RANDOM[6'h38][22:21];
        offsetRecord_33 = _RANDOM[6'h38][24:23];
        offsetRecord_34 = _RANDOM[6'h38][26:25];
        offsetRecord_35 = _RANDOM[6'h38][28:27];
        offsetRecord_36 = _RANDOM[6'h38][30:29];
        offsetRecord_37 = {_RANDOM[6'h38][31], _RANDOM[6'h39][0]};
        offsetRecord_38 = _RANDOM[6'h39][2:1];
        offsetRecord_39 = _RANDOM[6'h39][4:3];
        offsetRecord_40 = _RANDOM[6'h39][6:5];
        offsetRecord_41 = _RANDOM[6'h39][8:7];
        offsetRecord_42 = _RANDOM[6'h39][10:9];
        offsetRecord_43 = _RANDOM[6'h39][12:11];
        offsetRecord_44 = _RANDOM[6'h39][14:13];
        offsetRecord_45 = _RANDOM[6'h39][16:15];
        offsetRecord_46 = _RANDOM[6'h39][18:17];
        offsetRecord_47 = _RANDOM[6'h39][20:19];
        offsetRecord_48 = _RANDOM[6'h39][22:21];
        offsetRecord_49 = _RANDOM[6'h39][24:23];
        offsetRecord_50 = _RANDOM[6'h39][26:25];
        offsetRecord_51 = _RANDOM[6'h39][28:27];
        offsetRecord_52 = _RANDOM[6'h39][30:29];
        offsetRecord_53 = {_RANDOM[6'h39][31], _RANDOM[6'h3A][0]};
        offsetRecord_54 = _RANDOM[6'h3A][2:1];
        offsetRecord_55 = _RANDOM[6'h3A][4:3];
        offsetRecord_56 = _RANDOM[6'h3A][6:5];
        offsetRecord_57 = _RANDOM[6'h3A][8:7];
        offsetRecord_58 = _RANDOM[6'h3A][10:9];
        offsetRecord_59 = _RANDOM[6'h3A][12:11];
        offsetRecord_60 = _RANDOM[6'h3A][14:13];
        offsetRecord_61 = _RANDOM[6'h3A][16:15];
        offsetRecord_62 = _RANDOM[6'h3A][18:17];
        offsetRecord_63 = _RANDOM[6'h3A][20:19];
        offsetRecord_64 = _RANDOM[6'h3A][22:21];
        offsetRecord_65 = _RANDOM[6'h3A][24:23];
        offsetRecord_66 = _RANDOM[6'h3A][26:25];
        offsetRecord_67 = _RANDOM[6'h3A][28:27];
        offsetRecord_68 = _RANDOM[6'h3A][30:29];
        offsetRecord_69 = {_RANDOM[6'h3A][31], _RANDOM[6'h3B][0]};
        offsetRecord_70 = _RANDOM[6'h3B][2:1];
        offsetRecord_71 = _RANDOM[6'h3B][4:3];
        offsetRecord_72 = _RANDOM[6'h3B][6:5];
        offsetRecord_73 = _RANDOM[6'h3B][8:7];
        offsetRecord_74 = _RANDOM[6'h3B][10:9];
        offsetRecord_75 = _RANDOM[6'h3B][12:11];
        offsetRecord_76 = _RANDOM[6'h3B][14:13];
        offsetRecord_77 = _RANDOM[6'h3B][16:15];
        offsetRecord_78 = _RANDOM[6'h3B][18:17];
        offsetRecord_79 = _RANDOM[6'h3B][20:19];
        offsetRecord_80 = _RANDOM[6'h3B][22:21];
        offsetRecord_81 = _RANDOM[6'h3B][24:23];
        offsetRecord_82 = _RANDOM[6'h3B][26:25];
        offsetRecord_83 = _RANDOM[6'h3B][28:27];
        offsetRecord_84 = _RANDOM[6'h3B][30:29];
        offsetRecord_85 = {_RANDOM[6'h3B][31], _RANDOM[6'h3C][0]};
        offsetRecord_86 = _RANDOM[6'h3C][2:1];
        offsetRecord_87 = _RANDOM[6'h3C][4:3];
        offsetRecord_88 = _RANDOM[6'h3C][6:5];
        offsetRecord_89 = _RANDOM[6'h3C][8:7];
        offsetRecord_90 = _RANDOM[6'h3C][10:9];
        offsetRecord_91 = _RANDOM[6'h3C][12:11];
        offsetRecord_92 = _RANDOM[6'h3C][14:13];
        offsetRecord_93 = _RANDOM[6'h3C][16:15];
        offsetRecord_94 = _RANDOM[6'h3C][18:17];
        offsetRecord_95 = _RANDOM[6'h3C][20:19];
        offsetRecord_96 = _RANDOM[6'h3C][22:21];
        offsetRecord_97 = _RANDOM[6'h3C][24:23];
        offsetRecord_98 = _RANDOM[6'h3C][26:25];
        offsetRecord_99 = _RANDOM[6'h3C][28:27];
        offsetRecord_100 = _RANDOM[6'h3C][30:29];
        offsetRecord_101 = {_RANDOM[6'h3C][31], _RANDOM[6'h3D][0]};
        offsetRecord_102 = _RANDOM[6'h3D][2:1];
        offsetRecord_103 = _RANDOM[6'h3D][4:3];
        offsetRecord_104 = _RANDOM[6'h3D][6:5];
        offsetRecord_105 = _RANDOM[6'h3D][8:7];
        offsetRecord_106 = _RANDOM[6'h3D][10:9];
        offsetRecord_107 = _RANDOM[6'h3D][12:11];
        offsetRecord_108 = _RANDOM[6'h3D][14:13];
        offsetRecord_109 = _RANDOM[6'h3D][16:15];
        offsetRecord_110 = _RANDOM[6'h3D][18:17];
        offsetRecord_111 = _RANDOM[6'h3D][20:19];
        offsetRecord_112 = _RANDOM[6'h3D][22:21];
        offsetRecord_113 = _RANDOM[6'h3D][24:23];
        offsetRecord_114 = _RANDOM[6'h3D][26:25];
        offsetRecord_115 = _RANDOM[6'h3D][28:27];
        offsetRecord_116 = _RANDOM[6'h3D][30:29];
        offsetRecord_117 = {_RANDOM[6'h3D][31], _RANDOM[6'h3E][0]};
        offsetRecord_118 = _RANDOM[6'h3E][2:1];
        offsetRecord_119 = _RANDOM[6'h3E][4:3];
        offsetRecord_120 = _RANDOM[6'h3E][6:5];
        offsetRecord_121 = _RANDOM[6'h3E][8:7];
        offsetRecord_122 = _RANDOM[6'h3E][10:9];
        offsetRecord_123 = _RANDOM[6'h3E][12:11];
        offsetRecord_124 = _RANDOM[6'h3E][14:13];
        offsetRecord_125 = _RANDOM[6'h3E][16:15];
        offsetRecord_126 = _RANDOM[6'h3E][18:17];
        offsetRecord_127 = _RANDOM[6'h3E][20:19];
        invalidInstructionNext = _RANDOM[6'h3E][21];
        status_last_REG = _RANDOM[6'h3E][22];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  wire              offsetQueueVec_0_empty;
  assign offsetQueueVec_0_empty = _offsetQueueVec_queue_fifo_empty;
  wire              offsetQueueVec_0_full;
  assign offsetQueueVec_0_full = _offsetQueueVec_queue_fifo_full;
  wire              offsetQueueVec_1_empty;
  assign offsetQueueVec_1_empty = _offsetQueueVec_queue_fifo_1_empty;
  wire              offsetQueueVec_1_full;
  assign offsetQueueVec_1_full = _offsetQueueVec_queue_fifo_1_full;
  wire              offsetQueueVec_2_empty;
  assign offsetQueueVec_2_empty = _offsetQueueVec_queue_fifo_2_empty;
  wire              offsetQueueVec_2_full;
  assign offsetQueueVec_2_full = _offsetQueueVec_queue_fifo_2_full;
  wire              offsetQueueVec_3_empty;
  assign offsetQueueVec_3_empty = _offsetQueueVec_queue_fifo_3_empty;
  wire              offsetQueueVec_3_full;
  assign offsetQueueVec_3_full = _offsetQueueVec_queue_fifo_3_full;
  wire              offsetQueueVec_4_empty;
  assign offsetQueueVec_4_empty = _offsetQueueVec_queue_fifo_4_empty;
  wire              offsetQueueVec_4_full;
  assign offsetQueueVec_4_full = _offsetQueueVec_queue_fifo_4_full;
  wire              offsetQueueVec_5_empty;
  assign offsetQueueVec_5_empty = _offsetQueueVec_queue_fifo_5_empty;
  wire              offsetQueueVec_5_full;
  assign offsetQueueVec_5_full = _offsetQueueVec_queue_fifo_5_full;
  wire              offsetQueueVec_6_empty;
  assign offsetQueueVec_6_empty = _offsetQueueVec_queue_fifo_6_empty;
  wire              offsetQueueVec_6_full;
  assign offsetQueueVec_6_full = _offsetQueueVec_queue_fifo_6_full;
  wire              offsetQueueVec_7_empty;
  assign offsetQueueVec_7_empty = _offsetQueueVec_queue_fifo_7_empty;
  wire              offsetQueueVec_7_full;
  assign offsetQueueVec_7_full = _offsetQueueVec_queue_fifo_7_full;
  wire              offsetQueueVec_8_empty;
  assign offsetQueueVec_8_empty = _offsetQueueVec_queue_fifo_8_empty;
  wire              offsetQueueVec_8_full;
  assign offsetQueueVec_8_full = _offsetQueueVec_queue_fifo_8_full;
  wire              offsetQueueVec_9_empty;
  assign offsetQueueVec_9_empty = _offsetQueueVec_queue_fifo_9_empty;
  wire              offsetQueueVec_9_full;
  assign offsetQueueVec_9_full = _offsetQueueVec_queue_fifo_9_full;
  wire              offsetQueueVec_10_empty;
  assign offsetQueueVec_10_empty = _offsetQueueVec_queue_fifo_10_empty;
  wire              offsetQueueVec_10_full;
  assign offsetQueueVec_10_full = _offsetQueueVec_queue_fifo_10_full;
  wire              offsetQueueVec_11_empty;
  assign offsetQueueVec_11_empty = _offsetQueueVec_queue_fifo_11_empty;
  wire              offsetQueueVec_11_full;
  assign offsetQueueVec_11_full = _offsetQueueVec_queue_fifo_11_full;
  wire              offsetQueueVec_12_empty;
  assign offsetQueueVec_12_empty = _offsetQueueVec_queue_fifo_12_empty;
  wire              offsetQueueVec_12_full;
  assign offsetQueueVec_12_full = _offsetQueueVec_queue_fifo_12_full;
  wire              offsetQueueVec_13_empty;
  assign offsetQueueVec_13_empty = _offsetQueueVec_queue_fifo_13_empty;
  wire              offsetQueueVec_13_full;
  assign offsetQueueVec_13_full = _offsetQueueVec_queue_fifo_13_full;
  wire              offsetQueueVec_14_empty;
  assign offsetQueueVec_14_empty = _offsetQueueVec_queue_fifo_14_empty;
  wire              offsetQueueVec_14_full;
  assign offsetQueueVec_14_full = _offsetQueueVec_queue_fifo_14_full;
  wire              offsetQueueVec_15_empty;
  assign offsetQueueVec_15_empty = _offsetQueueVec_queue_fifo_15_empty;
  wire              offsetQueueVec_15_full;
  assign offsetQueueVec_15_full = _offsetQueueVec_queue_fifo_15_full;
  wire              offsetQueueVec_16_empty;
  assign offsetQueueVec_16_empty = _offsetQueueVec_queue_fifo_16_empty;
  wire              offsetQueueVec_16_full;
  assign offsetQueueVec_16_full = _offsetQueueVec_queue_fifo_16_full;
  wire              offsetQueueVec_17_empty;
  assign offsetQueueVec_17_empty = _offsetQueueVec_queue_fifo_17_empty;
  wire              offsetQueueVec_17_full;
  assign offsetQueueVec_17_full = _offsetQueueVec_queue_fifo_17_full;
  wire              offsetQueueVec_18_empty;
  assign offsetQueueVec_18_empty = _offsetQueueVec_queue_fifo_18_empty;
  wire              offsetQueueVec_18_full;
  assign offsetQueueVec_18_full = _offsetQueueVec_queue_fifo_18_full;
  wire              offsetQueueVec_19_empty;
  assign offsetQueueVec_19_empty = _offsetQueueVec_queue_fifo_19_empty;
  wire              offsetQueueVec_19_full;
  assign offsetQueueVec_19_full = _offsetQueueVec_queue_fifo_19_full;
  wire              offsetQueueVec_20_empty;
  assign offsetQueueVec_20_empty = _offsetQueueVec_queue_fifo_20_empty;
  wire              offsetQueueVec_20_full;
  assign offsetQueueVec_20_full = _offsetQueueVec_queue_fifo_20_full;
  wire              offsetQueueVec_21_empty;
  assign offsetQueueVec_21_empty = _offsetQueueVec_queue_fifo_21_empty;
  wire              offsetQueueVec_21_full;
  assign offsetQueueVec_21_full = _offsetQueueVec_queue_fifo_21_full;
  wire              offsetQueueVec_22_empty;
  assign offsetQueueVec_22_empty = _offsetQueueVec_queue_fifo_22_empty;
  wire              offsetQueueVec_22_full;
  assign offsetQueueVec_22_full = _offsetQueueVec_queue_fifo_22_full;
  wire              offsetQueueVec_23_empty;
  assign offsetQueueVec_23_empty = _offsetQueueVec_queue_fifo_23_empty;
  wire              offsetQueueVec_23_full;
  assign offsetQueueVec_23_full = _offsetQueueVec_queue_fifo_23_full;
  wire              offsetQueueVec_24_empty;
  assign offsetQueueVec_24_empty = _offsetQueueVec_queue_fifo_24_empty;
  wire              offsetQueueVec_24_full;
  assign offsetQueueVec_24_full = _offsetQueueVec_queue_fifo_24_full;
  wire              offsetQueueVec_25_empty;
  assign offsetQueueVec_25_empty = _offsetQueueVec_queue_fifo_25_empty;
  wire              offsetQueueVec_25_full;
  assign offsetQueueVec_25_full = _offsetQueueVec_queue_fifo_25_full;
  wire              offsetQueueVec_26_empty;
  assign offsetQueueVec_26_empty = _offsetQueueVec_queue_fifo_26_empty;
  wire              offsetQueueVec_26_full;
  assign offsetQueueVec_26_full = _offsetQueueVec_queue_fifo_26_full;
  wire              offsetQueueVec_27_empty;
  assign offsetQueueVec_27_empty = _offsetQueueVec_queue_fifo_27_empty;
  wire              offsetQueueVec_27_full;
  assign offsetQueueVec_27_full = _offsetQueueVec_queue_fifo_27_full;
  wire              offsetQueueVec_28_empty;
  assign offsetQueueVec_28_empty = _offsetQueueVec_queue_fifo_28_empty;
  wire              offsetQueueVec_28_full;
  assign offsetQueueVec_28_full = _offsetQueueVec_queue_fifo_28_full;
  wire              offsetQueueVec_29_empty;
  assign offsetQueueVec_29_empty = _offsetQueueVec_queue_fifo_29_empty;
  wire              offsetQueueVec_29_full;
  assign offsetQueueVec_29_full = _offsetQueueVec_queue_fifo_29_full;
  wire              offsetQueueVec_30_empty;
  assign offsetQueueVec_30_empty = _offsetQueueVec_queue_fifo_30_empty;
  wire              offsetQueueVec_30_full;
  assign offsetQueueVec_30_full = _offsetQueueVec_queue_fifo_30_full;
  wire              offsetQueueVec_31_empty;
  assign offsetQueueVec_31_empty = _offsetQueueVec_queue_fifo_31_empty;
  wire              offsetQueueVec_31_full;
  assign offsetQueueVec_31_full = _offsetQueueVec_queue_fifo_31_full;
  wire              s1EnqQueue_empty;
  assign s1EnqQueue_empty = _s1EnqQueue_fifo_empty;
  wire              s1EnqQueue_full;
  assign s1EnqQueue_full = _s1EnqQueue_fifo_full;
  wire              s1EnqDataQueue_empty;
  assign s1EnqDataQueue_empty = _s1EnqDataQueue_fifo_empty;
  wire              s1EnqDataQueue_full;
  assign s1EnqDataQueue_full = _s1EnqDataQueue_fifo_full;
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_0_enq_ready & offsetQueueVec_0_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_0_deq_ready & ~_offsetQueueVec_queue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_0_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_empty),
    .almost_empty (offsetQueueVec_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_0_almostFull),
    .full         (_offsetQueueVec_queue_fifo_full),
    .error        (_offsetQueueVec_queue_fifo_error),
    .data_out     (offsetQueueVec_0_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_1_enq_ready & offsetQueueVec_1_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_1_deq_ready & ~_offsetQueueVec_queue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_1_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_1_empty),
    .almost_empty (offsetQueueVec_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_1_almostFull),
    .full         (_offsetQueueVec_queue_fifo_1_full),
    .error        (_offsetQueueVec_queue_fifo_1_error),
    .data_out     (offsetQueueVec_1_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_2_enq_ready & offsetQueueVec_2_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_2_deq_ready & ~_offsetQueueVec_queue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_2_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_2_empty),
    .almost_empty (offsetQueueVec_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_2_almostFull),
    .full         (_offsetQueueVec_queue_fifo_2_full),
    .error        (_offsetQueueVec_queue_fifo_2_error),
    .data_out     (offsetQueueVec_2_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_3_enq_ready & offsetQueueVec_3_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_3_deq_ready & ~_offsetQueueVec_queue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_3_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_3_empty),
    .almost_empty (offsetQueueVec_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_3_almostFull),
    .full         (_offsetQueueVec_queue_fifo_3_full),
    .error        (_offsetQueueVec_queue_fifo_3_error),
    .data_out     (offsetQueueVec_3_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_4_enq_ready & offsetQueueVec_4_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_4_deq_ready & ~_offsetQueueVec_queue_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_4_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_4_empty),
    .almost_empty (offsetQueueVec_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_4_almostFull),
    .full         (_offsetQueueVec_queue_fifo_4_full),
    .error        (_offsetQueueVec_queue_fifo_4_error),
    .data_out     (offsetQueueVec_4_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_5_enq_ready & offsetQueueVec_5_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_5_deq_ready & ~_offsetQueueVec_queue_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_5_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_5_empty),
    .almost_empty (offsetQueueVec_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_5_almostFull),
    .full         (_offsetQueueVec_queue_fifo_5_full),
    .error        (_offsetQueueVec_queue_fifo_5_error),
    .data_out     (offsetQueueVec_5_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_6_enq_ready & offsetQueueVec_6_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_6_deq_ready & ~_offsetQueueVec_queue_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_6_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_6_empty),
    .almost_empty (offsetQueueVec_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_6_almostFull),
    .full         (_offsetQueueVec_queue_fifo_6_full),
    .error        (_offsetQueueVec_queue_fifo_6_error),
    .data_out     (offsetQueueVec_6_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_7_enq_ready & offsetQueueVec_7_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_7_deq_ready & ~_offsetQueueVec_queue_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_7_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_7_empty),
    .almost_empty (offsetQueueVec_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_7_almostFull),
    .full         (_offsetQueueVec_queue_fifo_7_full),
    .error        (_offsetQueueVec_queue_fifo_7_error),
    .data_out     (offsetQueueVec_7_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_8_enq_ready & offsetQueueVec_8_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_8_deq_ready & ~_offsetQueueVec_queue_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_8_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_8_empty),
    .almost_empty (offsetQueueVec_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_8_almostFull),
    .full         (_offsetQueueVec_queue_fifo_8_full),
    .error        (_offsetQueueVec_queue_fifo_8_error),
    .data_out     (offsetQueueVec_8_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_9_enq_ready & offsetQueueVec_9_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_9_deq_ready & ~_offsetQueueVec_queue_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_9_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_9_empty),
    .almost_empty (offsetQueueVec_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_9_almostFull),
    .full         (_offsetQueueVec_queue_fifo_9_full),
    .error        (_offsetQueueVec_queue_fifo_9_error),
    .data_out     (offsetQueueVec_9_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_10_enq_ready & offsetQueueVec_10_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_10_deq_ready & ~_offsetQueueVec_queue_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_10_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_10_empty),
    .almost_empty (offsetQueueVec_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_10_almostFull),
    .full         (_offsetQueueVec_queue_fifo_10_full),
    .error        (_offsetQueueVec_queue_fifo_10_error),
    .data_out     (offsetQueueVec_10_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_11_enq_ready & offsetQueueVec_11_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_11_deq_ready & ~_offsetQueueVec_queue_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_11_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_11_empty),
    .almost_empty (offsetQueueVec_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_11_almostFull),
    .full         (_offsetQueueVec_queue_fifo_11_full),
    .error        (_offsetQueueVec_queue_fifo_11_error),
    .data_out     (offsetQueueVec_11_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_12_enq_ready & offsetQueueVec_12_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_12_deq_ready & ~_offsetQueueVec_queue_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_12_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_12_empty),
    .almost_empty (offsetQueueVec_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_12_almostFull),
    .full         (_offsetQueueVec_queue_fifo_12_full),
    .error        (_offsetQueueVec_queue_fifo_12_error),
    .data_out     (offsetQueueVec_12_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_13_enq_ready & offsetQueueVec_13_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_13_deq_ready & ~_offsetQueueVec_queue_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_13_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_13_empty),
    .almost_empty (offsetQueueVec_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_13_almostFull),
    .full         (_offsetQueueVec_queue_fifo_13_full),
    .error        (_offsetQueueVec_queue_fifo_13_error),
    .data_out     (offsetQueueVec_13_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_14_enq_ready & offsetQueueVec_14_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_14_deq_ready & ~_offsetQueueVec_queue_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_14_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_14_empty),
    .almost_empty (offsetQueueVec_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_14_almostFull),
    .full         (_offsetQueueVec_queue_fifo_14_full),
    .error        (_offsetQueueVec_queue_fifo_14_error),
    .data_out     (offsetQueueVec_14_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_15_enq_ready & offsetQueueVec_15_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_15_deq_ready & ~_offsetQueueVec_queue_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_15_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_15_empty),
    .almost_empty (offsetQueueVec_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_15_almostFull),
    .full         (_offsetQueueVec_queue_fifo_15_full),
    .error        (_offsetQueueVec_queue_fifo_15_error),
    .data_out     (offsetQueueVec_15_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_16 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_16_enq_ready & offsetQueueVec_16_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_16_deq_ready & ~_offsetQueueVec_queue_fifo_16_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_16_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_16_empty),
    .almost_empty (offsetQueueVec_16_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_16_almostFull),
    .full         (_offsetQueueVec_queue_fifo_16_full),
    .error        (_offsetQueueVec_queue_fifo_16_error),
    .data_out     (offsetQueueVec_16_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_17 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_17_enq_ready & offsetQueueVec_17_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_17_deq_ready & ~_offsetQueueVec_queue_fifo_17_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_17_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_17_empty),
    .almost_empty (offsetQueueVec_17_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_17_almostFull),
    .full         (_offsetQueueVec_queue_fifo_17_full),
    .error        (_offsetQueueVec_queue_fifo_17_error),
    .data_out     (offsetQueueVec_17_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_18 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_18_enq_ready & offsetQueueVec_18_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_18_deq_ready & ~_offsetQueueVec_queue_fifo_18_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_18_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_18_empty),
    .almost_empty (offsetQueueVec_18_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_18_almostFull),
    .full         (_offsetQueueVec_queue_fifo_18_full),
    .error        (_offsetQueueVec_queue_fifo_18_error),
    .data_out     (offsetQueueVec_18_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_19 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_19_enq_ready & offsetQueueVec_19_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_19_deq_ready & ~_offsetQueueVec_queue_fifo_19_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_19_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_19_empty),
    .almost_empty (offsetQueueVec_19_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_19_almostFull),
    .full         (_offsetQueueVec_queue_fifo_19_full),
    .error        (_offsetQueueVec_queue_fifo_19_error),
    .data_out     (offsetQueueVec_19_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_20 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_20_enq_ready & offsetQueueVec_20_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_20_deq_ready & ~_offsetQueueVec_queue_fifo_20_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_20_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_20_empty),
    .almost_empty (offsetQueueVec_20_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_20_almostFull),
    .full         (_offsetQueueVec_queue_fifo_20_full),
    .error        (_offsetQueueVec_queue_fifo_20_error),
    .data_out     (offsetQueueVec_20_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_21 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_21_enq_ready & offsetQueueVec_21_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_21_deq_ready & ~_offsetQueueVec_queue_fifo_21_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_21_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_21_empty),
    .almost_empty (offsetQueueVec_21_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_21_almostFull),
    .full         (_offsetQueueVec_queue_fifo_21_full),
    .error        (_offsetQueueVec_queue_fifo_21_error),
    .data_out     (offsetQueueVec_21_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_22 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_22_enq_ready & offsetQueueVec_22_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_22_deq_ready & ~_offsetQueueVec_queue_fifo_22_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_22_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_22_empty),
    .almost_empty (offsetQueueVec_22_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_22_almostFull),
    .full         (_offsetQueueVec_queue_fifo_22_full),
    .error        (_offsetQueueVec_queue_fifo_22_error),
    .data_out     (offsetQueueVec_22_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_23 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_23_enq_ready & offsetQueueVec_23_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_23_deq_ready & ~_offsetQueueVec_queue_fifo_23_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_23_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_23_empty),
    .almost_empty (offsetQueueVec_23_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_23_almostFull),
    .full         (_offsetQueueVec_queue_fifo_23_full),
    .error        (_offsetQueueVec_queue_fifo_23_error),
    .data_out     (offsetQueueVec_23_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_24 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_24_enq_ready & offsetQueueVec_24_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_24_deq_ready & ~_offsetQueueVec_queue_fifo_24_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_24_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_24_empty),
    .almost_empty (offsetQueueVec_24_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_24_almostFull),
    .full         (_offsetQueueVec_queue_fifo_24_full),
    .error        (_offsetQueueVec_queue_fifo_24_error),
    .data_out     (offsetQueueVec_24_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_25 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_25_enq_ready & offsetQueueVec_25_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_25_deq_ready & ~_offsetQueueVec_queue_fifo_25_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_25_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_25_empty),
    .almost_empty (offsetQueueVec_25_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_25_almostFull),
    .full         (_offsetQueueVec_queue_fifo_25_full),
    .error        (_offsetQueueVec_queue_fifo_25_error),
    .data_out     (offsetQueueVec_25_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_26 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_26_enq_ready & offsetQueueVec_26_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_26_deq_ready & ~_offsetQueueVec_queue_fifo_26_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_26_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_26_empty),
    .almost_empty (offsetQueueVec_26_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_26_almostFull),
    .full         (_offsetQueueVec_queue_fifo_26_full),
    .error        (_offsetQueueVec_queue_fifo_26_error),
    .data_out     (offsetQueueVec_26_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_27 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_27_enq_ready & offsetQueueVec_27_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_27_deq_ready & ~_offsetQueueVec_queue_fifo_27_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_27_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_27_empty),
    .almost_empty (offsetQueueVec_27_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_27_almostFull),
    .full         (_offsetQueueVec_queue_fifo_27_full),
    .error        (_offsetQueueVec_queue_fifo_27_error),
    .data_out     (offsetQueueVec_27_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_28 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_28_enq_ready & offsetQueueVec_28_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_28_deq_ready & ~_offsetQueueVec_queue_fifo_28_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_28_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_28_empty),
    .almost_empty (offsetQueueVec_28_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_28_almostFull),
    .full         (_offsetQueueVec_queue_fifo_28_full),
    .error        (_offsetQueueVec_queue_fifo_28_error),
    .data_out     (offsetQueueVec_28_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_29 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_29_enq_ready & offsetQueueVec_29_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_29_deq_ready & ~_offsetQueueVec_queue_fifo_29_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_29_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_29_empty),
    .almost_empty (offsetQueueVec_29_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_29_almostFull),
    .full         (_offsetQueueVec_queue_fifo_29_full),
    .error        (_offsetQueueVec_queue_fifo_29_error),
    .data_out     (offsetQueueVec_29_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_30 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_30_enq_ready & offsetQueueVec_30_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_30_deq_ready & ~_offsetQueueVec_queue_fifo_30_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_30_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_30_empty),
    .almost_empty (offsetQueueVec_30_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_30_almostFull),
    .full         (_offsetQueueVec_queue_fifo_30_full),
    .error        (_offsetQueueVec_queue_fifo_30_error),
    .data_out     (offsetQueueVec_30_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) offsetQueueVec_queue_fifo_31 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(offsetQueueVec_31_enq_ready & offsetQueueVec_31_enq_valid)),
    .pop_req_n    (~(offsetQueueVec_31_deq_ready & ~_offsetQueueVec_queue_fifo_31_empty)),
    .diag_n       (1'h1),
    .data_in      (offsetQueueVec_31_enq_bits),
    .empty        (_offsetQueueVec_queue_fifo_31_empty),
    .almost_empty (offsetQueueVec_31_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (offsetQueueVec_31_almostFull),
    .full         (_offsetQueueVec_queue_fifo_31_full),
    .error        (_offsetQueueVec_queue_fifo_31_error),
    .data_out     (offsetQueueVec_31_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(6),
    .err_mode(2),
    .rst_mode(3),
    .width(74)
  ) s1EnqQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~s0DequeueFire),
    .pop_req_n    (~(s1EnqQueue_deq_ready & ~_s1EnqQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (s1EnqQueue_dataIn),
    .empty        (_s1EnqQueue_fifo_empty),
    .almost_empty (s1EnqQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (s1EnqQueue_almostFull),
    .full         (_s1EnqQueue_fifo_full),
    .error        (_s1EnqQueue_fifo_error),
    .data_out     (_s1EnqQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(6),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) s1EnqDataQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(s1EnqDataQueue_enq_ready & s1EnqDataQueue_enq_valid)),
    .pop_req_n    (~(s1EnqDataQueue_deq_ready & ~_s1EnqDataQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (s1EnqDataQueue_enq_bits),
    .empty        (_s1EnqDataQueue_fifo_empty),
    .almost_empty (s1EnqDataQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (s1EnqDataQueue_almostFull),
    .full         (_s1EnqDataQueue_fifo_full),
    .error        (_s1EnqDataQueue_fifo_error),
    .data_out     (s1EnqDataQueue_deq_bits)
  );
  assign vrfReadDataPorts_valid = vrfReadDataPorts_valid_0;
  assign vrfReadDataPorts_bits_vs = vrfReadDataPorts_bits_vs_0;
  assign vrfReadDataPorts_bits_offset = vrfReadDataPorts_bits_offset_0;
  assign vrfReadDataPorts_bits_instructionIndex = vrfReadDataPorts_bits_instructionIndex_0;
  assign maskSelect_valid = maskGroupEndAndRequestNewMask;
  assign maskSelect_bits = nextGroupIndex[3:0];
  assign memReadRequest_valid = memReadRequest_valid_0;
  assign memReadRequest_bits_address = memReadRequest_bits_address_0;
  assign memReadRequest_bits_source = memReadRequest_bits_source_0;
  assign memReadResponse_ready = memReadResponse_ready_0;
  assign memWriteRequest_valid = memWriteRequest_valid_0;
  assign memWriteRequest_bits_data = memWriteRequest_bits_data_0;
  assign memWriteRequest_bits_mask = memWriteRequest_bits_mask_0;
  assign memWriteRequest_bits_source = memWriteRequest_bits_source_0;
  assign memWriteRequest_bits_address = memWriteRequest_bits_address_0;
  assign memWriteRequest_bits_size = memWriteRequest_bits_size_0;
  assign vrfWritePort_valid = vrfWritePort_valid_0;
  assign vrfWritePort_bits_vd = vrfWritePort_bits_vd_0;
  assign vrfWritePort_bits_offset = vrfWritePort_bits_offset_0;
  assign vrfWritePort_bits_mask = vrfWritePort_bits_mask_0;
  assign vrfWritePort_bits_data = vrfWritePort_bits_data_0;
  assign vrfWritePort_bits_last = vrfWritePort_bits_last_0;
  assign vrfWritePort_bits_instructionIndex = vrfWritePort_bits_instructionIndex_0;
  assign status_idle = stateIdle;
  assign status_last = _status_last_output;
  assign status_instructionIndex = lsuRequestReg_instructionIndex;
  assign status_targetLane = 32'h1 << (lsuRequestReg_instructionInformation_isStore ? s0Reg_offsetForLane : loadBaseByteOffset[6:2]);
  assign status_isStore = lsuRequestReg_instructionInformation_isStore;
  assign offsetRelease_0 = _allElementsMasked_T_1;
  assign offsetRelease_1 = _allElementsMasked_T_2;
  assign offsetRelease_2 = _allElementsMasked_T_3;
  assign offsetRelease_3 = _allElementsMasked_T_4;
  assign offsetRelease_4 = _allElementsMasked_T_5;
  assign offsetRelease_5 = _allElementsMasked_T_6;
  assign offsetRelease_6 = _allElementsMasked_T_7;
  assign offsetRelease_7 = _allElementsMasked_T_8;
  assign offsetRelease_8 = _allElementsMasked_T_9;
  assign offsetRelease_9 = _allElementsMasked_T_10;
  assign offsetRelease_10 = _allElementsMasked_T_11;
  assign offsetRelease_11 = _allElementsMasked_T_12;
  assign offsetRelease_12 = _allElementsMasked_T_13;
  assign offsetRelease_13 = _allElementsMasked_T_14;
  assign offsetRelease_14 = _allElementsMasked_T_15;
  assign offsetRelease_15 = _allElementsMasked_T_16;
  assign offsetRelease_16 = _allElementsMasked_T_17;
  assign offsetRelease_17 = _allElementsMasked_T_18;
  assign offsetRelease_18 = _allElementsMasked_T_19;
  assign offsetRelease_19 = _allElementsMasked_T_20;
  assign offsetRelease_20 = _allElementsMasked_T_21;
  assign offsetRelease_21 = _allElementsMasked_T_22;
  assign offsetRelease_22 = _allElementsMasked_T_23;
  assign offsetRelease_23 = _allElementsMasked_T_24;
  assign offsetRelease_24 = _allElementsMasked_T_25;
  assign offsetRelease_25 = _allElementsMasked_T_26;
  assign offsetRelease_26 = _allElementsMasked_T_27;
  assign offsetRelease_27 = _allElementsMasked_T_28;
  assign offsetRelease_28 = _allElementsMasked_T_29;
  assign offsetRelease_29 = _allElementsMasked_T_30;
  assign offsetRelease_30 = _allElementsMasked_T_31;
  assign offsetRelease_31 = _allElementsMasked_T_32;
endmodule

