module VectorDecoder(
  input  [31:0] decodeInput,
  output        decodeResult_orderReduce,
                decodeResult_floatMul,
  output [1:0]  decodeResult_fpExecutionType,
  output        decodeResult_float,
                decodeResult_specialSlot,
  output [4:0]  decodeResult_topUop,
  output        decodeResult_popCount,
                decodeResult_ffo,
                decodeResult_average,
                decodeResult_reverse,
                decodeResult_dontNeedExecuteInLane,
                decodeResult_scheduler,
                decodeResult_sReadVD,
                decodeResult_vtype,
                decodeResult_sWrite,
                decodeResult_crossRead,
                decodeResult_crossWrite,
                decodeResult_maskUnit,
                decodeResult_special,
                decodeResult_saturate,
                decodeResult_vwmacc,
                decodeResult_readOnly,
                decodeResult_maskSource,
                decodeResult_maskDestination,
                decodeResult_maskLogic,
  output [3:0]  decodeResult_uop,
  output        decodeResult_iota,
                decodeResult_mv,
                decodeResult_extend,
                decodeResult_unOrderWrite,
                decodeResult_compress,
                decodeResult_gather16,
                decodeResult_gather,
                decodeResult_slid,
                decodeResult_targetRd,
                decodeResult_widenReduce,
                decodeResult_red,
                decodeResult_nr,
                decodeResult_itype,
                decodeResult_unsigned1,
                decodeResult_unsigned0,
                decodeResult_other,
                decodeResult_multiCycle,
                decodeResult_divider,
                decodeResult_multiplier,
                decodeResult_shift,
                decodeResult_adder,
                decodeResult_logic
);

  wire [31:0] decodeResult_plaInput = decodeInput;
  wire [31:0] decodeResult_invInputs = ~decodeResult_plaInput;
  wire [55:0] decodeResult_invMatrixOutputs;
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0 = decodeResult_invInputs[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_8 = decodeResult_invInputs[4];
  wire        decodeResult_andMatrixOutputs_96_2 = decodeResult_andMatrixOutputs_andMatrixInput_0;
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_1 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_2 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_4 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_5 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_6 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_7 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_11 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_13 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_15 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_16 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_17 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_38 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_39 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_41 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_42 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_44 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_46 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_60 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_61 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_66 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_73 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_74 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_79 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_99 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_101 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_103 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_104 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_107 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_110 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_111 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_112 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_113 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_114 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_115 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_116 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_117 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_118 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_122 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_128 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_129 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_130 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_131 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_133 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_134 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_135 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_136 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_142 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_143 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_144 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_145 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_147 = decodeResult_plaInput[4];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_1 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_4 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_10 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_12 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_19 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_20 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_21 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_22 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_23 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_34 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_37 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_40 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_40 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_45 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_49 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_51 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_53 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_56 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_58 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_59 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_60 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_64 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_65 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_65 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_68 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_72 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_73 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_86 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_87 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_95 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_96 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_98 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_98 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_102 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_102 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_105 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_109 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_109 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_110 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_111 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_115 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_121 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_123 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_126 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_127 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_127 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_132 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_134 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_135 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_137 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_138 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_140 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_141 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_146 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_148 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_149 = decodeResult_invInputs[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_2 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_7 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_8 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_16 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_28 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_38 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_48 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_53 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_54 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_57 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_60 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_61 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_62 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_63 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_65 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_66 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_67 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_69 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_70 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_73 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_74 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_75 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_76 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_79 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_80 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_80 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_82 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_83 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_106 = decodeResult_invInputs[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_117 = decodeResult_invInputs[14];
  wire [1:0]  decodeResult_andMatrixOutputs_hi = {decodeResult_andMatrixOutputs_andMatrixInput_0_1, decodeResult_andMatrixOutputs_andMatrixInput_1};
  wire        decodeResult_andMatrixOutputs_62_2 = &{decodeResult_andMatrixOutputs_hi, decodeResult_andMatrixOutputs_andMatrixInput_2};
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_1 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_2 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_3 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_8 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_11 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_13 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_17 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_21 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_29 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_37 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_36 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_37 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_42 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_42 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_47 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_49 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_54 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_59 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_59 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_61 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_62 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_68 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_69 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_70 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_74 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_76 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_77 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_77 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_81 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_84 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_85 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_86 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_94 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_95 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_96 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_97 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_97 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_99 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_99 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_104 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_106 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_109 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_110 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_111 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_118 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_119 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_122 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_123 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_126 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_126 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_127 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_130 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_131 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_133 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_136 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_139 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_140 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_144 = decodeResult_invInputs[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_1 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_2 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_3 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_4 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_8 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_11 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_14 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_19 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_20 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_23 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_36 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_36 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_40 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_44 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_49 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_55 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_52 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_56 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_57 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_61 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_62 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_64 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_68 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_63 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_75 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_76 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_78 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_42 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_84 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_86 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_88 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_88 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_91 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_100 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_105 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_108 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_106 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_112 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_113 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_112 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_118 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_124 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_141 = decodeResult_invInputs[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_1 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_2 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_3 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_4 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_5 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_7 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_7 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_10 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_11 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_8 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_13 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_15 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_17 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_18 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_19 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_20 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_23 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_21 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_18 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_25 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_31 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_28 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_29 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_53 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_54 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_55 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_56 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_23 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7_8 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_59 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_60 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7_9 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7_10 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_27 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_55 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_29 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_66 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_67 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_32 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_60 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_61 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_62 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_64 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_65 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_67 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_68 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_81 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_84 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_87 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_86 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_89 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_88 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_103 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_105 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_106 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_108 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_110 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_111 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_116 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_115 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_120 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_121 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_118 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_142 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_136 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_145 = decodeResult_invInputs[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_3 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_4 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_8 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7_2 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7_3 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_9 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_16 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_15 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_16 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_19 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_20 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_17 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_24 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_10 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_19 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_21 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_27 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_24 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_25 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_11 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_12 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_13 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_14 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7_5 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_32 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7_6 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_34 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_35 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_37 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_17 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_39 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_40 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_42 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_19 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_20 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_21 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_22 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_8_1 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_9 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_9_1 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_9_2 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_8_5 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7_12 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_8_6 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_30 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_31 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_8_7 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7_15 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7_16 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_8_8 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7_18 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7_19 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_9_3 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7_21 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7_22 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_9_4 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_43 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_71 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_44 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_45 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_74 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_46 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_77 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_47 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_79 = decodeResult_invInputs[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_49 = decodeResult_invInputs[31];
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi = {decodeResult_andMatrixOutputs_andMatrixInput_3, decodeResult_andMatrixOutputs_andMatrixInput_4};
  wire [2:0]  decodeResult_andMatrixOutputs_lo = {decodeResult_andMatrixOutputs_lo_hi, decodeResult_andMatrixOutputs_andMatrixInput_5};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi = {decodeResult_andMatrixOutputs_andMatrixInput_0_2, decodeResult_andMatrixOutputs_andMatrixInput_1_1};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_1 = {decodeResult_andMatrixOutputs_hi_hi, decodeResult_andMatrixOutputs_andMatrixInput_2_1};
  wire        decodeResult_andMatrixOutputs_15_2 = &{decodeResult_andMatrixOutputs_hi_1, decodeResult_andMatrixOutputs_lo};
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_3 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_3 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_5 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_9 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_12 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_14 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_14 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_16 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_18 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_24 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_26 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_27 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_30 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_31 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_32 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_35 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_36 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_38 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_41 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_43 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_43 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_48 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_50 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_62 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_63 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_67 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_69 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_70 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_71 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_75 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_76 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_77 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_78 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_78 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_82 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_85 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_90 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_91 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_92 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_97 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_100 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_100 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_103 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_106 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_108 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_112 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_116 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_117 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_119 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_120 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_121 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_124 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_125 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_128 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_129 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_132 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_133 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_139 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_141 = decodeResult_plaInput[12];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_142 = decodeResult_plaInput[12];
  wire [1:0]  decodeResult_andMatrixOutputs_hi_2 = {decodeResult_andMatrixOutputs_andMatrixInput_0_3, decodeResult_andMatrixOutputs_andMatrixInput_1_2};
  wire        decodeResult_andMatrixOutputs_89_2 = &{decodeResult_andMatrixOutputs_hi_2, decodeResult_andMatrixOutputs_andMatrixInput_2_2};
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_1 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_1 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_3 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_2 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_6 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_6 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_7 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7_4 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_14 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_17 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_18 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_21 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_22 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_20 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_29 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_22 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_23 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_30 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_31 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_26 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_27 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_28 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_29 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_30 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_16 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_43 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_44 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_46 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_49 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_51 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_104 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_88 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_89 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_90 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_112 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_116 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_117 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_100 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_122 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_103 = decodeResult_invInputs[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_107 = decodeResult_invInputs[30];
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_1 = {decodeResult_andMatrixOutputs_andMatrixInput_4_1, decodeResult_andMatrixOutputs_andMatrixInput_5_1};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_1 = {decodeResult_andMatrixOutputs_lo_hi_1, decodeResult_andMatrixOutputs_andMatrixInput_6};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo = {decodeResult_andMatrixOutputs_andMatrixInput_2_3, decodeResult_andMatrixOutputs_andMatrixInput_3_1};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_1 = {decodeResult_andMatrixOutputs_andMatrixInput_0_4, decodeResult_andMatrixOutputs_andMatrixInput_1_3};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_3 = {decodeResult_andMatrixOutputs_hi_hi_1, decodeResult_andMatrixOutputs_hi_lo};
  wire        decodeResult_andMatrixOutputs_110_2 = &{decodeResult_andMatrixOutputs_hi_3, decodeResult_andMatrixOutputs_lo_1};
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_4 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_5 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_6 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_9 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_15 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_15 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_18 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_25 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_25 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_26 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_28 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_29 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_33 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_34 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_35 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_39 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_39 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_40 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_45 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_44 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_50 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_52 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_55 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_63 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_64 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_64 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_66 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_67 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_71 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_75 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_80 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_81 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_83 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_84 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_89 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_90 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_91 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_94 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_101 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_101 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_102 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_105 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_107 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_108 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_113 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_114 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_114 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_115 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_116 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_120 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_120 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_125 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_128 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_131 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_132 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_134 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_137 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_138 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_140 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_143 = decodeResult_plaInput[13];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_2 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_18 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_22 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_24 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_25 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_25 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_28 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_35 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_37 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_47 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_51 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_49 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_55 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_58 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_48 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_24 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_85 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_89 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_96 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_98 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_97 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_100 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_101 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_110 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_121 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_123 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_125 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_127 = decodeResult_invInputs[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_124 = decodeResult_invInputs[27];
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo = {decodeResult_andMatrixOutputs_andMatrixInput_6_1, decodeResult_andMatrixOutputs_andMatrixInput_7};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_2 = {decodeResult_andMatrixOutputs_andMatrixInput_4_2, decodeResult_andMatrixOutputs_andMatrixInput_5_2};
  wire [3:0]  decodeResult_andMatrixOutputs_lo_2 = {decodeResult_andMatrixOutputs_lo_hi_2, decodeResult_andMatrixOutputs_lo_lo};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_1 = {decodeResult_andMatrixOutputs_andMatrixInput_2_4, decodeResult_andMatrixOutputs_andMatrixInput_3_2};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_2 = {decodeResult_andMatrixOutputs_andMatrixInput_0_5, decodeResult_andMatrixOutputs_andMatrixInput_1_4};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_4 = {decodeResult_andMatrixOutputs_hi_hi_2, decodeResult_andMatrixOutputs_hi_lo_1};
  wire        decodeResult_andMatrixOutputs_93_2 = &{decodeResult_andMatrixOutputs_hi_4, decodeResult_andMatrixOutputs_lo_2};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_3 = {decodeResult_andMatrixOutputs_andMatrixInput_3_3, decodeResult_andMatrixOutputs_andMatrixInput_4_3};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_3 = {decodeResult_andMatrixOutputs_andMatrixInput_0_6, decodeResult_andMatrixOutputs_andMatrixInput_1_5};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_5 = {decodeResult_andMatrixOutputs_hi_hi_3, decodeResult_andMatrixOutputs_andMatrixInput_2_5};
  wire        decodeResult_andMatrixOutputs_74_2 = &{decodeResult_andMatrixOutputs_hi_5, decodeResult_andMatrixOutputs_lo_3};
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_6 = decodeResult_plaInput[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_10 = decodeResult_plaInput[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_11 = decodeResult_plaInput[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_27 = decodeResult_plaInput[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_30 = decodeResult_plaInput[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_31 = decodeResult_plaInput[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_52 = decodeResult_plaInput[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_57 = decodeResult_plaInput[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_72 = decodeResult_plaInput[14];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_4 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_5 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_6 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_7 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_8 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_8 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7_1 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_9 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_11 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_12 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_12 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_14 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_35 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_34 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_38 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_39 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_31 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_41 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_40 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_43 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_44 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_25 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_56 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_69 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_69 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_77 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_93 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_95 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_99 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_100 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_105 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_107 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_108 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_111 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_113 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_114 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_124 = decodeResult_invInputs[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_126 = decodeResult_invInputs[28];
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_3 = {decodeResult_andMatrixOutputs_andMatrixInput_3_4, decodeResult_andMatrixOutputs_andMatrixInput_4_4};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_4 = {decodeResult_andMatrixOutputs_lo_hi_3, decodeResult_andMatrixOutputs_andMatrixInput_5_3};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_4 = {decodeResult_andMatrixOutputs_andMatrixInput_0_7, decodeResult_andMatrixOutputs_andMatrixInput_1_6};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_6 = {decodeResult_andMatrixOutputs_hi_hi_4, decodeResult_andMatrixOutputs_andMatrixInput_2_6};
  wire        decodeResult_andMatrixOutputs_16_2 = &{decodeResult_andMatrixOutputs_hi_6, decodeResult_andMatrixOutputs_lo_4};
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_7 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_5 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_6 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_9 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_10 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_14 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_17 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_26 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_29 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_30 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_41 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_46 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_47 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_51 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_56 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_72 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_59 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_71 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_70 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_71 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_93 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_93 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_103 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_104 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_107 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_114 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_129 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_130 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_128 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_129 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_143 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_148 = decodeResult_plaInput[26];
  wire        decodeResult_andMatrixOutputs_82_2 = &{decodeResult_andMatrixOutputs_andMatrixInput_0_8, decodeResult_andMatrixOutputs_andMatrixInput_1_7};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_4 = {decodeResult_andMatrixOutputs_andMatrixInput_4_5, decodeResult_andMatrixOutputs_andMatrixInput_5_4};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_5 = {decodeResult_andMatrixOutputs_lo_hi_4, decodeResult_andMatrixOutputs_andMatrixInput_6_2};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_2 = {decodeResult_andMatrixOutputs_andMatrixInput_2_7, decodeResult_andMatrixOutputs_andMatrixInput_3_5};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_5 = {decodeResult_andMatrixOutputs_andMatrixInput_0_9, decodeResult_andMatrixOutputs_andMatrixInput_1_8};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_7 = {decodeResult_andMatrixOutputs_hi_hi_5, decodeResult_andMatrixOutputs_hi_lo_2};
  wire        decodeResult_andMatrixOutputs_114_2 = &{decodeResult_andMatrixOutputs_hi_7, decodeResult_andMatrixOutputs_lo_5};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_5 = {decodeResult_andMatrixOutputs_andMatrixInput_4_6, decodeResult_andMatrixOutputs_andMatrixInput_5_5};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_6 = {decodeResult_andMatrixOutputs_lo_hi_5, decodeResult_andMatrixOutputs_andMatrixInput_6_3};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_3 = {decodeResult_andMatrixOutputs_andMatrixInput_2_8, decodeResult_andMatrixOutputs_andMatrixInput_3_6};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_6 = {decodeResult_andMatrixOutputs_andMatrixInput_0_10, decodeResult_andMatrixOutputs_andMatrixInput_1_9};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_8 = {decodeResult_andMatrixOutputs_hi_hi_6, decodeResult_andMatrixOutputs_hi_lo_3};
  wire        decodeResult_andMatrixOutputs_22_2 = &{decodeResult_andMatrixOutputs_hi_8, decodeResult_andMatrixOutputs_lo_6};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_6 = {decodeResult_andMatrixOutputs_andMatrixInput_4_7, decodeResult_andMatrixOutputs_andMatrixInput_5_6};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_7 = {decodeResult_andMatrixOutputs_lo_hi_6, decodeResult_andMatrixOutputs_andMatrixInput_6_4};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_4 = {decodeResult_andMatrixOutputs_andMatrixInput_2_9, decodeResult_andMatrixOutputs_andMatrixInput_3_7};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_7 = {decodeResult_andMatrixOutputs_andMatrixInput_0_11, decodeResult_andMatrixOutputs_andMatrixInput_1_10};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_9 = {decodeResult_andMatrixOutputs_hi_hi_7, decodeResult_andMatrixOutputs_hi_lo_4};
  wire        decodeResult_andMatrixOutputs_6_2 = &{decodeResult_andMatrixOutputs_hi_9, decodeResult_andMatrixOutputs_lo_7};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_8 = {decodeResult_andMatrixOutputs_andMatrixInput_2_10, decodeResult_andMatrixOutputs_andMatrixInput_3_8};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_10 = {decodeResult_andMatrixOutputs_andMatrixInput_0_12, decodeResult_andMatrixOutputs_andMatrixInput_1_11};
  wire        decodeResult_andMatrixOutputs_64_2 = &{decodeResult_andMatrixOutputs_hi_10, decodeResult_andMatrixOutputs_lo_8};
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_9 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_5 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_10 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_12 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_13 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_13 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_15 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_33 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_32 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_33 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_34 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_38 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_43 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_42 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_45 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_46 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_52 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_54 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_50 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_56 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_54 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_36 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_73 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_74 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7_20 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_76 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_79 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7_23 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_94 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_95 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_102 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_103 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_104 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_115 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_119 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_117 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_125 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_130 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_131 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_138 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_139 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_140 = decodeResult_plaInput[27];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_147 = decodeResult_plaInput[27];
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_7 = {decodeResult_andMatrixOutputs_andMatrixInput_3_9, decodeResult_andMatrixOutputs_andMatrixInput_4_8};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_9 = {decodeResult_andMatrixOutputs_lo_hi_7, decodeResult_andMatrixOutputs_andMatrixInput_5_7};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_8 = {decodeResult_andMatrixOutputs_andMatrixInput_0_13, decodeResult_andMatrixOutputs_andMatrixInput_1_12};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_11 = {decodeResult_andMatrixOutputs_hi_hi_8, decodeResult_andMatrixOutputs_andMatrixInput_2_11};
  wire        decodeResult_andMatrixOutputs_50_2 = &{decodeResult_andMatrixOutputs_hi_11, decodeResult_andMatrixOutputs_lo_9};
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_13 = decodeResult_invInputs[15];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_58 = decodeResult_invInputs[15];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_60 = decodeResult_invInputs[15];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_64 = decodeResult_invInputs[15];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_68 = decodeResult_invInputs[15];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_67 = decodeResult_invInputs[15];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_88 = decodeResult_invInputs[15];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_12 = decodeResult_invInputs[16];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_59 = decodeResult_invInputs[16];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_58 = decodeResult_invInputs[16];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_61 = decodeResult_invInputs[16];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_78 = decodeResult_invInputs[16];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_75 = decodeResult_invInputs[16];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_87 = decodeResult_invInputs[16];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_10 = decodeResult_invInputs[18];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_53 = decodeResult_invInputs[18];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_63 = decodeResult_invInputs[18];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_74 = decodeResult_invInputs[18];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_66 = decodeResult_invInputs[18];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_78 = decodeResult_invInputs[18];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_9 = decodeResult_invInputs[19];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_57 = decodeResult_invInputs[19];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_57 = decodeResult_invInputs[19];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_49 = decodeResult_invInputs[19];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_26 = decodeResult_invInputs[19];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_54 = decodeResult_invInputs[19];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_68 = decodeResult_invInputs[19];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_72 = decodeResult_invInputs[19];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_39 = decodeResult_invInputs[19];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_69 = decodeResult_invInputs[19];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_89 = decodeResult_invInputs[19];
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo_1 = {decodeResult_andMatrixOutputs_andMatrixInput_7_1, decodeResult_andMatrixOutputs_andMatrixInput_8};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_8 = {decodeResult_andMatrixOutputs_andMatrixInput_5_8, decodeResult_andMatrixOutputs_andMatrixInput_6_5};
  wire [3:0]  decodeResult_andMatrixOutputs_lo_10 = {decodeResult_andMatrixOutputs_lo_hi_8, decodeResult_andMatrixOutputs_lo_lo_1};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_5 = {decodeResult_andMatrixOutputs_andMatrixInput_3_10, decodeResult_andMatrixOutputs_andMatrixInput_4_9};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_hi = {decodeResult_andMatrixOutputs_andMatrixInput_0_14, decodeResult_andMatrixOutputs_andMatrixInput_1_13};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_hi_9 = {decodeResult_andMatrixOutputs_hi_hi_hi, decodeResult_andMatrixOutputs_andMatrixInput_2_12};
  wire [4:0]  decodeResult_andMatrixOutputs_hi_12 = {decodeResult_andMatrixOutputs_hi_hi_9, decodeResult_andMatrixOutputs_hi_lo_5};
  wire        decodeResult_andMatrixOutputs_44_2 = &{decodeResult_andMatrixOutputs_hi_12, decodeResult_andMatrixOutputs_lo_10};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo_2 = {decodeResult_andMatrixOutputs_andMatrixInput_6_6, decodeResult_andMatrixOutputs_andMatrixInput_7_2};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_9 = {decodeResult_andMatrixOutputs_andMatrixInput_4_10, decodeResult_andMatrixOutputs_andMatrixInput_5_9};
  wire [3:0]  decodeResult_andMatrixOutputs_lo_11 = {decodeResult_andMatrixOutputs_lo_hi_9, decodeResult_andMatrixOutputs_lo_lo_2};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_6 = {decodeResult_andMatrixOutputs_andMatrixInput_2_13, decodeResult_andMatrixOutputs_andMatrixInput_3_11};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_10 = {decodeResult_andMatrixOutputs_andMatrixInput_0_15, decodeResult_andMatrixOutputs_andMatrixInput_1_14};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_13 = {decodeResult_andMatrixOutputs_hi_hi_10, decodeResult_andMatrixOutputs_hi_lo_6};
  wire        decodeResult_andMatrixOutputs_138_2 = &{decodeResult_andMatrixOutputs_hi_13, decodeResult_andMatrixOutputs_lo_11};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo_3 = {decodeResult_andMatrixOutputs_andMatrixInput_6_7, decodeResult_andMatrixOutputs_andMatrixInput_7_3};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_10 = {decodeResult_andMatrixOutputs_andMatrixInput_4_11, decodeResult_andMatrixOutputs_andMatrixInput_5_10};
  wire [3:0]  decodeResult_andMatrixOutputs_lo_12 = {decodeResult_andMatrixOutputs_lo_hi_10, decodeResult_andMatrixOutputs_lo_lo_3};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_7 = {decodeResult_andMatrixOutputs_andMatrixInput_2_14, decodeResult_andMatrixOutputs_andMatrixInput_3_12};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_11 = {decodeResult_andMatrixOutputs_andMatrixInput_0_16, decodeResult_andMatrixOutputs_andMatrixInput_1_15};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_14 = {decodeResult_andMatrixOutputs_hi_hi_11, decodeResult_andMatrixOutputs_hi_lo_7};
  wire        decodeResult_andMatrixOutputs_30_2 = &{decodeResult_andMatrixOutputs_hi_14, decodeResult_andMatrixOutputs_lo_12};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_11 = {decodeResult_andMatrixOutputs_andMatrixInput_3_13, decodeResult_andMatrixOutputs_andMatrixInput_4_12};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_13 = {decodeResult_andMatrixOutputs_lo_hi_11, decodeResult_andMatrixOutputs_andMatrixInput_5_11};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_12 = {decodeResult_andMatrixOutputs_andMatrixInput_0_17, decodeResult_andMatrixOutputs_andMatrixInput_1_16};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_15 = {decodeResult_andMatrixOutputs_hi_hi_12, decodeResult_andMatrixOutputs_andMatrixInput_2_15};
  wire        decodeResult_andMatrixOutputs_25_2 = &{decodeResult_andMatrixOutputs_hi_15, decodeResult_andMatrixOutputs_lo_13};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo_4 = {decodeResult_andMatrixOutputs_andMatrixInput_6_8, decodeResult_andMatrixOutputs_andMatrixInput_7_4};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_12 = {decodeResult_andMatrixOutputs_andMatrixInput_4_13, decodeResult_andMatrixOutputs_andMatrixInput_5_12};
  wire [3:0]  decodeResult_andMatrixOutputs_lo_14 = {decodeResult_andMatrixOutputs_lo_hi_12, decodeResult_andMatrixOutputs_lo_lo_4};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_8 = {decodeResult_andMatrixOutputs_andMatrixInput_2_16, decodeResult_andMatrixOutputs_andMatrixInput_3_14};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_13 = {decodeResult_andMatrixOutputs_andMatrixInput_0_18, decodeResult_andMatrixOutputs_andMatrixInput_1_17};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_16 = {decodeResult_andMatrixOutputs_hi_hi_13, decodeResult_andMatrixOutputs_hi_lo_8};
  wire        decodeResult_andMatrixOutputs_0_2 = &{decodeResult_andMatrixOutputs_hi_16, decodeResult_andMatrixOutputs_lo_14};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_13 = {decodeResult_andMatrixOutputs_andMatrixInput_4_14, decodeResult_andMatrixOutputs_andMatrixInput_5_13};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_15 = {decodeResult_andMatrixOutputs_lo_hi_13, decodeResult_andMatrixOutputs_andMatrixInput_6_9};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_9 = {decodeResult_andMatrixOutputs_andMatrixInput_2_17, decodeResult_andMatrixOutputs_andMatrixInput_3_15};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_14 = {decodeResult_andMatrixOutputs_andMatrixInput_0_19, decodeResult_andMatrixOutputs_andMatrixInput_1_18};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_17 = {decodeResult_andMatrixOutputs_hi_hi_14, decodeResult_andMatrixOutputs_hi_lo_9};
  wire        decodeResult_andMatrixOutputs_92_2 = &{decodeResult_andMatrixOutputs_hi_17, decodeResult_andMatrixOutputs_lo_15};
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_16 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_19 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_20 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_21 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_22 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_24 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_22 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_23 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_26 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_23 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_24 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_27 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_26 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_32 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_30 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_31 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_32 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_47 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_48 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_45 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_50 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_47 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_50 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_53 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_41 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_55 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_52 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_81 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_82 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_83 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_87 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_85 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_86 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_90 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_88 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_92 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_90 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_91 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_92 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_118 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_122 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_123 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_124 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_122 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_135 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_136 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_137 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_135 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_136 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_146 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_147 = decodeResult_plaInput[28];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_144 = decodeResult_plaInput[28];
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_14 = {decodeResult_andMatrixOutputs_andMatrixInput_3_16, decodeResult_andMatrixOutputs_andMatrixInput_4_15};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_16 = {decodeResult_andMatrixOutputs_lo_hi_14, decodeResult_andMatrixOutputs_andMatrixInput_5_14};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_15 = {decodeResult_andMatrixOutputs_andMatrixInput_0_20, decodeResult_andMatrixOutputs_andMatrixInput_1_19};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_18 = {decodeResult_andMatrixOutputs_hi_hi_15, decodeResult_andMatrixOutputs_andMatrixInput_2_18};
  wire        decodeResult_andMatrixOutputs_24_2 = &{decodeResult_andMatrixOutputs_hi_18, decodeResult_andMatrixOutputs_lo_16};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_17 = {decodeResult_andMatrixOutputs_andMatrixInput_3_17, decodeResult_andMatrixOutputs_andMatrixInput_4_16};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_16 = {decodeResult_andMatrixOutputs_andMatrixInput_0_21, decodeResult_andMatrixOutputs_andMatrixInput_1_20};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_19 = {decodeResult_andMatrixOutputs_hi_hi_16, decodeResult_andMatrixOutputs_andMatrixInput_2_19};
  wire        decodeResult_andMatrixOutputs_23_2 = &{decodeResult_andMatrixOutputs_hi_19, decodeResult_andMatrixOutputs_lo_17};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_15 = {decodeResult_andMatrixOutputs_andMatrixInput_3_18, decodeResult_andMatrixOutputs_andMatrixInput_4_17};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_18 = {decodeResult_andMatrixOutputs_lo_hi_15, decodeResult_andMatrixOutputs_andMatrixInput_5_15};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_17 = {decodeResult_andMatrixOutputs_andMatrixInput_0_22, decodeResult_andMatrixOutputs_andMatrixInput_1_21};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_20 = {decodeResult_andMatrixOutputs_hi_hi_17, decodeResult_andMatrixOutputs_andMatrixInput_2_20};
  wire        decodeResult_andMatrixOutputs_58_2 = &{decodeResult_andMatrixOutputs_hi_20, decodeResult_andMatrixOutputs_lo_18};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_16 = {decodeResult_andMatrixOutputs_andMatrixInput_3_19, decodeResult_andMatrixOutputs_andMatrixInput_4_18};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_19 = {decodeResult_andMatrixOutputs_lo_hi_16, decodeResult_andMatrixOutputs_andMatrixInput_5_16};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_18 = {decodeResult_andMatrixOutputs_andMatrixInput_0_23, decodeResult_andMatrixOutputs_andMatrixInput_1_22};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_21 = {decodeResult_andMatrixOutputs_hi_hi_18, decodeResult_andMatrixOutputs_andMatrixInput_2_21};
  wire        decodeResult_andMatrixOutputs_45_2 = &{decodeResult_andMatrixOutputs_hi_21, decodeResult_andMatrixOutputs_lo_19};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_20 = {decodeResult_andMatrixOutputs_andMatrixInput_3_20, decodeResult_andMatrixOutputs_andMatrixInput_4_19};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_19 = {decodeResult_andMatrixOutputs_andMatrixInput_0_24, decodeResult_andMatrixOutputs_andMatrixInput_1_23};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_22 = {decodeResult_andMatrixOutputs_hi_hi_19, decodeResult_andMatrixOutputs_andMatrixInput_2_22};
  wire        decodeResult_andMatrixOutputs_10_2 = &{decodeResult_andMatrixOutputs_hi_22, decodeResult_andMatrixOutputs_lo_20};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_21 = {decodeResult_andMatrixOutputs_andMatrixInput_3_21, decodeResult_andMatrixOutputs_andMatrixInput_4_20};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_20 = {decodeResult_andMatrixOutputs_andMatrixInput_0_25, decodeResult_andMatrixOutputs_andMatrixInput_1_24};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_23 = {decodeResult_andMatrixOutputs_hi_hi_20, decodeResult_andMatrixOutputs_andMatrixInput_2_23};
  wire        decodeResult_andMatrixOutputs_123_2 = &{decodeResult_andMatrixOutputs_hi_23, decodeResult_andMatrixOutputs_lo_21};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_22 = {decodeResult_andMatrixOutputs_andMatrixInput_3_22, decodeResult_andMatrixOutputs_andMatrixInput_4_21};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_21 = {decodeResult_andMatrixOutputs_andMatrixInput_0_26, decodeResult_andMatrixOutputs_andMatrixInput_1_25};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_24 = {decodeResult_andMatrixOutputs_hi_hi_21, decodeResult_andMatrixOutputs_andMatrixInput_2_24};
  wire        decodeResult_andMatrixOutputs_128_2 = &{decodeResult_andMatrixOutputs_hi_24, decodeResult_andMatrixOutputs_lo_22};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_17 = {decodeResult_andMatrixOutputs_andMatrixInput_3_23, decodeResult_andMatrixOutputs_andMatrixInput_4_22};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_23 = {decodeResult_andMatrixOutputs_lo_hi_17, decodeResult_andMatrixOutputs_andMatrixInput_5_17};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_22 = {decodeResult_andMatrixOutputs_andMatrixInput_0_27, decodeResult_andMatrixOutputs_andMatrixInput_1_26};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_25 = {decodeResult_andMatrixOutputs_hi_hi_22, decodeResult_andMatrixOutputs_andMatrixInput_2_25};
  wire        decodeResult_andMatrixOutputs_83_2 = &{decodeResult_andMatrixOutputs_hi_25, decodeResult_andMatrixOutputs_lo_23};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_24 = {decodeResult_andMatrixOutputs_andMatrixInput_2_26, decodeResult_andMatrixOutputs_andMatrixInput_3_24};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_26 = {decodeResult_andMatrixOutputs_andMatrixInput_0_28, decodeResult_andMatrixOutputs_andMatrixInput_1_27};
  wire        decodeResult_andMatrixOutputs_149_2 = &{decodeResult_andMatrixOutputs_hi_26, decodeResult_andMatrixOutputs_lo_24};
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_28 = decodeResult_plaInput[15];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_63 = decodeResult_plaInput[15];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_77 = decodeResult_plaInput[15];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_81 = decodeResult_plaInput[15];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_83 = decodeResult_plaInput[15];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_0_93 = decodeResult_plaInput[15];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_27 = decodeResult_plaInput[16];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_62 = decodeResult_plaInput[16];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_82 = decodeResult_plaInput[16];
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_18 = {decodeResult_andMatrixOutputs_andMatrixInput_4_23, decodeResult_andMatrixOutputs_andMatrixInput_5_18};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_25 = {decodeResult_andMatrixOutputs_lo_hi_18, decodeResult_andMatrixOutputs_andMatrixInput_6_10};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_10 = {decodeResult_andMatrixOutputs_andMatrixInput_2_27, decodeResult_andMatrixOutputs_andMatrixInput_3_25};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_23 = {decodeResult_andMatrixOutputs_andMatrixInput_0_29, decodeResult_andMatrixOutputs_andMatrixInput_1_28};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_27 = {decodeResult_andMatrixOutputs_hi_hi_23, decodeResult_andMatrixOutputs_hi_lo_10};
  wire        decodeResult_andMatrixOutputs_32_2 = &{decodeResult_andMatrixOutputs_hi_27, decodeResult_andMatrixOutputs_lo_25};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_19 = {decodeResult_andMatrixOutputs_andMatrixInput_3_26, decodeResult_andMatrixOutputs_andMatrixInput_4_24};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_26 = {decodeResult_andMatrixOutputs_lo_hi_19, decodeResult_andMatrixOutputs_andMatrixInput_5_19};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_24 = {decodeResult_andMatrixOutputs_andMatrixInput_0_30, decodeResult_andMatrixOutputs_andMatrixInput_1_29};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_28 = {decodeResult_andMatrixOutputs_hi_hi_24, decodeResult_andMatrixOutputs_andMatrixInput_2_28};
  wire        decodeResult_andMatrixOutputs_53_2 = &{decodeResult_andMatrixOutputs_hi_28, decodeResult_andMatrixOutputs_lo_26};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_20 = {decodeResult_andMatrixOutputs_andMatrixInput_3_27, decodeResult_andMatrixOutputs_andMatrixInput_4_25};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_27 = {decodeResult_andMatrixOutputs_lo_hi_20, decodeResult_andMatrixOutputs_andMatrixInput_5_20};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_25 = {decodeResult_andMatrixOutputs_andMatrixInput_0_31, decodeResult_andMatrixOutputs_andMatrixInput_1_30};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_29 = {decodeResult_andMatrixOutputs_hi_hi_25, decodeResult_andMatrixOutputs_andMatrixInput_2_29};
  wire        decodeResult_andMatrixOutputs_40_2 = &{decodeResult_andMatrixOutputs_hi_29, decodeResult_andMatrixOutputs_lo_27};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_21 = {decodeResult_andMatrixOutputs_andMatrixInput_3_28, decodeResult_andMatrixOutputs_andMatrixInput_4_26};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_28 = {decodeResult_andMatrixOutputs_lo_hi_21, decodeResult_andMatrixOutputs_andMatrixInput_5_21};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_26 = {decodeResult_andMatrixOutputs_andMatrixInput_0_32, decodeResult_andMatrixOutputs_andMatrixInput_1_31};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_30 = {decodeResult_andMatrixOutputs_hi_hi_26, decodeResult_andMatrixOutputs_andMatrixInput_2_30};
  wire        decodeResult_andMatrixOutputs_78_2 = &{decodeResult_andMatrixOutputs_hi_30, decodeResult_andMatrixOutputs_lo_28};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_29 = {decodeResult_andMatrixOutputs_andMatrixInput_3_29, decodeResult_andMatrixOutputs_andMatrixInput_4_27};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_27 = {decodeResult_andMatrixOutputs_andMatrixInput_0_33, decodeResult_andMatrixOutputs_andMatrixInput_1_32};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_31 = {decodeResult_andMatrixOutputs_hi_hi_27, decodeResult_andMatrixOutputs_andMatrixInput_2_31};
  wire        decodeResult_andMatrixOutputs_107_2 = &{decodeResult_andMatrixOutputs_hi_31, decodeResult_andMatrixOutputs_lo_29};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_22 = {decodeResult_andMatrixOutputs_andMatrixInput_3_30, decodeResult_andMatrixOutputs_andMatrixInput_4_28};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_30 = {decodeResult_andMatrixOutputs_lo_hi_22, decodeResult_andMatrixOutputs_andMatrixInput_5_22};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_28 = {decodeResult_andMatrixOutputs_andMatrixInput_0_34, decodeResult_andMatrixOutputs_andMatrixInput_1_33};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_32 = {decodeResult_andMatrixOutputs_hi_hi_28, decodeResult_andMatrixOutputs_andMatrixInput_2_32};
  wire        decodeResult_andMatrixOutputs_84_2 = &{decodeResult_andMatrixOutputs_hi_32, decodeResult_andMatrixOutputs_lo_30};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_23 = {decodeResult_andMatrixOutputs_andMatrixInput_3_31, decodeResult_andMatrixOutputs_andMatrixInput_4_29};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_31 = {decodeResult_andMatrixOutputs_lo_hi_23, decodeResult_andMatrixOutputs_andMatrixInput_5_23};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_29 = {decodeResult_andMatrixOutputs_andMatrixInput_0_35, decodeResult_andMatrixOutputs_andMatrixInput_1_34};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_33 = {decodeResult_andMatrixOutputs_hi_hi_29, decodeResult_andMatrixOutputs_andMatrixInput_2_33};
  wire        decodeResult_andMatrixOutputs_56_2 = &{decodeResult_andMatrixOutputs_hi_33, decodeResult_andMatrixOutputs_lo_31};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_24 = {decodeResult_andMatrixOutputs_andMatrixInput_3_32, decodeResult_andMatrixOutputs_andMatrixInput_4_30};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_32 = {decodeResult_andMatrixOutputs_lo_hi_24, decodeResult_andMatrixOutputs_andMatrixInput_5_24};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_30 = {decodeResult_andMatrixOutputs_andMatrixInput_0_36, decodeResult_andMatrixOutputs_andMatrixInput_1_35};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_34 = {decodeResult_andMatrixOutputs_hi_hi_30, decodeResult_andMatrixOutputs_andMatrixInput_2_34};
  wire        decodeResult_andMatrixOutputs_71_2 = &{decodeResult_andMatrixOutputs_hi_34, decodeResult_andMatrixOutputs_lo_32};
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_33 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_32 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_33 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_34 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_35 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_36 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_37 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_15 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_39 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_33 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_41 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_42 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_45 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_46 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_36 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_48 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_38 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_48 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_51 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_18 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_53 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_43 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_91 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_94 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_93 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_96 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_95 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_98 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_97 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_98 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_99 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_83 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_101 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_102 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_119 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_120 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_121 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_126 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_123 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_104 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_125 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_106 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_127 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_132 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_133 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_134 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_131 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_132 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_145 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_146 = decodeResult_plaInput[29];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_139 = decodeResult_plaInput[29];
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_25 = {decodeResult_andMatrixOutputs_andMatrixInput_3_33, decodeResult_andMatrixOutputs_andMatrixInput_4_31};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_33 = {decodeResult_andMatrixOutputs_lo_hi_25, decodeResult_andMatrixOutputs_andMatrixInput_5_25};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_31 = {decodeResult_andMatrixOutputs_andMatrixInput_0_37, decodeResult_andMatrixOutputs_andMatrixInput_1_36};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_35 = {decodeResult_andMatrixOutputs_hi_hi_31, decodeResult_andMatrixOutputs_andMatrixInput_2_35};
  wire        decodeResult_andMatrixOutputs_7_2 = &{decodeResult_andMatrixOutputs_hi_35, decodeResult_andMatrixOutputs_lo_33};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_26 = {decodeResult_andMatrixOutputs_andMatrixInput_4_32, decodeResult_andMatrixOutputs_andMatrixInput_5_26};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_34 = {decodeResult_andMatrixOutputs_lo_hi_26, decodeResult_andMatrixOutputs_andMatrixInput_6_11};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_11 = {decodeResult_andMatrixOutputs_andMatrixInput_2_36, decodeResult_andMatrixOutputs_andMatrixInput_3_34};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_32 = {decodeResult_andMatrixOutputs_andMatrixInput_0_38, decodeResult_andMatrixOutputs_andMatrixInput_1_37};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_36 = {decodeResult_andMatrixOutputs_hi_hi_32, decodeResult_andMatrixOutputs_hi_lo_11};
  wire        decodeResult_andMatrixOutputs_75_2 = &{decodeResult_andMatrixOutputs_hi_36, decodeResult_andMatrixOutputs_lo_34};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_27 = {decodeResult_andMatrixOutputs_andMatrixInput_4_33, decodeResult_andMatrixOutputs_andMatrixInput_5_27};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_35 = {decodeResult_andMatrixOutputs_lo_hi_27, decodeResult_andMatrixOutputs_andMatrixInput_6_12};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_12 = {decodeResult_andMatrixOutputs_andMatrixInput_2_37, decodeResult_andMatrixOutputs_andMatrixInput_3_35};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_33 = {decodeResult_andMatrixOutputs_andMatrixInput_0_39, decodeResult_andMatrixOutputs_andMatrixInput_1_38};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_37 = {decodeResult_andMatrixOutputs_hi_hi_33, decodeResult_andMatrixOutputs_hi_lo_12};
  wire        decodeResult_andMatrixOutputs_68_2 = &{decodeResult_andMatrixOutputs_hi_37, decodeResult_andMatrixOutputs_lo_35};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_28 = {decodeResult_andMatrixOutputs_andMatrixInput_3_36, decodeResult_andMatrixOutputs_andMatrixInput_4_34};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_36 = {decodeResult_andMatrixOutputs_lo_hi_28, decodeResult_andMatrixOutputs_andMatrixInput_5_28};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_34 = {decodeResult_andMatrixOutputs_andMatrixInput_0_40, decodeResult_andMatrixOutputs_andMatrixInput_1_39};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_38 = {decodeResult_andMatrixOutputs_hi_hi_34, decodeResult_andMatrixOutputs_andMatrixInput_2_38};
  wire        decodeResult_andMatrixOutputs_48_2 = &{decodeResult_andMatrixOutputs_hi_38, decodeResult_andMatrixOutputs_lo_36};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_29 = {decodeResult_andMatrixOutputs_andMatrixInput_4_35, decodeResult_andMatrixOutputs_andMatrixInput_5_29};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_37 = {decodeResult_andMatrixOutputs_lo_hi_29, decodeResult_andMatrixOutputs_andMatrixInput_6_13};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_13 = {decodeResult_andMatrixOutputs_andMatrixInput_2_39, decodeResult_andMatrixOutputs_andMatrixInput_3_37};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_35 = {decodeResult_andMatrixOutputs_andMatrixInput_0_41, decodeResult_andMatrixOutputs_andMatrixInput_1_40};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_39 = {decodeResult_andMatrixOutputs_hi_hi_35, decodeResult_andMatrixOutputs_hi_lo_13};
  wire        decodeResult_andMatrixOutputs_73_2 = &{decodeResult_andMatrixOutputs_hi_39, decodeResult_andMatrixOutputs_lo_37};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_30 = {decodeResult_andMatrixOutputs_andMatrixInput_4_36, decodeResult_andMatrixOutputs_andMatrixInput_5_30};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_38 = {decodeResult_andMatrixOutputs_lo_hi_30, decodeResult_andMatrixOutputs_andMatrixInput_6_14};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_14 = {decodeResult_andMatrixOutputs_andMatrixInput_2_40, decodeResult_andMatrixOutputs_andMatrixInput_3_38};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_36 = {decodeResult_andMatrixOutputs_andMatrixInput_0_42, decodeResult_andMatrixOutputs_andMatrixInput_1_41};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_40 = {decodeResult_andMatrixOutputs_hi_hi_36, decodeResult_andMatrixOutputs_hi_lo_14};
  wire        decodeResult_andMatrixOutputs_130_2 = &{decodeResult_andMatrixOutputs_hi_40, decodeResult_andMatrixOutputs_lo_38};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_39 = {decodeResult_andMatrixOutputs_andMatrixInput_3_39, decodeResult_andMatrixOutputs_andMatrixInput_4_37};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_37 = {decodeResult_andMatrixOutputs_andMatrixInput_0_43, decodeResult_andMatrixOutputs_andMatrixInput_1_42};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_41 = {decodeResult_andMatrixOutputs_hi_hi_37, decodeResult_andMatrixOutputs_andMatrixInput_2_41};
  wire        decodeResult_andMatrixOutputs_120_2 = &{decodeResult_andMatrixOutputs_hi_41, decodeResult_andMatrixOutputs_lo_39};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo_5 = {decodeResult_andMatrixOutputs_andMatrixInput_6_15, decodeResult_andMatrixOutputs_andMatrixInput_7_5};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_31 = {decodeResult_andMatrixOutputs_andMatrixInput_4_38, decodeResult_andMatrixOutputs_andMatrixInput_5_31};
  wire [3:0]  decodeResult_andMatrixOutputs_lo_40 = {decodeResult_andMatrixOutputs_lo_hi_31, decodeResult_andMatrixOutputs_lo_lo_5};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_15 = {decodeResult_andMatrixOutputs_andMatrixInput_2_42, decodeResult_andMatrixOutputs_andMatrixInput_3_40};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_38 = {decodeResult_andMatrixOutputs_andMatrixInput_0_44, decodeResult_andMatrixOutputs_andMatrixInput_1_43};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_42 = {decodeResult_andMatrixOutputs_hi_hi_38, decodeResult_andMatrixOutputs_hi_lo_15};
  wire        decodeResult_andMatrixOutputs_136_2 = &{decodeResult_andMatrixOutputs_hi_42, decodeResult_andMatrixOutputs_lo_40};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_32 = {decodeResult_andMatrixOutputs_andMatrixInput_3_41, decodeResult_andMatrixOutputs_andMatrixInput_4_39};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_41 = {decodeResult_andMatrixOutputs_lo_hi_32, decodeResult_andMatrixOutputs_andMatrixInput_5_32};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_39 = {decodeResult_andMatrixOutputs_andMatrixInput_0_45, decodeResult_andMatrixOutputs_andMatrixInput_1_44};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_43 = {decodeResult_andMatrixOutputs_hi_hi_39, decodeResult_andMatrixOutputs_andMatrixInput_2_43};
  wire        decodeResult_andMatrixOutputs_34_2 = &{decodeResult_andMatrixOutputs_hi_43, decodeResult_andMatrixOutputs_lo_41};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo_6 = {decodeResult_andMatrixOutputs_andMatrixInput_6_16, decodeResult_andMatrixOutputs_andMatrixInput_7_6};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_33 = {decodeResult_andMatrixOutputs_andMatrixInput_4_40, decodeResult_andMatrixOutputs_andMatrixInput_5_33};
  wire [3:0]  decodeResult_andMatrixOutputs_lo_42 = {decodeResult_andMatrixOutputs_lo_hi_33, decodeResult_andMatrixOutputs_lo_lo_6};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_16 = {decodeResult_andMatrixOutputs_andMatrixInput_2_44, decodeResult_andMatrixOutputs_andMatrixInput_3_42};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_40 = {decodeResult_andMatrixOutputs_andMatrixInput_0_46, decodeResult_andMatrixOutputs_andMatrixInput_1_45};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_44 = {decodeResult_andMatrixOutputs_hi_hi_40, decodeResult_andMatrixOutputs_hi_lo_16};
  wire        decodeResult_andMatrixOutputs_57_2 = &{decodeResult_andMatrixOutputs_hi_44, decodeResult_andMatrixOutputs_lo_42};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_43 = {decodeResult_andMatrixOutputs_andMatrixInput_3_43, decodeResult_andMatrixOutputs_andMatrixInput_4_41};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_41 = {decodeResult_andMatrixOutputs_andMatrixInput_0_47, decodeResult_andMatrixOutputs_andMatrixInput_1_46};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_45 = {decodeResult_andMatrixOutputs_hi_hi_41, decodeResult_andMatrixOutputs_andMatrixInput_2_45};
  wire        decodeResult_andMatrixOutputs_66_2 = &{decodeResult_andMatrixOutputs_hi_45, decodeResult_andMatrixOutputs_lo_43};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_44 = {decodeResult_andMatrixOutputs_andMatrixInput_3_44, decodeResult_andMatrixOutputs_andMatrixInput_4_42};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_42 = {decodeResult_andMatrixOutputs_andMatrixInput_0_48, decodeResult_andMatrixOutputs_andMatrixInput_1_47};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_46 = {decodeResult_andMatrixOutputs_hi_hi_42, decodeResult_andMatrixOutputs_andMatrixInput_2_46};
  wire        decodeResult_andMatrixOutputs_9_2 = &{decodeResult_andMatrixOutputs_hi_46, decodeResult_andMatrixOutputs_lo_44};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_34 = {decodeResult_andMatrixOutputs_andMatrixInput_3_45, decodeResult_andMatrixOutputs_andMatrixInput_4_43};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_45 = {decodeResult_andMatrixOutputs_lo_hi_34, decodeResult_andMatrixOutputs_andMatrixInput_5_34};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_43 = {decodeResult_andMatrixOutputs_andMatrixInput_0_49, decodeResult_andMatrixOutputs_andMatrixInput_1_48};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_47 = {decodeResult_andMatrixOutputs_hi_hi_43, decodeResult_andMatrixOutputs_andMatrixInput_2_47};
  wire        decodeResult_andMatrixOutputs_18_2 = &{decodeResult_andMatrixOutputs_hi_47, decodeResult_andMatrixOutputs_lo_45};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_35 = {decodeResult_andMatrixOutputs_andMatrixInput_3_46, decodeResult_andMatrixOutputs_andMatrixInput_4_44};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_46 = {decodeResult_andMatrixOutputs_lo_hi_35, decodeResult_andMatrixOutputs_andMatrixInput_5_35};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_44 = {decodeResult_andMatrixOutputs_andMatrixInput_0_50, decodeResult_andMatrixOutputs_andMatrixInput_1_49};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_48 = {decodeResult_andMatrixOutputs_hi_hi_44, decodeResult_andMatrixOutputs_andMatrixInput_2_48};
  wire        decodeResult_andMatrixOutputs_4_2 = &{decodeResult_andMatrixOutputs_hi_48, decodeResult_andMatrixOutputs_lo_46};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_36 = {decodeResult_andMatrixOutputs_andMatrixInput_3_47, decodeResult_andMatrixOutputs_andMatrixInput_4_45};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_47 = {decodeResult_andMatrixOutputs_lo_hi_36, decodeResult_andMatrixOutputs_andMatrixInput_5_36};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_45 = {decodeResult_andMatrixOutputs_andMatrixInput_0_51, decodeResult_andMatrixOutputs_andMatrixInput_1_50};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_49 = {decodeResult_andMatrixOutputs_hi_hi_45, decodeResult_andMatrixOutputs_andMatrixInput_2_49};
  wire        decodeResult_andMatrixOutputs_146_2 = &{decodeResult_andMatrixOutputs_hi_49, decodeResult_andMatrixOutputs_lo_47};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_37 = {decodeResult_andMatrixOutputs_andMatrixInput_3_48, decodeResult_andMatrixOutputs_andMatrixInput_4_46};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_48 = {decodeResult_andMatrixOutputs_lo_hi_37, decodeResult_andMatrixOutputs_andMatrixInput_5_37};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_46 = {decodeResult_andMatrixOutputs_andMatrixInput_0_52, decodeResult_andMatrixOutputs_andMatrixInput_1_51};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_50 = {decodeResult_andMatrixOutputs_hi_hi_46, decodeResult_andMatrixOutputs_andMatrixInput_2_50};
  wire        decodeResult_andMatrixOutputs_55_2 = &{decodeResult_andMatrixOutputs_hi_50, decodeResult_andMatrixOutputs_lo_48};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_38 = {decodeResult_andMatrixOutputs_andMatrixInput_4_47, decodeResult_andMatrixOutputs_andMatrixInput_5_38};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_49 = {decodeResult_andMatrixOutputs_lo_hi_38, decodeResult_andMatrixOutputs_andMatrixInput_6_17};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_17 = {decodeResult_andMatrixOutputs_andMatrixInput_2_51, decodeResult_andMatrixOutputs_andMatrixInput_3_49};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_47 = {decodeResult_andMatrixOutputs_andMatrixInput_0_53, decodeResult_andMatrixOutputs_andMatrixInput_1_52};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_51 = {decodeResult_andMatrixOutputs_hi_hi_47, decodeResult_andMatrixOutputs_hi_lo_17};
  wire        decodeResult_andMatrixOutputs_137_2 = &{decodeResult_andMatrixOutputs_hi_51, decodeResult_andMatrixOutputs_lo_49};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_39 = {decodeResult_andMatrixOutputs_andMatrixInput_3_50, decodeResult_andMatrixOutputs_andMatrixInput_4_48};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_50 = {decodeResult_andMatrixOutputs_lo_hi_39, decodeResult_andMatrixOutputs_andMatrixInput_5_39};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_48 = {decodeResult_andMatrixOutputs_andMatrixInput_0_54, decodeResult_andMatrixOutputs_andMatrixInput_1_53};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_52 = {decodeResult_andMatrixOutputs_hi_hi_48, decodeResult_andMatrixOutputs_andMatrixInput_2_52};
  wire        decodeResult_andMatrixOutputs_108_2 = &{decodeResult_andMatrixOutputs_hi_52, decodeResult_andMatrixOutputs_lo_50};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_40 = {decodeResult_andMatrixOutputs_andMatrixInput_3_51, decodeResult_andMatrixOutputs_andMatrixInput_4_49};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_51 = {decodeResult_andMatrixOutputs_lo_hi_40, decodeResult_andMatrixOutputs_andMatrixInput_5_40};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_49 = {decodeResult_andMatrixOutputs_andMatrixInput_0_55, decodeResult_andMatrixOutputs_andMatrixInput_1_54};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_53 = {decodeResult_andMatrixOutputs_hi_hi_49, decodeResult_andMatrixOutputs_andMatrixInput_2_53};
  wire        decodeResult_andMatrixOutputs_69_2 = &{decodeResult_andMatrixOutputs_hi_53, decodeResult_andMatrixOutputs_lo_51};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_41 = {decodeResult_andMatrixOutputs_andMatrixInput_4_50, decodeResult_andMatrixOutputs_andMatrixInput_5_41};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_52 = {decodeResult_andMatrixOutputs_lo_hi_41, decodeResult_andMatrixOutputs_andMatrixInput_6_18};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_18 = {decodeResult_andMatrixOutputs_andMatrixInput_2_54, decodeResult_andMatrixOutputs_andMatrixInput_3_52};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_50 = {decodeResult_andMatrixOutputs_andMatrixInput_0_56, decodeResult_andMatrixOutputs_andMatrixInput_1_55};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_54 = {decodeResult_andMatrixOutputs_hi_hi_50, decodeResult_andMatrixOutputs_hi_lo_18};
  wire        decodeResult_andMatrixOutputs_117_2 = &{decodeResult_andMatrixOutputs_hi_54, decodeResult_andMatrixOutputs_lo_52};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_42 = {decodeResult_andMatrixOutputs_andMatrixInput_3_53, decodeResult_andMatrixOutputs_andMatrixInput_4_51};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_53 = {decodeResult_andMatrixOutputs_lo_hi_42, decodeResult_andMatrixOutputs_andMatrixInput_5_42};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_51 = {decodeResult_andMatrixOutputs_andMatrixInput_0_57, decodeResult_andMatrixOutputs_andMatrixInput_1_56};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_55 = {decodeResult_andMatrixOutputs_hi_hi_51, decodeResult_andMatrixOutputs_andMatrixInput_2_55};
  wire        decodeResult_andMatrixOutputs_106_2 = &{decodeResult_andMatrixOutputs_hi_55, decodeResult_andMatrixOutputs_lo_53};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_43 = {decodeResult_andMatrixOutputs_andMatrixInput_3_54, decodeResult_andMatrixOutputs_andMatrixInput_4_52};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_54 = {decodeResult_andMatrixOutputs_lo_hi_43, decodeResult_andMatrixOutputs_andMatrixInput_5_43};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_52 = {decodeResult_andMatrixOutputs_andMatrixInput_0_58, decodeResult_andMatrixOutputs_andMatrixInput_1_57};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_56 = {decodeResult_andMatrixOutputs_hi_hi_52, decodeResult_andMatrixOutputs_andMatrixInput_2_56};
  wire        decodeResult_andMatrixOutputs_141_2 = &{decodeResult_andMatrixOutputs_hi_56, decodeResult_andMatrixOutputs_lo_54};
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_44 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_58 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_45 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_46 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_47 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7_7 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_8_2 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_50 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_51 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_8_3 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_8_4 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7_11 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_28 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7_13 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_57 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_58 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7_14 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_33 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_34 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_35 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_7_17 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_37 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_38 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_8_9 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_40 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_41 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_8_10 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_79 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_80 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_70 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_82 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_83 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_84 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_85 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_72 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_87 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_73 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_89 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_90 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_75 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_92 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_76 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_94 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_78 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_96 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_80 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_81 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_82 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_48 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_84 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_85 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_137 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_138 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_139 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_110 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_144 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_142 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_143 = decodeResult_plaInput[30];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_111 = decodeResult_plaInput[30];
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_44 = {decodeResult_andMatrixOutputs_andMatrixInput_4_53, decodeResult_andMatrixOutputs_andMatrixInput_5_44};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_55 = {decodeResult_andMatrixOutputs_lo_hi_44, decodeResult_andMatrixOutputs_andMatrixInput_6_19};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_19 = {decodeResult_andMatrixOutputs_andMatrixInput_2_57, decodeResult_andMatrixOutputs_andMatrixInput_3_55};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_53 = {decodeResult_andMatrixOutputs_andMatrixInput_0_59, decodeResult_andMatrixOutputs_andMatrixInput_1_58};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_57 = {decodeResult_andMatrixOutputs_hi_hi_53, decodeResult_andMatrixOutputs_hi_lo_19};
  wire        decodeResult_andMatrixOutputs_148_2 = &{decodeResult_andMatrixOutputs_hi_57, decodeResult_andMatrixOutputs_lo_55};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_58 = {decodeResult_andMatrixOutputs_andMatrixInput_0_60, decodeResult_andMatrixOutputs_andMatrixInput_1_59};
  wire        decodeResult_andMatrixOutputs_90_2 = &{decodeResult_andMatrixOutputs_hi_58, decodeResult_andMatrixOutputs_andMatrixInput_2_58};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_45 = {decodeResult_andMatrixOutputs_andMatrixInput_4_54, decodeResult_andMatrixOutputs_andMatrixInput_5_45};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_56 = {decodeResult_andMatrixOutputs_lo_hi_45, decodeResult_andMatrixOutputs_andMatrixInput_6_20};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_20 = {decodeResult_andMatrixOutputs_andMatrixInput_2_59, decodeResult_andMatrixOutputs_andMatrixInput_3_56};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_54 = {decodeResult_andMatrixOutputs_andMatrixInput_0_61, decodeResult_andMatrixOutputs_andMatrixInput_1_60};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_59 = {decodeResult_andMatrixOutputs_hi_hi_54, decodeResult_andMatrixOutputs_hi_lo_20};
  wire        decodeResult_andMatrixOutputs_20_2 = &{decodeResult_andMatrixOutputs_hi_59, decodeResult_andMatrixOutputs_lo_56};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_46 = {decodeResult_andMatrixOutputs_andMatrixInput_4_55, decodeResult_andMatrixOutputs_andMatrixInput_5_46};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_57 = {decodeResult_andMatrixOutputs_lo_hi_46, decodeResult_andMatrixOutputs_andMatrixInput_6_21};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_21 = {decodeResult_andMatrixOutputs_andMatrixInput_2_60, decodeResult_andMatrixOutputs_andMatrixInput_3_57};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_55 = {decodeResult_andMatrixOutputs_andMatrixInput_0_62, decodeResult_andMatrixOutputs_andMatrixInput_1_61};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_60 = {decodeResult_andMatrixOutputs_hi_hi_55, decodeResult_andMatrixOutputs_hi_lo_21};
  wire        decodeResult_andMatrixOutputs_133_2 = &{decodeResult_andMatrixOutputs_hi_60, decodeResult_andMatrixOutputs_lo_57};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_47 = {decodeResult_andMatrixOutputs_andMatrixInput_4_56, decodeResult_andMatrixOutputs_andMatrixInput_5_47};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_58 = {decodeResult_andMatrixOutputs_lo_hi_47, decodeResult_andMatrixOutputs_andMatrixInput_6_22};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_22 = {decodeResult_andMatrixOutputs_andMatrixInput_2_61, decodeResult_andMatrixOutputs_andMatrixInput_3_58};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_56 = {decodeResult_andMatrixOutputs_andMatrixInput_0_63, decodeResult_andMatrixOutputs_andMatrixInput_1_62};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_61 = {decodeResult_andMatrixOutputs_hi_hi_56, decodeResult_andMatrixOutputs_hi_lo_22};
  wire        decodeResult_andMatrixOutputs_21_2 = &{decodeResult_andMatrixOutputs_hi_61, decodeResult_andMatrixOutputs_lo_58};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo_7 = {decodeResult_andMatrixOutputs_andMatrixInput_7_7, decodeResult_andMatrixOutputs_andMatrixInput_8_1};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_48 = {decodeResult_andMatrixOutputs_andMatrixInput_5_48, decodeResult_andMatrixOutputs_andMatrixInput_6_23};
  wire [3:0]  decodeResult_andMatrixOutputs_lo_59 = {decodeResult_andMatrixOutputs_lo_hi_48, decodeResult_andMatrixOutputs_lo_lo_7};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_23 = {decodeResult_andMatrixOutputs_andMatrixInput_3_59, decodeResult_andMatrixOutputs_andMatrixInput_4_57};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_hi_1 = {decodeResult_andMatrixOutputs_andMatrixInput_0_64, decodeResult_andMatrixOutputs_andMatrixInput_1_63};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_hi_57 = {decodeResult_andMatrixOutputs_hi_hi_hi_1, decodeResult_andMatrixOutputs_andMatrixInput_2_62};
  wire [4:0]  decodeResult_andMatrixOutputs_hi_62 = {decodeResult_andMatrixOutputs_hi_hi_57, decodeResult_andMatrixOutputs_hi_lo_23};
  wire        decodeResult_andMatrixOutputs_121_2 = &{decodeResult_andMatrixOutputs_hi_62, decodeResult_andMatrixOutputs_lo_59};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo_8 = {decodeResult_andMatrixOutputs_andMatrixInput_8_2, decodeResult_andMatrixOutputs_andMatrixInput_9};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_hi = {decodeResult_andMatrixOutputs_andMatrixInput_5_49, decodeResult_andMatrixOutputs_andMatrixInput_6_24};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_hi_49 = {decodeResult_andMatrixOutputs_lo_hi_hi, decodeResult_andMatrixOutputs_andMatrixInput_7_8};
  wire [4:0]  decodeResult_andMatrixOutputs_lo_60 = {decodeResult_andMatrixOutputs_lo_hi_49, decodeResult_andMatrixOutputs_lo_lo_8};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_24 = {decodeResult_andMatrixOutputs_andMatrixInput_3_60, decodeResult_andMatrixOutputs_andMatrixInput_4_58};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_hi_2 = {decodeResult_andMatrixOutputs_andMatrixInput_0_65, decodeResult_andMatrixOutputs_andMatrixInput_1_64};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_hi_58 = {decodeResult_andMatrixOutputs_hi_hi_hi_2, decodeResult_andMatrixOutputs_andMatrixInput_2_63};
  wire [4:0]  decodeResult_andMatrixOutputs_hi_63 = {decodeResult_andMatrixOutputs_hi_hi_58, decodeResult_andMatrixOutputs_hi_lo_24};
  wire        decodeResult_andMatrixOutputs_63_2 = &{decodeResult_andMatrixOutputs_hi_63, decodeResult_andMatrixOutputs_lo_60};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_50 = {decodeResult_andMatrixOutputs_andMatrixInput_3_61, decodeResult_andMatrixOutputs_andMatrixInput_4_59};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_61 = {decodeResult_andMatrixOutputs_lo_hi_50, decodeResult_andMatrixOutputs_andMatrixInput_5_50};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_59 = {decodeResult_andMatrixOutputs_andMatrixInput_0_66, decodeResult_andMatrixOutputs_andMatrixInput_1_65};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_64 = {decodeResult_andMatrixOutputs_hi_hi_59, decodeResult_andMatrixOutputs_andMatrixInput_2_64};
  wire        decodeResult_andMatrixOutputs_11_2 = &{decodeResult_andMatrixOutputs_hi_64, decodeResult_andMatrixOutputs_lo_61};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_51 = {decodeResult_andMatrixOutputs_andMatrixInput_3_62, decodeResult_andMatrixOutputs_andMatrixInput_4_60};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_62 = {decodeResult_andMatrixOutputs_lo_hi_51, decodeResult_andMatrixOutputs_andMatrixInput_5_51};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_60 = {decodeResult_andMatrixOutputs_andMatrixInput_0_67, decodeResult_andMatrixOutputs_andMatrixInput_1_66};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_65 = {decodeResult_andMatrixOutputs_hi_hi_60, decodeResult_andMatrixOutputs_andMatrixInput_2_65};
  wire        decodeResult_andMatrixOutputs_94_2 = &{decodeResult_andMatrixOutputs_hi_65, decodeResult_andMatrixOutputs_lo_62};
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_52 = decodeResult_invInputs[17];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_70 = decodeResult_invInputs[17];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_79 = decodeResult_invInputs[17];
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo_9 = {decodeResult_andMatrixOutputs_andMatrixInput_8_3, decodeResult_andMatrixOutputs_andMatrixInput_9_1};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_hi_1 = {decodeResult_andMatrixOutputs_andMatrixInput_5_52, decodeResult_andMatrixOutputs_andMatrixInput_6_25};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_hi_52 = {decodeResult_andMatrixOutputs_lo_hi_hi_1, decodeResult_andMatrixOutputs_andMatrixInput_7_9};
  wire [4:0]  decodeResult_andMatrixOutputs_lo_63 = {decodeResult_andMatrixOutputs_lo_hi_52, decodeResult_andMatrixOutputs_lo_lo_9};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_25 = {decodeResult_andMatrixOutputs_andMatrixInput_3_63, decodeResult_andMatrixOutputs_andMatrixInput_4_61};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_hi_3 = {decodeResult_andMatrixOutputs_andMatrixInput_0_68, decodeResult_andMatrixOutputs_andMatrixInput_1_67};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_hi_61 = {decodeResult_andMatrixOutputs_hi_hi_hi_3, decodeResult_andMatrixOutputs_andMatrixInput_2_66};
  wire [4:0]  decodeResult_andMatrixOutputs_hi_66 = {decodeResult_andMatrixOutputs_hi_hi_61, decodeResult_andMatrixOutputs_hi_lo_25};
  wire        decodeResult_andMatrixOutputs_144_2 = &{decodeResult_andMatrixOutputs_hi_66, decodeResult_andMatrixOutputs_lo_63};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo_10 = {decodeResult_andMatrixOutputs_andMatrixInput_8_4, decodeResult_andMatrixOutputs_andMatrixInput_9_2};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_hi_2 = {decodeResult_andMatrixOutputs_andMatrixInput_5_53, decodeResult_andMatrixOutputs_andMatrixInput_6_26};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_hi_53 = {decodeResult_andMatrixOutputs_lo_hi_hi_2, decodeResult_andMatrixOutputs_andMatrixInput_7_10};
  wire [4:0]  decodeResult_andMatrixOutputs_lo_64 = {decodeResult_andMatrixOutputs_lo_hi_53, decodeResult_andMatrixOutputs_lo_lo_10};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_26 = {decodeResult_andMatrixOutputs_andMatrixInput_3_64, decodeResult_andMatrixOutputs_andMatrixInput_4_62};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_hi_4 = {decodeResult_andMatrixOutputs_andMatrixInput_0_69, decodeResult_andMatrixOutputs_andMatrixInput_1_68};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_hi_62 = {decodeResult_andMatrixOutputs_hi_hi_hi_4, decodeResult_andMatrixOutputs_andMatrixInput_2_67};
  wire [4:0]  decodeResult_andMatrixOutputs_hi_67 = {decodeResult_andMatrixOutputs_hi_hi_62, decodeResult_andMatrixOutputs_hi_lo_26};
  wire        decodeResult_andMatrixOutputs_77_2 = &{decodeResult_andMatrixOutputs_hi_67, decodeResult_andMatrixOutputs_lo_64};
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_65 = decodeResult_plaInput[17];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_72 = decodeResult_plaInput[17];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_80 = decodeResult_plaInput[17];
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo_11 = {decodeResult_andMatrixOutputs_andMatrixInput_7_11, decodeResult_andMatrixOutputs_andMatrixInput_8_5};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_54 = {decodeResult_andMatrixOutputs_andMatrixInput_5_54, decodeResult_andMatrixOutputs_andMatrixInput_6_27};
  wire [3:0]  decodeResult_andMatrixOutputs_lo_65 = {decodeResult_andMatrixOutputs_lo_hi_54, decodeResult_andMatrixOutputs_lo_lo_11};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_27 = {decodeResult_andMatrixOutputs_andMatrixInput_3_65, decodeResult_andMatrixOutputs_andMatrixInput_4_63};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_hi_5 = {decodeResult_andMatrixOutputs_andMatrixInput_0_70, decodeResult_andMatrixOutputs_andMatrixInput_1_69};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_hi_63 = {decodeResult_andMatrixOutputs_hi_hi_hi_5, decodeResult_andMatrixOutputs_andMatrixInput_2_68};
  wire [4:0]  decodeResult_andMatrixOutputs_hi_68 = {decodeResult_andMatrixOutputs_hi_hi_63, decodeResult_andMatrixOutputs_hi_lo_27};
  wire        decodeResult_andMatrixOutputs_54_2 = &{decodeResult_andMatrixOutputs_hi_68, decodeResult_andMatrixOutputs_lo_65};
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_66 = decodeResult_plaInput[19];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_65 = decodeResult_plaInput[19];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_73 = decodeResult_plaInput[19];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_1_92 = decodeResult_plaInput[19];
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo_12 = {decodeResult_andMatrixOutputs_andMatrixInput_6_28, decodeResult_andMatrixOutputs_andMatrixInput_7_12};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_55 = {decodeResult_andMatrixOutputs_andMatrixInput_4_64, decodeResult_andMatrixOutputs_andMatrixInput_5_55};
  wire [3:0]  decodeResult_andMatrixOutputs_lo_66 = {decodeResult_andMatrixOutputs_lo_hi_55, decodeResult_andMatrixOutputs_lo_lo_12};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_28 = {decodeResult_andMatrixOutputs_andMatrixInput_2_69, decodeResult_andMatrixOutputs_andMatrixInput_3_66};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_64 = {decodeResult_andMatrixOutputs_andMatrixInput_0_71, decodeResult_andMatrixOutputs_andMatrixInput_1_70};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_69 = {decodeResult_andMatrixOutputs_hi_hi_64, decodeResult_andMatrixOutputs_hi_lo_28};
  wire        decodeResult_andMatrixOutputs_140_2 = &{decodeResult_andMatrixOutputs_hi_69, decodeResult_andMatrixOutputs_lo_66};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo_13 = {decodeResult_andMatrixOutputs_andMatrixInput_7_13, decodeResult_andMatrixOutputs_andMatrixInput_8_6};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_56 = {decodeResult_andMatrixOutputs_andMatrixInput_5_56, decodeResult_andMatrixOutputs_andMatrixInput_6_29};
  wire [3:0]  decodeResult_andMatrixOutputs_lo_67 = {decodeResult_andMatrixOutputs_lo_hi_56, decodeResult_andMatrixOutputs_lo_lo_13};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_29 = {decodeResult_andMatrixOutputs_andMatrixInput_3_67, decodeResult_andMatrixOutputs_andMatrixInput_4_65};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_hi_6 = {decodeResult_andMatrixOutputs_andMatrixInput_0_72, decodeResult_andMatrixOutputs_andMatrixInput_1_71};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_hi_65 = {decodeResult_andMatrixOutputs_hi_hi_hi_6, decodeResult_andMatrixOutputs_andMatrixInput_2_70};
  wire [4:0]  decodeResult_andMatrixOutputs_hi_70 = {decodeResult_andMatrixOutputs_hi_hi_65, decodeResult_andMatrixOutputs_hi_lo_29};
  wire        decodeResult_andMatrixOutputs_33_2 = &{decodeResult_andMatrixOutputs_hi_70, decodeResult_andMatrixOutputs_lo_67};
  wire        decodeResult_andMatrixOutputs_andMatrixInput_2_71 = decodeResult_plaInput[25];
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_57 = {decodeResult_andMatrixOutputs_andMatrixInput_4_66, decodeResult_andMatrixOutputs_andMatrixInput_5_57};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_68 = {decodeResult_andMatrixOutputs_lo_hi_57, decodeResult_andMatrixOutputs_andMatrixInput_6_30};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_30 = {decodeResult_andMatrixOutputs_andMatrixInput_2_71, decodeResult_andMatrixOutputs_andMatrixInput_3_68};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_66 = {decodeResult_andMatrixOutputs_andMatrixInput_0_73, decodeResult_andMatrixOutputs_andMatrixInput_1_72};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_71 = {decodeResult_andMatrixOutputs_hi_hi_66, decodeResult_andMatrixOutputs_hi_lo_30};
  wire        decodeResult_andMatrixOutputs_67_2 = &{decodeResult_andMatrixOutputs_hi_71, decodeResult_andMatrixOutputs_lo_68};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_58 = {decodeResult_andMatrixOutputs_andMatrixInput_4_67, decodeResult_andMatrixOutputs_andMatrixInput_5_58};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_69 = {decodeResult_andMatrixOutputs_lo_hi_58, decodeResult_andMatrixOutputs_andMatrixInput_6_31};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_31 = {decodeResult_andMatrixOutputs_andMatrixInput_2_72, decodeResult_andMatrixOutputs_andMatrixInput_3_69};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_67 = {decodeResult_andMatrixOutputs_andMatrixInput_0_74, decodeResult_andMatrixOutputs_andMatrixInput_1_73};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_72 = {decodeResult_andMatrixOutputs_hi_hi_67, decodeResult_andMatrixOutputs_hi_lo_31};
  wire        decodeResult_andMatrixOutputs_14_2 = &{decodeResult_andMatrixOutputs_hi_72, decodeResult_andMatrixOutputs_lo_69};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo_14 = {decodeResult_andMatrixOutputs_andMatrixInput_7_14, decodeResult_andMatrixOutputs_andMatrixInput_8_7};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_59 = {decodeResult_andMatrixOutputs_andMatrixInput_5_59, decodeResult_andMatrixOutputs_andMatrixInput_6_32};
  wire [3:0]  decodeResult_andMatrixOutputs_lo_70 = {decodeResult_andMatrixOutputs_lo_hi_59, decodeResult_andMatrixOutputs_lo_lo_14};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_32 = {decodeResult_andMatrixOutputs_andMatrixInput_3_70, decodeResult_andMatrixOutputs_andMatrixInput_4_68};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_hi_7 = {decodeResult_andMatrixOutputs_andMatrixInput_0_75, decodeResult_andMatrixOutputs_andMatrixInput_1_74};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_hi_68 = {decodeResult_andMatrixOutputs_hi_hi_hi_7, decodeResult_andMatrixOutputs_andMatrixInput_2_73};
  wire [4:0]  decodeResult_andMatrixOutputs_hi_73 = {decodeResult_andMatrixOutputs_hi_hi_68, decodeResult_andMatrixOutputs_hi_lo_32};
  wire        decodeResult_andMatrixOutputs_13_2 = &{decodeResult_andMatrixOutputs_hi_73, decodeResult_andMatrixOutputs_lo_70};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_60 = {decodeResult_andMatrixOutputs_andMatrixInput_4_69, decodeResult_andMatrixOutputs_andMatrixInput_5_60};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_71 = {decodeResult_andMatrixOutputs_lo_hi_60, decodeResult_andMatrixOutputs_andMatrixInput_6_33};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_33 = {decodeResult_andMatrixOutputs_andMatrixInput_2_74, decodeResult_andMatrixOutputs_andMatrixInput_3_71};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_69 = {decodeResult_andMatrixOutputs_andMatrixInput_0_76, decodeResult_andMatrixOutputs_andMatrixInput_1_75};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_74 = {decodeResult_andMatrixOutputs_hi_hi_69, decodeResult_andMatrixOutputs_hi_lo_33};
  wire        decodeResult_andMatrixOutputs_98_2 = &{decodeResult_andMatrixOutputs_hi_74, decodeResult_andMatrixOutputs_lo_71};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo_15 = {decodeResult_andMatrixOutputs_andMatrixInput_6_34, decodeResult_andMatrixOutputs_andMatrixInput_7_15};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_61 = {decodeResult_andMatrixOutputs_andMatrixInput_4_70, decodeResult_andMatrixOutputs_andMatrixInput_5_61};
  wire [3:0]  decodeResult_andMatrixOutputs_lo_72 = {decodeResult_andMatrixOutputs_lo_hi_61, decodeResult_andMatrixOutputs_lo_lo_15};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_34 = {decodeResult_andMatrixOutputs_andMatrixInput_2_75, decodeResult_andMatrixOutputs_andMatrixInput_3_72};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_70 = {decodeResult_andMatrixOutputs_andMatrixInput_0_77, decodeResult_andMatrixOutputs_andMatrixInput_1_76};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_75 = {decodeResult_andMatrixOutputs_hi_hi_70, decodeResult_andMatrixOutputs_hi_lo_34};
  wire        decodeResult_andMatrixOutputs_46_2 = &{decodeResult_andMatrixOutputs_hi_75, decodeResult_andMatrixOutputs_lo_72};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo_16 = {decodeResult_andMatrixOutputs_andMatrixInput_6_35, decodeResult_andMatrixOutputs_andMatrixInput_7_16};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_62 = {decodeResult_andMatrixOutputs_andMatrixInput_4_71, decodeResult_andMatrixOutputs_andMatrixInput_5_62};
  wire [3:0]  decodeResult_andMatrixOutputs_lo_73 = {decodeResult_andMatrixOutputs_lo_hi_62, decodeResult_andMatrixOutputs_lo_lo_16};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_35 = {decodeResult_andMatrixOutputs_andMatrixInput_2_76, decodeResult_andMatrixOutputs_andMatrixInput_3_73};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_71 = {decodeResult_andMatrixOutputs_andMatrixInput_0_78, decodeResult_andMatrixOutputs_andMatrixInput_1_77};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_76 = {decodeResult_andMatrixOutputs_hi_hi_71, decodeResult_andMatrixOutputs_hi_lo_35};
  wire        decodeResult_andMatrixOutputs_101_2 = &{decodeResult_andMatrixOutputs_hi_76, decodeResult_andMatrixOutputs_lo_73};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo_17 = {decodeResult_andMatrixOutputs_andMatrixInput_7_17, decodeResult_andMatrixOutputs_andMatrixInput_8_8};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_63 = {decodeResult_andMatrixOutputs_andMatrixInput_5_63, decodeResult_andMatrixOutputs_andMatrixInput_6_36};
  wire [3:0]  decodeResult_andMatrixOutputs_lo_74 = {decodeResult_andMatrixOutputs_lo_hi_63, decodeResult_andMatrixOutputs_lo_lo_17};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_36 = {decodeResult_andMatrixOutputs_andMatrixInput_3_74, decodeResult_andMatrixOutputs_andMatrixInput_4_72};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_hi_8 = {decodeResult_andMatrixOutputs_andMatrixInput_0_79, decodeResult_andMatrixOutputs_andMatrixInput_1_78};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_hi_72 = {decodeResult_andMatrixOutputs_hi_hi_hi_8, decodeResult_andMatrixOutputs_andMatrixInput_2_77};
  wire [4:0]  decodeResult_andMatrixOutputs_hi_77 = {decodeResult_andMatrixOutputs_hi_hi_72, decodeResult_andMatrixOutputs_hi_lo_36};
  wire        decodeResult_andMatrixOutputs_142_2 = &{decodeResult_andMatrixOutputs_hi_77, decodeResult_andMatrixOutputs_lo_74};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo_18 = {decodeResult_andMatrixOutputs_andMatrixInput_6_37, decodeResult_andMatrixOutputs_andMatrixInput_7_18};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_64 = {decodeResult_andMatrixOutputs_andMatrixInput_4_73, decodeResult_andMatrixOutputs_andMatrixInput_5_64};
  wire [3:0]  decodeResult_andMatrixOutputs_lo_75 = {decodeResult_andMatrixOutputs_lo_hi_64, decodeResult_andMatrixOutputs_lo_lo_18};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_37 = {decodeResult_andMatrixOutputs_andMatrixInput_2_78, decodeResult_andMatrixOutputs_andMatrixInput_3_75};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_73 = {decodeResult_andMatrixOutputs_andMatrixInput_0_80, decodeResult_andMatrixOutputs_andMatrixInput_1_79};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_78 = {decodeResult_andMatrixOutputs_hi_hi_73, decodeResult_andMatrixOutputs_hi_lo_37};
  wire        decodeResult_andMatrixOutputs_19_2 = &{decodeResult_andMatrixOutputs_hi_78, decodeResult_andMatrixOutputs_lo_75};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo_19 = {decodeResult_andMatrixOutputs_andMatrixInput_6_38, decodeResult_andMatrixOutputs_andMatrixInput_7_19};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_65 = {decodeResult_andMatrixOutputs_andMatrixInput_4_74, decodeResult_andMatrixOutputs_andMatrixInput_5_65};
  wire [3:0]  decodeResult_andMatrixOutputs_lo_76 = {decodeResult_andMatrixOutputs_lo_hi_65, decodeResult_andMatrixOutputs_lo_lo_19};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_38 = {decodeResult_andMatrixOutputs_andMatrixInput_2_79, decodeResult_andMatrixOutputs_andMatrixInput_3_76};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_74 = {decodeResult_andMatrixOutputs_andMatrixInput_0_81, decodeResult_andMatrixOutputs_andMatrixInput_1_80};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_79 = {decodeResult_andMatrixOutputs_hi_hi_74, decodeResult_andMatrixOutputs_hi_lo_38};
  wire        decodeResult_andMatrixOutputs_17_2 = &{decodeResult_andMatrixOutputs_hi_79, decodeResult_andMatrixOutputs_lo_76};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo_20 = {decodeResult_andMatrixOutputs_andMatrixInput_8_9, decodeResult_andMatrixOutputs_andMatrixInput_9_3};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_hi_3 = {decodeResult_andMatrixOutputs_andMatrixInput_5_66, decodeResult_andMatrixOutputs_andMatrixInput_6_39};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_hi_66 = {decodeResult_andMatrixOutputs_lo_hi_hi_3, decodeResult_andMatrixOutputs_andMatrixInput_7_20};
  wire [4:0]  decodeResult_andMatrixOutputs_lo_77 = {decodeResult_andMatrixOutputs_lo_hi_66, decodeResult_andMatrixOutputs_lo_lo_20};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_39 = {decodeResult_andMatrixOutputs_andMatrixInput_3_77, decodeResult_andMatrixOutputs_andMatrixInput_4_75};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_hi_9 = {decodeResult_andMatrixOutputs_andMatrixInput_0_82, decodeResult_andMatrixOutputs_andMatrixInput_1_81};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_hi_75 = {decodeResult_andMatrixOutputs_hi_hi_hi_9, decodeResult_andMatrixOutputs_andMatrixInput_2_80};
  wire [4:0]  decodeResult_andMatrixOutputs_hi_80 = {decodeResult_andMatrixOutputs_hi_hi_75, decodeResult_andMatrixOutputs_hi_lo_39};
  wire        decodeResult_andMatrixOutputs_8_2 = &{decodeResult_andMatrixOutputs_hi_80, decodeResult_andMatrixOutputs_lo_77};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo_21 = {decodeResult_andMatrixOutputs_andMatrixInput_6_40, decodeResult_andMatrixOutputs_andMatrixInput_7_21};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_67 = {decodeResult_andMatrixOutputs_andMatrixInput_4_76, decodeResult_andMatrixOutputs_andMatrixInput_5_67};
  wire [3:0]  decodeResult_andMatrixOutputs_lo_78 = {decodeResult_andMatrixOutputs_lo_hi_67, decodeResult_andMatrixOutputs_lo_lo_21};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_40 = {decodeResult_andMatrixOutputs_andMatrixInput_2_81, decodeResult_andMatrixOutputs_andMatrixInput_3_78};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_76 = {decodeResult_andMatrixOutputs_andMatrixInput_0_83, decodeResult_andMatrixOutputs_andMatrixInput_1_82};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_81 = {decodeResult_andMatrixOutputs_hi_hi_76, decodeResult_andMatrixOutputs_hi_lo_40};
  wire        decodeResult_andMatrixOutputs_61_2 = &{decodeResult_andMatrixOutputs_hi_81, decodeResult_andMatrixOutputs_lo_78};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo_22 = {decodeResult_andMatrixOutputs_andMatrixInput_6_41, decodeResult_andMatrixOutputs_andMatrixInput_7_22};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_68 = {decodeResult_andMatrixOutputs_andMatrixInput_4_77, decodeResult_andMatrixOutputs_andMatrixInput_5_68};
  wire [3:0]  decodeResult_andMatrixOutputs_lo_79 = {decodeResult_andMatrixOutputs_lo_hi_68, decodeResult_andMatrixOutputs_lo_lo_22};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_41 = {decodeResult_andMatrixOutputs_andMatrixInput_2_82, decodeResult_andMatrixOutputs_andMatrixInput_3_79};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_77 = {decodeResult_andMatrixOutputs_andMatrixInput_0_84, decodeResult_andMatrixOutputs_andMatrixInput_1_83};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_82 = {decodeResult_andMatrixOutputs_hi_hi_77, decodeResult_andMatrixOutputs_hi_lo_41};
  wire        decodeResult_andMatrixOutputs_36_2 = &{decodeResult_andMatrixOutputs_hi_82, decodeResult_andMatrixOutputs_lo_79};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_lo_23 = {decodeResult_andMatrixOutputs_andMatrixInput_8_10, decodeResult_andMatrixOutputs_andMatrixInput_9_4};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_hi_4 = {decodeResult_andMatrixOutputs_andMatrixInput_5_69, decodeResult_andMatrixOutputs_andMatrixInput_6_42};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_hi_69 = {decodeResult_andMatrixOutputs_lo_hi_hi_4, decodeResult_andMatrixOutputs_andMatrixInput_7_23};
  wire [4:0]  decodeResult_andMatrixOutputs_lo_80 = {decodeResult_andMatrixOutputs_lo_hi_69, decodeResult_andMatrixOutputs_lo_lo_23};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_42 = {decodeResult_andMatrixOutputs_andMatrixInput_3_80, decodeResult_andMatrixOutputs_andMatrixInput_4_78};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_hi_10 = {decodeResult_andMatrixOutputs_andMatrixInput_0_85, decodeResult_andMatrixOutputs_andMatrixInput_1_84};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_hi_78 = {decodeResult_andMatrixOutputs_hi_hi_hi_10, decodeResult_andMatrixOutputs_andMatrixInput_2_83};
  wire [4:0]  decodeResult_andMatrixOutputs_hi_83 = {decodeResult_andMatrixOutputs_hi_hi_78, decodeResult_andMatrixOutputs_hi_lo_42};
  wire        decodeResult_andMatrixOutputs_86_2 = &{decodeResult_andMatrixOutputs_hi_83, decodeResult_andMatrixOutputs_lo_80};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_81 = {decodeResult_andMatrixOutputs_andMatrixInput_3_81, decodeResult_andMatrixOutputs_andMatrixInput_4_79};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_79 = {decodeResult_andMatrixOutputs_andMatrixInput_0_86, decodeResult_andMatrixOutputs_andMatrixInput_1_85};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_84 = {decodeResult_andMatrixOutputs_hi_hi_79, decodeResult_andMatrixOutputs_andMatrixInput_2_84};
  wire        decodeResult_andMatrixOutputs_145_2 = &{decodeResult_andMatrixOutputs_hi_84, decodeResult_andMatrixOutputs_lo_81};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_82 = {decodeResult_andMatrixOutputs_andMatrixInput_3_82, decodeResult_andMatrixOutputs_andMatrixInput_4_80};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_80 = {decodeResult_andMatrixOutputs_andMatrixInput_0_87, decodeResult_andMatrixOutputs_andMatrixInput_1_86};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_85 = {decodeResult_andMatrixOutputs_hi_hi_80, decodeResult_andMatrixOutputs_andMatrixInput_2_85};
  wire        decodeResult_andMatrixOutputs_2_2 = &{decodeResult_andMatrixOutputs_hi_85, decodeResult_andMatrixOutputs_lo_82};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_70 = {decodeResult_andMatrixOutputs_andMatrixInput_4_81, decodeResult_andMatrixOutputs_andMatrixInput_5_70};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_83 = {decodeResult_andMatrixOutputs_lo_hi_70, decodeResult_andMatrixOutputs_andMatrixInput_6_43};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_43 = {decodeResult_andMatrixOutputs_andMatrixInput_2_86, decodeResult_andMatrixOutputs_andMatrixInput_3_83};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_81 = {decodeResult_andMatrixOutputs_andMatrixInput_0_88, decodeResult_andMatrixOutputs_andMatrixInput_1_87};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_86 = {decodeResult_andMatrixOutputs_hi_hi_81, decodeResult_andMatrixOutputs_hi_lo_43};
  wire        decodeResult_andMatrixOutputs_113_2 = &{decodeResult_andMatrixOutputs_hi_86, decodeResult_andMatrixOutputs_lo_83};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_71 = {decodeResult_andMatrixOutputs_andMatrixInput_3_84, decodeResult_andMatrixOutputs_andMatrixInput_4_82};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_84 = {decodeResult_andMatrixOutputs_lo_hi_71, decodeResult_andMatrixOutputs_andMatrixInput_5_71};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_82 = {decodeResult_andMatrixOutputs_andMatrixInput_0_89, decodeResult_andMatrixOutputs_andMatrixInput_1_88};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_87 = {decodeResult_andMatrixOutputs_hi_hi_82, decodeResult_andMatrixOutputs_andMatrixInput_2_87};
  wire        decodeResult_andMatrixOutputs_147_2 = &{decodeResult_andMatrixOutputs_hi_87, decodeResult_andMatrixOutputs_lo_84};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_85 = {decodeResult_andMatrixOutputs_andMatrixInput_3_85, decodeResult_andMatrixOutputs_andMatrixInput_4_83};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_83 = {decodeResult_andMatrixOutputs_andMatrixInput_0_90, decodeResult_andMatrixOutputs_andMatrixInput_1_89};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_88 = {decodeResult_andMatrixOutputs_hi_hi_83, decodeResult_andMatrixOutputs_andMatrixInput_2_88};
  wire        decodeResult_andMatrixOutputs_59_2 = &{decodeResult_andMatrixOutputs_hi_88, decodeResult_andMatrixOutputs_lo_85};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_86 = {decodeResult_andMatrixOutputs_andMatrixInput_3_86, decodeResult_andMatrixOutputs_andMatrixInput_4_84};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_84 = {decodeResult_andMatrixOutputs_andMatrixInput_0_91, decodeResult_andMatrixOutputs_andMatrixInput_1_90};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_89 = {decodeResult_andMatrixOutputs_hi_hi_84, decodeResult_andMatrixOutputs_andMatrixInput_2_89};
  wire        decodeResult_andMatrixOutputs_60_2 = &{decodeResult_andMatrixOutputs_hi_89, decodeResult_andMatrixOutputs_lo_86};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_87 = {decodeResult_andMatrixOutputs_andMatrixInput_3_87, decodeResult_andMatrixOutputs_andMatrixInput_4_85};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_85 = {decodeResult_andMatrixOutputs_andMatrixInput_0_92, decodeResult_andMatrixOutputs_andMatrixInput_1_91};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_90 = {decodeResult_andMatrixOutputs_hi_hi_85, decodeResult_andMatrixOutputs_andMatrixInput_2_90};
  wire        decodeResult_andMatrixOutputs_39_2 = &{decodeResult_andMatrixOutputs_hi_90, decodeResult_andMatrixOutputs_lo_87};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_72 = {decodeResult_andMatrixOutputs_andMatrixInput_4_86, decodeResult_andMatrixOutputs_andMatrixInput_5_72};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_88 = {decodeResult_andMatrixOutputs_lo_hi_72, decodeResult_andMatrixOutputs_andMatrixInput_6_44};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_44 = {decodeResult_andMatrixOutputs_andMatrixInput_2_91, decodeResult_andMatrixOutputs_andMatrixInput_3_88};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_86 = {decodeResult_andMatrixOutputs_andMatrixInput_0_93, decodeResult_andMatrixOutputs_andMatrixInput_1_92};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_91 = {decodeResult_andMatrixOutputs_hi_hi_86, decodeResult_andMatrixOutputs_hi_lo_44};
  wire        decodeResult_andMatrixOutputs_80_2 = &{decodeResult_andMatrixOutputs_hi_91, decodeResult_andMatrixOutputs_lo_88};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_89 = {decodeResult_andMatrixOutputs_andMatrixInput_3_89, decodeResult_andMatrixOutputs_andMatrixInput_4_87};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_87 = {decodeResult_andMatrixOutputs_andMatrixInput_0_94, decodeResult_andMatrixOutputs_andMatrixInput_1_93};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_92 = {decodeResult_andMatrixOutputs_hi_hi_87, decodeResult_andMatrixOutputs_andMatrixInput_2_92};
  wire        decodeResult_andMatrixOutputs_29_2 = &{decodeResult_andMatrixOutputs_hi_92, decodeResult_andMatrixOutputs_lo_89};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_73 = {decodeResult_andMatrixOutputs_andMatrixInput_4_88, decodeResult_andMatrixOutputs_andMatrixInput_5_73};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_90 = {decodeResult_andMatrixOutputs_lo_hi_73, decodeResult_andMatrixOutputs_andMatrixInput_6_45};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_45 = {decodeResult_andMatrixOutputs_andMatrixInput_2_93, decodeResult_andMatrixOutputs_andMatrixInput_3_90};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_88 = {decodeResult_andMatrixOutputs_andMatrixInput_0_95, decodeResult_andMatrixOutputs_andMatrixInput_1_94};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_93 = {decodeResult_andMatrixOutputs_hi_hi_88, decodeResult_andMatrixOutputs_hi_lo_45};
  wire        decodeResult_andMatrixOutputs_132_2 = &{decodeResult_andMatrixOutputs_hi_93, decodeResult_andMatrixOutputs_lo_90};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_91 = {decodeResult_andMatrixOutputs_andMatrixInput_3_91, decodeResult_andMatrixOutputs_andMatrixInput_4_89};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_89 = {decodeResult_andMatrixOutputs_andMatrixInput_0_96, decodeResult_andMatrixOutputs_andMatrixInput_1_95};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_94 = {decodeResult_andMatrixOutputs_hi_hi_89, decodeResult_andMatrixOutputs_andMatrixInput_2_94};
  wire        decodeResult_andMatrixOutputs_87_2 = &{decodeResult_andMatrixOutputs_hi_94, decodeResult_andMatrixOutputs_lo_91};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_74 = {decodeResult_andMatrixOutputs_andMatrixInput_3_92, decodeResult_andMatrixOutputs_andMatrixInput_4_90};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_92 = {decodeResult_andMatrixOutputs_lo_hi_74, decodeResult_andMatrixOutputs_andMatrixInput_5_74};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_90 = {decodeResult_andMatrixOutputs_andMatrixInput_0_97, decodeResult_andMatrixOutputs_andMatrixInput_1_96};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_95 = {decodeResult_andMatrixOutputs_hi_hi_90, decodeResult_andMatrixOutputs_andMatrixInput_2_95};
  wire        decodeResult_andMatrixOutputs_70_2 = &{decodeResult_andMatrixOutputs_hi_95, decodeResult_andMatrixOutputs_lo_92};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_75 = {decodeResult_andMatrixOutputs_andMatrixInput_3_93, decodeResult_andMatrixOutputs_andMatrixInput_4_91};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_93 = {decodeResult_andMatrixOutputs_lo_hi_75, decodeResult_andMatrixOutputs_andMatrixInput_5_75};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_91 = {decodeResult_andMatrixOutputs_andMatrixInput_0_98, decodeResult_andMatrixOutputs_andMatrixInput_1_97};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_96 = {decodeResult_andMatrixOutputs_hi_hi_91, decodeResult_andMatrixOutputs_andMatrixInput_2_96};
  wire        decodeResult_andMatrixOutputs_135_2 = &{decodeResult_andMatrixOutputs_hi_96, decodeResult_andMatrixOutputs_lo_93};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_94 = {decodeResult_andMatrixOutputs_andMatrixInput_3_94, decodeResult_andMatrixOutputs_andMatrixInput_4_92};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_92 = {decodeResult_andMatrixOutputs_andMatrixInput_0_99, decodeResult_andMatrixOutputs_andMatrixInput_1_98};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_97 = {decodeResult_andMatrixOutputs_hi_hi_92, decodeResult_andMatrixOutputs_andMatrixInput_2_97};
  wire        decodeResult_andMatrixOutputs_49_2 = &{decodeResult_andMatrixOutputs_hi_97, decodeResult_andMatrixOutputs_lo_94};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_76 = {decodeResult_andMatrixOutputs_andMatrixInput_4_93, decodeResult_andMatrixOutputs_andMatrixInput_5_76};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_95 = {decodeResult_andMatrixOutputs_lo_hi_76, decodeResult_andMatrixOutputs_andMatrixInput_6_46};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_46 = {decodeResult_andMatrixOutputs_andMatrixInput_2_98, decodeResult_andMatrixOutputs_andMatrixInput_3_95};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_93 = {decodeResult_andMatrixOutputs_andMatrixInput_0_100, decodeResult_andMatrixOutputs_andMatrixInput_1_99};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_98 = {decodeResult_andMatrixOutputs_hi_hi_93, decodeResult_andMatrixOutputs_hi_lo_46};
  wire        decodeResult_andMatrixOutputs_79_2 = &{decodeResult_andMatrixOutputs_hi_98, decodeResult_andMatrixOutputs_lo_95};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_77 = {decodeResult_andMatrixOutputs_andMatrixInput_3_96, decodeResult_andMatrixOutputs_andMatrixInput_4_94};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_96 = {decodeResult_andMatrixOutputs_lo_hi_77, decodeResult_andMatrixOutputs_andMatrixInput_5_77};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_94 = {decodeResult_andMatrixOutputs_andMatrixInput_0_101, decodeResult_andMatrixOutputs_andMatrixInput_1_100};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_99 = {decodeResult_andMatrixOutputs_hi_hi_94, decodeResult_andMatrixOutputs_andMatrixInput_2_99};
  wire        decodeResult_andMatrixOutputs_47_2 = &{decodeResult_andMatrixOutputs_hi_99, decodeResult_andMatrixOutputs_lo_96};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_78 = {decodeResult_andMatrixOutputs_andMatrixInput_4_95, decodeResult_andMatrixOutputs_andMatrixInput_5_78};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_97 = {decodeResult_andMatrixOutputs_lo_hi_78, decodeResult_andMatrixOutputs_andMatrixInput_6_47};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_47 = {decodeResult_andMatrixOutputs_andMatrixInput_2_100, decodeResult_andMatrixOutputs_andMatrixInput_3_97};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_95 = {decodeResult_andMatrixOutputs_andMatrixInput_0_102, decodeResult_andMatrixOutputs_andMatrixInput_1_101};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_100 = {decodeResult_andMatrixOutputs_hi_hi_95, decodeResult_andMatrixOutputs_hi_lo_47};
  wire        decodeResult_andMatrixOutputs_99_2 = &{decodeResult_andMatrixOutputs_hi_100, decodeResult_andMatrixOutputs_lo_97};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_79 = {decodeResult_andMatrixOutputs_andMatrixInput_3_98, decodeResult_andMatrixOutputs_andMatrixInput_4_96};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_98 = {decodeResult_andMatrixOutputs_lo_hi_79, decodeResult_andMatrixOutputs_andMatrixInput_5_79};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_96 = {decodeResult_andMatrixOutputs_andMatrixInput_0_103, decodeResult_andMatrixOutputs_andMatrixInput_1_102};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_101 = {decodeResult_andMatrixOutputs_hi_hi_96, decodeResult_andMatrixOutputs_andMatrixInput_2_101};
  wire        decodeResult_andMatrixOutputs_127_2 = &{decodeResult_andMatrixOutputs_hi_101, decodeResult_andMatrixOutputs_lo_98};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_80 = {decodeResult_andMatrixOutputs_andMatrixInput_3_99, decodeResult_andMatrixOutputs_andMatrixInput_4_97};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_99 = {decodeResult_andMatrixOutputs_lo_hi_80, decodeResult_andMatrixOutputs_andMatrixInput_5_80};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_97 = {decodeResult_andMatrixOutputs_andMatrixInput_0_104, decodeResult_andMatrixOutputs_andMatrixInput_1_103};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_102 = {decodeResult_andMatrixOutputs_hi_hi_97, decodeResult_andMatrixOutputs_andMatrixInput_2_102};
  wire        decodeResult_andMatrixOutputs_122_2 = &{decodeResult_andMatrixOutputs_hi_102, decodeResult_andMatrixOutputs_lo_99};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_81 = {decodeResult_andMatrixOutputs_andMatrixInput_3_100, decodeResult_andMatrixOutputs_andMatrixInput_4_98};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_100 = {decodeResult_andMatrixOutputs_lo_hi_81, decodeResult_andMatrixOutputs_andMatrixInput_5_81};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_98 = {decodeResult_andMatrixOutputs_andMatrixInput_0_105, decodeResult_andMatrixOutputs_andMatrixInput_1_104};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_103 = {decodeResult_andMatrixOutputs_hi_hi_98, decodeResult_andMatrixOutputs_andMatrixInput_2_103};
  wire        decodeResult_andMatrixOutputs_134_2 = &{decodeResult_andMatrixOutputs_hi_103, decodeResult_andMatrixOutputs_lo_100};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_82 = {decodeResult_andMatrixOutputs_andMatrixInput_3_101, decodeResult_andMatrixOutputs_andMatrixInput_4_99};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_101 = {decodeResult_andMatrixOutputs_lo_hi_82, decodeResult_andMatrixOutputs_andMatrixInput_5_82};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_99 = {decodeResult_andMatrixOutputs_andMatrixInput_0_106, decodeResult_andMatrixOutputs_andMatrixInput_1_105};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_104 = {decodeResult_andMatrixOutputs_hi_hi_99, decodeResult_andMatrixOutputs_andMatrixInput_2_104};
  wire        decodeResult_andMatrixOutputs_35_2 = &{decodeResult_andMatrixOutputs_hi_104, decodeResult_andMatrixOutputs_lo_101};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_83 = {decodeResult_andMatrixOutputs_andMatrixInput_4_100, decodeResult_andMatrixOutputs_andMatrixInput_5_83};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_102 = {decodeResult_andMatrixOutputs_lo_hi_83, decodeResult_andMatrixOutputs_andMatrixInput_6_48};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_48 = {decodeResult_andMatrixOutputs_andMatrixInput_2_105, decodeResult_andMatrixOutputs_andMatrixInput_3_102};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_100 = {decodeResult_andMatrixOutputs_andMatrixInput_0_107, decodeResult_andMatrixOutputs_andMatrixInput_1_106};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_105 = {decodeResult_andMatrixOutputs_hi_hi_100, decodeResult_andMatrixOutputs_hi_lo_48};
  wire        decodeResult_andMatrixOutputs_131_2 = &{decodeResult_andMatrixOutputs_hi_105, decodeResult_andMatrixOutputs_lo_102};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_84 = {decodeResult_andMatrixOutputs_andMatrixInput_3_103, decodeResult_andMatrixOutputs_andMatrixInput_4_101};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_103 = {decodeResult_andMatrixOutputs_lo_hi_84, decodeResult_andMatrixOutputs_andMatrixInput_5_84};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_101 = {decodeResult_andMatrixOutputs_andMatrixInput_0_108, decodeResult_andMatrixOutputs_andMatrixInput_1_107};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_106 = {decodeResult_andMatrixOutputs_hi_hi_101, decodeResult_andMatrixOutputs_andMatrixInput_2_106};
  wire        decodeResult_andMatrixOutputs_125_2 = &{decodeResult_andMatrixOutputs_hi_106, decodeResult_andMatrixOutputs_lo_103};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_85 = {decodeResult_andMatrixOutputs_andMatrixInput_4_102, decodeResult_andMatrixOutputs_andMatrixInput_5_85};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_104 = {decodeResult_andMatrixOutputs_lo_hi_85, decodeResult_andMatrixOutputs_andMatrixInput_6_49};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_49 = {decodeResult_andMatrixOutputs_andMatrixInput_2_107, decodeResult_andMatrixOutputs_andMatrixInput_3_104};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_102 = {decodeResult_andMatrixOutputs_andMatrixInput_0_109, decodeResult_andMatrixOutputs_andMatrixInput_1_108};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_107 = {decodeResult_andMatrixOutputs_hi_hi_102, decodeResult_andMatrixOutputs_hi_lo_49};
  wire        decodeResult_andMatrixOutputs_43_2 = &{decodeResult_andMatrixOutputs_hi_107, decodeResult_andMatrixOutputs_lo_104};
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_86 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_87 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_50 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_51 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_109 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_107 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_52 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_109 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_91 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_92 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_93 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_113 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_94 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_95 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_119 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_96 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_97 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_98 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_99 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_53 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_101 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_102 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_54 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_55 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_105 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_56 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_57 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_128 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_129 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_130 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_108 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_5_109 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_133 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_134 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_135 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_58 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_3_141 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_137 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_4_138 = decodeResult_plaInput[31];
  wire        decodeResult_andMatrixOutputs_andMatrixInput_6_59 = decodeResult_plaInput[31];
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_86 = {decodeResult_andMatrixOutputs_andMatrixInput_3_105, decodeResult_andMatrixOutputs_andMatrixInput_4_103};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_105 = {decodeResult_andMatrixOutputs_lo_hi_86, decodeResult_andMatrixOutputs_andMatrixInput_5_86};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_103 = {decodeResult_andMatrixOutputs_andMatrixInput_0_110, decodeResult_andMatrixOutputs_andMatrixInput_1_109};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_108 = {decodeResult_andMatrixOutputs_hi_hi_103, decodeResult_andMatrixOutputs_andMatrixInput_2_108};
  wire        decodeResult_andMatrixOutputs_100_2 = &{decodeResult_andMatrixOutputs_hi_108, decodeResult_andMatrixOutputs_lo_105};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_87 = {decodeResult_andMatrixOutputs_andMatrixInput_3_106, decodeResult_andMatrixOutputs_andMatrixInput_4_104};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_106 = {decodeResult_andMatrixOutputs_lo_hi_87, decodeResult_andMatrixOutputs_andMatrixInput_5_87};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_104 = {decodeResult_andMatrixOutputs_andMatrixInput_0_111, decodeResult_andMatrixOutputs_andMatrixInput_1_110};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_109 = {decodeResult_andMatrixOutputs_hi_hi_104, decodeResult_andMatrixOutputs_andMatrixInput_2_109};
  wire        decodeResult_andMatrixOutputs_119_2 = &{decodeResult_andMatrixOutputs_hi_109, decodeResult_andMatrixOutputs_lo_106};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_88 = {decodeResult_andMatrixOutputs_andMatrixInput_4_105, decodeResult_andMatrixOutputs_andMatrixInput_5_88};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_107 = {decodeResult_andMatrixOutputs_lo_hi_88, decodeResult_andMatrixOutputs_andMatrixInput_6_50};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_50 = {decodeResult_andMatrixOutputs_andMatrixInput_2_110, decodeResult_andMatrixOutputs_andMatrixInput_3_107};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_105 = {decodeResult_andMatrixOutputs_andMatrixInput_0_112, decodeResult_andMatrixOutputs_andMatrixInput_1_111};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_110 = {decodeResult_andMatrixOutputs_hi_hi_105, decodeResult_andMatrixOutputs_hi_lo_50};
  wire        decodeResult_andMatrixOutputs_27_2 = &{decodeResult_andMatrixOutputs_hi_110, decodeResult_andMatrixOutputs_lo_107};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_89 = {decodeResult_andMatrixOutputs_andMatrixInput_4_106, decodeResult_andMatrixOutputs_andMatrixInput_5_89};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_108 = {decodeResult_andMatrixOutputs_lo_hi_89, decodeResult_andMatrixOutputs_andMatrixInput_6_51};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_51 = {decodeResult_andMatrixOutputs_andMatrixInput_2_111, decodeResult_andMatrixOutputs_andMatrixInput_3_108};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_106 = {decodeResult_andMatrixOutputs_andMatrixInput_0_113, decodeResult_andMatrixOutputs_andMatrixInput_1_112};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_111 = {decodeResult_andMatrixOutputs_hi_hi_106, decodeResult_andMatrixOutputs_hi_lo_51};
  wire        decodeResult_andMatrixOutputs_105_2 = &{decodeResult_andMatrixOutputs_hi_111, decodeResult_andMatrixOutputs_lo_108};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_109 = {decodeResult_andMatrixOutputs_andMatrixInput_2_112, decodeResult_andMatrixOutputs_andMatrixInput_3_109};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_112 = {decodeResult_andMatrixOutputs_andMatrixInput_0_114, decodeResult_andMatrixOutputs_andMatrixInput_1_113};
  wire        decodeResult_andMatrixOutputs_51_2 = &{decodeResult_andMatrixOutputs_hi_112, decodeResult_andMatrixOutputs_lo_109};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_110 = {decodeResult_andMatrixOutputs_andMatrixInput_3_110, decodeResult_andMatrixOutputs_andMatrixInput_4_107};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_107 = {decodeResult_andMatrixOutputs_andMatrixInput_0_115, decodeResult_andMatrixOutputs_andMatrixInput_1_114};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_113 = {decodeResult_andMatrixOutputs_hi_hi_107, decodeResult_andMatrixOutputs_andMatrixInput_2_113};
  wire        decodeResult_andMatrixOutputs_118_2 = &{decodeResult_andMatrixOutputs_hi_113, decodeResult_andMatrixOutputs_lo_110};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_90 = {decodeResult_andMatrixOutputs_andMatrixInput_4_108, decodeResult_andMatrixOutputs_andMatrixInput_5_90};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_111 = {decodeResult_andMatrixOutputs_lo_hi_90, decodeResult_andMatrixOutputs_andMatrixInput_6_52};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_52 = {decodeResult_andMatrixOutputs_andMatrixInput_2_114, decodeResult_andMatrixOutputs_andMatrixInput_3_111};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_108 = {decodeResult_andMatrixOutputs_andMatrixInput_0_116, decodeResult_andMatrixOutputs_andMatrixInput_1_115};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_114 = {decodeResult_andMatrixOutputs_hi_hi_108, decodeResult_andMatrixOutputs_hi_lo_52};
  wire        decodeResult_andMatrixOutputs_38_2 = &{decodeResult_andMatrixOutputs_hi_114, decodeResult_andMatrixOutputs_lo_111};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_112 = {decodeResult_andMatrixOutputs_andMatrixInput_3_112, decodeResult_andMatrixOutputs_andMatrixInput_4_109};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_109 = {decodeResult_andMatrixOutputs_andMatrixInput_0_117, decodeResult_andMatrixOutputs_andMatrixInput_1_116};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_115 = {decodeResult_andMatrixOutputs_hi_hi_109, decodeResult_andMatrixOutputs_andMatrixInput_2_115};
  wire        decodeResult_andMatrixOutputs_115_2 = &{decodeResult_andMatrixOutputs_hi_115, decodeResult_andMatrixOutputs_lo_112};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_91 = {decodeResult_andMatrixOutputs_andMatrixInput_3_113, decodeResult_andMatrixOutputs_andMatrixInput_4_110};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_113 = {decodeResult_andMatrixOutputs_lo_hi_91, decodeResult_andMatrixOutputs_andMatrixInput_5_91};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_110 = {decodeResult_andMatrixOutputs_andMatrixInput_0_118, decodeResult_andMatrixOutputs_andMatrixInput_1_117};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_116 = {decodeResult_andMatrixOutputs_hi_hi_110, decodeResult_andMatrixOutputs_andMatrixInput_2_116};
  wire        decodeResult_andMatrixOutputs_31_2 = &{decodeResult_andMatrixOutputs_hi_116, decodeResult_andMatrixOutputs_lo_113};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_92 = {decodeResult_andMatrixOutputs_andMatrixInput_3_114, decodeResult_andMatrixOutputs_andMatrixInput_4_111};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_114 = {decodeResult_andMatrixOutputs_lo_hi_92, decodeResult_andMatrixOutputs_andMatrixInput_5_92};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_111 = {decodeResult_andMatrixOutputs_andMatrixInput_0_119, decodeResult_andMatrixOutputs_andMatrixInput_1_118};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_117 = {decodeResult_andMatrixOutputs_hi_hi_111, decodeResult_andMatrixOutputs_andMatrixInput_2_117};
  wire        decodeResult_andMatrixOutputs_1_2 = &{decodeResult_andMatrixOutputs_hi_117, decodeResult_andMatrixOutputs_lo_114};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_93 = {decodeResult_andMatrixOutputs_andMatrixInput_3_115, decodeResult_andMatrixOutputs_andMatrixInput_4_112};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_115 = {decodeResult_andMatrixOutputs_lo_hi_93, decodeResult_andMatrixOutputs_andMatrixInput_5_93};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_112 = {decodeResult_andMatrixOutputs_andMatrixInput_0_120, decodeResult_andMatrixOutputs_andMatrixInput_1_119};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_118 = {decodeResult_andMatrixOutputs_hi_hi_112, decodeResult_andMatrixOutputs_andMatrixInput_2_118};
  wire        decodeResult_andMatrixOutputs_102_2 = &{decodeResult_andMatrixOutputs_hi_118, decodeResult_andMatrixOutputs_lo_115};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_116 = {decodeResult_andMatrixOutputs_andMatrixInput_3_116, decodeResult_andMatrixOutputs_andMatrixInput_4_113};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_113 = {decodeResult_andMatrixOutputs_andMatrixInput_0_121, decodeResult_andMatrixOutputs_andMatrixInput_1_120};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_119 = {decodeResult_andMatrixOutputs_hi_hi_113, decodeResult_andMatrixOutputs_andMatrixInput_2_119};
  wire        decodeResult_andMatrixOutputs_112_2 = &{decodeResult_andMatrixOutputs_hi_119, decodeResult_andMatrixOutputs_lo_116};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_94 = {decodeResult_andMatrixOutputs_andMatrixInput_3_117, decodeResult_andMatrixOutputs_andMatrixInput_4_114};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_117 = {decodeResult_andMatrixOutputs_lo_hi_94, decodeResult_andMatrixOutputs_andMatrixInput_5_94};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_114 = {decodeResult_andMatrixOutputs_andMatrixInput_0_122, decodeResult_andMatrixOutputs_andMatrixInput_1_121};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_120 = {decodeResult_andMatrixOutputs_hi_hi_114, decodeResult_andMatrixOutputs_andMatrixInput_2_120};
  wire        decodeResult_andMatrixOutputs_91_2 = &{decodeResult_andMatrixOutputs_hi_120, decodeResult_andMatrixOutputs_lo_117};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_95 = {decodeResult_andMatrixOutputs_andMatrixInput_3_118, decodeResult_andMatrixOutputs_andMatrixInput_4_115};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_118 = {decodeResult_andMatrixOutputs_lo_hi_95, decodeResult_andMatrixOutputs_andMatrixInput_5_95};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_115 = {decodeResult_andMatrixOutputs_andMatrixInput_0_123, decodeResult_andMatrixOutputs_andMatrixInput_1_122};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_121 = {decodeResult_andMatrixOutputs_hi_hi_115, decodeResult_andMatrixOutputs_andMatrixInput_2_121};
  wire        decodeResult_andMatrixOutputs_81_2 = &{decodeResult_andMatrixOutputs_hi_121, decodeResult_andMatrixOutputs_lo_118};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_119 = {decodeResult_andMatrixOutputs_andMatrixInput_2_122, decodeResult_andMatrixOutputs_andMatrixInput_3_119};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_122 = {decodeResult_andMatrixOutputs_andMatrixInput_0_124, decodeResult_andMatrixOutputs_andMatrixInput_1_123};
  wire        decodeResult_andMatrixOutputs_42_2 = &{decodeResult_andMatrixOutputs_hi_122, decodeResult_andMatrixOutputs_lo_119};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_96 = {decodeResult_andMatrixOutputs_andMatrixInput_3_120, decodeResult_andMatrixOutputs_andMatrixInput_4_116};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_120 = {decodeResult_andMatrixOutputs_lo_hi_96, decodeResult_andMatrixOutputs_andMatrixInput_5_96};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_116 = {decodeResult_andMatrixOutputs_andMatrixInput_0_125, decodeResult_andMatrixOutputs_andMatrixInput_1_124};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_123 = {decodeResult_andMatrixOutputs_hi_hi_116, decodeResult_andMatrixOutputs_andMatrixInput_2_123};
  wire        decodeResult_andMatrixOutputs_109_2 = &{decodeResult_andMatrixOutputs_hi_123, decodeResult_andMatrixOutputs_lo_120};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_97 = {decodeResult_andMatrixOutputs_andMatrixInput_3_121, decodeResult_andMatrixOutputs_andMatrixInput_4_117};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_121 = {decodeResult_andMatrixOutputs_lo_hi_97, decodeResult_andMatrixOutputs_andMatrixInput_5_97};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_117 = {decodeResult_andMatrixOutputs_andMatrixInput_0_126, decodeResult_andMatrixOutputs_andMatrixInput_1_125};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_124 = {decodeResult_andMatrixOutputs_hi_hi_117, decodeResult_andMatrixOutputs_andMatrixInput_2_124};
  wire        decodeResult_andMatrixOutputs_124_2 = &{decodeResult_andMatrixOutputs_hi_124, decodeResult_andMatrixOutputs_lo_121};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_98 = {decodeResult_andMatrixOutputs_andMatrixInput_3_122, decodeResult_andMatrixOutputs_andMatrixInput_4_118};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_122 = {decodeResult_andMatrixOutputs_lo_hi_98, decodeResult_andMatrixOutputs_andMatrixInput_5_98};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_118 = {decodeResult_andMatrixOutputs_andMatrixInput_0_127, decodeResult_andMatrixOutputs_andMatrixInput_1_126};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_125 = {decodeResult_andMatrixOutputs_hi_hi_118, decodeResult_andMatrixOutputs_andMatrixInput_2_125};
  wire        decodeResult_andMatrixOutputs_5_2 = &{decodeResult_andMatrixOutputs_hi_125, decodeResult_andMatrixOutputs_lo_122};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_99 = {decodeResult_andMatrixOutputs_andMatrixInput_3_123, decodeResult_andMatrixOutputs_andMatrixInput_4_119};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_123 = {decodeResult_andMatrixOutputs_lo_hi_99, decodeResult_andMatrixOutputs_andMatrixInput_5_99};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_119 = {decodeResult_andMatrixOutputs_andMatrixInput_0_128, decodeResult_andMatrixOutputs_andMatrixInput_1_127};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_126 = {decodeResult_andMatrixOutputs_hi_hi_119, decodeResult_andMatrixOutputs_andMatrixInput_2_126};
  wire        decodeResult_andMatrixOutputs_72_2 = &{decodeResult_andMatrixOutputs_hi_126, decodeResult_andMatrixOutputs_lo_123};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_100 = {decodeResult_andMatrixOutputs_andMatrixInput_4_120, decodeResult_andMatrixOutputs_andMatrixInput_5_100};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_124 = {decodeResult_andMatrixOutputs_lo_hi_100, decodeResult_andMatrixOutputs_andMatrixInput_6_53};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_53 = {decodeResult_andMatrixOutputs_andMatrixInput_2_127, decodeResult_andMatrixOutputs_andMatrixInput_3_124};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_120 = {decodeResult_andMatrixOutputs_andMatrixInput_0_129, decodeResult_andMatrixOutputs_andMatrixInput_1_128};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_127 = {decodeResult_andMatrixOutputs_hi_hi_120, decodeResult_andMatrixOutputs_hi_lo_53};
  wire        decodeResult_andMatrixOutputs_111_2 = &{decodeResult_andMatrixOutputs_hi_127, decodeResult_andMatrixOutputs_lo_124};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_101 = {decodeResult_andMatrixOutputs_andMatrixInput_3_125, decodeResult_andMatrixOutputs_andMatrixInput_4_121};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_125 = {decodeResult_andMatrixOutputs_lo_hi_101, decodeResult_andMatrixOutputs_andMatrixInput_5_101};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_121 = {decodeResult_andMatrixOutputs_andMatrixInput_0_130, decodeResult_andMatrixOutputs_andMatrixInput_1_129};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_128 = {decodeResult_andMatrixOutputs_hi_hi_121, decodeResult_andMatrixOutputs_andMatrixInput_2_128};
  wire        decodeResult_andMatrixOutputs_3_2 = &{decodeResult_andMatrixOutputs_hi_128, decodeResult_andMatrixOutputs_lo_125};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_102 = {decodeResult_andMatrixOutputs_andMatrixInput_3_126, decodeResult_andMatrixOutputs_andMatrixInput_4_122};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_126 = {decodeResult_andMatrixOutputs_lo_hi_102, decodeResult_andMatrixOutputs_andMatrixInput_5_102};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_122 = {decodeResult_andMatrixOutputs_andMatrixInput_0_131, decodeResult_andMatrixOutputs_andMatrixInput_1_130};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_129 = {decodeResult_andMatrixOutputs_hi_hi_122, decodeResult_andMatrixOutputs_andMatrixInput_2_129};
  wire        decodeResult_andMatrixOutputs_37_2 = &{decodeResult_andMatrixOutputs_hi_129, decodeResult_andMatrixOutputs_lo_126};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_103 = {decodeResult_andMatrixOutputs_andMatrixInput_4_123, decodeResult_andMatrixOutputs_andMatrixInput_5_103};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_127 = {decodeResult_andMatrixOutputs_lo_hi_103, decodeResult_andMatrixOutputs_andMatrixInput_6_54};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_54 = {decodeResult_andMatrixOutputs_andMatrixInput_2_130, decodeResult_andMatrixOutputs_andMatrixInput_3_127};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_123 = {decodeResult_andMatrixOutputs_andMatrixInput_0_132, decodeResult_andMatrixOutputs_andMatrixInput_1_131};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_130 = {decodeResult_andMatrixOutputs_hi_hi_123, decodeResult_andMatrixOutputs_hi_lo_54};
  wire        decodeResult_andMatrixOutputs_26_2 = &{decodeResult_andMatrixOutputs_hi_130, decodeResult_andMatrixOutputs_lo_127};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_104 = {decodeResult_andMatrixOutputs_andMatrixInput_4_124, decodeResult_andMatrixOutputs_andMatrixInput_5_104};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_128 = {decodeResult_andMatrixOutputs_lo_hi_104, decodeResult_andMatrixOutputs_andMatrixInput_6_55};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_55 = {decodeResult_andMatrixOutputs_andMatrixInput_2_131, decodeResult_andMatrixOutputs_andMatrixInput_3_128};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_124 = {decodeResult_andMatrixOutputs_andMatrixInput_0_133, decodeResult_andMatrixOutputs_andMatrixInput_1_132};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_131 = {decodeResult_andMatrixOutputs_hi_hi_124, decodeResult_andMatrixOutputs_hi_lo_55};
  wire        decodeResult_andMatrixOutputs_52_2 = &{decodeResult_andMatrixOutputs_hi_131, decodeResult_andMatrixOutputs_lo_128};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_105 = {decodeResult_andMatrixOutputs_andMatrixInput_3_129, decodeResult_andMatrixOutputs_andMatrixInput_4_125};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_129 = {decodeResult_andMatrixOutputs_lo_hi_105, decodeResult_andMatrixOutputs_andMatrixInput_5_105};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_125 = {decodeResult_andMatrixOutputs_andMatrixInput_0_134, decodeResult_andMatrixOutputs_andMatrixInput_1_133};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_132 = {decodeResult_andMatrixOutputs_hi_hi_125, decodeResult_andMatrixOutputs_andMatrixInput_2_132};
  wire        decodeResult_andMatrixOutputs_41_2 = &{decodeResult_andMatrixOutputs_hi_132, decodeResult_andMatrixOutputs_lo_129};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_106 = {decodeResult_andMatrixOutputs_andMatrixInput_4_126, decodeResult_andMatrixOutputs_andMatrixInput_5_106};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_130 = {decodeResult_andMatrixOutputs_lo_hi_106, decodeResult_andMatrixOutputs_andMatrixInput_6_56};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_56 = {decodeResult_andMatrixOutputs_andMatrixInput_2_133, decodeResult_andMatrixOutputs_andMatrixInput_3_130};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_126 = {decodeResult_andMatrixOutputs_andMatrixInput_0_135, decodeResult_andMatrixOutputs_andMatrixInput_1_134};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_133 = {decodeResult_andMatrixOutputs_hi_hi_126, decodeResult_andMatrixOutputs_hi_lo_56};
  wire        decodeResult_andMatrixOutputs_28_2 = &{decodeResult_andMatrixOutputs_hi_133, decodeResult_andMatrixOutputs_lo_130};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_107 = {decodeResult_andMatrixOutputs_andMatrixInput_4_127, decodeResult_andMatrixOutputs_andMatrixInput_5_107};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_131 = {decodeResult_andMatrixOutputs_lo_hi_107, decodeResult_andMatrixOutputs_andMatrixInput_6_57};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_57 = {decodeResult_andMatrixOutputs_andMatrixInput_2_134, decodeResult_andMatrixOutputs_andMatrixInput_3_131};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_127 = {decodeResult_andMatrixOutputs_andMatrixInput_0_136, decodeResult_andMatrixOutputs_andMatrixInput_1_135};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_134 = {decodeResult_andMatrixOutputs_hi_hi_127, decodeResult_andMatrixOutputs_hi_lo_57};
  wire        decodeResult_andMatrixOutputs_116_2 = &{decodeResult_andMatrixOutputs_hi_134, decodeResult_andMatrixOutputs_lo_131};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_132 = {decodeResult_andMatrixOutputs_andMatrixInput_3_132, decodeResult_andMatrixOutputs_andMatrixInput_4_128};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_128 = {decodeResult_andMatrixOutputs_andMatrixInput_0_137, decodeResult_andMatrixOutputs_andMatrixInput_1_136};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_135 = {decodeResult_andMatrixOutputs_hi_hi_128, decodeResult_andMatrixOutputs_andMatrixInput_2_135};
  wire        decodeResult_andMatrixOutputs_129_2 = &{decodeResult_andMatrixOutputs_hi_135, decodeResult_andMatrixOutputs_lo_132};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_133 = {decodeResult_andMatrixOutputs_andMatrixInput_3_133, decodeResult_andMatrixOutputs_andMatrixInput_4_129};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_129 = {decodeResult_andMatrixOutputs_andMatrixInput_0_138, decodeResult_andMatrixOutputs_andMatrixInput_1_137};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_136 = {decodeResult_andMatrixOutputs_hi_hi_129, decodeResult_andMatrixOutputs_andMatrixInput_2_136};
  wire        decodeResult_andMatrixOutputs_97_2 = &{decodeResult_andMatrixOutputs_hi_136, decodeResult_andMatrixOutputs_lo_133};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_134 = {decodeResult_andMatrixOutputs_andMatrixInput_3_134, decodeResult_andMatrixOutputs_andMatrixInput_4_130};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_130 = {decodeResult_andMatrixOutputs_andMatrixInput_0_139, decodeResult_andMatrixOutputs_andMatrixInput_1_138};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_137 = {decodeResult_andMatrixOutputs_hi_hi_130, decodeResult_andMatrixOutputs_andMatrixInput_2_137};
  wire        decodeResult_andMatrixOutputs_65_2 = &{decodeResult_andMatrixOutputs_hi_137, decodeResult_andMatrixOutputs_lo_134};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_108 = {decodeResult_andMatrixOutputs_andMatrixInput_3_135, decodeResult_andMatrixOutputs_andMatrixInput_4_131};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_135 = {decodeResult_andMatrixOutputs_lo_hi_108, decodeResult_andMatrixOutputs_andMatrixInput_5_108};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_131 = {decodeResult_andMatrixOutputs_andMatrixInput_0_140, decodeResult_andMatrixOutputs_andMatrixInput_1_139};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_138 = {decodeResult_andMatrixOutputs_hi_hi_131, decodeResult_andMatrixOutputs_andMatrixInput_2_138};
  wire        decodeResult_andMatrixOutputs_95_2 = &{decodeResult_andMatrixOutputs_hi_138, decodeResult_andMatrixOutputs_lo_135};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_109 = {decodeResult_andMatrixOutputs_andMatrixInput_3_136, decodeResult_andMatrixOutputs_andMatrixInput_4_132};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_136 = {decodeResult_andMatrixOutputs_lo_hi_109, decodeResult_andMatrixOutputs_andMatrixInput_5_109};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_132 = {decodeResult_andMatrixOutputs_andMatrixInput_0_141, decodeResult_andMatrixOutputs_andMatrixInput_1_140};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_139 = {decodeResult_andMatrixOutputs_hi_hi_132, decodeResult_andMatrixOutputs_andMatrixInput_2_139};
  wire        decodeResult_andMatrixOutputs_12_2 = &{decodeResult_andMatrixOutputs_hi_139, decodeResult_andMatrixOutputs_lo_136};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_137 = {decodeResult_andMatrixOutputs_andMatrixInput_3_137, decodeResult_andMatrixOutputs_andMatrixInput_4_133};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_133 = {decodeResult_andMatrixOutputs_andMatrixInput_0_142, decodeResult_andMatrixOutputs_andMatrixInput_1_141};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_140 = {decodeResult_andMatrixOutputs_hi_hi_133, decodeResult_andMatrixOutputs_andMatrixInput_2_140};
  wire        decodeResult_andMatrixOutputs_103_2 = &{decodeResult_andMatrixOutputs_hi_140, decodeResult_andMatrixOutputs_lo_137};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_138 = {decodeResult_andMatrixOutputs_andMatrixInput_3_138, decodeResult_andMatrixOutputs_andMatrixInput_4_134};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_134 = {decodeResult_andMatrixOutputs_andMatrixInput_0_143, decodeResult_andMatrixOutputs_andMatrixInput_1_142};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_141 = {decodeResult_andMatrixOutputs_hi_hi_134, decodeResult_andMatrixOutputs_andMatrixInput_2_141};
  wire        decodeResult_andMatrixOutputs_139_2 = &{decodeResult_andMatrixOutputs_hi_141, decodeResult_andMatrixOutputs_lo_138};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_139 = {decodeResult_andMatrixOutputs_andMatrixInput_3_139, decodeResult_andMatrixOutputs_andMatrixInput_4_135};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_135 = {decodeResult_andMatrixOutputs_andMatrixInput_0_144, decodeResult_andMatrixOutputs_andMatrixInput_1_143};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_142 = {decodeResult_andMatrixOutputs_hi_hi_135, decodeResult_andMatrixOutputs_andMatrixInput_2_142};
  wire        decodeResult_andMatrixOutputs_104_2 = &{decodeResult_andMatrixOutputs_hi_142, decodeResult_andMatrixOutputs_lo_139};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_110 = {decodeResult_andMatrixOutputs_andMatrixInput_4_136, decodeResult_andMatrixOutputs_andMatrixInput_5_110};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_140 = {decodeResult_andMatrixOutputs_lo_hi_110, decodeResult_andMatrixOutputs_andMatrixInput_6_58};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_58 = {decodeResult_andMatrixOutputs_andMatrixInput_2_143, decodeResult_andMatrixOutputs_andMatrixInput_3_140};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_136 = {decodeResult_andMatrixOutputs_andMatrixInput_0_145, decodeResult_andMatrixOutputs_andMatrixInput_1_144};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_143 = {decodeResult_andMatrixOutputs_hi_hi_136, decodeResult_andMatrixOutputs_hi_lo_58};
  wire        decodeResult_andMatrixOutputs_126_2 = &{decodeResult_andMatrixOutputs_hi_143, decodeResult_andMatrixOutputs_lo_140};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_141 = {decodeResult_andMatrixOutputs_andMatrixInput_2_144, decodeResult_andMatrixOutputs_andMatrixInput_3_141};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_144 = {decodeResult_andMatrixOutputs_andMatrixInput_0_146, decodeResult_andMatrixOutputs_andMatrixInput_1_145};
  wire        decodeResult_andMatrixOutputs_143_2 = &{decodeResult_andMatrixOutputs_hi_144, decodeResult_andMatrixOutputs_lo_141};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_142 = {decodeResult_andMatrixOutputs_andMatrixInput_3_142, decodeResult_andMatrixOutputs_andMatrixInput_4_137};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_137 = {decodeResult_andMatrixOutputs_andMatrixInput_0_147, decodeResult_andMatrixOutputs_andMatrixInput_1_146};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_145 = {decodeResult_andMatrixOutputs_hi_hi_137, decodeResult_andMatrixOutputs_andMatrixInput_2_145};
  wire        decodeResult_andMatrixOutputs_88_2 = &{decodeResult_andMatrixOutputs_hi_145, decodeResult_andMatrixOutputs_lo_142};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_143 = {decodeResult_andMatrixOutputs_andMatrixInput_3_143, decodeResult_andMatrixOutputs_andMatrixInput_4_138};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_138 = {decodeResult_andMatrixOutputs_andMatrixInput_0_148, decodeResult_andMatrixOutputs_andMatrixInput_1_147};
  wire [2:0]  decodeResult_andMatrixOutputs_hi_146 = {decodeResult_andMatrixOutputs_hi_hi_138, decodeResult_andMatrixOutputs_andMatrixInput_2_146};
  wire        decodeResult_andMatrixOutputs_85_2 = &{decodeResult_andMatrixOutputs_hi_146, decodeResult_andMatrixOutputs_lo_143};
  wire [1:0]  decodeResult_andMatrixOutputs_lo_hi_111 = {decodeResult_andMatrixOutputs_andMatrixInput_4_139, decodeResult_andMatrixOutputs_andMatrixInput_5_111};
  wire [2:0]  decodeResult_andMatrixOutputs_lo_144 = {decodeResult_andMatrixOutputs_lo_hi_111, decodeResult_andMatrixOutputs_andMatrixInput_6_59};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_lo_59 = {decodeResult_andMatrixOutputs_andMatrixInput_2_147, decodeResult_andMatrixOutputs_andMatrixInput_3_144};
  wire [1:0]  decodeResult_andMatrixOutputs_hi_hi_139 = {decodeResult_andMatrixOutputs_andMatrixInput_0_149, decodeResult_andMatrixOutputs_andMatrixInput_1_148};
  wire [3:0]  decodeResult_andMatrixOutputs_hi_147 = {decodeResult_andMatrixOutputs_hi_hi_139, decodeResult_andMatrixOutputs_hi_lo_59};
  wire        decodeResult_andMatrixOutputs_76_2 = &{decodeResult_andMatrixOutputs_hi_147, decodeResult_andMatrixOutputs_lo_144};
  wire [1:0]  decodeResult_orMatrixOutputs_lo = {decodeResult_andMatrixOutputs_130_2, decodeResult_andMatrixOutputs_127_2};
  wire [1:0]  _GEN = {decodeResult_andMatrixOutputs_22_2, decodeResult_andMatrixOutputs_30_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi;
  assign decodeResult_orMatrixOutputs_hi_hi = _GEN;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_lo_4;
  assign decodeResult_orMatrixOutputs_hi_hi_hi_lo_4 = _GEN;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_16;
  assign decodeResult_orMatrixOutputs_hi_hi_hi_16 = _GEN;
  wire [2:0]  decodeResult_orMatrixOutputs_hi = {decodeResult_orMatrixOutputs_hi_hi, decodeResult_andMatrixOutputs_75_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_lo = {decodeResult_andMatrixOutputs_103_2, decodeResult_andMatrixOutputs_104_2};
  wire [1:0]  _GEN_0 = {decodeResult_andMatrixOutputs_27_2, decodeResult_andMatrixOutputs_31_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi;
  assign decodeResult_orMatrixOutputs_lo_lo_hi = _GEN_0;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_19;
  assign decodeResult_orMatrixOutputs_hi_hi_19 = _GEN_0;
  wire [3:0]  decodeResult_orMatrixOutputs_lo_lo = {decodeResult_orMatrixOutputs_lo_lo_hi, decodeResult_orMatrixOutputs_lo_lo_lo};
  wire [1:0]  _GEN_1 = {decodeResult_andMatrixOutputs_122_2, decodeResult_andMatrixOutputs_125_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_lo;
  assign decodeResult_orMatrixOutputs_lo_hi_lo = _GEN_1;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_lo_3;
  assign decodeResult_orMatrixOutputs_lo_hi_lo_3 = _GEN_1;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_lo_12;
  assign decodeResult_orMatrixOutputs_lo_lo_lo_12 = _GEN_1;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_15;
  assign decodeResult_orMatrixOutputs_lo_lo_hi_15 = _GEN_1;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_hi = {decodeResult_andMatrixOutputs_98_2, decodeResult_andMatrixOutputs_60_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_hi = {decodeResult_orMatrixOutputs_lo_hi_hi_hi, decodeResult_andMatrixOutputs_49_2};
  wire [4:0]  decodeResult_orMatrixOutputs_lo_hi = {decodeResult_orMatrixOutputs_lo_hi_hi, decodeResult_orMatrixOutputs_lo_hi_lo};
  wire [8:0]  decodeResult_orMatrixOutputs_lo_1 = {decodeResult_orMatrixOutputs_lo_hi, decodeResult_orMatrixOutputs_lo_lo};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_lo = {decodeResult_andMatrixOutputs_57_2, decodeResult_andMatrixOutputs_14_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_hi = {decodeResult_andMatrixOutputs_58_2, decodeResult_andMatrixOutputs_123_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_lo_hi = {decodeResult_orMatrixOutputs_hi_lo_hi_hi, decodeResult_andMatrixOutputs_73_2};
  wire [4:0]  decodeResult_orMatrixOutputs_hi_lo = {decodeResult_orMatrixOutputs_hi_lo_hi, decodeResult_orMatrixOutputs_hi_lo_lo};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo = {decodeResult_andMatrixOutputs_50_2, decodeResult_andMatrixOutputs_25_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_hi = {decodeResult_andMatrixOutputs_15_2, decodeResult_andMatrixOutputs_93_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_hi_hi = {decodeResult_orMatrixOutputs_hi_hi_hi_hi, decodeResult_andMatrixOutputs_74_2};
  wire [4:0]  decodeResult_orMatrixOutputs_hi_hi_1 = {decodeResult_orMatrixOutputs_hi_hi_hi, decodeResult_orMatrixOutputs_hi_hi_lo};
  wire [9:0]  decodeResult_orMatrixOutputs_hi_1 = {decodeResult_orMatrixOutputs_hi_hi_1, decodeResult_orMatrixOutputs_hi_lo};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_1 = {decodeResult_andMatrixOutputs_72_2, decodeResult_andMatrixOutputs_3_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_2 = {decodeResult_orMatrixOutputs_lo_hi_1, decodeResult_andMatrixOutputs_28_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_2 = {decodeResult_andMatrixOutputs_128_2, decodeResult_andMatrixOutputs_91_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_2 = {decodeResult_orMatrixOutputs_hi_hi_2, decodeResult_andMatrixOutputs_81_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_3 = {decodeResult_andMatrixOutputs_116_2, decodeResult_andMatrixOutputs_88_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_3 = {decodeResult_andMatrixOutputs_124_2, decodeResult_andMatrixOutputs_5_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_3 = {decodeResult_orMatrixOutputs_hi_hi_3, decodeResult_andMatrixOutputs_52_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_4 = {decodeResult_andMatrixOutputs_13_2, decodeResult_andMatrixOutputs_105_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_1 = {decodeResult_andMatrixOutputs_111_2, decodeResult_andMatrixOutputs_139_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_1 = {decodeResult_andMatrixOutputs_105_2, decodeResult_andMatrixOutputs_38_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_2 = {decodeResult_orMatrixOutputs_lo_hi_hi_1, decodeResult_andMatrixOutputs_42_2};
  wire [4:0]  decodeResult_orMatrixOutputs_lo_4 = {decodeResult_orMatrixOutputs_lo_hi_2, decodeResult_orMatrixOutputs_lo_lo_1};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_1 = {decodeResult_andMatrixOutputs_68_2, decodeResult_andMatrixOutputs_47_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_1 = {decodeResult_andMatrixOutputs_89_2, decodeResult_andMatrixOutputs_110_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_hi_4 = {decodeResult_orMatrixOutputs_hi_hi_hi_1, decodeResult_andMatrixOutputs_138_2};
  wire [4:0]  decodeResult_orMatrixOutputs_hi_5 = {decodeResult_orMatrixOutputs_hi_hi_4, decodeResult_orMatrixOutputs_hi_lo_1};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_1 = {decodeResult_andMatrixOutputs_29_2, decodeResult_andMatrixOutputs_95_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_lo_2 = {decodeResult_orMatrixOutputs_lo_lo_hi_1, decodeResult_andMatrixOutputs_12_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_2 = {decodeResult_andMatrixOutputs_147_2, decodeResult_andMatrixOutputs_39_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_3 = {decodeResult_orMatrixOutputs_lo_hi_hi_2, decodeResult_andMatrixOutputs_80_2};
  wire [5:0]  decodeResult_orMatrixOutputs_lo_5 = {decodeResult_orMatrixOutputs_lo_hi_3, decodeResult_orMatrixOutputs_lo_lo_2};
  wire [1:0]  _GEN_2 = {decodeResult_andMatrixOutputs_144_2, decodeResult_andMatrixOutputs_33_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_1;
  assign decodeResult_orMatrixOutputs_hi_lo_hi_1 = _GEN_2;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_10;
  assign decodeResult_orMatrixOutputs_lo_10 = _GEN_2;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_15;
  assign decodeResult_orMatrixOutputs_hi_hi_15 = _GEN_2;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_lo_hi_3;
  assign decodeResult_orMatrixOutputs_hi_lo_lo_hi_3 = _GEN_2;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_lo_hi_4;
  assign decodeResult_orMatrixOutputs_hi_lo_lo_hi_4 = _GEN_2;
  wire [2:0]  decodeResult_orMatrixOutputs_hi_lo_2 = {decodeResult_orMatrixOutputs_hi_lo_hi_1, decodeResult_andMatrixOutputs_67_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_1 = {decodeResult_andMatrixOutputs_55_2, decodeResult_andMatrixOutputs_121_2};
  wire [1:0]  _GEN_3 = {decodeResult_andMatrixOutputs_83_2, decodeResult_andMatrixOutputs_18_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_2;
  assign decodeResult_orMatrixOutputs_hi_hi_hi_2 = _GEN_3;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_12;
  assign decodeResult_orMatrixOutputs_hi_12 = _GEN_3;
  wire [3:0]  decodeResult_orMatrixOutputs_hi_hi_5 = {decodeResult_orMatrixOutputs_hi_hi_hi_2, decodeResult_orMatrixOutputs_hi_hi_lo_1};
  wire [6:0]  decodeResult_orMatrixOutputs_hi_6 = {decodeResult_orMatrixOutputs_hi_hi_5, decodeResult_orMatrixOutputs_hi_lo_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_lo_1 = {decodeResult_andMatrixOutputs_51_2, decodeResult_andMatrixOutputs_81_2};
  wire [1:0]  _GEN_4 = {decodeResult_andMatrixOutputs_100_2, decodeResult_andMatrixOutputs_119_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_2;
  assign decodeResult_orMatrixOutputs_lo_lo_hi_2 = _GEN_4;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_lo_2;
  assign decodeResult_orMatrixOutputs_lo_hi_lo_2 = _GEN_4;
  wire [3:0]  decodeResult_orMatrixOutputs_lo_lo_3 = {decodeResult_orMatrixOutputs_lo_lo_hi_2, decodeResult_orMatrixOutputs_lo_lo_lo_1};
  wire [1:0]  _GEN_5 = {decodeResult_andMatrixOutputs_59_2, decodeResult_andMatrixOutputs_131_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_lo_1;
  assign decodeResult_orMatrixOutputs_lo_hi_lo_1 = _GEN_5;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_4;
  assign decodeResult_orMatrixOutputs_lo_hi_hi_4 = _GEN_5;
  wire [1:0]  _GEN_6 = {decodeResult_andMatrixOutputs_46_2, decodeResult_andMatrixOutputs_101_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_hi_1;
  assign decodeResult_orMatrixOutputs_lo_hi_hi_hi_1 = _GEN_6;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_28;
  assign decodeResult_orMatrixOutputs_lo_hi_28 = _GEN_6;
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_hi_3 = {decodeResult_orMatrixOutputs_lo_hi_hi_hi_1, decodeResult_andMatrixOutputs_145_2};
  wire [4:0]  decodeResult_orMatrixOutputs_lo_hi_4 = {decodeResult_orMatrixOutputs_lo_hi_hi_3, decodeResult_orMatrixOutputs_lo_hi_lo_1};
  wire [8:0]  decodeResult_orMatrixOutputs_lo_6 = {decodeResult_orMatrixOutputs_lo_hi_4, decodeResult_orMatrixOutputs_lo_lo_3};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_lo_1 = {decodeResult_andMatrixOutputs_13_2, decodeResult_andMatrixOutputs_98_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_hi_1 = {decodeResult_andMatrixOutputs_11_2, decodeResult_andMatrixOutputs_67_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_lo_hi_2 = {decodeResult_orMatrixOutputs_hi_lo_hi_hi_1, decodeResult_andMatrixOutputs_14_2};
  wire [4:0]  decodeResult_orMatrixOutputs_hi_lo_3 = {decodeResult_orMatrixOutputs_hi_lo_hi_2, decodeResult_orMatrixOutputs_hi_lo_lo_1};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_2 = {decodeResult_andMatrixOutputs_48_2, decodeResult_andMatrixOutputs_133_2};
  wire [1:0]  _GEN_7 = {decodeResult_andMatrixOutputs_16_2, decodeResult_andMatrixOutputs_23_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_hi_1;
  assign decodeResult_orMatrixOutputs_hi_hi_hi_hi_1 = _GEN_7;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_hi_2;
  assign decodeResult_orMatrixOutputs_hi_hi_hi_hi_2 = _GEN_7;
  wire [2:0]  decodeResult_orMatrixOutputs_hi_hi_hi_3 = {decodeResult_orMatrixOutputs_hi_hi_hi_hi_1, decodeResult_andMatrixOutputs_128_2};
  wire [4:0]  decodeResult_orMatrixOutputs_hi_hi_6 = {decodeResult_orMatrixOutputs_hi_hi_hi_3, decodeResult_orMatrixOutputs_hi_hi_lo_2};
  wire [9:0]  decodeResult_orMatrixOutputs_hi_7 = {decodeResult_orMatrixOutputs_hi_hi_6, decodeResult_orMatrixOutputs_hi_lo_3};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_lo_2 = {decodeResult_andMatrixOutputs_81_2, decodeResult_andMatrixOutputs_76_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_3 = {decodeResult_andMatrixOutputs_118_2, decodeResult_andMatrixOutputs_115_2};
  wire [3:0]  decodeResult_orMatrixOutputs_lo_lo_4 = {decodeResult_orMatrixOutputs_lo_lo_hi_3, decodeResult_orMatrixOutputs_lo_lo_lo_2};
  wire [3:0]  decodeResult_orMatrixOutputs_lo_hi_5 = {decodeResult_orMatrixOutputs_lo_hi_hi_4, decodeResult_orMatrixOutputs_lo_hi_lo_2};
  wire [7:0]  decodeResult_orMatrixOutputs_lo_7 = {decodeResult_orMatrixOutputs_lo_hi_5, decodeResult_orMatrixOutputs_lo_lo_4};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_lo_2 = {decodeResult_andMatrixOutputs_98_2, decodeResult_andMatrixOutputs_145_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_3 = {decodeResult_andMatrixOutputs_77_2, decodeResult_andMatrixOutputs_14_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_lo_4 = {decodeResult_orMatrixOutputs_hi_lo_hi_3, decodeResult_orMatrixOutputs_hi_lo_lo_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_3 = {decodeResult_andMatrixOutputs_48_2, decodeResult_andMatrixOutputs_11_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_hi_hi_4 = {decodeResult_orMatrixOutputs_hi_hi_hi_hi_2, decodeResult_andMatrixOutputs_128_2};
  wire [4:0]  decodeResult_orMatrixOutputs_hi_hi_7 = {decodeResult_orMatrixOutputs_hi_hi_hi_4, decodeResult_orMatrixOutputs_hi_hi_lo_3};
  wire [8:0]  decodeResult_orMatrixOutputs_hi_8 = {decodeResult_orMatrixOutputs_hi_hi_7, decodeResult_orMatrixOutputs_hi_lo_4};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_lo_3 = {decodeResult_andMatrixOutputs_3_2, decodeResult_andMatrixOutputs_12_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_4 = {decodeResult_andMatrixOutputs_31_2, decodeResult_andMatrixOutputs_91_2};
  wire [3:0]  decodeResult_orMatrixOutputs_lo_lo_5 = {decodeResult_orMatrixOutputs_lo_lo_hi_4, decodeResult_orMatrixOutputs_lo_lo_lo_3};
  wire [1:0]  _GEN_8 = {decodeResult_andMatrixOutputs_60_2, decodeResult_andMatrixOutputs_39_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_5;
  assign decodeResult_orMatrixOutputs_lo_hi_hi_5 = _GEN_8;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_lo;
  assign decodeResult_orMatrixOutputs_lo_hi_hi_lo = _GEN_8;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_lo_14;
  assign decodeResult_orMatrixOutputs_hi_lo_lo_14 = _GEN_8;
  wire [3:0]  decodeResult_orMatrixOutputs_lo_hi_6 = {decodeResult_orMatrixOutputs_lo_hi_hi_5, decodeResult_orMatrixOutputs_lo_hi_lo_3};
  wire [7:0]  decodeResult_orMatrixOutputs_lo_8 = {decodeResult_orMatrixOutputs_lo_hi_6, decodeResult_orMatrixOutputs_lo_lo_5};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_lo_3 = {decodeResult_andMatrixOutputs_130_2, decodeResult_andMatrixOutputs_98_2};
  wire [1:0]  _GEN_9 = {decodeResult_andMatrixOutputs_56_2, decodeResult_andMatrixOutputs_71_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_4;
  assign decodeResult_orMatrixOutputs_hi_lo_hi_4 = _GEN_9;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_hi_lo;
  assign decodeResult_orMatrixOutputs_hi_lo_hi_hi_lo = _GEN_9;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_lo_hi_1;
  assign decodeResult_orMatrixOutputs_hi_hi_lo_lo_hi_1 = _GEN_9;
  wire [3:0]  decodeResult_orMatrixOutputs_hi_lo_5 = {decodeResult_orMatrixOutputs_hi_lo_hi_4, decodeResult_orMatrixOutputs_hi_lo_lo_3};
  wire [1:0]  _GEN_10 = {decodeResult_andMatrixOutputs_128_2, decodeResult_andMatrixOutputs_83_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_4;
  assign decodeResult_orMatrixOutputs_hi_hi_lo_4 = _GEN_10;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_lo_hi;
  assign decodeResult_orMatrixOutputs_hi_hi_lo_lo_hi = _GEN_10;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_5 = {decodeResult_andMatrixOutputs_74_2, decodeResult_andMatrixOutputs_25_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_hi_8 = {decodeResult_orMatrixOutputs_hi_hi_hi_5, decodeResult_orMatrixOutputs_hi_hi_lo_4};
  wire [7:0]  decodeResult_orMatrixOutputs_hi_9 = {decodeResult_orMatrixOutputs_hi_hi_8, decodeResult_orMatrixOutputs_hi_lo_5};
  wire [1:0]  _GEN_11 = {decodeResult_andMatrixOutputs_1_2, decodeResult_andMatrixOutputs_103_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_6;
  assign decodeResult_orMatrixOutputs_lo_lo_6 = _GEN_11;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_lo_13;
  assign decodeResult_orMatrixOutputs_lo_lo_lo_13 = _GEN_11;
  wire [1:0]  _GEN_12 = {decodeResult_andMatrixOutputs_53_2, decodeResult_andMatrixOutputs_33_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_7;
  assign decodeResult_orMatrixOutputs_lo_hi_7 = _GEN_12;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_15;
  assign decodeResult_orMatrixOutputs_hi_lo_hi_15 = _GEN_12;
  wire [3:0]  decodeResult_orMatrixOutputs_lo_9 = {decodeResult_orMatrixOutputs_lo_hi_7, decodeResult_orMatrixOutputs_lo_lo_6};
  wire [1:0]  _GEN_13 = {decodeResult_andMatrixOutputs_30_2, decodeResult_andMatrixOutputs_123_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_6;
  assign decodeResult_orMatrixOutputs_hi_lo_6 = _GEN_13;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_hi_3;
  assign decodeResult_orMatrixOutputs_hi_hi_lo_hi_3 = _GEN_13;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_14;
  assign decodeResult_orMatrixOutputs_hi_hi_lo_14 = _GEN_13;
  wire [1:0]  _GEN_14 = {decodeResult_andMatrixOutputs_93_2, decodeResult_andMatrixOutputs_114_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_6;
  assign decodeResult_orMatrixOutputs_hi_hi_hi_6 = _GEN_14;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_hi_8;
  assign decodeResult_orMatrixOutputs_hi_hi_hi_hi_8 = _GEN_14;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_hi_11;
  assign decodeResult_orMatrixOutputs_hi_hi_hi_hi_11 = _GEN_14;
  wire [2:0]  decodeResult_orMatrixOutputs_hi_hi_9 = {decodeResult_orMatrixOutputs_hi_hi_hi_6, decodeResult_andMatrixOutputs_22_2};
  wire [4:0]  decodeResult_orMatrixOutputs_hi_10 = {decodeResult_orMatrixOutputs_hi_hi_9, decodeResult_orMatrixOutputs_hi_lo_6};
  wire [1:0]  _GEN_15 = {decodeResult_andMatrixOutputs_21_2, decodeResult_andMatrixOutputs_63_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_11;
  assign decodeResult_orMatrixOutputs_hi_11 = _GEN_15;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_14;
  assign decodeResult_orMatrixOutputs_hi_14 = _GEN_15;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_19;
  assign decodeResult_orMatrixOutputs_hi_lo_19 = _GEN_15;
  wire [1:0]  _GEN_16 = {decodeResult_andMatrixOutputs_63_2, decodeResult_andMatrixOutputs_67_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_8;
  assign decodeResult_orMatrixOutputs_lo_hi_8 = _GEN_16;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_hi_hi_1;
  assign decodeResult_orMatrixOutputs_lo_hi_hi_hi_hi_1 = _GEN_16;
  wire [2:0]  decodeResult_orMatrixOutputs_lo_11 = {decodeResult_orMatrixOutputs_lo_hi_8, decodeResult_andMatrixOutputs_113_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_7 = {decodeResult_andMatrixOutputs_106_2, decodeResult_andMatrixOutputs_21_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_10 = {decodeResult_andMatrixOutputs_0_2, decodeResult_andMatrixOutputs_71_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_13 = {decodeResult_orMatrixOutputs_hi_hi_10, decodeResult_orMatrixOutputs_hi_lo_7};
  wire [1:0]  _decodeResult_orMatrixOutputs_T_34 = {decodeResult_andMatrixOutputs_19_2, decodeResult_andMatrixOutputs_36_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_lo_2;
  assign decodeResult_orMatrixOutputs_lo_hi_hi_lo_2 = _decodeResult_orMatrixOutputs_T_34;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_lo_3;
  assign decodeResult_orMatrixOutputs_lo_hi_hi_lo_3 = _decodeResult_orMatrixOutputs_T_34;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_lo_12;
  assign decodeResult_orMatrixOutputs_hi_lo_lo_12 = _decodeResult_orMatrixOutputs_T_34;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_hi_10;
  assign decodeResult_orMatrixOutputs_lo_hi_hi_hi_10 = _decodeResult_orMatrixOutputs_T_34;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_lo_lo = {decodeResult_andMatrixOutputs_52_2, decodeResult_andMatrixOutputs_85_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_lo_hi = {decodeResult_andMatrixOutputs_81_2, decodeResult_andMatrixOutputs_26_2};
  wire [3:0]  decodeResult_orMatrixOutputs_lo_lo_lo_4 = {decodeResult_orMatrixOutputs_lo_lo_lo_hi, decodeResult_orMatrixOutputs_lo_lo_lo_lo};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_lo = {decodeResult_andMatrixOutputs_102_2, decodeResult_andMatrixOutputs_112_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_hi = {decodeResult_andMatrixOutputs_134_2, decodeResult_andMatrixOutputs_35_2};
  wire [3:0]  decodeResult_orMatrixOutputs_lo_lo_hi_5 = {decodeResult_orMatrixOutputs_lo_lo_hi_hi, decodeResult_orMatrixOutputs_lo_lo_hi_lo};
  wire [7:0]  decodeResult_orMatrixOutputs_lo_lo_7 = {decodeResult_orMatrixOutputs_lo_lo_hi_5, decodeResult_orMatrixOutputs_lo_lo_lo_4};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_lo_lo = {decodeResult_andMatrixOutputs_70_2, decodeResult_andMatrixOutputs_79_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_lo_hi = {decodeResult_andMatrixOutputs_80_2, decodeResult_andMatrixOutputs_29_2};
  wire [3:0]  decodeResult_orMatrixOutputs_lo_hi_lo_4 = {decodeResult_orMatrixOutputs_lo_hi_lo_hi, decodeResult_orMatrixOutputs_lo_hi_lo_lo};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_hi_hi = {decodeResult_andMatrixOutputs_67_2, decodeResult_andMatrixOutputs_13_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_hi_hi_2 = {decodeResult_orMatrixOutputs_lo_hi_hi_hi_hi, decodeResult_andMatrixOutputs_2_2};
  wire [4:0]  decodeResult_orMatrixOutputs_lo_hi_hi_6 = {decodeResult_orMatrixOutputs_lo_hi_hi_hi_2, decodeResult_orMatrixOutputs_lo_hi_hi_lo};
  wire [8:0]  decodeResult_orMatrixOutputs_lo_hi_9 = {decodeResult_orMatrixOutputs_lo_hi_hi_6, decodeResult_orMatrixOutputs_lo_hi_lo_4};
  wire [16:0] decodeResult_orMatrixOutputs_lo_12 = {decodeResult_orMatrixOutputs_lo_hi_9, decodeResult_orMatrixOutputs_lo_lo_7};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_lo_lo = {decodeResult_andMatrixOutputs_121_2, decodeResult_andMatrixOutputs_54_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_lo_hi = {decodeResult_andMatrixOutputs_146_2, decodeResult_andMatrixOutputs_117_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_lo_lo_4 = {decodeResult_orMatrixOutputs_hi_lo_lo_hi, decodeResult_orMatrixOutputs_hi_lo_lo_lo};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_lo = {decodeResult_andMatrixOutputs_34_2, decodeResult_andMatrixOutputs_57_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_hi_2 = {decodeResult_andMatrixOutputs_40_2, decodeResult_andMatrixOutputs_7_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_lo_hi_5 = {decodeResult_orMatrixOutputs_hi_lo_hi_hi_2, decodeResult_orMatrixOutputs_hi_lo_hi_lo};
  wire [7:0]  decodeResult_orMatrixOutputs_hi_lo_8 = {decodeResult_orMatrixOutputs_hi_lo_hi_5, decodeResult_orMatrixOutputs_hi_lo_lo_4};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_lo = {decodeResult_andMatrixOutputs_128_2, decodeResult_andMatrixOutputs_32_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_hi = {decodeResult_andMatrixOutputs_24_2, decodeResult_andMatrixOutputs_45_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_hi_lo_5 = {decodeResult_orMatrixOutputs_hi_hi_lo_hi, decodeResult_orMatrixOutputs_hi_hi_lo_lo};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_lo = {decodeResult_andMatrixOutputs_30_2, decodeResult_andMatrixOutputs_25_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_hi_hi = {decodeResult_andMatrixOutputs_50_2, decodeResult_andMatrixOutputs_44_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_hi_hi_hi_3 = {decodeResult_orMatrixOutputs_hi_hi_hi_hi_hi, decodeResult_andMatrixOutputs_138_2};
  wire [4:0]  decodeResult_orMatrixOutputs_hi_hi_hi_7 = {decodeResult_orMatrixOutputs_hi_hi_hi_hi_3, decodeResult_orMatrixOutputs_hi_hi_hi_lo};
  wire [8:0]  decodeResult_orMatrixOutputs_hi_hi_11 = {decodeResult_orMatrixOutputs_hi_hi_hi_7, decodeResult_orMatrixOutputs_hi_hi_lo_5};
  wire [16:0] decodeResult_orMatrixOutputs_hi_15 = {decodeResult_orMatrixOutputs_hi_hi_11, decodeResult_orMatrixOutputs_hi_lo_8};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_lo_hi_1 = {decodeResult_andMatrixOutputs_116_2, decodeResult_andMatrixOutputs_95_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_lo_lo_5 = {decodeResult_orMatrixOutputs_lo_lo_lo_hi_1, decodeResult_andMatrixOutputs_12_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_lo_1 = {decodeResult_andMatrixOutputs_37_2, decodeResult_andMatrixOutputs_41_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_hi_1 = {decodeResult_andMatrixOutputs_131_2, decodeResult_andMatrixOutputs_43_2};
  wire [3:0]  decodeResult_orMatrixOutputs_lo_lo_hi_6 = {decodeResult_orMatrixOutputs_lo_lo_hi_hi_1, decodeResult_orMatrixOutputs_lo_lo_hi_lo_1};
  wire [6:0]  decodeResult_orMatrixOutputs_lo_lo_8 = {decodeResult_orMatrixOutputs_lo_lo_hi_6, decodeResult_orMatrixOutputs_lo_lo_lo_5};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_lo_hi_1 = {decodeResult_andMatrixOutputs_86_2, decodeResult_andMatrixOutputs_2_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_lo_5 = {decodeResult_orMatrixOutputs_lo_hi_lo_hi_1, decodeResult_andMatrixOutputs_60_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_lo_1 = {decodeResult_andMatrixOutputs_46_2, decodeResult_andMatrixOutputs_8_2};
  wire [1:0]  _GEN_17 = {decodeResult_andMatrixOutputs_14_2, decodeResult_andMatrixOutputs_98_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_hi_3;
  assign decodeResult_orMatrixOutputs_lo_hi_hi_hi_3 = _GEN_17;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_16;
  assign decodeResult_orMatrixOutputs_hi_hi_16 = _GEN_17;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_hi_6;
  assign decodeResult_orMatrixOutputs_lo_hi_hi_hi_6 = _GEN_17;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_hi_7;
  assign decodeResult_orMatrixOutputs_lo_hi_hi_hi_7 = _GEN_17;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_14;
  assign decodeResult_orMatrixOutputs_hi_lo_hi_14 = _GEN_17;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_lo_13;
  assign decodeResult_orMatrixOutputs_hi_lo_lo_13 = _GEN_17;
  wire [3:0]  decodeResult_orMatrixOutputs_lo_hi_hi_7 = {decodeResult_orMatrixOutputs_lo_hi_hi_hi_3, decodeResult_orMatrixOutputs_lo_hi_hi_lo_1};
  wire [6:0]  decodeResult_orMatrixOutputs_lo_hi_10 = {decodeResult_orMatrixOutputs_lo_hi_hi_7, decodeResult_orMatrixOutputs_lo_hi_lo_5};
  wire [13:0] decodeResult_orMatrixOutputs_lo_13 = {decodeResult_orMatrixOutputs_lo_hi_10, decodeResult_orMatrixOutputs_lo_lo_8};
  wire [1:0]  _GEN_18 = {decodeResult_andMatrixOutputs_20_2, decodeResult_andMatrixOutputs_94_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_lo_hi_1;
  assign decodeResult_orMatrixOutputs_hi_lo_lo_hi_1 = _GEN_18;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_17;
  assign decodeResult_orMatrixOutputs_hi_hi_17 = _GEN_18;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_hi_12;
  assign decodeResult_orMatrixOutputs_hi_hi_hi_hi_12 = _GEN_18;
  wire [2:0]  decodeResult_orMatrixOutputs_hi_lo_lo_5 = {decodeResult_orMatrixOutputs_hi_lo_lo_hi_1, decodeResult_andMatrixOutputs_67_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_lo_1 = {decodeResult_andMatrixOutputs_9_2, decodeResult_andMatrixOutputs_148_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_hi_3 = {decodeResult_andMatrixOutputs_136_2, decodeResult_andMatrixOutputs_66_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_lo_hi_6 = {decodeResult_orMatrixOutputs_hi_lo_hi_hi_3, decodeResult_orMatrixOutputs_hi_lo_hi_lo_1};
  wire [6:0]  decodeResult_orMatrixOutputs_hi_lo_9 = {decodeResult_orMatrixOutputs_hi_lo_hi_6, decodeResult_orMatrixOutputs_hi_lo_lo_5};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_lo_1 = {decodeResult_andMatrixOutputs_84_2, decodeResult_andMatrixOutputs_120_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_hi_1 = {decodeResult_andMatrixOutputs_123_2, decodeResult_andMatrixOutputs_32_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_hi_lo_6 = {decodeResult_orMatrixOutputs_hi_hi_lo_hi_1, decodeResult_orMatrixOutputs_hi_hi_lo_lo_1};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_lo_1 = {decodeResult_andMatrixOutputs_24_2, decodeResult_andMatrixOutputs_58_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_hi_4 = {decodeResult_andMatrixOutputs_64_2, decodeResult_andMatrixOutputs_92_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_hi_hi_8 = {decodeResult_orMatrixOutputs_hi_hi_hi_hi_4, decodeResult_orMatrixOutputs_hi_hi_hi_lo_1};
  wire [7:0]  decodeResult_orMatrixOutputs_hi_hi_12 = {decodeResult_orMatrixOutputs_hi_hi_hi_8, decodeResult_orMatrixOutputs_hi_hi_lo_6};
  wire [14:0] decodeResult_orMatrixOutputs_hi_16 = {decodeResult_orMatrixOutputs_hi_hi_12, decodeResult_orMatrixOutputs_hi_lo_9};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_lo_hi_2 = {decodeResult_andMatrixOutputs_97_2, decodeResult_andMatrixOutputs_95_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_lo_lo_6 = {decodeResult_orMatrixOutputs_lo_lo_lo_hi_2, decodeResult_andMatrixOutputs_12_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_hi_2 = {decodeResult_andMatrixOutputs_91_2, decodeResult_andMatrixOutputs_111_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_lo_hi_7 = {decodeResult_orMatrixOutputs_lo_lo_hi_hi_2, decodeResult_andMatrixOutputs_28_2};
  wire [5:0]  decodeResult_orMatrixOutputs_lo_lo_9 = {decodeResult_orMatrixOutputs_lo_lo_hi_7, decodeResult_orMatrixOutputs_lo_lo_lo_6};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_lo_hi_2 = {decodeResult_andMatrixOutputs_70_2, decodeResult_andMatrixOutputs_99_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_lo_6 = {decodeResult_orMatrixOutputs_lo_hi_lo_hi_2, decodeResult_andMatrixOutputs_125_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_hi_4 = {decodeResult_andMatrixOutputs_86_2, decodeResult_andMatrixOutputs_39_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_hi_8 = {decodeResult_orMatrixOutputs_lo_hi_hi_hi_4, decodeResult_andMatrixOutputs_87_2};
  wire [5:0]  decodeResult_orMatrixOutputs_lo_hi_11 = {decodeResult_orMatrixOutputs_lo_hi_hi_8, decodeResult_orMatrixOutputs_lo_hi_lo_6};
  wire [11:0] decodeResult_orMatrixOutputs_lo_14 = {decodeResult_orMatrixOutputs_lo_hi_11, decodeResult_orMatrixOutputs_lo_lo_9};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_lo_hi_2 = {decodeResult_andMatrixOutputs_67_2, decodeResult_andMatrixOutputs_46_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_lo_lo_6 = {decodeResult_orMatrixOutputs_hi_lo_lo_hi_2, decodeResult_andMatrixOutputs_101_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_hi_4 = {decodeResult_andMatrixOutputs_141_2, decodeResult_andMatrixOutputs_63_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_lo_hi_7 = {decodeResult_orMatrixOutputs_hi_lo_hi_hi_4, decodeResult_andMatrixOutputs_54_2};
  wire [5:0]  decodeResult_orMatrixOutputs_hi_lo_10 = {decodeResult_orMatrixOutputs_hi_lo_hi_7, decodeResult_orMatrixOutputs_hi_lo_lo_6};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_hi_2 = {decodeResult_andMatrixOutputs_107_2, decodeResult_andMatrixOutputs_18_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_hi_lo_7 = {decodeResult_orMatrixOutputs_hi_hi_lo_hi_2, decodeResult_andMatrixOutputs_55_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_lo_2 = {decodeResult_andMatrixOutputs_40_2, decodeResult_andMatrixOutputs_78_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_hi_5 = {decodeResult_andMatrixOutputs_45_2, decodeResult_andMatrixOutputs_83_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_hi_hi_9 = {decodeResult_orMatrixOutputs_hi_hi_hi_hi_5, decodeResult_orMatrixOutputs_hi_hi_hi_lo_2};
  wire [6:0]  decodeResult_orMatrixOutputs_hi_hi_13 = {decodeResult_orMatrixOutputs_hi_hi_hi_9, decodeResult_orMatrixOutputs_hi_hi_lo_7};
  wire [12:0] decodeResult_orMatrixOutputs_hi_17 = {decodeResult_orMatrixOutputs_hi_hi_13, decodeResult_orMatrixOutputs_hi_lo_10};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_lo_7 = {decodeResult_andMatrixOutputs_105_2, decodeResult_andMatrixOutputs_116_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_8 = {decodeResult_andMatrixOutputs_135_2, decodeResult_andMatrixOutputs_122_2};
  wire [3:0]  decodeResult_orMatrixOutputs_lo_lo_10 = {decodeResult_orMatrixOutputs_lo_lo_hi_8, decodeResult_orMatrixOutputs_lo_lo_lo_7};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_lo_7 = {decodeResult_andMatrixOutputs_142_2, decodeResult_andMatrixOutputs_80_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_hi_5 = {decodeResult_andMatrixOutputs_14_2, decodeResult_andMatrixOutputs_13_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_hi_9 = {decodeResult_orMatrixOutputs_lo_hi_hi_hi_5, decodeResult_andMatrixOutputs_98_2};
  wire [4:0]  decodeResult_orMatrixOutputs_lo_hi_12 = {decodeResult_orMatrixOutputs_lo_hi_hi_9, decodeResult_orMatrixOutputs_lo_hi_lo_7};
  wire [8:0]  decodeResult_orMatrixOutputs_lo_15 = {decodeResult_orMatrixOutputs_lo_hi_12, decodeResult_orMatrixOutputs_lo_lo_10};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_lo_7 = {decodeResult_andMatrixOutputs_94_2, decodeResult_andMatrixOutputs_33_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_8 = {decodeResult_andMatrixOutputs_117_2, decodeResult_andMatrixOutputs_20_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_lo_11 = {decodeResult_orMatrixOutputs_hi_lo_hi_8, decodeResult_orMatrixOutputs_hi_lo_lo_7};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_8 = {decodeResult_andMatrixOutputs_40_2, decodeResult_andMatrixOutputs_137_2};
  wire [1:0]  _GEN_19 = {decodeResult_andMatrixOutputs_110_2, decodeResult_andMatrixOutputs_114_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_hi_6;
  assign decodeResult_orMatrixOutputs_hi_hi_hi_hi_6 = _GEN_19;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_20;
  assign decodeResult_orMatrixOutputs_hi_hi_hi_20 = _GEN_19;
  wire [2:0]  decodeResult_orMatrixOutputs_hi_hi_hi_10 = {decodeResult_orMatrixOutputs_hi_hi_hi_hi_6, decodeResult_andMatrixOutputs_53_2};
  wire [4:0]  decodeResult_orMatrixOutputs_hi_hi_14 = {decodeResult_orMatrixOutputs_hi_hi_hi_10, decodeResult_orMatrixOutputs_hi_hi_lo_8};
  wire [8:0]  decodeResult_orMatrixOutputs_hi_18 = {decodeResult_orMatrixOutputs_hi_hi_14, decodeResult_orMatrixOutputs_hi_lo_11};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_16 = {decodeResult_andMatrixOutputs_147_2, decodeResult_andMatrixOutputs_127_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_19 = {decodeResult_orMatrixOutputs_hi_hi_15, decodeResult_andMatrixOutputs_113_2};
  wire [1:0]  _GEN_20 = {decodeResult_andMatrixOutputs_47_2, decodeResult_andMatrixOutputs_122_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_13;
  assign decodeResult_orMatrixOutputs_lo_hi_13 = _GEN_20;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_lo_2;
  assign decodeResult_orMatrixOutputs_lo_lo_hi_lo_2 = _GEN_20;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_lo_3;
  assign decodeResult_orMatrixOutputs_lo_lo_hi_lo_3 = _GEN_20;
  wire [2:0]  decodeResult_orMatrixOutputs_lo_17 = {decodeResult_orMatrixOutputs_lo_hi_13, decodeResult_andMatrixOutputs_125_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_12 = {decodeResult_andMatrixOutputs_60_2, decodeResult_andMatrixOutputs_49_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_20 = {decodeResult_orMatrixOutputs_hi_hi_16, decodeResult_orMatrixOutputs_hi_lo_12};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_14 = {decodeResult_andMatrixOutputs_98_2, decodeResult_andMatrixOutputs_39_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_18 = {decodeResult_orMatrixOutputs_lo_hi_14, decodeResult_andMatrixOutputs_29_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_21 = {decodeResult_orMatrixOutputs_hi_hi_17, decodeResult_andMatrixOutputs_14_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_19 = {decodeResult_andMatrixOutputs_113_2, decodeResult_andMatrixOutputs_132_2};
  wire [1:0]  _GEN_21 = {decodeResult_andMatrixOutputs_18_2, decodeResult_andMatrixOutputs_19_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_18;
  assign decodeResult_orMatrixOutputs_hi_hi_18 = _GEN_21;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_18;
  assign decodeResult_orMatrixOutputs_hi_lo_18 = _GEN_21;
  wire [2:0]  decodeResult_orMatrixOutputs_hi_22 = {decodeResult_orMatrixOutputs_hi_hi_18, decodeResult_andMatrixOutputs_36_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_20 = {decodeResult_andMatrixOutputs_5_2, decodeResult_andMatrixOutputs_28_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_23 = {decodeResult_orMatrixOutputs_hi_hi_19, decodeResult_andMatrixOutputs_91_2};
  wire [1:0]  _GEN_22 = {decodeResult_andMatrixOutputs_125_2, decodeResult_andMatrixOutputs_1_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_lo_hi_3;
  assign decodeResult_orMatrixOutputs_lo_lo_lo_hi_3 = _GEN_22;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_lo_hi_4;
  assign decodeResult_orMatrixOutputs_lo_lo_lo_hi_4 = _GEN_22;
  wire [2:0]  decodeResult_orMatrixOutputs_lo_lo_lo_8 = {decodeResult_orMatrixOutputs_lo_lo_lo_hi_3, decodeResult_andMatrixOutputs_103_2};
  wire [1:0]  _GEN_23 = {decodeResult_andMatrixOutputs_132_2, decodeResult_andMatrixOutputs_49_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_hi_3;
  assign decodeResult_orMatrixOutputs_lo_lo_hi_hi_3 = _GEN_23;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_hi_4;
  assign decodeResult_orMatrixOutputs_lo_lo_hi_hi_4 = _GEN_23;
  wire [3:0]  decodeResult_orMatrixOutputs_lo_lo_hi_9 = {decodeResult_orMatrixOutputs_lo_lo_hi_hi_3, decodeResult_orMatrixOutputs_lo_lo_hi_lo_2};
  wire [6:0]  decodeResult_orMatrixOutputs_lo_lo_11 = {decodeResult_orMatrixOutputs_lo_lo_hi_9, decodeResult_orMatrixOutputs_lo_lo_lo_8};
  wire [1:0]  _GEN_24 = {decodeResult_andMatrixOutputs_113_2, decodeResult_andMatrixOutputs_147_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_lo_hi_3;
  assign decodeResult_orMatrixOutputs_lo_hi_lo_hi_3 = _GEN_24;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_lo_hi_4;
  assign decodeResult_orMatrixOutputs_lo_hi_lo_hi_4 = _GEN_24;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_16;
  assign decodeResult_orMatrixOutputs_lo_hi_hi_16 = _GEN_24;
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_lo_8 = {decodeResult_orMatrixOutputs_lo_hi_lo_hi_3, decodeResult_andMatrixOutputs_60_2};
  wire [3:0]  decodeResult_orMatrixOutputs_lo_hi_hi_10 = {decodeResult_orMatrixOutputs_lo_hi_hi_hi_6, decodeResult_orMatrixOutputs_lo_hi_hi_lo_2};
  wire [6:0]  decodeResult_orMatrixOutputs_lo_hi_15 = {decodeResult_orMatrixOutputs_lo_hi_hi_10, decodeResult_orMatrixOutputs_lo_hi_lo_8};
  wire [13:0] decodeResult_orMatrixOutputs_lo_21 = {decodeResult_orMatrixOutputs_lo_hi_15, decodeResult_orMatrixOutputs_lo_lo_11};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_lo_lo_8 = {decodeResult_orMatrixOutputs_hi_lo_lo_hi_3, decodeResult_andMatrixOutputs_67_2};
  wire [1:0]  _GEN_25 = {decodeResult_andMatrixOutputs_21_2, decodeResult_andMatrixOutputs_121_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_lo_2;
  assign decodeResult_orMatrixOutputs_hi_lo_hi_lo_2 = _GEN_25;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_lo_3;
  assign decodeResult_orMatrixOutputs_hi_lo_hi_lo_3 = _GEN_25;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_17;
  assign decodeResult_orMatrixOutputs_hi_hi_hi_17 = _GEN_25;
  wire [1:0]  _GEN_26 = {decodeResult_andMatrixOutputs_18_2, decodeResult_andMatrixOutputs_106_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_hi_5;
  assign decodeResult_orMatrixOutputs_hi_lo_hi_hi_5 = _GEN_26;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_hi_6;
  assign decodeResult_orMatrixOutputs_hi_lo_hi_hi_6 = _GEN_26;
  wire [3:0]  decodeResult_orMatrixOutputs_hi_lo_hi_9 = {decodeResult_orMatrixOutputs_hi_lo_hi_hi_5, decodeResult_orMatrixOutputs_hi_lo_hi_lo_2};
  wire [6:0]  decodeResult_orMatrixOutputs_hi_lo_13 = {decodeResult_orMatrixOutputs_hi_lo_hi_9, decodeResult_orMatrixOutputs_hi_lo_lo_8};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_lo_2 = {decodeResult_andMatrixOutputs_53_2, decodeResult_andMatrixOutputs_71_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_hi_lo_9 = {decodeResult_orMatrixOutputs_hi_hi_lo_hi_3, decodeResult_orMatrixOutputs_hi_hi_lo_lo_2};
  wire [1:0]  _GEN_27 = {decodeResult_andMatrixOutputs_114_2, decodeResult_andMatrixOutputs_22_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_lo_3;
  assign decodeResult_orMatrixOutputs_hi_hi_hi_lo_3 = _GEN_27;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_lo_hi;
  assign decodeResult_orMatrixOutputs_hi_hi_hi_lo_hi = _GEN_27;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_hi_7 = {decodeResult_andMatrixOutputs_93_2, decodeResult_andMatrixOutputs_82_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_hi_hi_11 = {decodeResult_orMatrixOutputs_hi_hi_hi_hi_7, decodeResult_orMatrixOutputs_hi_hi_hi_lo_3};
  wire [7:0]  decodeResult_orMatrixOutputs_hi_hi_20 = {decodeResult_orMatrixOutputs_hi_hi_hi_11, decodeResult_orMatrixOutputs_hi_hi_lo_9};
  wire [14:0] decodeResult_orMatrixOutputs_hi_24 = {decodeResult_orMatrixOutputs_hi_hi_20, decodeResult_orMatrixOutputs_hi_lo_13};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_lo_lo_9 = {decodeResult_orMatrixOutputs_lo_lo_lo_hi_4, decodeResult_andMatrixOutputs_103_2};
  wire [3:0]  decodeResult_orMatrixOutputs_lo_lo_hi_10 = {decodeResult_orMatrixOutputs_lo_lo_hi_hi_4, decodeResult_orMatrixOutputs_lo_lo_hi_lo_3};
  wire [6:0]  decodeResult_orMatrixOutputs_lo_lo_12 = {decodeResult_orMatrixOutputs_lo_lo_hi_10, decodeResult_orMatrixOutputs_lo_lo_lo_9};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_lo_9 = {decodeResult_orMatrixOutputs_lo_hi_lo_hi_4, decodeResult_andMatrixOutputs_60_2};
  wire [3:0]  decodeResult_orMatrixOutputs_lo_hi_hi_11 = {decodeResult_orMatrixOutputs_lo_hi_hi_hi_7, decodeResult_orMatrixOutputs_lo_hi_hi_lo_3};
  wire [6:0]  decodeResult_orMatrixOutputs_lo_hi_16 = {decodeResult_orMatrixOutputs_lo_hi_hi_11, decodeResult_orMatrixOutputs_lo_hi_lo_9};
  wire [13:0] decodeResult_orMatrixOutputs_lo_22 = {decodeResult_orMatrixOutputs_lo_hi_16, decodeResult_orMatrixOutputs_lo_lo_12};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_lo_lo_9 = {decodeResult_orMatrixOutputs_hi_lo_lo_hi_4, decodeResult_andMatrixOutputs_67_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_lo_hi_10 = {decodeResult_orMatrixOutputs_hi_lo_hi_hi_6, decodeResult_orMatrixOutputs_hi_lo_hi_lo_3};
  wire [6:0]  decodeResult_orMatrixOutputs_hi_lo_14 = {decodeResult_orMatrixOutputs_hi_lo_hi_10, decodeResult_orMatrixOutputs_hi_lo_lo_9};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_hi_4 = {decodeResult_andMatrixOutputs_123_2, decodeResult_andMatrixOutputs_53_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_hi_lo_10 = {decodeResult_orMatrixOutputs_hi_hi_lo_hi_4, decodeResult_andMatrixOutputs_71_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_hi_hi_12 = {decodeResult_orMatrixOutputs_hi_hi_hi_hi_8, decodeResult_orMatrixOutputs_hi_hi_hi_lo_4};
  wire [6:0]  decodeResult_orMatrixOutputs_hi_hi_21 = {decodeResult_orMatrixOutputs_hi_hi_hi_12, decodeResult_orMatrixOutputs_hi_hi_lo_10};
  wire [13:0] decodeResult_orMatrixOutputs_hi_25 = {decodeResult_orMatrixOutputs_hi_hi_21, decodeResult_orMatrixOutputs_hi_lo_14};
  wire [1:0]  _decodeResult_orMatrixOutputs_T_62 = {decodeResult_andMatrixOutputs_104_2, decodeResult_andMatrixOutputs_88_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_13;
  assign decodeResult_orMatrixOutputs_lo_lo_13 = _decodeResult_orMatrixOutputs_T_62;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_lo_lo_2;
  assign decodeResult_orMatrixOutputs_lo_lo_lo_lo_2 = _decodeResult_orMatrixOutputs_T_62;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_23 = {decodeResult_andMatrixOutputs_143_2, decodeResult_andMatrixOutputs_85_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_22 = {decodeResult_andMatrixOutputs_140_2, decodeResult_andMatrixOutputs_129_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_26 = {decodeResult_orMatrixOutputs_hi_hi_22, decodeResult_andMatrixOutputs_65_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_17 = {decodeResult_andMatrixOutputs_33_2, decodeResult_andMatrixOutputs_103_2};
  wire [3:0]  decodeResult_orMatrixOutputs_lo_24 = {decodeResult_orMatrixOutputs_lo_hi_17, decodeResult_orMatrixOutputs_lo_lo_13};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_15 = {decodeResult_andMatrixOutputs_63_2, decodeResult_andMatrixOutputs_144_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_23 = {decodeResult_andMatrixOutputs_96_2, decodeResult_andMatrixOutputs_21_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_27 = {decodeResult_orMatrixOutputs_hi_hi_23, decodeResult_orMatrixOutputs_hi_lo_15};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_lo_lo_hi = {decodeResult_andMatrixOutputs_95_2, decodeResult_andMatrixOutputs_104_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_lo_lo_lo_1 = {decodeResult_orMatrixOutputs_lo_lo_lo_lo_hi, decodeResult_andMatrixOutputs_88_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_lo_hi_hi = {decodeResult_andMatrixOutputs_72_2, decodeResult_andMatrixOutputs_41_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_lo_lo_hi_5 = {decodeResult_orMatrixOutputs_lo_lo_lo_hi_hi, decodeResult_andMatrixOutputs_28_2};
  wire [5:0]  decodeResult_orMatrixOutputs_lo_lo_lo_10 = {decodeResult_orMatrixOutputs_lo_lo_lo_hi_5, decodeResult_orMatrixOutputs_lo_lo_lo_lo_1};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_lo_hi = {decodeResult_andMatrixOutputs_109_2, decodeResult_andMatrixOutputs_124_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_lo_hi_lo_4 = {decodeResult_orMatrixOutputs_lo_lo_hi_lo_hi, decodeResult_andMatrixOutputs_5_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_hi_lo = {decodeResult_andMatrixOutputs_31_2, decodeResult_andMatrixOutputs_81_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_hi_hi = {decodeResult_andMatrixOutputs_51_2, decodeResult_andMatrixOutputs_38_2};
  wire [3:0]  decodeResult_orMatrixOutputs_lo_lo_hi_hi_5 = {decodeResult_orMatrixOutputs_lo_lo_hi_hi_hi, decodeResult_orMatrixOutputs_lo_lo_hi_hi_lo};
  wire [6:0]  decodeResult_orMatrixOutputs_lo_lo_hi_11 = {decodeResult_orMatrixOutputs_lo_lo_hi_hi_5, decodeResult_orMatrixOutputs_lo_lo_hi_lo_4};
  wire [12:0] decodeResult_orMatrixOutputs_lo_lo_14 = {decodeResult_orMatrixOutputs_lo_lo_hi_11, decodeResult_orMatrixOutputs_lo_lo_lo_10};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_lo_lo_hi = {decodeResult_andMatrixOutputs_125_2, decodeResult_andMatrixOutputs_27_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_lo_lo_1 = {decodeResult_orMatrixOutputs_lo_hi_lo_lo_hi, decodeResult_andMatrixOutputs_105_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_lo_hi_hi = {decodeResult_andMatrixOutputs_80_2, decodeResult_andMatrixOutputs_132_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_lo_hi_5 = {decodeResult_orMatrixOutputs_lo_hi_lo_hi_hi, decodeResult_andMatrixOutputs_122_2};
  wire [5:0]  decodeResult_orMatrixOutputs_lo_hi_lo_10 = {decodeResult_orMatrixOutputs_lo_hi_lo_hi_5, decodeResult_orMatrixOutputs_lo_hi_lo_lo_1};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_lo_hi = {decodeResult_andMatrixOutputs_36_2, decodeResult_andMatrixOutputs_60_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_hi_lo_4 = {decodeResult_orMatrixOutputs_lo_hi_hi_lo_hi, decodeResult_andMatrixOutputs_39_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_hi_lo = {decodeResult_andMatrixOutputs_98_2, decodeResult_andMatrixOutputs_19_2};
  wire [3:0]  decodeResult_orMatrixOutputs_lo_hi_hi_hi_8 = {decodeResult_orMatrixOutputs_lo_hi_hi_hi_hi_1, decodeResult_orMatrixOutputs_lo_hi_hi_hi_lo};
  wire [6:0]  decodeResult_orMatrixOutputs_lo_hi_hi_12 = {decodeResult_orMatrixOutputs_lo_hi_hi_hi_8, decodeResult_orMatrixOutputs_lo_hi_hi_lo_4};
  wire [12:0] decodeResult_orMatrixOutputs_lo_hi_18 = {decodeResult_orMatrixOutputs_lo_hi_hi_12, decodeResult_orMatrixOutputs_lo_hi_lo_10};
  wire [25:0] decodeResult_orMatrixOutputs_lo_25 = {decodeResult_orMatrixOutputs_lo_hi_18, decodeResult_orMatrixOutputs_lo_lo_14};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_lo_lo_hi = {decodeResult_andMatrixOutputs_55_2, decodeResult_andMatrixOutputs_106_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_lo_lo_lo_1 = {decodeResult_orMatrixOutputs_hi_lo_lo_lo_hi, decodeResult_andMatrixOutputs_90_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_lo_hi_hi = {decodeResult_andMatrixOutputs_130_2, decodeResult_andMatrixOutputs_57_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_lo_lo_hi_5 = {decodeResult_orMatrixOutputs_hi_lo_lo_hi_hi, decodeResult_andMatrixOutputs_18_2};
  wire [5:0]  decodeResult_orMatrixOutputs_hi_lo_lo_10 = {decodeResult_orMatrixOutputs_hi_lo_lo_hi_5, decodeResult_orMatrixOutputs_hi_lo_lo_lo_1};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_lo_hi = {decodeResult_andMatrixOutputs_75_2, decodeResult_andMatrixOutputs_68_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_lo_hi_lo_4 = {decodeResult_orMatrixOutputs_hi_lo_hi_lo_hi, decodeResult_andMatrixOutputs_73_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_hi_hi = {decodeResult_andMatrixOutputs_40_2, decodeResult_andMatrixOutputs_107_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_lo_hi_hi_7 = {decodeResult_orMatrixOutputs_hi_lo_hi_hi_hi, decodeResult_orMatrixOutputs_hi_lo_hi_hi_lo};
  wire [6:0]  decodeResult_orMatrixOutputs_hi_lo_hi_11 = {decodeResult_orMatrixOutputs_hi_lo_hi_hi_7, decodeResult_orMatrixOutputs_hi_lo_hi_lo_4};
  wire [12:0] decodeResult_orMatrixOutputs_hi_lo_16 = {decodeResult_orMatrixOutputs_hi_lo_hi_11, decodeResult_orMatrixOutputs_hi_lo_lo_10};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_hi_lo_lo_3 = {decodeResult_orMatrixOutputs_hi_hi_lo_lo_hi, decodeResult_andMatrixOutputs_53_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_hi_lo = {decodeResult_andMatrixOutputs_25_2, decodeResult_andMatrixOutputs_45_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_hi_hi = {decodeResult_andMatrixOutputs_138_2, decodeResult_andMatrixOutputs_30_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_hi_lo_hi_5 = {decodeResult_orMatrixOutputs_hi_hi_lo_hi_hi, decodeResult_orMatrixOutputs_hi_hi_lo_hi_lo};
  wire [6:0]  decodeResult_orMatrixOutputs_hi_hi_lo_11 = {decodeResult_orMatrixOutputs_hi_hi_lo_hi_5, decodeResult_orMatrixOutputs_hi_hi_lo_lo_3};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_hi_hi_lo_5 = {decodeResult_orMatrixOutputs_hi_hi_hi_lo_hi, decodeResult_andMatrixOutputs_50_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_hi_lo = {decodeResult_andMatrixOutputs_93_2, decodeResult_andMatrixOutputs_74_2};
  wire [1:0]  _GEN_28 = {decodeResult_andMatrixOutputs_15_2, decodeResult_andMatrixOutputs_110_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_hi_hi_1;
  assign decodeResult_orMatrixOutputs_hi_hi_hi_hi_hi_1 = _GEN_28;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_hi_hi_2;
  assign decodeResult_orMatrixOutputs_hi_hi_hi_hi_hi_2 = _GEN_28;
  wire [3:0]  decodeResult_orMatrixOutputs_hi_hi_hi_hi_9 = {decodeResult_orMatrixOutputs_hi_hi_hi_hi_hi_1, decodeResult_orMatrixOutputs_hi_hi_hi_hi_lo};
  wire [6:0]  decodeResult_orMatrixOutputs_hi_hi_hi_13 = {decodeResult_orMatrixOutputs_hi_hi_hi_hi_9, decodeResult_orMatrixOutputs_hi_hi_hi_lo_5};
  wire [13:0] decodeResult_orMatrixOutputs_hi_hi_24 = {decodeResult_orMatrixOutputs_hi_hi_hi_13, decodeResult_orMatrixOutputs_hi_hi_lo_11};
  wire [26:0] decodeResult_orMatrixOutputs_hi_28 = {decodeResult_orMatrixOutputs_hi_hi_24, decodeResult_orMatrixOutputs_hi_lo_16};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_lo_hi_hi_1 = {decodeResult_andMatrixOutputs_41_2, decodeResult_andMatrixOutputs_116_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_lo_lo_hi_6 = {decodeResult_orMatrixOutputs_lo_lo_lo_hi_hi_1, decodeResult_andMatrixOutputs_139_2};
  wire [4:0]  decodeResult_orMatrixOutputs_lo_lo_lo_11 = {decodeResult_orMatrixOutputs_lo_lo_lo_hi_6, decodeResult_orMatrixOutputs_lo_lo_lo_lo_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_lo_hi_1 = {decodeResult_andMatrixOutputs_111_2, decodeResult_andMatrixOutputs_37_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_lo_hi_lo_5 = {decodeResult_orMatrixOutputs_lo_lo_hi_lo_hi_1, decodeResult_andMatrixOutputs_52_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_hi_hi_1 = {decodeResult_andMatrixOutputs_42_2, decodeResult_andMatrixOutputs_124_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_lo_hi_hi_6 = {decodeResult_orMatrixOutputs_lo_lo_hi_hi_hi_1, decodeResult_andMatrixOutputs_5_2};
  wire [5:0]  decodeResult_orMatrixOutputs_lo_lo_hi_12 = {decodeResult_orMatrixOutputs_lo_lo_hi_hi_6, decodeResult_orMatrixOutputs_lo_lo_hi_lo_5};
  wire [10:0] decodeResult_orMatrixOutputs_lo_lo_15 = {decodeResult_orMatrixOutputs_lo_lo_hi_12, decodeResult_orMatrixOutputs_lo_lo_lo_11};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_lo_lo_hi_1 = {decodeResult_andMatrixOutputs_38_2, decodeResult_andMatrixOutputs_31_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_lo_lo_2 = {decodeResult_orMatrixOutputs_lo_hi_lo_lo_hi_1, decodeResult_andMatrixOutputs_81_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_lo_hi_hi_1 = {decodeResult_andMatrixOutputs_27_2, decodeResult_andMatrixOutputs_105_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_lo_hi_6 = {decodeResult_orMatrixOutputs_lo_hi_lo_hi_hi_1, decodeResult_andMatrixOutputs_51_2};
  wire [5:0]  decodeResult_orMatrixOutputs_lo_hi_lo_11 = {decodeResult_orMatrixOutputs_lo_hi_lo_hi_6, decodeResult_orMatrixOutputs_lo_hi_lo_lo_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_lo_hi_1 = {decodeResult_andMatrixOutputs_29_2, decodeResult_andMatrixOutputs_127_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_hi_lo_5 = {decodeResult_orMatrixOutputs_lo_hi_hi_lo_hi_1, decodeResult_andMatrixOutputs_119_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_hi_hi_2 = {decodeResult_andMatrixOutputs_101_2, decodeResult_andMatrixOutputs_39_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_hi_hi_9 = {decodeResult_orMatrixOutputs_lo_hi_hi_hi_hi_2, decodeResult_andMatrixOutputs_80_2};
  wire [5:0]  decodeResult_orMatrixOutputs_lo_hi_hi_13 = {decodeResult_orMatrixOutputs_lo_hi_hi_hi_9, decodeResult_orMatrixOutputs_lo_hi_hi_lo_5};
  wire [11:0] decodeResult_orMatrixOutputs_lo_hi_19 = {decodeResult_orMatrixOutputs_lo_hi_hi_13, decodeResult_orMatrixOutputs_lo_hi_lo_11};
  wire [22:0] decodeResult_orMatrixOutputs_lo_26 = {decodeResult_orMatrixOutputs_lo_hi_19, decodeResult_orMatrixOutputs_lo_lo_15};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_lo_lo_2 = {decodeResult_andMatrixOutputs_13_2, decodeResult_andMatrixOutputs_46_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_lo_hi_hi_1 = {decodeResult_andMatrixOutputs_133_2, decodeResult_andMatrixOutputs_63_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_lo_lo_hi_6 = {decodeResult_orMatrixOutputs_hi_lo_lo_hi_hi_1, decodeResult_andMatrixOutputs_67_2};
  wire [4:0]  decodeResult_orMatrixOutputs_hi_lo_lo_11 = {decodeResult_orMatrixOutputs_hi_lo_lo_hi_6, decodeResult_orMatrixOutputs_hi_lo_lo_lo_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_lo_hi_1 = {decodeResult_andMatrixOutputs_57_2, decodeResult_andMatrixOutputs_55_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_lo_hi_lo_5 = {decodeResult_orMatrixOutputs_hi_lo_hi_lo_hi_1, decodeResult_andMatrixOutputs_106_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_hi_hi_1 = {decodeResult_andMatrixOutputs_68_2, decodeResult_andMatrixOutputs_73_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_lo_hi_hi_8 = {decodeResult_orMatrixOutputs_hi_lo_hi_hi_hi_1, decodeResult_andMatrixOutputs_130_2};
  wire [5:0]  decodeResult_orMatrixOutputs_hi_lo_hi_12 = {decodeResult_orMatrixOutputs_hi_lo_hi_hi_8, decodeResult_orMatrixOutputs_hi_lo_hi_lo_5};
  wire [10:0] decodeResult_orMatrixOutputs_hi_lo_17 = {decodeResult_orMatrixOutputs_hi_lo_hi_12, decodeResult_orMatrixOutputs_hi_lo_lo_11};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_hi_lo_lo_4 = {decodeResult_orMatrixOutputs_hi_hi_lo_lo_hi_1, decodeResult_andMatrixOutputs_75_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_hi_hi_1 = {decodeResult_andMatrixOutputs_58_2, decodeResult_andMatrixOutputs_128_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_hi_lo_hi_6 = {decodeResult_orMatrixOutputs_hi_hi_lo_hi_hi_1, decodeResult_andMatrixOutputs_83_2};
  wire [5:0]  decodeResult_orMatrixOutputs_hi_hi_lo_12 = {decodeResult_orMatrixOutputs_hi_hi_lo_hi_6, decodeResult_orMatrixOutputs_hi_hi_lo_lo_4};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_lo_hi_1 = {decodeResult_andMatrixOutputs_6_2, decodeResult_andMatrixOutputs_138_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_hi_hi_lo_6 = {decodeResult_orMatrixOutputs_hi_hi_hi_lo_hi_1, decodeResult_andMatrixOutputs_25_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_hi_hi_hi_10 = {decodeResult_orMatrixOutputs_hi_hi_hi_hi_hi_2, decodeResult_andMatrixOutputs_74_2};
  wire [5:0]  decodeResult_orMatrixOutputs_hi_hi_hi_14 = {decodeResult_orMatrixOutputs_hi_hi_hi_hi_10, decodeResult_orMatrixOutputs_hi_hi_hi_lo_6};
  wire [11:0] decodeResult_orMatrixOutputs_hi_hi_25 = {decodeResult_orMatrixOutputs_hi_hi_hi_14, decodeResult_orMatrixOutputs_hi_hi_lo_12};
  wire [22:0] decodeResult_orMatrixOutputs_hi_29 = {decodeResult_orMatrixOutputs_hi_hi_25, decodeResult_orMatrixOutputs_hi_lo_17};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_20 = {decodeResult_andMatrixOutputs_36_2, decodeResult_andMatrixOutputs_113_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_27 = {decodeResult_orMatrixOutputs_lo_hi_20, decodeResult_andMatrixOutputs_132_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_26 = {decodeResult_andMatrixOutputs_96_2, decodeResult_andMatrixOutputs_56_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_30 = {decodeResult_orMatrixOutputs_hi_hi_26, decodeResult_orMatrixOutputs_hi_lo_18};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_16 = {decodeResult_andMatrixOutputs_103_2, decodeResult_andMatrixOutputs_126_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_14 = {decodeResult_andMatrixOutputs_144_2, decodeResult_andMatrixOutputs_61_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_21 = {decodeResult_orMatrixOutputs_lo_hi_hi_14, decodeResult_andMatrixOutputs_132_2};
  wire [4:0]  decodeResult_orMatrixOutputs_lo_28 = {decodeResult_orMatrixOutputs_lo_hi_21, decodeResult_orMatrixOutputs_lo_lo_16};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_15 = {decodeResult_andMatrixOutputs_0_2, decodeResult_andMatrixOutputs_53_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_hi_27 = {decodeResult_orMatrixOutputs_hi_hi_hi_15, decodeResult_andMatrixOutputs_69_2};
  wire [4:0]  decodeResult_orMatrixOutputs_hi_31 = {decodeResult_orMatrixOutputs_hi_hi_27, decodeResult_orMatrixOutputs_hi_lo_19};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_13 = {decodeResult_andMatrixOutputs_36_2, decodeResult_andMatrixOutputs_147_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_lo_17 = {decodeResult_orMatrixOutputs_lo_lo_hi_13, decodeResult_andMatrixOutputs_1_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_15 = {decodeResult_andMatrixOutputs_121_2, decodeResult_andMatrixOutputs_144_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_22 = {decodeResult_orMatrixOutputs_lo_hi_hi_15, decodeResult_andMatrixOutputs_67_2};
  wire [5:0]  decodeResult_orMatrixOutputs_lo_29 = {decodeResult_orMatrixOutputs_lo_hi_22, decodeResult_orMatrixOutputs_lo_lo_17};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_13 = {decodeResult_andMatrixOutputs_53_2, decodeResult_andMatrixOutputs_4_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_lo_20 = {decodeResult_orMatrixOutputs_hi_lo_hi_13, decodeResult_andMatrixOutputs_21_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_hi_28 = {decodeResult_orMatrixOutputs_hi_hi_hi_16, decodeResult_andMatrixOutputs_149_2};
  wire [5:0]  decodeResult_orMatrixOutputs_hi_32 = {decodeResult_orMatrixOutputs_hi_hi_28, decodeResult_orMatrixOutputs_hi_lo_20};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_23 = {decodeResult_andMatrixOutputs_17_2, decodeResult_andMatrixOutputs_147_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_30 = {decodeResult_orMatrixOutputs_lo_hi_23, decodeResult_andMatrixOutputs_1_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_21 = {decodeResult_andMatrixOutputs_144_2, decodeResult_andMatrixOutputs_19_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_29 = {decodeResult_andMatrixOutputs_114_2, decodeResult_andMatrixOutputs_18_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_33 = {decodeResult_orMatrixOutputs_hi_hi_29, decodeResult_orMatrixOutputs_hi_lo_21};
  wire [1:0]  _GEN_29 = {decodeResult_andMatrixOutputs_49_2, decodeResult_andMatrixOutputs_47_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_14;
  assign decodeResult_orMatrixOutputs_lo_lo_hi_14 = _GEN_29;
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_lo_13;
  assign decodeResult_orMatrixOutputs_lo_hi_lo_13 = _GEN_29;
  wire [3:0]  decodeResult_orMatrixOutputs_lo_lo_18 = {decodeResult_orMatrixOutputs_lo_lo_hi_14, decodeResult_orMatrixOutputs_lo_lo_lo_12};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_lo_12 = {decodeResult_andMatrixOutputs_60_2, decodeResult_andMatrixOutputs_132_2};
  wire [3:0]  decodeResult_orMatrixOutputs_lo_hi_24 = {decodeResult_orMatrixOutputs_lo_hi_hi_16, decodeResult_orMatrixOutputs_lo_hi_lo_12};
  wire [7:0]  decodeResult_orMatrixOutputs_lo_31 = {decodeResult_orMatrixOutputs_lo_hi_24, decodeResult_orMatrixOutputs_lo_lo_18};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_lo_22 = {decodeResult_orMatrixOutputs_hi_lo_hi_14, decodeResult_orMatrixOutputs_hi_lo_lo_12};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_13 = {decodeResult_andMatrixOutputs_144_2, decodeResult_andMatrixOutputs_67_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_hi_30 = {decodeResult_orMatrixOutputs_hi_hi_hi_17, decodeResult_orMatrixOutputs_hi_hi_lo_13};
  wire [7:0]  decodeResult_orMatrixOutputs_hi_34 = {decodeResult_orMatrixOutputs_hi_hi_30, decodeResult_orMatrixOutputs_hi_lo_22};
  wire [3:0]  decodeResult_orMatrixOutputs_lo_lo_19 = {decodeResult_orMatrixOutputs_lo_lo_hi_15, decodeResult_orMatrixOutputs_lo_lo_lo_13};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_hi_17 = {decodeResult_orMatrixOutputs_lo_hi_hi_hi_10, decodeResult_andMatrixOutputs_60_2};
  wire [4:0]  decodeResult_orMatrixOutputs_lo_hi_25 = {decodeResult_orMatrixOutputs_lo_hi_hi_17, decodeResult_orMatrixOutputs_lo_hi_lo_13};
  wire [8:0]  decodeResult_orMatrixOutputs_lo_32 = {decodeResult_orMatrixOutputs_lo_hi_25, decodeResult_orMatrixOutputs_lo_lo_19};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_lo_23 = {decodeResult_orMatrixOutputs_hi_lo_hi_15, decodeResult_orMatrixOutputs_hi_lo_lo_13};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_hi_hi_18 = {decodeResult_orMatrixOutputs_hi_hi_hi_hi_11, decodeResult_andMatrixOutputs_22_2};
  wire [4:0]  decodeResult_orMatrixOutputs_hi_hi_31 = {decodeResult_orMatrixOutputs_hi_hi_hi_18, decodeResult_orMatrixOutputs_hi_hi_lo_14};
  wire [8:0]  decodeResult_orMatrixOutputs_hi_35 = {decodeResult_orMatrixOutputs_hi_hi_31, decodeResult_orMatrixOutputs_hi_lo_23};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_lo_14 = {decodeResult_andMatrixOutputs_143_2, decodeResult_andMatrixOutputs_88_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_hi_7 = {decodeResult_andMatrixOutputs_129_2, decodeResult_andMatrixOutputs_65_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_lo_hi_16 = {decodeResult_orMatrixOutputs_lo_lo_hi_hi_7, decodeResult_andMatrixOutputs_104_2};
  wire [4:0]  decodeResult_orMatrixOutputs_lo_lo_20 = {decodeResult_orMatrixOutputs_lo_lo_hi_16, decodeResult_orMatrixOutputs_lo_lo_lo_14};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_lo_hi_7 = {decodeResult_andMatrixOutputs_127_2, decodeResult_andMatrixOutputs_122_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_lo_14 = {decodeResult_orMatrixOutputs_lo_hi_lo_hi_7, decodeResult_andMatrixOutputs_125_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_hi_11 = {decodeResult_andMatrixOutputs_29_2, decodeResult_andMatrixOutputs_49_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_hi_18 = {decodeResult_orMatrixOutputs_lo_hi_hi_hi_11, decodeResult_andMatrixOutputs_47_2};
  wire [5:0]  decodeResult_orMatrixOutputs_lo_hi_26 = {decodeResult_orMatrixOutputs_lo_hi_hi_18, decodeResult_orMatrixOutputs_lo_hi_lo_14};
  wire [10:0] decodeResult_orMatrixOutputs_lo_33 = {decodeResult_orMatrixOutputs_lo_hi_26, decodeResult_orMatrixOutputs_lo_lo_20};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_hi_9 = {decodeResult_andMatrixOutputs_98_2, decodeResult_andMatrixOutputs_113_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_lo_hi_16 = {decodeResult_orMatrixOutputs_hi_lo_hi_hi_9, decodeResult_andMatrixOutputs_147_2};
  wire [4:0]  decodeResult_orMatrixOutputs_hi_lo_24 = {decodeResult_orMatrixOutputs_hi_lo_hi_16, decodeResult_orMatrixOutputs_hi_lo_lo_14};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_hi_7 = {decodeResult_andMatrixOutputs_140_2, decodeResult_andMatrixOutputs_33_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_hi_lo_15 = {decodeResult_orMatrixOutputs_hi_hi_lo_hi_7, decodeResult_andMatrixOutputs_14_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_hi_hi_19 = {decodeResult_orMatrixOutputs_hi_hi_hi_hi_12, decodeResult_andMatrixOutputs_144_2};
  wire [5:0]  decodeResult_orMatrixOutputs_hi_hi_32 = {decodeResult_orMatrixOutputs_hi_hi_hi_19, decodeResult_orMatrixOutputs_hi_hi_lo_15};
  wire [10:0] decodeResult_orMatrixOutputs_hi_36 = {decodeResult_orMatrixOutputs_hi_hi_32, decodeResult_orMatrixOutputs_hi_lo_24};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_17 = {decodeResult_andMatrixOutputs_42_2, decodeResult_andMatrixOutputs_111_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_lo_21 = {decodeResult_orMatrixOutputs_lo_lo_hi_17, decodeResult_andMatrixOutputs_139_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_19 = {decodeResult_andMatrixOutputs_101_2, decodeResult_andMatrixOutputs_47_2};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_27 = {decodeResult_orMatrixOutputs_lo_hi_hi_19, decodeResult_andMatrixOutputs_1_2};
  wire [5:0]  decodeResult_orMatrixOutputs_lo_34 = {decodeResult_orMatrixOutputs_lo_hi_27, decodeResult_orMatrixOutputs_lo_lo_21};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_17 = {decodeResult_andMatrixOutputs_68_2, decodeResult_andMatrixOutputs_133_2};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_lo_25 = {decodeResult_orMatrixOutputs_hi_lo_hi_17, decodeResult_andMatrixOutputs_46_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_16 = {decodeResult_andMatrixOutputs_138_2, decodeResult_andMatrixOutputs_53_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_hi_33 = {decodeResult_orMatrixOutputs_hi_hi_hi_20, decodeResult_orMatrixOutputs_hi_hi_lo_16};
  wire [6:0]  decodeResult_orMatrixOutputs_hi_37 = {decodeResult_orMatrixOutputs_hi_hi_33, decodeResult_orMatrixOutputs_hi_lo_25};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_35 = {decodeResult_andMatrixOutputs_101_2, decodeResult_andMatrixOutputs_142_2};
  wire [1:0]  _GEN_30 = {decodeResult_andMatrixOutputs_68_2, decodeResult_andMatrixOutputs_136_2};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_34;
  assign decodeResult_orMatrixOutputs_hi_hi_34 = _GEN_30;
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_26;
  assign decodeResult_orMatrixOutputs_hi_lo_26 = _GEN_30;
  wire [2:0]  decodeResult_orMatrixOutputs_hi_38 = {decodeResult_orMatrixOutputs_hi_hi_34, decodeResult_andMatrixOutputs_46_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_22 = {decodeResult_andMatrixOutputs_142_2, decodeResult_andMatrixOutputs_47_2};
  wire [3:0]  decodeResult_orMatrixOutputs_lo_36 = {decodeResult_orMatrixOutputs_lo_hi_28, decodeResult_orMatrixOutputs_lo_lo_22};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_35 = {decodeResult_andMatrixOutputs_10_2, decodeResult_andMatrixOutputs_53_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_39 = {decodeResult_orMatrixOutputs_hi_hi_35, decodeResult_orMatrixOutputs_hi_lo_26};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_lo_lo_hi_1 = {|{decodeResult_orMatrixOutputs_hi_2, decodeResult_orMatrixOutputs_lo_2}, |{decodeResult_orMatrixOutputs_hi_1, decodeResult_orMatrixOutputs_lo_1}};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_lo_lo_lo_3 = {decodeResult_orMatrixOutputs_lo_lo_lo_lo_hi_1, |{decodeResult_orMatrixOutputs_hi, decodeResult_orMatrixOutputs_lo}};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_lo_hi_lo = {|{decodeResult_orMatrixOutputs_hi_4, decodeResult_andMatrixOutputs_38_2}, |{decodeResult_orMatrixOutputs_hi_3, decodeResult_orMatrixOutputs_lo_3}};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_lo_hi_hi_2 = {|{decodeResult_orMatrixOutputs_hi_6, decodeResult_orMatrixOutputs_lo_5}, |{decodeResult_orMatrixOutputs_hi_5, decodeResult_orMatrixOutputs_lo_4}};
  wire [3:0]  decodeResult_orMatrixOutputs_lo_lo_lo_hi_7 = {decodeResult_orMatrixOutputs_lo_lo_lo_hi_hi_2, decodeResult_orMatrixOutputs_lo_lo_lo_hi_lo};
  wire [6:0]  decodeResult_orMatrixOutputs_lo_lo_lo_15 = {decodeResult_orMatrixOutputs_lo_lo_lo_hi_7, decodeResult_orMatrixOutputs_lo_lo_lo_lo_3};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_lo_hi_2 = {|{decodeResult_orMatrixOutputs_hi_9, decodeResult_orMatrixOutputs_lo_8}, |{decodeResult_orMatrixOutputs_hi_8, decodeResult_orMatrixOutputs_lo_7}};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_lo_hi_lo_6 = {decodeResult_orMatrixOutputs_lo_lo_hi_lo_hi_2, |{decodeResult_orMatrixOutputs_hi_7, decodeResult_orMatrixOutputs_lo_6}};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_hi_lo_1 = {|{decodeResult_orMatrixOutputs_hi_10, decodeResult_orMatrixOutputs_lo_9}, decodeResult_andMatrixOutputs_56_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_lo_hi_hi_hi_2 = {|{decodeResult_orMatrixOutputs_hi_11, decodeResult_orMatrixOutputs_lo_10}, decodeResult_andMatrixOutputs_103_2};
  wire [3:0]  decodeResult_orMatrixOutputs_lo_lo_hi_hi_8 = {decodeResult_orMatrixOutputs_lo_lo_hi_hi_hi_2, decodeResult_orMatrixOutputs_lo_lo_hi_hi_lo_1};
  wire [6:0]  decodeResult_orMatrixOutputs_lo_lo_hi_18 = {decodeResult_orMatrixOutputs_lo_lo_hi_hi_8, decodeResult_orMatrixOutputs_lo_lo_hi_lo_6};
  wire [13:0] decodeResult_orMatrixOutputs_lo_lo_23 = {decodeResult_orMatrixOutputs_lo_lo_hi_18, decodeResult_orMatrixOutputs_lo_lo_lo_15};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_lo_lo_hi_2 = {decodeResult_andMatrixOutputs_108_2, |{decodeResult_orMatrixOutputs_hi_12, decodeResult_andMatrixOutputs_55_2}};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_lo_lo_3 = {decodeResult_orMatrixOutputs_lo_hi_lo_lo_hi_2, |{decodeResult_andMatrixOutputs_71_2, decodeResult_andMatrixOutputs_106_2}};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_lo_hi_lo = {|{decodeResult_orMatrixOutputs_hi_13, decodeResult_orMatrixOutputs_lo_11}, decodeResult_andMatrixOutputs_132_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_lo_hi_hi_2 = {|{decodeResult_orMatrixOutputs_hi_14, decodeResult_andMatrixOutputs_67_2}, |_decodeResult_orMatrixOutputs_T_34};
  wire [3:0]  decodeResult_orMatrixOutputs_lo_hi_lo_hi_8 = {decodeResult_orMatrixOutputs_lo_hi_lo_hi_hi_2, decodeResult_orMatrixOutputs_lo_hi_lo_hi_lo};
  wire [6:0]  decodeResult_orMatrixOutputs_lo_hi_lo_15 = {decodeResult_orMatrixOutputs_lo_hi_lo_hi_8, decodeResult_orMatrixOutputs_lo_hi_lo_lo_3};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_lo_hi_2 = {|{decodeResult_orMatrixOutputs_hi_16, decodeResult_orMatrixOutputs_lo_13}, |{decodeResult_orMatrixOutputs_hi_15, decodeResult_orMatrixOutputs_lo_12}};
  wire [2:0]  decodeResult_orMatrixOutputs_lo_hi_hi_lo_6 = {decodeResult_orMatrixOutputs_lo_hi_hi_lo_hi_2, decodeResult_andMatrixOutputs_113_2};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_hi_lo_1 = {|{decodeResult_orMatrixOutputs_hi_18, decodeResult_orMatrixOutputs_lo_15}, |{decodeResult_orMatrixOutputs_hi_17, decodeResult_orMatrixOutputs_lo_14}};
  wire [1:0]  decodeResult_orMatrixOutputs_lo_hi_hi_hi_hi_3 = {|{decodeResult_orMatrixOutputs_hi_20, decodeResult_orMatrixOutputs_lo_17}, |{decodeResult_orMatrixOutputs_hi_19, decodeResult_orMatrixOutputs_lo_16}};
  wire [3:0]  decodeResult_orMatrixOutputs_lo_hi_hi_hi_12 = {decodeResult_orMatrixOutputs_lo_hi_hi_hi_hi_3, decodeResult_orMatrixOutputs_lo_hi_hi_hi_lo_1};
  wire [6:0]  decodeResult_orMatrixOutputs_lo_hi_hi_20 = {decodeResult_orMatrixOutputs_lo_hi_hi_hi_12, decodeResult_orMatrixOutputs_lo_hi_hi_lo_6};
  wire [13:0] decodeResult_orMatrixOutputs_lo_hi_29 = {decodeResult_orMatrixOutputs_lo_hi_hi_20, decodeResult_orMatrixOutputs_lo_hi_lo_15};
  wire [27:0] decodeResult_orMatrixOutputs_lo_37 = {decodeResult_orMatrixOutputs_lo_hi_29, decodeResult_orMatrixOutputs_lo_lo_23};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_lo_lo_hi_1 = {decodeResult_andMatrixOutputs_85_2, |{decodeResult_orMatrixOutputs_hi_22, decodeResult_orMatrixOutputs_lo_19}};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_lo_lo_lo_3 = {decodeResult_orMatrixOutputs_hi_lo_lo_lo_hi_1, |{decodeResult_orMatrixOutputs_hi_21, decodeResult_orMatrixOutputs_lo_18}};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_lo_hi_lo = {|{decodeResult_orMatrixOutputs_hi_24, decodeResult_orMatrixOutputs_lo_21}, |{decodeResult_orMatrixOutputs_hi_23, decodeResult_orMatrixOutputs_lo_20}};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_lo_hi_hi_2 = {|_decodeResult_orMatrixOutputs_T_62, |{decodeResult_orMatrixOutputs_hi_25, decodeResult_orMatrixOutputs_lo_22}};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_lo_lo_hi_7 = {decodeResult_orMatrixOutputs_hi_lo_lo_hi_hi_2, decodeResult_orMatrixOutputs_hi_lo_lo_hi_lo};
  wire [6:0]  decodeResult_orMatrixOutputs_hi_lo_lo_15 = {decodeResult_orMatrixOutputs_hi_lo_lo_hi_7, decodeResult_orMatrixOutputs_hi_lo_lo_lo_3};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_lo_hi_2 = {|{decodeResult_andMatrixOutputs_62_2, decodeResult_andMatrixOutputs_89_2}, |{decodeResult_orMatrixOutputs_hi_27, decodeResult_orMatrixOutputs_lo_24}};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_lo_hi_lo_6 = {decodeResult_orMatrixOutputs_hi_lo_hi_lo_hi_2, |{decodeResult_orMatrixOutputs_hi_26, decodeResult_orMatrixOutputs_lo_23}};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_hi_lo_1 = {|{decodeResult_orMatrixOutputs_hi_29, decodeResult_orMatrixOutputs_lo_26}, |{decodeResult_orMatrixOutputs_hi_28, decodeResult_orMatrixOutputs_lo_25}};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_lo_hi_hi_hi_2 = {|{decodeResult_andMatrixOutputs_6_2, decodeResult_andMatrixOutputs_25_2}, |{decodeResult_orMatrixOutputs_hi_30, decodeResult_orMatrixOutputs_lo_27}};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_lo_hi_hi_10 = {decodeResult_orMatrixOutputs_hi_lo_hi_hi_hi_2, decodeResult_orMatrixOutputs_hi_lo_hi_hi_lo_1};
  wire [6:0]  decodeResult_orMatrixOutputs_hi_lo_hi_18 = {decodeResult_orMatrixOutputs_hi_lo_hi_hi_10, decodeResult_orMatrixOutputs_hi_lo_hi_lo_6};
  wire [13:0] decodeResult_orMatrixOutputs_hi_lo_27 = {decodeResult_orMatrixOutputs_hi_lo_hi_18, decodeResult_orMatrixOutputs_hi_lo_lo_15};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_lo_hi_2 = {decodeResult_andMatrixOutputs_33_2, |{decodeResult_andMatrixOutputs_144_2, decodeResult_andMatrixOutputs_147_2}};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_hi_lo_lo_5 = {decodeResult_orMatrixOutputs_hi_hi_lo_lo_hi_2, |{decodeResult_andMatrixOutputs_73_2, decodeResult_andMatrixOutputs_57_2}};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_hi_lo_1 = {|{decodeResult_orMatrixOutputs_hi_32, decodeResult_orMatrixOutputs_lo_29}, |{decodeResult_orMatrixOutputs_hi_31, decodeResult_orMatrixOutputs_lo_28}};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_lo_hi_hi_2 = {|{decodeResult_orMatrixOutputs_hi_34, decodeResult_orMatrixOutputs_lo_31}, |{decodeResult_orMatrixOutputs_hi_33, decodeResult_orMatrixOutputs_lo_30}};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_hi_lo_hi_8 = {decodeResult_orMatrixOutputs_hi_hi_lo_hi_hi_2, decodeResult_orMatrixOutputs_hi_hi_lo_hi_lo_1};
  wire [6:0]  decodeResult_orMatrixOutputs_hi_hi_lo_17 = {decodeResult_orMatrixOutputs_hi_hi_lo_hi_8, decodeResult_orMatrixOutputs_hi_hi_lo_lo_5};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_lo_hi_2 = {|{decodeResult_orMatrixOutputs_hi_37, decodeResult_orMatrixOutputs_lo_34}, |{decodeResult_orMatrixOutputs_hi_36, decodeResult_orMatrixOutputs_lo_33}};
  wire [2:0]  decodeResult_orMatrixOutputs_hi_hi_hi_lo_7 = {decodeResult_orMatrixOutputs_hi_hi_hi_lo_hi_2, |{decodeResult_orMatrixOutputs_hi_35, decodeResult_orMatrixOutputs_lo_32}};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_hi_lo_1 = {|{decodeResult_orMatrixOutputs_hi_39, decodeResult_orMatrixOutputs_lo_36}, |{decodeResult_orMatrixOutputs_hi_38, decodeResult_orMatrixOutputs_lo_35}};
  wire [1:0]  decodeResult_orMatrixOutputs_hi_hi_hi_hi_hi_3 = {decodeResult_andMatrixOutputs_0_2, decodeResult_andMatrixOutputs_109_2};
  wire [3:0]  decodeResult_orMatrixOutputs_hi_hi_hi_hi_13 = {decodeResult_orMatrixOutputs_hi_hi_hi_hi_hi_3, decodeResult_orMatrixOutputs_hi_hi_hi_hi_lo_1};
  wire [6:0]  decodeResult_orMatrixOutputs_hi_hi_hi_21 = {decodeResult_orMatrixOutputs_hi_hi_hi_hi_13, decodeResult_orMatrixOutputs_hi_hi_hi_lo_7};
  wire [13:0] decodeResult_orMatrixOutputs_hi_hi_36 = {decodeResult_orMatrixOutputs_hi_hi_hi_21, decodeResult_orMatrixOutputs_hi_hi_lo_17};
  wire [27:0] decodeResult_orMatrixOutputs_hi_40 = {decodeResult_orMatrixOutputs_hi_hi_36, decodeResult_orMatrixOutputs_hi_lo_27};
  wire [55:0] decodeResult_orMatrixOutputs = {decodeResult_orMatrixOutputs_hi_40, decodeResult_orMatrixOutputs_lo_37};
  wire [1:0]  decodeResult_invMatrixOutputs_lo_lo_lo_lo_hi = decodeResult_orMatrixOutputs[2:1];
  wire [2:0]  decodeResult_invMatrixOutputs_lo_lo_lo_lo = {decodeResult_invMatrixOutputs_lo_lo_lo_lo_hi, decodeResult_orMatrixOutputs[0]};
  wire [1:0]  decodeResult_invMatrixOutputs_lo_lo_lo_hi_lo = decodeResult_orMatrixOutputs[4:3];
  wire [1:0]  decodeResult_invMatrixOutputs_lo_lo_lo_hi_hi = decodeResult_orMatrixOutputs[6:5];
  wire [3:0]  decodeResult_invMatrixOutputs_lo_lo_lo_hi = {decodeResult_invMatrixOutputs_lo_lo_lo_hi_hi, decodeResult_invMatrixOutputs_lo_lo_lo_hi_lo};
  wire [6:0]  decodeResult_invMatrixOutputs_lo_lo_lo = {decodeResult_invMatrixOutputs_lo_lo_lo_hi, decodeResult_invMatrixOutputs_lo_lo_lo_lo};
  wire [1:0]  decodeResult_invMatrixOutputs_lo_lo_hi_lo_hi = decodeResult_orMatrixOutputs[9:8];
  wire [2:0]  decodeResult_invMatrixOutputs_lo_lo_hi_lo = {decodeResult_invMatrixOutputs_lo_lo_hi_lo_hi, decodeResult_orMatrixOutputs[7]};
  wire [1:0]  decodeResult_invMatrixOutputs_lo_lo_hi_hi_lo = decodeResult_orMatrixOutputs[11:10];
  wire [1:0]  decodeResult_invMatrixOutputs_lo_lo_hi_hi_hi = decodeResult_orMatrixOutputs[13:12];
  wire [3:0]  decodeResult_invMatrixOutputs_lo_lo_hi_hi = {decodeResult_invMatrixOutputs_lo_lo_hi_hi_hi, decodeResult_invMatrixOutputs_lo_lo_hi_hi_lo};
  wire [6:0]  decodeResult_invMatrixOutputs_lo_lo_hi = {decodeResult_invMatrixOutputs_lo_lo_hi_hi, decodeResult_invMatrixOutputs_lo_lo_hi_lo};
  wire [13:0] decodeResult_invMatrixOutputs_lo_lo = {decodeResult_invMatrixOutputs_lo_lo_hi, decodeResult_invMatrixOutputs_lo_lo_lo};
  wire [1:0]  decodeResult_invMatrixOutputs_lo_hi_lo_lo_hi = decodeResult_orMatrixOutputs[16:15];
  wire [2:0]  decodeResult_invMatrixOutputs_lo_hi_lo_lo = {decodeResult_invMatrixOutputs_lo_hi_lo_lo_hi, decodeResult_orMatrixOutputs[14]};
  wire [1:0]  decodeResult_invMatrixOutputs_lo_hi_lo_hi_lo = decodeResult_orMatrixOutputs[18:17];
  wire [1:0]  decodeResult_invMatrixOutputs_lo_hi_lo_hi_hi = decodeResult_orMatrixOutputs[20:19];
  wire [3:0]  decodeResult_invMatrixOutputs_lo_hi_lo_hi = {decodeResult_invMatrixOutputs_lo_hi_lo_hi_hi, decodeResult_invMatrixOutputs_lo_hi_lo_hi_lo};
  wire [6:0]  decodeResult_invMatrixOutputs_lo_hi_lo = {decodeResult_invMatrixOutputs_lo_hi_lo_hi, decodeResult_invMatrixOutputs_lo_hi_lo_lo};
  wire [1:0]  decodeResult_invMatrixOutputs_lo_hi_hi_lo_hi = decodeResult_orMatrixOutputs[23:22];
  wire [2:0]  decodeResult_invMatrixOutputs_lo_hi_hi_lo = {decodeResult_invMatrixOutputs_lo_hi_hi_lo_hi, decodeResult_orMatrixOutputs[21]};
  wire [1:0]  decodeResult_invMatrixOutputs_lo_hi_hi_hi_lo = decodeResult_orMatrixOutputs[25:24];
  wire [1:0]  decodeResult_invMatrixOutputs_lo_hi_hi_hi_hi = decodeResult_orMatrixOutputs[27:26];
  wire [3:0]  decodeResult_invMatrixOutputs_lo_hi_hi_hi = {decodeResult_invMatrixOutputs_lo_hi_hi_hi_hi, decodeResult_invMatrixOutputs_lo_hi_hi_hi_lo};
  wire [6:0]  decodeResult_invMatrixOutputs_lo_hi_hi = {decodeResult_invMatrixOutputs_lo_hi_hi_hi, decodeResult_invMatrixOutputs_lo_hi_hi_lo};
  wire [13:0] decodeResult_invMatrixOutputs_lo_hi = {decodeResult_invMatrixOutputs_lo_hi_hi, decodeResult_invMatrixOutputs_lo_hi_lo};
  wire [27:0] decodeResult_invMatrixOutputs_lo = {decodeResult_invMatrixOutputs_lo_hi, decodeResult_invMatrixOutputs_lo_lo};
  wire [1:0]  decodeResult_invMatrixOutputs_hi_lo_lo_lo_hi = decodeResult_orMatrixOutputs[30:29];
  wire [2:0]  decodeResult_invMatrixOutputs_hi_lo_lo_lo = {decodeResult_invMatrixOutputs_hi_lo_lo_lo_hi, decodeResult_orMatrixOutputs[28]};
  wire [1:0]  decodeResult_invMatrixOutputs_hi_lo_lo_hi_lo = decodeResult_orMatrixOutputs[32:31];
  wire [1:0]  decodeResult_invMatrixOutputs_hi_lo_lo_hi_hi = decodeResult_orMatrixOutputs[34:33];
  wire [3:0]  decodeResult_invMatrixOutputs_hi_lo_lo_hi = {decodeResult_invMatrixOutputs_hi_lo_lo_hi_hi, decodeResult_invMatrixOutputs_hi_lo_lo_hi_lo};
  wire [6:0]  decodeResult_invMatrixOutputs_hi_lo_lo = {decodeResult_invMatrixOutputs_hi_lo_lo_hi, decodeResult_invMatrixOutputs_hi_lo_lo_lo};
  wire [1:0]  decodeResult_invMatrixOutputs_hi_lo_hi_lo_hi = decodeResult_orMatrixOutputs[37:36];
  wire [2:0]  decodeResult_invMatrixOutputs_hi_lo_hi_lo = {decodeResult_invMatrixOutputs_hi_lo_hi_lo_hi, decodeResult_orMatrixOutputs[35]};
  wire [1:0]  decodeResult_invMatrixOutputs_hi_lo_hi_hi_lo = decodeResult_orMatrixOutputs[39:38];
  wire [1:0]  decodeResult_invMatrixOutputs_hi_lo_hi_hi_hi = decodeResult_orMatrixOutputs[41:40];
  wire [3:0]  decodeResult_invMatrixOutputs_hi_lo_hi_hi = {decodeResult_invMatrixOutputs_hi_lo_hi_hi_hi, decodeResult_invMatrixOutputs_hi_lo_hi_hi_lo};
  wire [6:0]  decodeResult_invMatrixOutputs_hi_lo_hi = {decodeResult_invMatrixOutputs_hi_lo_hi_hi, decodeResult_invMatrixOutputs_hi_lo_hi_lo};
  wire [13:0] decodeResult_invMatrixOutputs_hi_lo = {decodeResult_invMatrixOutputs_hi_lo_hi, decodeResult_invMatrixOutputs_hi_lo_lo};
  wire [1:0]  decodeResult_invMatrixOutputs_hi_hi_lo_lo_hi = decodeResult_orMatrixOutputs[44:43];
  wire [2:0]  decodeResult_invMatrixOutputs_hi_hi_lo_lo = {decodeResult_invMatrixOutputs_hi_hi_lo_lo_hi, decodeResult_orMatrixOutputs[42]};
  wire [1:0]  decodeResult_invMatrixOutputs_hi_hi_lo_hi_lo = decodeResult_orMatrixOutputs[46:45];
  wire [1:0]  decodeResult_invMatrixOutputs_hi_hi_lo_hi_hi = decodeResult_orMatrixOutputs[48:47];
  wire [3:0]  decodeResult_invMatrixOutputs_hi_hi_lo_hi = {decodeResult_invMatrixOutputs_hi_hi_lo_hi_hi, decodeResult_invMatrixOutputs_hi_hi_lo_hi_lo};
  wire [6:0]  decodeResult_invMatrixOutputs_hi_hi_lo = {decodeResult_invMatrixOutputs_hi_hi_lo_hi, decodeResult_invMatrixOutputs_hi_hi_lo_lo};
  wire [1:0]  decodeResult_invMatrixOutputs_hi_hi_hi_lo_hi = decodeResult_orMatrixOutputs[51:50];
  wire [2:0]  decodeResult_invMatrixOutputs_hi_hi_hi_lo = {decodeResult_invMatrixOutputs_hi_hi_hi_lo_hi, decodeResult_orMatrixOutputs[49]};
  wire [1:0]  decodeResult_invMatrixOutputs_hi_hi_hi_hi_lo = decodeResult_orMatrixOutputs[53:52];
  wire [1:0]  decodeResult_invMatrixOutputs_hi_hi_hi_hi_hi = decodeResult_orMatrixOutputs[55:54];
  wire [3:0]  decodeResult_invMatrixOutputs_hi_hi_hi_hi = {decodeResult_invMatrixOutputs_hi_hi_hi_hi_hi, decodeResult_invMatrixOutputs_hi_hi_hi_hi_lo};
  wire [6:0]  decodeResult_invMatrixOutputs_hi_hi_hi = {decodeResult_invMatrixOutputs_hi_hi_hi_hi, decodeResult_invMatrixOutputs_hi_hi_hi_lo};
  wire [13:0] decodeResult_invMatrixOutputs_hi_hi = {decodeResult_invMatrixOutputs_hi_hi_hi, decodeResult_invMatrixOutputs_hi_hi_lo};
  wire [27:0] decodeResult_invMatrixOutputs_hi = {decodeResult_invMatrixOutputs_hi_hi, decodeResult_invMatrixOutputs_hi_lo};
  assign decodeResult_invMatrixOutputs = {decodeResult_invMatrixOutputs_hi, decodeResult_invMatrixOutputs_lo};
  wire [55:0] decodeResult_plaOutput = decodeResult_invMatrixOutputs;
  assign decodeResult_orderReduce = decodeResult_plaOutput[55];
  assign decodeResult_floatMul = decodeResult_plaOutput[54];
  assign decodeResult_fpExecutionType = decodeResult_plaOutput[53:52];
  assign decodeResult_float = decodeResult_plaOutput[51];
  assign decodeResult_specialSlot = decodeResult_plaOutput[50];
  assign decodeResult_topUop = decodeResult_plaOutput[49:45];
  assign decodeResult_popCount = decodeResult_plaOutput[44];
  assign decodeResult_ffo = decodeResult_plaOutput[43];
  assign decodeResult_average = decodeResult_plaOutput[42];
  assign decodeResult_reverse = decodeResult_plaOutput[41];
  assign decodeResult_dontNeedExecuteInLane = decodeResult_plaOutput[40];
  assign decodeResult_scheduler = decodeResult_plaOutput[39];
  assign decodeResult_sReadVD = decodeResult_plaOutput[38];
  assign decodeResult_vtype = decodeResult_plaOutput[37];
  assign decodeResult_sWrite = decodeResult_plaOutput[36];
  assign decodeResult_crossRead = decodeResult_plaOutput[35];
  assign decodeResult_crossWrite = decodeResult_plaOutput[34];
  assign decodeResult_maskUnit = decodeResult_plaOutput[33];
  assign decodeResult_special = decodeResult_plaOutput[32];
  assign decodeResult_saturate = decodeResult_plaOutput[31];
  assign decodeResult_vwmacc = decodeResult_plaOutput[30];
  assign decodeResult_readOnly = decodeResult_plaOutput[29];
  assign decodeResult_maskSource = decodeResult_plaOutput[28];
  assign decodeResult_maskDestination = decodeResult_plaOutput[27];
  assign decodeResult_maskLogic = decodeResult_plaOutput[26];
  assign decodeResult_uop = decodeResult_plaOutput[25:22];
  assign decodeResult_iota = decodeResult_plaOutput[21];
  assign decodeResult_mv = decodeResult_plaOutput[20];
  assign decodeResult_extend = decodeResult_plaOutput[19];
  assign decodeResult_unOrderWrite = decodeResult_plaOutput[18];
  assign decodeResult_compress = decodeResult_plaOutput[17];
  assign decodeResult_gather16 = decodeResult_plaOutput[16];
  assign decodeResult_gather = decodeResult_plaOutput[15];
  assign decodeResult_slid = decodeResult_plaOutput[14];
  assign decodeResult_targetRd = decodeResult_plaOutput[13];
  assign decodeResult_widenReduce = decodeResult_plaOutput[12];
  assign decodeResult_red = decodeResult_plaOutput[11];
  assign decodeResult_nr = decodeResult_plaOutput[10];
  assign decodeResult_itype = decodeResult_plaOutput[9];
  assign decodeResult_unsigned1 = decodeResult_plaOutput[8];
  assign decodeResult_unsigned0 = decodeResult_plaOutput[7];
  assign decodeResult_other = decodeResult_plaOutput[6];
  assign decodeResult_multiCycle = decodeResult_plaOutput[5];
  assign decodeResult_divider = decodeResult_plaOutput[4];
  assign decodeResult_multiplier = decodeResult_plaOutput[3];
  assign decodeResult_shift = decodeResult_plaOutput[2];
  assign decodeResult_adder = decodeResult_plaOutput[1];
  assign decodeResult_logic = decodeResult_plaOutput[0];
endmodule

