`define ref_T1_t1Probe_instructionCounter verification.probeWire_instructionCounter_probe
`define ref_T1_t1Probe_instructionIssue verification.probeWire_instructionIssue_probe
`define ref_T1_t1Probe_issueTag verification.probeWire_issueTag_probe
`define ref_T1_t1Probe_retireValid verification.probeWire_retireValid_probe
`define ref_T1_t1Probe_requestReg_valid verification.probeWire_requestReg_valid_probe
`define ref_T1_t1Probe_requestReg_bits_issue_instruction verification.probeWire_requestReg_bits_issue_instruction_probe
`define ref_T1_t1Probe_requestReg_bits_issue_rs1Data verification.probeWire_requestReg_bits_issue_rs1Data_probe
`define ref_T1_t1Probe_requestReg_bits_issue_rs2Data verification.probeWire_requestReg_bits_issue_rs2Data_probe
`define ref_T1_t1Probe_requestReg_bits_issue_vtype verification.probeWire_requestReg_bits_issue_vtype_probe
`define ref_T1_t1Probe_requestReg_bits_issue_vl verification.probeWire_requestReg_bits_issue_vl_probe
`define ref_T1_t1Probe_requestReg_bits_issue_vstart verification.probeWire_requestReg_bits_issue_vstart_probe
`define ref_T1_t1Probe_requestReg_bits_issue_vcsr verification.probeWire_requestReg_bits_issue_vcsr_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_specialSlot verification.probeWire_requestReg_bits_decodeResult_specialSlot_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_topUop verification.probeWire_requestReg_bits_decodeResult_topUop_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_popCount verification.probeWire_requestReg_bits_decodeResult_popCount_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_ffo verification.probeWire_requestReg_bits_decodeResult_ffo_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_average verification.probeWire_requestReg_bits_decodeResult_average_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_reverse verification.probeWire_requestReg_bits_decodeResult_reverse_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_dontNeedExecuteInLane verification.probeWire_requestReg_bits_decodeResult_dontNeedExecuteInLane_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_scheduler verification.probeWire_requestReg_bits_decodeResult_scheduler_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_sReadVD verification.probeWire_requestReg_bits_decodeResult_sReadVD_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_vtype verification.probeWire_requestReg_bits_decodeResult_vtype_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_sWrite verification.probeWire_requestReg_bits_decodeResult_sWrite_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_crossRead verification.probeWire_requestReg_bits_decodeResult_crossRead_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_crossWrite verification.probeWire_requestReg_bits_decodeResult_crossWrite_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_maskUnit verification.probeWire_requestReg_bits_decodeResult_maskUnit_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_special verification.probeWire_requestReg_bits_decodeResult_special_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_saturate verification.probeWire_requestReg_bits_decodeResult_saturate_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_vwmacc verification.probeWire_requestReg_bits_decodeResult_vwmacc_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_readOnly verification.probeWire_requestReg_bits_decodeResult_readOnly_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_maskSource verification.probeWire_requestReg_bits_decodeResult_maskSource_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_maskDestination verification.probeWire_requestReg_bits_decodeResult_maskDestination_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_maskLogic verification.probeWire_requestReg_bits_decodeResult_maskLogic_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_uop verification.probeWire_requestReg_bits_decodeResult_uop_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_iota verification.probeWire_requestReg_bits_decodeResult_iota_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_mv verification.probeWire_requestReg_bits_decodeResult_mv_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_extend verification.probeWire_requestReg_bits_decodeResult_extend_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_unOrderWrite verification.probeWire_requestReg_bits_decodeResult_unOrderWrite_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_compress verification.probeWire_requestReg_bits_decodeResult_compress_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_gather16 verification.probeWire_requestReg_bits_decodeResult_gather16_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_gather verification.probeWire_requestReg_bits_decodeResult_gather_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_slid verification.probeWire_requestReg_bits_decodeResult_slid_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_targetRd verification.probeWire_requestReg_bits_decodeResult_targetRd_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_widenReduce verification.probeWire_requestReg_bits_decodeResult_widenReduce_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_red verification.probeWire_requestReg_bits_decodeResult_red_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_nr verification.probeWire_requestReg_bits_decodeResult_nr_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_itype verification.probeWire_requestReg_bits_decodeResult_itype_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_unsigned1 verification.probeWire_requestReg_bits_decodeResult_unsigned1_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_unsigned0 verification.probeWire_requestReg_bits_decodeResult_unsigned0_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_other verification.probeWire_requestReg_bits_decodeResult_other_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_multiCycle verification.probeWire_requestReg_bits_decodeResult_multiCycle_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_divider verification.probeWire_requestReg_bits_decodeResult_divider_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_multiplier verification.probeWire_requestReg_bits_decodeResult_multiplier_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_shift verification.probeWire_requestReg_bits_decodeResult_shift_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_adder verification.probeWire_requestReg_bits_decodeResult_adder_probe
`define ref_T1_t1Probe_requestReg_bits_decodeResult_logic verification.probeWire_requestReg_bits_decodeResult_logic_probe
`define ref_T1_t1Probe_requestReg_bits_instructionIndex verification.probeWire_requestReg_bits_instructionIndex_probe
`define ref_T1_t1Probe_requestReg_bits_vdIsV0 verification.probeWire_requestReg_bits_vdIsV0_probe
`define ref_T1_t1Probe_requestReg_bits_writeByte verification.probeWire_requestReg_bits_writeByte_probe
`define ref_T1_t1Probe_requestRegReady verification.probeWire_requestRegReady_probe
`define ref_T1_t1Probe_writeQueueEnqVec_0_valid verification.probeWire_writeQueueEnqVec_0_valid_probe
`define ref_T1_t1Probe_writeQueueEnqVec_0_bits verification.probeWire_writeQueueEnqVec_0_bits_probe
`define ref_T1_t1Probe_writeQueueEnqVec_1_valid verification.probeWire_writeQueueEnqVec_1_valid_probe
`define ref_T1_t1Probe_writeQueueEnqVec_1_bits verification.probeWire_writeQueueEnqVec_1_bits_probe
`define ref_T1_t1Probe_writeQueueEnqVec_2_valid verification.probeWire_writeQueueEnqVec_2_valid_probe
`define ref_T1_t1Probe_writeQueueEnqVec_2_bits verification.probeWire_writeQueueEnqVec_2_bits_probe
`define ref_T1_t1Probe_writeQueueEnqVec_3_valid verification.probeWire_writeQueueEnqVec_3_valid_probe
`define ref_T1_t1Probe_writeQueueEnqVec_3_bits verification.probeWire_writeQueueEnqVec_3_bits_probe
`define ref_T1_t1Probe_writeQueueEnqVec_4_valid verification.probeWire_writeQueueEnqVec_4_valid_probe
`define ref_T1_t1Probe_writeQueueEnqVec_4_bits verification.probeWire_writeQueueEnqVec_4_bits_probe
`define ref_T1_t1Probe_writeQueueEnqVec_5_valid verification.probeWire_writeQueueEnqVec_5_valid_probe
`define ref_T1_t1Probe_writeQueueEnqVec_5_bits verification.probeWire_writeQueueEnqVec_5_bits_probe
`define ref_T1_t1Probe_writeQueueEnqVec_6_valid verification.probeWire_writeQueueEnqVec_6_valid_probe
`define ref_T1_t1Probe_writeQueueEnqVec_6_bits verification.probeWire_writeQueueEnqVec_6_bits_probe
`define ref_T1_t1Probe_writeQueueEnqVec_7_valid verification.probeWire_writeQueueEnqVec_7_valid_probe
`define ref_T1_t1Probe_writeQueueEnqVec_7_bits verification.probeWire_writeQueueEnqVec_7_bits_probe
`define ref_T1_t1Probe_writeQueueEnqVec_8_valid verification.probeWire_writeQueueEnqVec_8_valid_probe
`define ref_T1_t1Probe_writeQueueEnqVec_8_bits verification.probeWire_writeQueueEnqVec_8_bits_probe
`define ref_T1_t1Probe_writeQueueEnqVec_9_valid verification.probeWire_writeQueueEnqVec_9_valid_probe
`define ref_T1_t1Probe_writeQueueEnqVec_9_bits verification.probeWire_writeQueueEnqVec_9_bits_probe
`define ref_T1_t1Probe_writeQueueEnqVec_10_valid verification.probeWire_writeQueueEnqVec_10_valid_probe
`define ref_T1_t1Probe_writeQueueEnqVec_10_bits verification.probeWire_writeQueueEnqVec_10_bits_probe
`define ref_T1_t1Probe_writeQueueEnqVec_11_valid verification.probeWire_writeQueueEnqVec_11_valid_probe
`define ref_T1_t1Probe_writeQueueEnqVec_11_bits verification.probeWire_writeQueueEnqVec_11_bits_probe
`define ref_T1_t1Probe_writeQueueEnqVec_12_valid verification.probeWire_writeQueueEnqVec_12_valid_probe
`define ref_T1_t1Probe_writeQueueEnqVec_12_bits verification.probeWire_writeQueueEnqVec_12_bits_probe
`define ref_T1_t1Probe_writeQueueEnqVec_13_valid verification.probeWire_writeQueueEnqVec_13_valid_probe
`define ref_T1_t1Probe_writeQueueEnqVec_13_bits verification.probeWire_writeQueueEnqVec_13_bits_probe
`define ref_T1_t1Probe_writeQueueEnqVec_14_valid verification.probeWire_writeQueueEnqVec_14_valid_probe
`define ref_T1_t1Probe_writeQueueEnqVec_14_bits verification.probeWire_writeQueueEnqVec_14_bits_probe
`define ref_T1_t1Probe_writeQueueEnqVec_15_valid verification.probeWire_writeQueueEnqVec_15_valid_probe
`define ref_T1_t1Probe_writeQueueEnqVec_15_bits verification.probeWire_writeQueueEnqVec_15_bits_probe
`define ref_T1_t1Probe_instructionValid verification.probeWire_instructionValid_probe
`define ref_T1_t1Probe_responseCounter verification.probeWire_responseCounter_probe
`define ref_T1_t1Probe_lsuProbe_slots_0_dataVd verification.probeWire_lsuProbe_slots_0_dataVd_probe
`define ref_T1_t1Probe_lsuProbe_slots_0_dataOffset verification.probeWire_lsuProbe_slots_0_dataOffset_probe
`define ref_T1_t1Probe_lsuProbe_slots_0_dataMask verification.probeWire_lsuProbe_slots_0_dataMask_probe
`define ref_T1_t1Probe_lsuProbe_slots_0_dataData verification.probeWire_lsuProbe_slots_0_dataData_probe
`define ref_T1_t1Probe_lsuProbe_slots_0_dataInstruction verification.probeWire_lsuProbe_slots_0_dataInstruction_probe
`define ref_T1_t1Probe_lsuProbe_slots_0_writeValid verification.probeWire_lsuProbe_slots_0_writeValid_probe
`define ref_T1_t1Probe_lsuProbe_slots_0_targetLane verification.probeWire_lsuProbe_slots_0_targetLane_probe
`define ref_T1_t1Probe_lsuProbe_slots_1_dataVd verification.probeWire_lsuProbe_slots_1_dataVd_probe
`define ref_T1_t1Probe_lsuProbe_slots_1_dataOffset verification.probeWire_lsuProbe_slots_1_dataOffset_probe
`define ref_T1_t1Probe_lsuProbe_slots_1_dataMask verification.probeWire_lsuProbe_slots_1_dataMask_probe
`define ref_T1_t1Probe_lsuProbe_slots_1_dataData verification.probeWire_lsuProbe_slots_1_dataData_probe
`define ref_T1_t1Probe_lsuProbe_slots_1_dataInstruction verification.probeWire_lsuProbe_slots_1_dataInstruction_probe
`define ref_T1_t1Probe_lsuProbe_slots_1_writeValid verification.probeWire_lsuProbe_slots_1_writeValid_probe
`define ref_T1_t1Probe_lsuProbe_slots_1_targetLane verification.probeWire_lsuProbe_slots_1_targetLane_probe
`define ref_T1_t1Probe_lsuProbe_slots_2_dataVd verification.probeWire_lsuProbe_slots_2_dataVd_probe
`define ref_T1_t1Probe_lsuProbe_slots_2_dataOffset verification.probeWire_lsuProbe_slots_2_dataOffset_probe
`define ref_T1_t1Probe_lsuProbe_slots_2_dataMask verification.probeWire_lsuProbe_slots_2_dataMask_probe
`define ref_T1_t1Probe_lsuProbe_slots_2_dataData verification.probeWire_lsuProbe_slots_2_dataData_probe
`define ref_T1_t1Probe_lsuProbe_slots_2_dataInstruction verification.probeWire_lsuProbe_slots_2_dataInstruction_probe
`define ref_T1_t1Probe_lsuProbe_slots_2_writeValid verification.probeWire_lsuProbe_slots_2_writeValid_probe
`define ref_T1_t1Probe_lsuProbe_slots_2_targetLane verification.probeWire_lsuProbe_slots_2_targetLane_probe
`define ref_T1_t1Probe_lsuProbe_slots_3_dataVd verification.probeWire_lsuProbe_slots_3_dataVd_probe
`define ref_T1_t1Probe_lsuProbe_slots_3_dataOffset verification.probeWire_lsuProbe_slots_3_dataOffset_probe
`define ref_T1_t1Probe_lsuProbe_slots_3_dataMask verification.probeWire_lsuProbe_slots_3_dataMask_probe
`define ref_T1_t1Probe_lsuProbe_slots_3_dataData verification.probeWire_lsuProbe_slots_3_dataData_probe
`define ref_T1_t1Probe_lsuProbe_slots_3_dataInstruction verification.probeWire_lsuProbe_slots_3_dataInstruction_probe
`define ref_T1_t1Probe_lsuProbe_slots_3_writeValid verification.probeWire_lsuProbe_slots_3_writeValid_probe
`define ref_T1_t1Probe_lsuProbe_slots_3_targetLane verification.probeWire_lsuProbe_slots_3_targetLane_probe
`define ref_T1_t1Probe_lsuProbe_slots_4_dataVd verification.probeWire_lsuProbe_slots_4_dataVd_probe
`define ref_T1_t1Probe_lsuProbe_slots_4_dataOffset verification.probeWire_lsuProbe_slots_4_dataOffset_probe
`define ref_T1_t1Probe_lsuProbe_slots_4_dataMask verification.probeWire_lsuProbe_slots_4_dataMask_probe
`define ref_T1_t1Probe_lsuProbe_slots_4_dataData verification.probeWire_lsuProbe_slots_4_dataData_probe
`define ref_T1_t1Probe_lsuProbe_slots_4_dataInstruction verification.probeWire_lsuProbe_slots_4_dataInstruction_probe
`define ref_T1_t1Probe_lsuProbe_slots_4_writeValid verification.probeWire_lsuProbe_slots_4_writeValid_probe
`define ref_T1_t1Probe_lsuProbe_slots_4_targetLane verification.probeWire_lsuProbe_slots_4_targetLane_probe
`define ref_T1_t1Probe_lsuProbe_slots_5_dataVd verification.probeWire_lsuProbe_slots_5_dataVd_probe
`define ref_T1_t1Probe_lsuProbe_slots_5_dataOffset verification.probeWire_lsuProbe_slots_5_dataOffset_probe
`define ref_T1_t1Probe_lsuProbe_slots_5_dataMask verification.probeWire_lsuProbe_slots_5_dataMask_probe
`define ref_T1_t1Probe_lsuProbe_slots_5_dataData verification.probeWire_lsuProbe_slots_5_dataData_probe
`define ref_T1_t1Probe_lsuProbe_slots_5_dataInstruction verification.probeWire_lsuProbe_slots_5_dataInstruction_probe
`define ref_T1_t1Probe_lsuProbe_slots_5_writeValid verification.probeWire_lsuProbe_slots_5_writeValid_probe
`define ref_T1_t1Probe_lsuProbe_slots_5_targetLane verification.probeWire_lsuProbe_slots_5_targetLane_probe
`define ref_T1_t1Probe_lsuProbe_slots_6_dataVd verification.probeWire_lsuProbe_slots_6_dataVd_probe
`define ref_T1_t1Probe_lsuProbe_slots_6_dataOffset verification.probeWire_lsuProbe_slots_6_dataOffset_probe
`define ref_T1_t1Probe_lsuProbe_slots_6_dataMask verification.probeWire_lsuProbe_slots_6_dataMask_probe
`define ref_T1_t1Probe_lsuProbe_slots_6_dataData verification.probeWire_lsuProbe_slots_6_dataData_probe
`define ref_T1_t1Probe_lsuProbe_slots_6_dataInstruction verification.probeWire_lsuProbe_slots_6_dataInstruction_probe
`define ref_T1_t1Probe_lsuProbe_slots_6_writeValid verification.probeWire_lsuProbe_slots_6_writeValid_probe
`define ref_T1_t1Probe_lsuProbe_slots_6_targetLane verification.probeWire_lsuProbe_slots_6_targetLane_probe
`define ref_T1_t1Probe_lsuProbe_slots_7_dataVd verification.probeWire_lsuProbe_slots_7_dataVd_probe
`define ref_T1_t1Probe_lsuProbe_slots_7_dataOffset verification.probeWire_lsuProbe_slots_7_dataOffset_probe
`define ref_T1_t1Probe_lsuProbe_slots_7_dataMask verification.probeWire_lsuProbe_slots_7_dataMask_probe
`define ref_T1_t1Probe_lsuProbe_slots_7_dataData verification.probeWire_lsuProbe_slots_7_dataData_probe
`define ref_T1_t1Probe_lsuProbe_slots_7_dataInstruction verification.probeWire_lsuProbe_slots_7_dataInstruction_probe
`define ref_T1_t1Probe_lsuProbe_slots_7_writeValid verification.probeWire_lsuProbe_slots_7_writeValid_probe
`define ref_T1_t1Probe_lsuProbe_slots_7_targetLane verification.probeWire_lsuProbe_slots_7_targetLane_probe
`define ref_T1_t1Probe_lsuProbe_slots_8_dataVd verification.probeWire_lsuProbe_slots_8_dataVd_probe
`define ref_T1_t1Probe_lsuProbe_slots_8_dataOffset verification.probeWire_lsuProbe_slots_8_dataOffset_probe
`define ref_T1_t1Probe_lsuProbe_slots_8_dataMask verification.probeWire_lsuProbe_slots_8_dataMask_probe
`define ref_T1_t1Probe_lsuProbe_slots_8_dataData verification.probeWire_lsuProbe_slots_8_dataData_probe
`define ref_T1_t1Probe_lsuProbe_slots_8_dataInstruction verification.probeWire_lsuProbe_slots_8_dataInstruction_probe
`define ref_T1_t1Probe_lsuProbe_slots_8_writeValid verification.probeWire_lsuProbe_slots_8_writeValid_probe
`define ref_T1_t1Probe_lsuProbe_slots_8_targetLane verification.probeWire_lsuProbe_slots_8_targetLane_probe
`define ref_T1_t1Probe_lsuProbe_slots_9_dataVd verification.probeWire_lsuProbe_slots_9_dataVd_probe
`define ref_T1_t1Probe_lsuProbe_slots_9_dataOffset verification.probeWire_lsuProbe_slots_9_dataOffset_probe
`define ref_T1_t1Probe_lsuProbe_slots_9_dataMask verification.probeWire_lsuProbe_slots_9_dataMask_probe
`define ref_T1_t1Probe_lsuProbe_slots_9_dataData verification.probeWire_lsuProbe_slots_9_dataData_probe
`define ref_T1_t1Probe_lsuProbe_slots_9_dataInstruction verification.probeWire_lsuProbe_slots_9_dataInstruction_probe
`define ref_T1_t1Probe_lsuProbe_slots_9_writeValid verification.probeWire_lsuProbe_slots_9_writeValid_probe
`define ref_T1_t1Probe_lsuProbe_slots_9_targetLane verification.probeWire_lsuProbe_slots_9_targetLane_probe
`define ref_T1_t1Probe_lsuProbe_slots_10_dataVd verification.probeWire_lsuProbe_slots_10_dataVd_probe
`define ref_T1_t1Probe_lsuProbe_slots_10_dataOffset verification.probeWire_lsuProbe_slots_10_dataOffset_probe
`define ref_T1_t1Probe_lsuProbe_slots_10_dataMask verification.probeWire_lsuProbe_slots_10_dataMask_probe
`define ref_T1_t1Probe_lsuProbe_slots_10_dataData verification.probeWire_lsuProbe_slots_10_dataData_probe
`define ref_T1_t1Probe_lsuProbe_slots_10_dataInstruction verification.probeWire_lsuProbe_slots_10_dataInstruction_probe
`define ref_T1_t1Probe_lsuProbe_slots_10_writeValid verification.probeWire_lsuProbe_slots_10_writeValid_probe
`define ref_T1_t1Probe_lsuProbe_slots_10_targetLane verification.probeWire_lsuProbe_slots_10_targetLane_probe
`define ref_T1_t1Probe_lsuProbe_slots_11_dataVd verification.probeWire_lsuProbe_slots_11_dataVd_probe
`define ref_T1_t1Probe_lsuProbe_slots_11_dataOffset verification.probeWire_lsuProbe_slots_11_dataOffset_probe
`define ref_T1_t1Probe_lsuProbe_slots_11_dataMask verification.probeWire_lsuProbe_slots_11_dataMask_probe
`define ref_T1_t1Probe_lsuProbe_slots_11_dataData verification.probeWire_lsuProbe_slots_11_dataData_probe
`define ref_T1_t1Probe_lsuProbe_slots_11_dataInstruction verification.probeWire_lsuProbe_slots_11_dataInstruction_probe
`define ref_T1_t1Probe_lsuProbe_slots_11_writeValid verification.probeWire_lsuProbe_slots_11_writeValid_probe
`define ref_T1_t1Probe_lsuProbe_slots_11_targetLane verification.probeWire_lsuProbe_slots_11_targetLane_probe
`define ref_T1_t1Probe_lsuProbe_slots_12_dataVd verification.probeWire_lsuProbe_slots_12_dataVd_probe
`define ref_T1_t1Probe_lsuProbe_slots_12_dataOffset verification.probeWire_lsuProbe_slots_12_dataOffset_probe
`define ref_T1_t1Probe_lsuProbe_slots_12_dataMask verification.probeWire_lsuProbe_slots_12_dataMask_probe
`define ref_T1_t1Probe_lsuProbe_slots_12_dataData verification.probeWire_lsuProbe_slots_12_dataData_probe
`define ref_T1_t1Probe_lsuProbe_slots_12_dataInstruction verification.probeWire_lsuProbe_slots_12_dataInstruction_probe
`define ref_T1_t1Probe_lsuProbe_slots_12_writeValid verification.probeWire_lsuProbe_slots_12_writeValid_probe
`define ref_T1_t1Probe_lsuProbe_slots_12_targetLane verification.probeWire_lsuProbe_slots_12_targetLane_probe
`define ref_T1_t1Probe_lsuProbe_slots_13_dataVd verification.probeWire_lsuProbe_slots_13_dataVd_probe
`define ref_T1_t1Probe_lsuProbe_slots_13_dataOffset verification.probeWire_lsuProbe_slots_13_dataOffset_probe
`define ref_T1_t1Probe_lsuProbe_slots_13_dataMask verification.probeWire_lsuProbe_slots_13_dataMask_probe
`define ref_T1_t1Probe_lsuProbe_slots_13_dataData verification.probeWire_lsuProbe_slots_13_dataData_probe
`define ref_T1_t1Probe_lsuProbe_slots_13_dataInstruction verification.probeWire_lsuProbe_slots_13_dataInstruction_probe
`define ref_T1_t1Probe_lsuProbe_slots_13_writeValid verification.probeWire_lsuProbe_slots_13_writeValid_probe
`define ref_T1_t1Probe_lsuProbe_slots_13_targetLane verification.probeWire_lsuProbe_slots_13_targetLane_probe
`define ref_T1_t1Probe_lsuProbe_slots_14_dataVd verification.probeWire_lsuProbe_slots_14_dataVd_probe
`define ref_T1_t1Probe_lsuProbe_slots_14_dataOffset verification.probeWire_lsuProbe_slots_14_dataOffset_probe
`define ref_T1_t1Probe_lsuProbe_slots_14_dataMask verification.probeWire_lsuProbe_slots_14_dataMask_probe
`define ref_T1_t1Probe_lsuProbe_slots_14_dataData verification.probeWire_lsuProbe_slots_14_dataData_probe
`define ref_T1_t1Probe_lsuProbe_slots_14_dataInstruction verification.probeWire_lsuProbe_slots_14_dataInstruction_probe
`define ref_T1_t1Probe_lsuProbe_slots_14_writeValid verification.probeWire_lsuProbe_slots_14_writeValid_probe
`define ref_T1_t1Probe_lsuProbe_slots_14_targetLane verification.probeWire_lsuProbe_slots_14_targetLane_probe
`define ref_T1_t1Probe_lsuProbe_slots_15_dataVd verification.probeWire_lsuProbe_slots_15_dataVd_probe
`define ref_T1_t1Probe_lsuProbe_slots_15_dataOffset verification.probeWire_lsuProbe_slots_15_dataOffset_probe
`define ref_T1_t1Probe_lsuProbe_slots_15_dataMask verification.probeWire_lsuProbe_slots_15_dataMask_probe
`define ref_T1_t1Probe_lsuProbe_slots_15_dataData verification.probeWire_lsuProbe_slots_15_dataData_probe
`define ref_T1_t1Probe_lsuProbe_slots_15_dataInstruction verification.probeWire_lsuProbe_slots_15_dataInstruction_probe
`define ref_T1_t1Probe_lsuProbe_slots_15_writeValid verification.probeWire_lsuProbe_slots_15_writeValid_probe
`define ref_T1_t1Probe_lsuProbe_slots_15_targetLane verification.probeWire_lsuProbe_slots_15_targetLane_probe
`define ref_T1_t1Probe_lsuProbe_storeUnitProbe_valid verification.probeWire_lsuProbe_storeUnitProbe_valid_probe
`define ref_T1_t1Probe_lsuProbe_storeUnitProbe_data verification.probeWire_lsuProbe_storeUnitProbe_data_probe
`define ref_T1_t1Probe_lsuProbe_storeUnitProbe_mask verification.probeWire_lsuProbe_storeUnitProbe_mask_probe
`define ref_T1_t1Probe_lsuProbe_storeUnitProbe_index verification.probeWire_lsuProbe_storeUnitProbe_index_probe
`define ref_T1_t1Probe_lsuProbe_storeUnitProbe_address verification.probeWire_lsuProbe_storeUnitProbe_address_probe
`define ref_T1_t1Probe_lsuProbe_otherUnitProbe_valid verification.probeWire_lsuProbe_otherUnitProbe_valid_probe
`define ref_T1_t1Probe_lsuProbe_otherUnitProbe_data verification.probeWire_lsuProbe_otherUnitProbe_data_probe
`define ref_T1_t1Probe_lsuProbe_otherUnitProbe_mask verification.probeWire_lsuProbe_otherUnitProbe_mask_probe
`define ref_T1_t1Probe_lsuProbe_otherUnitProbe_index verification.probeWire_lsuProbe_otherUnitProbe_index_probe
`define ref_T1_t1Probe_lsuProbe_otherUnitProbe_address verification.probeWire_lsuProbe_otherUnitProbe_address_probe
`define ref_T1_t1Probe_lsuProbe_reqEnq verification.probeWire_lsuProbe_reqEnq_probe
`define ref_T1_t1Probe_lsuProbe_lsuInstructionValid verification.probeWire_lsuProbe_lsuInstructionValid_probe
`define ref_T1_t1Probe_laneProbes_0_slots_0_stage0EnqueueReady verification.probeWire_laneProbes_0_slots_0_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_0_slots_0_stage0EnqueueValid verification.probeWire_laneProbes_0_slots_0_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_0_slots_0_changingMaskSet verification.probeWire_laneProbes_0_slots_0_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_0_slots_0_slotActive verification.probeWire_laneProbes_0_slots_0_slotActive_probe
`define ref_T1_t1Probe_laneProbes_0_slots_0_slotOccupied verification.probeWire_laneProbes_0_slots_0_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_0_slots_0_pipeFinish verification.probeWire_laneProbes_0_slots_0_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_0_slots_0_slotShiftValid verification.probeWire_laneProbes_0_slots_0_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_0_slots_0_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_0_slots_0_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_0_slots_0_decodeResultIsScheduler verification.probeWire_laneProbes_0_slots_0_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_0_slots_0_executionUnitVfuRequestReady verification.probeWire_laneProbes_0_slots_0_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_0_slots_0_executionUnitVfuRequestValid verification.probeWire_laneProbes_0_slots_0_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_0_slots_0_stage3VrfWriteReady verification.probeWire_laneProbes_0_slots_0_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_0_slots_0_stage3VrfWriteValid verification.probeWire_laneProbes_0_slots_0_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_0_slots_0_writeQueueEnq verification.probeWire_laneProbes_0_slots_0_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_0_slots_0_writeTag verification.probeWire_laneProbes_0_slots_0_writeTag_probe
`define ref_T1_t1Probe_laneProbes_0_slots_0_writeMask verification.probeWire_laneProbes_0_slots_0_writeMask_probe
`define ref_T1_t1Probe_laneProbes_0_slots_1_stage0EnqueueReady verification.probeWire_laneProbes_0_slots_1_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_0_slots_1_stage0EnqueueValid verification.probeWire_laneProbes_0_slots_1_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_0_slots_1_changingMaskSet verification.probeWire_laneProbes_0_slots_1_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_0_slots_1_slotActive verification.probeWire_laneProbes_0_slots_1_slotActive_probe
`define ref_T1_t1Probe_laneProbes_0_slots_1_slotOccupied verification.probeWire_laneProbes_0_slots_1_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_0_slots_1_pipeFinish verification.probeWire_laneProbes_0_slots_1_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_0_slots_1_slotShiftValid verification.probeWire_laneProbes_0_slots_1_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_0_slots_1_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_0_slots_1_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_0_slots_1_decodeResultIsScheduler verification.probeWire_laneProbes_0_slots_1_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_0_slots_1_executionUnitVfuRequestReady verification.probeWire_laneProbes_0_slots_1_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_0_slots_1_executionUnitVfuRequestValid verification.probeWire_laneProbes_0_slots_1_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_0_slots_1_stage3VrfWriteReady verification.probeWire_laneProbes_0_slots_1_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_0_slots_1_stage3VrfWriteValid verification.probeWire_laneProbes_0_slots_1_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_0_slots_1_writeQueueEnq verification.probeWire_laneProbes_0_slots_1_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_0_slots_1_writeTag verification.probeWire_laneProbes_0_slots_1_writeTag_probe
`define ref_T1_t1Probe_laneProbes_0_slots_1_writeMask verification.probeWire_laneProbes_0_slots_1_writeMask_probe
`define ref_T1_t1Probe_laneProbes_0_slots_2_stage0EnqueueReady verification.probeWire_laneProbes_0_slots_2_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_0_slots_2_stage0EnqueueValid verification.probeWire_laneProbes_0_slots_2_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_0_slots_2_changingMaskSet verification.probeWire_laneProbes_0_slots_2_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_0_slots_2_slotActive verification.probeWire_laneProbes_0_slots_2_slotActive_probe
`define ref_T1_t1Probe_laneProbes_0_slots_2_slotOccupied verification.probeWire_laneProbes_0_slots_2_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_0_slots_2_pipeFinish verification.probeWire_laneProbes_0_slots_2_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_0_slots_2_slotShiftValid verification.probeWire_laneProbes_0_slots_2_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_0_slots_2_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_0_slots_2_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_0_slots_2_decodeResultIsScheduler verification.probeWire_laneProbes_0_slots_2_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_0_slots_2_executionUnitVfuRequestReady verification.probeWire_laneProbes_0_slots_2_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_0_slots_2_executionUnitVfuRequestValid verification.probeWire_laneProbes_0_slots_2_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_0_slots_2_stage3VrfWriteReady verification.probeWire_laneProbes_0_slots_2_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_0_slots_2_stage3VrfWriteValid verification.probeWire_laneProbes_0_slots_2_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_0_slots_2_writeQueueEnq verification.probeWire_laneProbes_0_slots_2_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_0_slots_2_writeTag verification.probeWire_laneProbes_0_slots_2_writeTag_probe
`define ref_T1_t1Probe_laneProbes_0_slots_2_writeMask verification.probeWire_laneProbes_0_slots_2_writeMask_probe
`define ref_T1_t1Probe_laneProbes_0_slots_3_stage0EnqueueReady verification.probeWire_laneProbes_0_slots_3_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_0_slots_3_stage0EnqueueValid verification.probeWire_laneProbes_0_slots_3_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_0_slots_3_changingMaskSet verification.probeWire_laneProbes_0_slots_3_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_0_slots_3_slotActive verification.probeWire_laneProbes_0_slots_3_slotActive_probe
`define ref_T1_t1Probe_laneProbes_0_slots_3_slotOccupied verification.probeWire_laneProbes_0_slots_3_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_0_slots_3_pipeFinish verification.probeWire_laneProbes_0_slots_3_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_0_slots_3_slotShiftValid verification.probeWire_laneProbes_0_slots_3_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_0_slots_3_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_0_slots_3_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_0_slots_3_decodeResultIsScheduler verification.probeWire_laneProbes_0_slots_3_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_0_slots_3_executionUnitVfuRequestReady verification.probeWire_laneProbes_0_slots_3_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_0_slots_3_executionUnitVfuRequestValid verification.probeWire_laneProbes_0_slots_3_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_0_slots_3_stage3VrfWriteReady verification.probeWire_laneProbes_0_slots_3_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_0_slots_3_stage3VrfWriteValid verification.probeWire_laneProbes_0_slots_3_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_0_slots_3_writeQueueEnq verification.probeWire_laneProbes_0_slots_3_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_0_slots_3_writeTag verification.probeWire_laneProbes_0_slots_3_writeTag_probe
`define ref_T1_t1Probe_laneProbes_0_slots_3_writeMask verification.probeWire_laneProbes_0_slots_3_writeMask_probe
`define ref_T1_t1Probe_laneProbes_0_laneRequestStall verification.probeWire_laneProbes_0_laneRequestStall_probe
`define ref_T1_t1Probe_laneProbes_0_lastSlotOccupied verification.probeWire_laneProbes_0_lastSlotOccupied_probe
`define ref_T1_t1Probe_laneProbes_0_instructionFinished verification.probeWire_laneProbes_0_instructionFinished_probe
`define ref_T1_t1Probe_laneProbes_0_instructionValid verification.probeWire_laneProbes_0_instructionValid_probe
`define ref_T1_t1Probe_laneProbes_0_crossWriteProbe_0_valid verification.probeWire_laneProbes_0_crossWriteProbe_0_valid_probe
`define ref_T1_t1Probe_laneProbes_0_crossWriteProbe_0_bits_writeTag verification.probeWire_laneProbes_0_crossWriteProbe_0_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_0_crossWriteProbe_0_bits_writeMask verification.probeWire_laneProbes_0_crossWriteProbe_0_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_0_crossWriteProbe_1_valid verification.probeWire_laneProbes_0_crossWriteProbe_1_valid_probe
`define ref_T1_t1Probe_laneProbes_0_crossWriteProbe_1_bits_writeTag verification.probeWire_laneProbes_0_crossWriteProbe_1_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_0_crossWriteProbe_1_bits_writeMask verification.probeWire_laneProbes_0_crossWriteProbe_1_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_0_vrfProbe_valid verification.probeWire_laneProbes_0_vrfProbe_valid_probe
`define ref_T1_t1Probe_laneProbes_0_vrfProbe_requestVd verification.probeWire_laneProbes_0_vrfProbe_requestVd_probe
`define ref_T1_t1Probe_laneProbes_0_vrfProbe_requestOffset verification.probeWire_laneProbes_0_vrfProbe_requestOffset_probe
`define ref_T1_t1Probe_laneProbes_0_vrfProbe_requestMask verification.probeWire_laneProbes_0_vrfProbe_requestMask_probe
`define ref_T1_t1Probe_laneProbes_0_vrfProbe_requestData verification.probeWire_laneProbes_0_vrfProbe_requestData_probe
`define ref_T1_t1Probe_laneProbes_0_vrfProbe_requestInstruction verification.probeWire_laneProbes_0_vrfProbe_requestInstruction_probe
`define ref_T1_t1Probe_laneProbes_1_slots_0_stage0EnqueueReady verification.probeWire_laneProbes_1_slots_0_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_1_slots_0_stage0EnqueueValid verification.probeWire_laneProbes_1_slots_0_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_1_slots_0_changingMaskSet verification.probeWire_laneProbes_1_slots_0_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_1_slots_0_slotActive verification.probeWire_laneProbes_1_slots_0_slotActive_probe
`define ref_T1_t1Probe_laneProbes_1_slots_0_slotOccupied verification.probeWire_laneProbes_1_slots_0_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_1_slots_0_pipeFinish verification.probeWire_laneProbes_1_slots_0_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_1_slots_0_slotShiftValid verification.probeWire_laneProbes_1_slots_0_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_1_slots_0_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_1_slots_0_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_1_slots_0_decodeResultIsScheduler verification.probeWire_laneProbes_1_slots_0_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_1_slots_0_executionUnitVfuRequestReady verification.probeWire_laneProbes_1_slots_0_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_1_slots_0_executionUnitVfuRequestValid verification.probeWire_laneProbes_1_slots_0_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_1_slots_0_stage3VrfWriteReady verification.probeWire_laneProbes_1_slots_0_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_1_slots_0_stage3VrfWriteValid verification.probeWire_laneProbes_1_slots_0_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_1_slots_0_writeQueueEnq verification.probeWire_laneProbes_1_slots_0_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_1_slots_0_writeTag verification.probeWire_laneProbes_1_slots_0_writeTag_probe
`define ref_T1_t1Probe_laneProbes_1_slots_0_writeMask verification.probeWire_laneProbes_1_slots_0_writeMask_probe
`define ref_T1_t1Probe_laneProbes_1_slots_1_stage0EnqueueReady verification.probeWire_laneProbes_1_slots_1_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_1_slots_1_stage0EnqueueValid verification.probeWire_laneProbes_1_slots_1_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_1_slots_1_changingMaskSet verification.probeWire_laneProbes_1_slots_1_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_1_slots_1_slotActive verification.probeWire_laneProbes_1_slots_1_slotActive_probe
`define ref_T1_t1Probe_laneProbes_1_slots_1_slotOccupied verification.probeWire_laneProbes_1_slots_1_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_1_slots_1_pipeFinish verification.probeWire_laneProbes_1_slots_1_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_1_slots_1_slotShiftValid verification.probeWire_laneProbes_1_slots_1_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_1_slots_1_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_1_slots_1_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_1_slots_1_decodeResultIsScheduler verification.probeWire_laneProbes_1_slots_1_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_1_slots_1_executionUnitVfuRequestReady verification.probeWire_laneProbes_1_slots_1_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_1_slots_1_executionUnitVfuRequestValid verification.probeWire_laneProbes_1_slots_1_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_1_slots_1_stage3VrfWriteReady verification.probeWire_laneProbes_1_slots_1_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_1_slots_1_stage3VrfWriteValid verification.probeWire_laneProbes_1_slots_1_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_1_slots_1_writeQueueEnq verification.probeWire_laneProbes_1_slots_1_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_1_slots_1_writeTag verification.probeWire_laneProbes_1_slots_1_writeTag_probe
`define ref_T1_t1Probe_laneProbes_1_slots_1_writeMask verification.probeWire_laneProbes_1_slots_1_writeMask_probe
`define ref_T1_t1Probe_laneProbes_1_slots_2_stage0EnqueueReady verification.probeWire_laneProbes_1_slots_2_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_1_slots_2_stage0EnqueueValid verification.probeWire_laneProbes_1_slots_2_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_1_slots_2_changingMaskSet verification.probeWire_laneProbes_1_slots_2_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_1_slots_2_slotActive verification.probeWire_laneProbes_1_slots_2_slotActive_probe
`define ref_T1_t1Probe_laneProbes_1_slots_2_slotOccupied verification.probeWire_laneProbes_1_slots_2_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_1_slots_2_pipeFinish verification.probeWire_laneProbes_1_slots_2_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_1_slots_2_slotShiftValid verification.probeWire_laneProbes_1_slots_2_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_1_slots_2_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_1_slots_2_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_1_slots_2_decodeResultIsScheduler verification.probeWire_laneProbes_1_slots_2_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_1_slots_2_executionUnitVfuRequestReady verification.probeWire_laneProbes_1_slots_2_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_1_slots_2_executionUnitVfuRequestValid verification.probeWire_laneProbes_1_slots_2_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_1_slots_2_stage3VrfWriteReady verification.probeWire_laneProbes_1_slots_2_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_1_slots_2_stage3VrfWriteValid verification.probeWire_laneProbes_1_slots_2_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_1_slots_2_writeQueueEnq verification.probeWire_laneProbes_1_slots_2_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_1_slots_2_writeTag verification.probeWire_laneProbes_1_slots_2_writeTag_probe
`define ref_T1_t1Probe_laneProbes_1_slots_2_writeMask verification.probeWire_laneProbes_1_slots_2_writeMask_probe
`define ref_T1_t1Probe_laneProbes_1_slots_3_stage0EnqueueReady verification.probeWire_laneProbes_1_slots_3_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_1_slots_3_stage0EnqueueValid verification.probeWire_laneProbes_1_slots_3_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_1_slots_3_changingMaskSet verification.probeWire_laneProbes_1_slots_3_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_1_slots_3_slotActive verification.probeWire_laneProbes_1_slots_3_slotActive_probe
`define ref_T1_t1Probe_laneProbes_1_slots_3_slotOccupied verification.probeWire_laneProbes_1_slots_3_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_1_slots_3_pipeFinish verification.probeWire_laneProbes_1_slots_3_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_1_slots_3_slotShiftValid verification.probeWire_laneProbes_1_slots_3_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_1_slots_3_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_1_slots_3_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_1_slots_3_decodeResultIsScheduler verification.probeWire_laneProbes_1_slots_3_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_1_slots_3_executionUnitVfuRequestReady verification.probeWire_laneProbes_1_slots_3_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_1_slots_3_executionUnitVfuRequestValid verification.probeWire_laneProbes_1_slots_3_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_1_slots_3_stage3VrfWriteReady verification.probeWire_laneProbes_1_slots_3_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_1_slots_3_stage3VrfWriteValid verification.probeWire_laneProbes_1_slots_3_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_1_slots_3_writeQueueEnq verification.probeWire_laneProbes_1_slots_3_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_1_slots_3_writeTag verification.probeWire_laneProbes_1_slots_3_writeTag_probe
`define ref_T1_t1Probe_laneProbes_1_slots_3_writeMask verification.probeWire_laneProbes_1_slots_3_writeMask_probe
`define ref_T1_t1Probe_laneProbes_1_laneRequestStall verification.probeWire_laneProbes_1_laneRequestStall_probe
`define ref_T1_t1Probe_laneProbes_1_lastSlotOccupied verification.probeWire_laneProbes_1_lastSlotOccupied_probe
`define ref_T1_t1Probe_laneProbes_1_instructionFinished verification.probeWire_laneProbes_1_instructionFinished_probe
`define ref_T1_t1Probe_laneProbes_1_instructionValid verification.probeWire_laneProbes_1_instructionValid_probe
`define ref_T1_t1Probe_laneProbes_1_crossWriteProbe_0_valid verification.probeWire_laneProbes_1_crossWriteProbe_0_valid_probe
`define ref_T1_t1Probe_laneProbes_1_crossWriteProbe_0_bits_writeTag verification.probeWire_laneProbes_1_crossWriteProbe_0_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_1_crossWriteProbe_0_bits_writeMask verification.probeWire_laneProbes_1_crossWriteProbe_0_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_1_crossWriteProbe_1_valid verification.probeWire_laneProbes_1_crossWriteProbe_1_valid_probe
`define ref_T1_t1Probe_laneProbes_1_crossWriteProbe_1_bits_writeTag verification.probeWire_laneProbes_1_crossWriteProbe_1_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_1_crossWriteProbe_1_bits_writeMask verification.probeWire_laneProbes_1_crossWriteProbe_1_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_1_vrfProbe_valid verification.probeWire_laneProbes_1_vrfProbe_valid_probe
`define ref_T1_t1Probe_laneProbes_1_vrfProbe_requestVd verification.probeWire_laneProbes_1_vrfProbe_requestVd_probe
`define ref_T1_t1Probe_laneProbes_1_vrfProbe_requestOffset verification.probeWire_laneProbes_1_vrfProbe_requestOffset_probe
`define ref_T1_t1Probe_laneProbes_1_vrfProbe_requestMask verification.probeWire_laneProbes_1_vrfProbe_requestMask_probe
`define ref_T1_t1Probe_laneProbes_1_vrfProbe_requestData verification.probeWire_laneProbes_1_vrfProbe_requestData_probe
`define ref_T1_t1Probe_laneProbes_1_vrfProbe_requestInstruction verification.probeWire_laneProbes_1_vrfProbe_requestInstruction_probe
`define ref_T1_t1Probe_laneProbes_2_slots_0_stage0EnqueueReady verification.probeWire_laneProbes_2_slots_0_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_2_slots_0_stage0EnqueueValid verification.probeWire_laneProbes_2_slots_0_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_2_slots_0_changingMaskSet verification.probeWire_laneProbes_2_slots_0_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_2_slots_0_slotActive verification.probeWire_laneProbes_2_slots_0_slotActive_probe
`define ref_T1_t1Probe_laneProbes_2_slots_0_slotOccupied verification.probeWire_laneProbes_2_slots_0_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_2_slots_0_pipeFinish verification.probeWire_laneProbes_2_slots_0_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_2_slots_0_slotShiftValid verification.probeWire_laneProbes_2_slots_0_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_2_slots_0_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_2_slots_0_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_2_slots_0_decodeResultIsScheduler verification.probeWire_laneProbes_2_slots_0_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_2_slots_0_executionUnitVfuRequestReady verification.probeWire_laneProbes_2_slots_0_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_2_slots_0_executionUnitVfuRequestValid verification.probeWire_laneProbes_2_slots_0_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_2_slots_0_stage3VrfWriteReady verification.probeWire_laneProbes_2_slots_0_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_2_slots_0_stage3VrfWriteValid verification.probeWire_laneProbes_2_slots_0_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_2_slots_0_writeQueueEnq verification.probeWire_laneProbes_2_slots_0_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_2_slots_0_writeTag verification.probeWire_laneProbes_2_slots_0_writeTag_probe
`define ref_T1_t1Probe_laneProbes_2_slots_0_writeMask verification.probeWire_laneProbes_2_slots_0_writeMask_probe
`define ref_T1_t1Probe_laneProbes_2_slots_1_stage0EnqueueReady verification.probeWire_laneProbes_2_slots_1_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_2_slots_1_stage0EnqueueValid verification.probeWire_laneProbes_2_slots_1_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_2_slots_1_changingMaskSet verification.probeWire_laneProbes_2_slots_1_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_2_slots_1_slotActive verification.probeWire_laneProbes_2_slots_1_slotActive_probe
`define ref_T1_t1Probe_laneProbes_2_slots_1_slotOccupied verification.probeWire_laneProbes_2_slots_1_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_2_slots_1_pipeFinish verification.probeWire_laneProbes_2_slots_1_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_2_slots_1_slotShiftValid verification.probeWire_laneProbes_2_slots_1_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_2_slots_1_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_2_slots_1_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_2_slots_1_decodeResultIsScheduler verification.probeWire_laneProbes_2_slots_1_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_2_slots_1_executionUnitVfuRequestReady verification.probeWire_laneProbes_2_slots_1_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_2_slots_1_executionUnitVfuRequestValid verification.probeWire_laneProbes_2_slots_1_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_2_slots_1_stage3VrfWriteReady verification.probeWire_laneProbes_2_slots_1_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_2_slots_1_stage3VrfWriteValid verification.probeWire_laneProbes_2_slots_1_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_2_slots_1_writeQueueEnq verification.probeWire_laneProbes_2_slots_1_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_2_slots_1_writeTag verification.probeWire_laneProbes_2_slots_1_writeTag_probe
`define ref_T1_t1Probe_laneProbes_2_slots_1_writeMask verification.probeWire_laneProbes_2_slots_1_writeMask_probe
`define ref_T1_t1Probe_laneProbes_2_slots_2_stage0EnqueueReady verification.probeWire_laneProbes_2_slots_2_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_2_slots_2_stage0EnqueueValid verification.probeWire_laneProbes_2_slots_2_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_2_slots_2_changingMaskSet verification.probeWire_laneProbes_2_slots_2_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_2_slots_2_slotActive verification.probeWire_laneProbes_2_slots_2_slotActive_probe
`define ref_T1_t1Probe_laneProbes_2_slots_2_slotOccupied verification.probeWire_laneProbes_2_slots_2_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_2_slots_2_pipeFinish verification.probeWire_laneProbes_2_slots_2_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_2_slots_2_slotShiftValid verification.probeWire_laneProbes_2_slots_2_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_2_slots_2_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_2_slots_2_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_2_slots_2_decodeResultIsScheduler verification.probeWire_laneProbes_2_slots_2_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_2_slots_2_executionUnitVfuRequestReady verification.probeWire_laneProbes_2_slots_2_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_2_slots_2_executionUnitVfuRequestValid verification.probeWire_laneProbes_2_slots_2_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_2_slots_2_stage3VrfWriteReady verification.probeWire_laneProbes_2_slots_2_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_2_slots_2_stage3VrfWriteValid verification.probeWire_laneProbes_2_slots_2_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_2_slots_2_writeQueueEnq verification.probeWire_laneProbes_2_slots_2_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_2_slots_2_writeTag verification.probeWire_laneProbes_2_slots_2_writeTag_probe
`define ref_T1_t1Probe_laneProbes_2_slots_2_writeMask verification.probeWire_laneProbes_2_slots_2_writeMask_probe
`define ref_T1_t1Probe_laneProbes_2_slots_3_stage0EnqueueReady verification.probeWire_laneProbes_2_slots_3_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_2_slots_3_stage0EnqueueValid verification.probeWire_laneProbes_2_slots_3_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_2_slots_3_changingMaskSet verification.probeWire_laneProbes_2_slots_3_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_2_slots_3_slotActive verification.probeWire_laneProbes_2_slots_3_slotActive_probe
`define ref_T1_t1Probe_laneProbes_2_slots_3_slotOccupied verification.probeWire_laneProbes_2_slots_3_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_2_slots_3_pipeFinish verification.probeWire_laneProbes_2_slots_3_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_2_slots_3_slotShiftValid verification.probeWire_laneProbes_2_slots_3_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_2_slots_3_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_2_slots_3_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_2_slots_3_decodeResultIsScheduler verification.probeWire_laneProbes_2_slots_3_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_2_slots_3_executionUnitVfuRequestReady verification.probeWire_laneProbes_2_slots_3_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_2_slots_3_executionUnitVfuRequestValid verification.probeWire_laneProbes_2_slots_3_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_2_slots_3_stage3VrfWriteReady verification.probeWire_laneProbes_2_slots_3_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_2_slots_3_stage3VrfWriteValid verification.probeWire_laneProbes_2_slots_3_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_2_slots_3_writeQueueEnq verification.probeWire_laneProbes_2_slots_3_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_2_slots_3_writeTag verification.probeWire_laneProbes_2_slots_3_writeTag_probe
`define ref_T1_t1Probe_laneProbes_2_slots_3_writeMask verification.probeWire_laneProbes_2_slots_3_writeMask_probe
`define ref_T1_t1Probe_laneProbes_2_laneRequestStall verification.probeWire_laneProbes_2_laneRequestStall_probe
`define ref_T1_t1Probe_laneProbes_2_lastSlotOccupied verification.probeWire_laneProbes_2_lastSlotOccupied_probe
`define ref_T1_t1Probe_laneProbes_2_instructionFinished verification.probeWire_laneProbes_2_instructionFinished_probe
`define ref_T1_t1Probe_laneProbes_2_instructionValid verification.probeWire_laneProbes_2_instructionValid_probe
`define ref_T1_t1Probe_laneProbes_2_crossWriteProbe_0_valid verification.probeWire_laneProbes_2_crossWriteProbe_0_valid_probe
`define ref_T1_t1Probe_laneProbes_2_crossWriteProbe_0_bits_writeTag verification.probeWire_laneProbes_2_crossWriteProbe_0_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_2_crossWriteProbe_0_bits_writeMask verification.probeWire_laneProbes_2_crossWriteProbe_0_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_2_crossWriteProbe_1_valid verification.probeWire_laneProbes_2_crossWriteProbe_1_valid_probe
`define ref_T1_t1Probe_laneProbes_2_crossWriteProbe_1_bits_writeTag verification.probeWire_laneProbes_2_crossWriteProbe_1_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_2_crossWriteProbe_1_bits_writeMask verification.probeWire_laneProbes_2_crossWriteProbe_1_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_2_vrfProbe_valid verification.probeWire_laneProbes_2_vrfProbe_valid_probe
`define ref_T1_t1Probe_laneProbes_2_vrfProbe_requestVd verification.probeWire_laneProbes_2_vrfProbe_requestVd_probe
`define ref_T1_t1Probe_laneProbes_2_vrfProbe_requestOffset verification.probeWire_laneProbes_2_vrfProbe_requestOffset_probe
`define ref_T1_t1Probe_laneProbes_2_vrfProbe_requestMask verification.probeWire_laneProbes_2_vrfProbe_requestMask_probe
`define ref_T1_t1Probe_laneProbes_2_vrfProbe_requestData verification.probeWire_laneProbes_2_vrfProbe_requestData_probe
`define ref_T1_t1Probe_laneProbes_2_vrfProbe_requestInstruction verification.probeWire_laneProbes_2_vrfProbe_requestInstruction_probe
`define ref_T1_t1Probe_laneProbes_3_slots_0_stage0EnqueueReady verification.probeWire_laneProbes_3_slots_0_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_3_slots_0_stage0EnqueueValid verification.probeWire_laneProbes_3_slots_0_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_3_slots_0_changingMaskSet verification.probeWire_laneProbes_3_slots_0_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_3_slots_0_slotActive verification.probeWire_laneProbes_3_slots_0_slotActive_probe
`define ref_T1_t1Probe_laneProbes_3_slots_0_slotOccupied verification.probeWire_laneProbes_3_slots_0_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_3_slots_0_pipeFinish verification.probeWire_laneProbes_3_slots_0_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_3_slots_0_slotShiftValid verification.probeWire_laneProbes_3_slots_0_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_3_slots_0_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_3_slots_0_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_3_slots_0_decodeResultIsScheduler verification.probeWire_laneProbes_3_slots_0_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_3_slots_0_executionUnitVfuRequestReady verification.probeWire_laneProbes_3_slots_0_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_3_slots_0_executionUnitVfuRequestValid verification.probeWire_laneProbes_3_slots_0_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_3_slots_0_stage3VrfWriteReady verification.probeWire_laneProbes_3_slots_0_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_3_slots_0_stage3VrfWriteValid verification.probeWire_laneProbes_3_slots_0_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_3_slots_0_writeQueueEnq verification.probeWire_laneProbes_3_slots_0_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_3_slots_0_writeTag verification.probeWire_laneProbes_3_slots_0_writeTag_probe
`define ref_T1_t1Probe_laneProbes_3_slots_0_writeMask verification.probeWire_laneProbes_3_slots_0_writeMask_probe
`define ref_T1_t1Probe_laneProbes_3_slots_1_stage0EnqueueReady verification.probeWire_laneProbes_3_slots_1_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_3_slots_1_stage0EnqueueValid verification.probeWire_laneProbes_3_slots_1_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_3_slots_1_changingMaskSet verification.probeWire_laneProbes_3_slots_1_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_3_slots_1_slotActive verification.probeWire_laneProbes_3_slots_1_slotActive_probe
`define ref_T1_t1Probe_laneProbes_3_slots_1_slotOccupied verification.probeWire_laneProbes_3_slots_1_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_3_slots_1_pipeFinish verification.probeWire_laneProbes_3_slots_1_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_3_slots_1_slotShiftValid verification.probeWire_laneProbes_3_slots_1_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_3_slots_1_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_3_slots_1_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_3_slots_1_decodeResultIsScheduler verification.probeWire_laneProbes_3_slots_1_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_3_slots_1_executionUnitVfuRequestReady verification.probeWire_laneProbes_3_slots_1_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_3_slots_1_executionUnitVfuRequestValid verification.probeWire_laneProbes_3_slots_1_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_3_slots_1_stage3VrfWriteReady verification.probeWire_laneProbes_3_slots_1_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_3_slots_1_stage3VrfWriteValid verification.probeWire_laneProbes_3_slots_1_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_3_slots_1_writeQueueEnq verification.probeWire_laneProbes_3_slots_1_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_3_slots_1_writeTag verification.probeWire_laneProbes_3_slots_1_writeTag_probe
`define ref_T1_t1Probe_laneProbes_3_slots_1_writeMask verification.probeWire_laneProbes_3_slots_1_writeMask_probe
`define ref_T1_t1Probe_laneProbes_3_slots_2_stage0EnqueueReady verification.probeWire_laneProbes_3_slots_2_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_3_slots_2_stage0EnqueueValid verification.probeWire_laneProbes_3_slots_2_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_3_slots_2_changingMaskSet verification.probeWire_laneProbes_3_slots_2_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_3_slots_2_slotActive verification.probeWire_laneProbes_3_slots_2_slotActive_probe
`define ref_T1_t1Probe_laneProbes_3_slots_2_slotOccupied verification.probeWire_laneProbes_3_slots_2_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_3_slots_2_pipeFinish verification.probeWire_laneProbes_3_slots_2_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_3_slots_2_slotShiftValid verification.probeWire_laneProbes_3_slots_2_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_3_slots_2_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_3_slots_2_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_3_slots_2_decodeResultIsScheduler verification.probeWire_laneProbes_3_slots_2_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_3_slots_2_executionUnitVfuRequestReady verification.probeWire_laneProbes_3_slots_2_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_3_slots_2_executionUnitVfuRequestValid verification.probeWire_laneProbes_3_slots_2_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_3_slots_2_stage3VrfWriteReady verification.probeWire_laneProbes_3_slots_2_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_3_slots_2_stage3VrfWriteValid verification.probeWire_laneProbes_3_slots_2_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_3_slots_2_writeQueueEnq verification.probeWire_laneProbes_3_slots_2_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_3_slots_2_writeTag verification.probeWire_laneProbes_3_slots_2_writeTag_probe
`define ref_T1_t1Probe_laneProbes_3_slots_2_writeMask verification.probeWire_laneProbes_3_slots_2_writeMask_probe
`define ref_T1_t1Probe_laneProbes_3_slots_3_stage0EnqueueReady verification.probeWire_laneProbes_3_slots_3_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_3_slots_3_stage0EnqueueValid verification.probeWire_laneProbes_3_slots_3_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_3_slots_3_changingMaskSet verification.probeWire_laneProbes_3_slots_3_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_3_slots_3_slotActive verification.probeWire_laneProbes_3_slots_3_slotActive_probe
`define ref_T1_t1Probe_laneProbes_3_slots_3_slotOccupied verification.probeWire_laneProbes_3_slots_3_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_3_slots_3_pipeFinish verification.probeWire_laneProbes_3_slots_3_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_3_slots_3_slotShiftValid verification.probeWire_laneProbes_3_slots_3_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_3_slots_3_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_3_slots_3_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_3_slots_3_decodeResultIsScheduler verification.probeWire_laneProbes_3_slots_3_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_3_slots_3_executionUnitVfuRequestReady verification.probeWire_laneProbes_3_slots_3_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_3_slots_3_executionUnitVfuRequestValid verification.probeWire_laneProbes_3_slots_3_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_3_slots_3_stage3VrfWriteReady verification.probeWire_laneProbes_3_slots_3_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_3_slots_3_stage3VrfWriteValid verification.probeWire_laneProbes_3_slots_3_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_3_slots_3_writeQueueEnq verification.probeWire_laneProbes_3_slots_3_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_3_slots_3_writeTag verification.probeWire_laneProbes_3_slots_3_writeTag_probe
`define ref_T1_t1Probe_laneProbes_3_slots_3_writeMask verification.probeWire_laneProbes_3_slots_3_writeMask_probe
`define ref_T1_t1Probe_laneProbes_3_laneRequestStall verification.probeWire_laneProbes_3_laneRequestStall_probe
`define ref_T1_t1Probe_laneProbes_3_lastSlotOccupied verification.probeWire_laneProbes_3_lastSlotOccupied_probe
`define ref_T1_t1Probe_laneProbes_3_instructionFinished verification.probeWire_laneProbes_3_instructionFinished_probe
`define ref_T1_t1Probe_laneProbes_3_instructionValid verification.probeWire_laneProbes_3_instructionValid_probe
`define ref_T1_t1Probe_laneProbes_3_crossWriteProbe_0_valid verification.probeWire_laneProbes_3_crossWriteProbe_0_valid_probe
`define ref_T1_t1Probe_laneProbes_3_crossWriteProbe_0_bits_writeTag verification.probeWire_laneProbes_3_crossWriteProbe_0_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_3_crossWriteProbe_0_bits_writeMask verification.probeWire_laneProbes_3_crossWriteProbe_0_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_3_crossWriteProbe_1_valid verification.probeWire_laneProbes_3_crossWriteProbe_1_valid_probe
`define ref_T1_t1Probe_laneProbes_3_crossWriteProbe_1_bits_writeTag verification.probeWire_laneProbes_3_crossWriteProbe_1_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_3_crossWriteProbe_1_bits_writeMask verification.probeWire_laneProbes_3_crossWriteProbe_1_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_3_vrfProbe_valid verification.probeWire_laneProbes_3_vrfProbe_valid_probe
`define ref_T1_t1Probe_laneProbes_3_vrfProbe_requestVd verification.probeWire_laneProbes_3_vrfProbe_requestVd_probe
`define ref_T1_t1Probe_laneProbes_3_vrfProbe_requestOffset verification.probeWire_laneProbes_3_vrfProbe_requestOffset_probe
`define ref_T1_t1Probe_laneProbes_3_vrfProbe_requestMask verification.probeWire_laneProbes_3_vrfProbe_requestMask_probe
`define ref_T1_t1Probe_laneProbes_3_vrfProbe_requestData verification.probeWire_laneProbes_3_vrfProbe_requestData_probe
`define ref_T1_t1Probe_laneProbes_3_vrfProbe_requestInstruction verification.probeWire_laneProbes_3_vrfProbe_requestInstruction_probe
`define ref_T1_t1Probe_laneProbes_4_slots_0_stage0EnqueueReady verification.probeWire_laneProbes_4_slots_0_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_4_slots_0_stage0EnqueueValid verification.probeWire_laneProbes_4_slots_0_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_4_slots_0_changingMaskSet verification.probeWire_laneProbes_4_slots_0_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_4_slots_0_slotActive verification.probeWire_laneProbes_4_slots_0_slotActive_probe
`define ref_T1_t1Probe_laneProbes_4_slots_0_slotOccupied verification.probeWire_laneProbes_4_slots_0_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_4_slots_0_pipeFinish verification.probeWire_laneProbes_4_slots_0_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_4_slots_0_slotShiftValid verification.probeWire_laneProbes_4_slots_0_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_4_slots_0_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_4_slots_0_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_4_slots_0_decodeResultIsScheduler verification.probeWire_laneProbes_4_slots_0_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_4_slots_0_executionUnitVfuRequestReady verification.probeWire_laneProbes_4_slots_0_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_4_slots_0_executionUnitVfuRequestValid verification.probeWire_laneProbes_4_slots_0_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_4_slots_0_stage3VrfWriteReady verification.probeWire_laneProbes_4_slots_0_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_4_slots_0_stage3VrfWriteValid verification.probeWire_laneProbes_4_slots_0_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_4_slots_0_writeQueueEnq verification.probeWire_laneProbes_4_slots_0_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_4_slots_0_writeTag verification.probeWire_laneProbes_4_slots_0_writeTag_probe
`define ref_T1_t1Probe_laneProbes_4_slots_0_writeMask verification.probeWire_laneProbes_4_slots_0_writeMask_probe
`define ref_T1_t1Probe_laneProbes_4_slots_1_stage0EnqueueReady verification.probeWire_laneProbes_4_slots_1_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_4_slots_1_stage0EnqueueValid verification.probeWire_laneProbes_4_slots_1_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_4_slots_1_changingMaskSet verification.probeWire_laneProbes_4_slots_1_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_4_slots_1_slotActive verification.probeWire_laneProbes_4_slots_1_slotActive_probe
`define ref_T1_t1Probe_laneProbes_4_slots_1_slotOccupied verification.probeWire_laneProbes_4_slots_1_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_4_slots_1_pipeFinish verification.probeWire_laneProbes_4_slots_1_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_4_slots_1_slotShiftValid verification.probeWire_laneProbes_4_slots_1_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_4_slots_1_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_4_slots_1_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_4_slots_1_decodeResultIsScheduler verification.probeWire_laneProbes_4_slots_1_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_4_slots_1_executionUnitVfuRequestReady verification.probeWire_laneProbes_4_slots_1_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_4_slots_1_executionUnitVfuRequestValid verification.probeWire_laneProbes_4_slots_1_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_4_slots_1_stage3VrfWriteReady verification.probeWire_laneProbes_4_slots_1_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_4_slots_1_stage3VrfWriteValid verification.probeWire_laneProbes_4_slots_1_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_4_slots_1_writeQueueEnq verification.probeWire_laneProbes_4_slots_1_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_4_slots_1_writeTag verification.probeWire_laneProbes_4_slots_1_writeTag_probe
`define ref_T1_t1Probe_laneProbes_4_slots_1_writeMask verification.probeWire_laneProbes_4_slots_1_writeMask_probe
`define ref_T1_t1Probe_laneProbes_4_slots_2_stage0EnqueueReady verification.probeWire_laneProbes_4_slots_2_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_4_slots_2_stage0EnqueueValid verification.probeWire_laneProbes_4_slots_2_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_4_slots_2_changingMaskSet verification.probeWire_laneProbes_4_slots_2_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_4_slots_2_slotActive verification.probeWire_laneProbes_4_slots_2_slotActive_probe
`define ref_T1_t1Probe_laneProbes_4_slots_2_slotOccupied verification.probeWire_laneProbes_4_slots_2_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_4_slots_2_pipeFinish verification.probeWire_laneProbes_4_slots_2_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_4_slots_2_slotShiftValid verification.probeWire_laneProbes_4_slots_2_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_4_slots_2_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_4_slots_2_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_4_slots_2_decodeResultIsScheduler verification.probeWire_laneProbes_4_slots_2_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_4_slots_2_executionUnitVfuRequestReady verification.probeWire_laneProbes_4_slots_2_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_4_slots_2_executionUnitVfuRequestValid verification.probeWire_laneProbes_4_slots_2_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_4_slots_2_stage3VrfWriteReady verification.probeWire_laneProbes_4_slots_2_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_4_slots_2_stage3VrfWriteValid verification.probeWire_laneProbes_4_slots_2_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_4_slots_2_writeQueueEnq verification.probeWire_laneProbes_4_slots_2_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_4_slots_2_writeTag verification.probeWire_laneProbes_4_slots_2_writeTag_probe
`define ref_T1_t1Probe_laneProbes_4_slots_2_writeMask verification.probeWire_laneProbes_4_slots_2_writeMask_probe
`define ref_T1_t1Probe_laneProbes_4_slots_3_stage0EnqueueReady verification.probeWire_laneProbes_4_slots_3_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_4_slots_3_stage0EnqueueValid verification.probeWire_laneProbes_4_slots_3_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_4_slots_3_changingMaskSet verification.probeWire_laneProbes_4_slots_3_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_4_slots_3_slotActive verification.probeWire_laneProbes_4_slots_3_slotActive_probe
`define ref_T1_t1Probe_laneProbes_4_slots_3_slotOccupied verification.probeWire_laneProbes_4_slots_3_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_4_slots_3_pipeFinish verification.probeWire_laneProbes_4_slots_3_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_4_slots_3_slotShiftValid verification.probeWire_laneProbes_4_slots_3_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_4_slots_3_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_4_slots_3_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_4_slots_3_decodeResultIsScheduler verification.probeWire_laneProbes_4_slots_3_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_4_slots_3_executionUnitVfuRequestReady verification.probeWire_laneProbes_4_slots_3_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_4_slots_3_executionUnitVfuRequestValid verification.probeWire_laneProbes_4_slots_3_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_4_slots_3_stage3VrfWriteReady verification.probeWire_laneProbes_4_slots_3_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_4_slots_3_stage3VrfWriteValid verification.probeWire_laneProbes_4_slots_3_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_4_slots_3_writeQueueEnq verification.probeWire_laneProbes_4_slots_3_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_4_slots_3_writeTag verification.probeWire_laneProbes_4_slots_3_writeTag_probe
`define ref_T1_t1Probe_laneProbes_4_slots_3_writeMask verification.probeWire_laneProbes_4_slots_3_writeMask_probe
`define ref_T1_t1Probe_laneProbes_4_laneRequestStall verification.probeWire_laneProbes_4_laneRequestStall_probe
`define ref_T1_t1Probe_laneProbes_4_lastSlotOccupied verification.probeWire_laneProbes_4_lastSlotOccupied_probe
`define ref_T1_t1Probe_laneProbes_4_instructionFinished verification.probeWire_laneProbes_4_instructionFinished_probe
`define ref_T1_t1Probe_laneProbes_4_instructionValid verification.probeWire_laneProbes_4_instructionValid_probe
`define ref_T1_t1Probe_laneProbes_4_crossWriteProbe_0_valid verification.probeWire_laneProbes_4_crossWriteProbe_0_valid_probe
`define ref_T1_t1Probe_laneProbes_4_crossWriteProbe_0_bits_writeTag verification.probeWire_laneProbes_4_crossWriteProbe_0_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_4_crossWriteProbe_0_bits_writeMask verification.probeWire_laneProbes_4_crossWriteProbe_0_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_4_crossWriteProbe_1_valid verification.probeWire_laneProbes_4_crossWriteProbe_1_valid_probe
`define ref_T1_t1Probe_laneProbes_4_crossWriteProbe_1_bits_writeTag verification.probeWire_laneProbes_4_crossWriteProbe_1_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_4_crossWriteProbe_1_bits_writeMask verification.probeWire_laneProbes_4_crossWriteProbe_1_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_4_vrfProbe_valid verification.probeWire_laneProbes_4_vrfProbe_valid_probe
`define ref_T1_t1Probe_laneProbes_4_vrfProbe_requestVd verification.probeWire_laneProbes_4_vrfProbe_requestVd_probe
`define ref_T1_t1Probe_laneProbes_4_vrfProbe_requestOffset verification.probeWire_laneProbes_4_vrfProbe_requestOffset_probe
`define ref_T1_t1Probe_laneProbes_4_vrfProbe_requestMask verification.probeWire_laneProbes_4_vrfProbe_requestMask_probe
`define ref_T1_t1Probe_laneProbes_4_vrfProbe_requestData verification.probeWire_laneProbes_4_vrfProbe_requestData_probe
`define ref_T1_t1Probe_laneProbes_4_vrfProbe_requestInstruction verification.probeWire_laneProbes_4_vrfProbe_requestInstruction_probe
`define ref_T1_t1Probe_laneProbes_5_slots_0_stage0EnqueueReady verification.probeWire_laneProbes_5_slots_0_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_5_slots_0_stage0EnqueueValid verification.probeWire_laneProbes_5_slots_0_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_5_slots_0_changingMaskSet verification.probeWire_laneProbes_5_slots_0_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_5_slots_0_slotActive verification.probeWire_laneProbes_5_slots_0_slotActive_probe
`define ref_T1_t1Probe_laneProbes_5_slots_0_slotOccupied verification.probeWire_laneProbes_5_slots_0_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_5_slots_0_pipeFinish verification.probeWire_laneProbes_5_slots_0_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_5_slots_0_slotShiftValid verification.probeWire_laneProbes_5_slots_0_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_5_slots_0_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_5_slots_0_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_5_slots_0_decodeResultIsScheduler verification.probeWire_laneProbes_5_slots_0_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_5_slots_0_executionUnitVfuRequestReady verification.probeWire_laneProbes_5_slots_0_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_5_slots_0_executionUnitVfuRequestValid verification.probeWire_laneProbes_5_slots_0_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_5_slots_0_stage3VrfWriteReady verification.probeWire_laneProbes_5_slots_0_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_5_slots_0_stage3VrfWriteValid verification.probeWire_laneProbes_5_slots_0_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_5_slots_0_writeQueueEnq verification.probeWire_laneProbes_5_slots_0_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_5_slots_0_writeTag verification.probeWire_laneProbes_5_slots_0_writeTag_probe
`define ref_T1_t1Probe_laneProbes_5_slots_0_writeMask verification.probeWire_laneProbes_5_slots_0_writeMask_probe
`define ref_T1_t1Probe_laneProbes_5_slots_1_stage0EnqueueReady verification.probeWire_laneProbes_5_slots_1_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_5_slots_1_stage0EnqueueValid verification.probeWire_laneProbes_5_slots_1_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_5_slots_1_changingMaskSet verification.probeWire_laneProbes_5_slots_1_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_5_slots_1_slotActive verification.probeWire_laneProbes_5_slots_1_slotActive_probe
`define ref_T1_t1Probe_laneProbes_5_slots_1_slotOccupied verification.probeWire_laneProbes_5_slots_1_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_5_slots_1_pipeFinish verification.probeWire_laneProbes_5_slots_1_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_5_slots_1_slotShiftValid verification.probeWire_laneProbes_5_slots_1_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_5_slots_1_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_5_slots_1_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_5_slots_1_decodeResultIsScheduler verification.probeWire_laneProbes_5_slots_1_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_5_slots_1_executionUnitVfuRequestReady verification.probeWire_laneProbes_5_slots_1_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_5_slots_1_executionUnitVfuRequestValid verification.probeWire_laneProbes_5_slots_1_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_5_slots_1_stage3VrfWriteReady verification.probeWire_laneProbes_5_slots_1_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_5_slots_1_stage3VrfWriteValid verification.probeWire_laneProbes_5_slots_1_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_5_slots_1_writeQueueEnq verification.probeWire_laneProbes_5_slots_1_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_5_slots_1_writeTag verification.probeWire_laneProbes_5_slots_1_writeTag_probe
`define ref_T1_t1Probe_laneProbes_5_slots_1_writeMask verification.probeWire_laneProbes_5_slots_1_writeMask_probe
`define ref_T1_t1Probe_laneProbes_5_slots_2_stage0EnqueueReady verification.probeWire_laneProbes_5_slots_2_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_5_slots_2_stage0EnqueueValid verification.probeWire_laneProbes_5_slots_2_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_5_slots_2_changingMaskSet verification.probeWire_laneProbes_5_slots_2_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_5_slots_2_slotActive verification.probeWire_laneProbes_5_slots_2_slotActive_probe
`define ref_T1_t1Probe_laneProbes_5_slots_2_slotOccupied verification.probeWire_laneProbes_5_slots_2_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_5_slots_2_pipeFinish verification.probeWire_laneProbes_5_slots_2_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_5_slots_2_slotShiftValid verification.probeWire_laneProbes_5_slots_2_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_5_slots_2_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_5_slots_2_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_5_slots_2_decodeResultIsScheduler verification.probeWire_laneProbes_5_slots_2_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_5_slots_2_executionUnitVfuRequestReady verification.probeWire_laneProbes_5_slots_2_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_5_slots_2_executionUnitVfuRequestValid verification.probeWire_laneProbes_5_slots_2_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_5_slots_2_stage3VrfWriteReady verification.probeWire_laneProbes_5_slots_2_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_5_slots_2_stage3VrfWriteValid verification.probeWire_laneProbes_5_slots_2_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_5_slots_2_writeQueueEnq verification.probeWire_laneProbes_5_slots_2_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_5_slots_2_writeTag verification.probeWire_laneProbes_5_slots_2_writeTag_probe
`define ref_T1_t1Probe_laneProbes_5_slots_2_writeMask verification.probeWire_laneProbes_5_slots_2_writeMask_probe
`define ref_T1_t1Probe_laneProbes_5_slots_3_stage0EnqueueReady verification.probeWire_laneProbes_5_slots_3_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_5_slots_3_stage0EnqueueValid verification.probeWire_laneProbes_5_slots_3_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_5_slots_3_changingMaskSet verification.probeWire_laneProbes_5_slots_3_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_5_slots_3_slotActive verification.probeWire_laneProbes_5_slots_3_slotActive_probe
`define ref_T1_t1Probe_laneProbes_5_slots_3_slotOccupied verification.probeWire_laneProbes_5_slots_3_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_5_slots_3_pipeFinish verification.probeWire_laneProbes_5_slots_3_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_5_slots_3_slotShiftValid verification.probeWire_laneProbes_5_slots_3_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_5_slots_3_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_5_slots_3_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_5_slots_3_decodeResultIsScheduler verification.probeWire_laneProbes_5_slots_3_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_5_slots_3_executionUnitVfuRequestReady verification.probeWire_laneProbes_5_slots_3_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_5_slots_3_executionUnitVfuRequestValid verification.probeWire_laneProbes_5_slots_3_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_5_slots_3_stage3VrfWriteReady verification.probeWire_laneProbes_5_slots_3_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_5_slots_3_stage3VrfWriteValid verification.probeWire_laneProbes_5_slots_3_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_5_slots_3_writeQueueEnq verification.probeWire_laneProbes_5_slots_3_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_5_slots_3_writeTag verification.probeWire_laneProbes_5_slots_3_writeTag_probe
`define ref_T1_t1Probe_laneProbes_5_slots_3_writeMask verification.probeWire_laneProbes_5_slots_3_writeMask_probe
`define ref_T1_t1Probe_laneProbes_5_laneRequestStall verification.probeWire_laneProbes_5_laneRequestStall_probe
`define ref_T1_t1Probe_laneProbes_5_lastSlotOccupied verification.probeWire_laneProbes_5_lastSlotOccupied_probe
`define ref_T1_t1Probe_laneProbes_5_instructionFinished verification.probeWire_laneProbes_5_instructionFinished_probe
`define ref_T1_t1Probe_laneProbes_5_instructionValid verification.probeWire_laneProbes_5_instructionValid_probe
`define ref_T1_t1Probe_laneProbes_5_crossWriteProbe_0_valid verification.probeWire_laneProbes_5_crossWriteProbe_0_valid_probe
`define ref_T1_t1Probe_laneProbes_5_crossWriteProbe_0_bits_writeTag verification.probeWire_laneProbes_5_crossWriteProbe_0_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_5_crossWriteProbe_0_bits_writeMask verification.probeWire_laneProbes_5_crossWriteProbe_0_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_5_crossWriteProbe_1_valid verification.probeWire_laneProbes_5_crossWriteProbe_1_valid_probe
`define ref_T1_t1Probe_laneProbes_5_crossWriteProbe_1_bits_writeTag verification.probeWire_laneProbes_5_crossWriteProbe_1_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_5_crossWriteProbe_1_bits_writeMask verification.probeWire_laneProbes_5_crossWriteProbe_1_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_5_vrfProbe_valid verification.probeWire_laneProbes_5_vrfProbe_valid_probe
`define ref_T1_t1Probe_laneProbes_5_vrfProbe_requestVd verification.probeWire_laneProbes_5_vrfProbe_requestVd_probe
`define ref_T1_t1Probe_laneProbes_5_vrfProbe_requestOffset verification.probeWire_laneProbes_5_vrfProbe_requestOffset_probe
`define ref_T1_t1Probe_laneProbes_5_vrfProbe_requestMask verification.probeWire_laneProbes_5_vrfProbe_requestMask_probe
`define ref_T1_t1Probe_laneProbes_5_vrfProbe_requestData verification.probeWire_laneProbes_5_vrfProbe_requestData_probe
`define ref_T1_t1Probe_laneProbes_5_vrfProbe_requestInstruction verification.probeWire_laneProbes_5_vrfProbe_requestInstruction_probe
`define ref_T1_t1Probe_laneProbes_6_slots_0_stage0EnqueueReady verification.probeWire_laneProbes_6_slots_0_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_6_slots_0_stage0EnqueueValid verification.probeWire_laneProbes_6_slots_0_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_6_slots_0_changingMaskSet verification.probeWire_laneProbes_6_slots_0_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_6_slots_0_slotActive verification.probeWire_laneProbes_6_slots_0_slotActive_probe
`define ref_T1_t1Probe_laneProbes_6_slots_0_slotOccupied verification.probeWire_laneProbes_6_slots_0_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_6_slots_0_pipeFinish verification.probeWire_laneProbes_6_slots_0_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_6_slots_0_slotShiftValid verification.probeWire_laneProbes_6_slots_0_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_6_slots_0_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_6_slots_0_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_6_slots_0_decodeResultIsScheduler verification.probeWire_laneProbes_6_slots_0_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_6_slots_0_executionUnitVfuRequestReady verification.probeWire_laneProbes_6_slots_0_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_6_slots_0_executionUnitVfuRequestValid verification.probeWire_laneProbes_6_slots_0_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_6_slots_0_stage3VrfWriteReady verification.probeWire_laneProbes_6_slots_0_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_6_slots_0_stage3VrfWriteValid verification.probeWire_laneProbes_6_slots_0_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_6_slots_0_writeQueueEnq verification.probeWire_laneProbes_6_slots_0_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_6_slots_0_writeTag verification.probeWire_laneProbes_6_slots_0_writeTag_probe
`define ref_T1_t1Probe_laneProbes_6_slots_0_writeMask verification.probeWire_laneProbes_6_slots_0_writeMask_probe
`define ref_T1_t1Probe_laneProbes_6_slots_1_stage0EnqueueReady verification.probeWire_laneProbes_6_slots_1_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_6_slots_1_stage0EnqueueValid verification.probeWire_laneProbes_6_slots_1_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_6_slots_1_changingMaskSet verification.probeWire_laneProbes_6_slots_1_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_6_slots_1_slotActive verification.probeWire_laneProbes_6_slots_1_slotActive_probe
`define ref_T1_t1Probe_laneProbes_6_slots_1_slotOccupied verification.probeWire_laneProbes_6_slots_1_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_6_slots_1_pipeFinish verification.probeWire_laneProbes_6_slots_1_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_6_slots_1_slotShiftValid verification.probeWire_laneProbes_6_slots_1_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_6_slots_1_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_6_slots_1_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_6_slots_1_decodeResultIsScheduler verification.probeWire_laneProbes_6_slots_1_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_6_slots_1_executionUnitVfuRequestReady verification.probeWire_laneProbes_6_slots_1_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_6_slots_1_executionUnitVfuRequestValid verification.probeWire_laneProbes_6_slots_1_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_6_slots_1_stage3VrfWriteReady verification.probeWire_laneProbes_6_slots_1_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_6_slots_1_stage3VrfWriteValid verification.probeWire_laneProbes_6_slots_1_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_6_slots_1_writeQueueEnq verification.probeWire_laneProbes_6_slots_1_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_6_slots_1_writeTag verification.probeWire_laneProbes_6_slots_1_writeTag_probe
`define ref_T1_t1Probe_laneProbes_6_slots_1_writeMask verification.probeWire_laneProbes_6_slots_1_writeMask_probe
`define ref_T1_t1Probe_laneProbes_6_slots_2_stage0EnqueueReady verification.probeWire_laneProbes_6_slots_2_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_6_slots_2_stage0EnqueueValid verification.probeWire_laneProbes_6_slots_2_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_6_slots_2_changingMaskSet verification.probeWire_laneProbes_6_slots_2_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_6_slots_2_slotActive verification.probeWire_laneProbes_6_slots_2_slotActive_probe
`define ref_T1_t1Probe_laneProbes_6_slots_2_slotOccupied verification.probeWire_laneProbes_6_slots_2_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_6_slots_2_pipeFinish verification.probeWire_laneProbes_6_slots_2_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_6_slots_2_slotShiftValid verification.probeWire_laneProbes_6_slots_2_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_6_slots_2_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_6_slots_2_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_6_slots_2_decodeResultIsScheduler verification.probeWire_laneProbes_6_slots_2_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_6_slots_2_executionUnitVfuRequestReady verification.probeWire_laneProbes_6_slots_2_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_6_slots_2_executionUnitVfuRequestValid verification.probeWire_laneProbes_6_slots_2_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_6_slots_2_stage3VrfWriteReady verification.probeWire_laneProbes_6_slots_2_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_6_slots_2_stage3VrfWriteValid verification.probeWire_laneProbes_6_slots_2_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_6_slots_2_writeQueueEnq verification.probeWire_laneProbes_6_slots_2_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_6_slots_2_writeTag verification.probeWire_laneProbes_6_slots_2_writeTag_probe
`define ref_T1_t1Probe_laneProbes_6_slots_2_writeMask verification.probeWire_laneProbes_6_slots_2_writeMask_probe
`define ref_T1_t1Probe_laneProbes_6_slots_3_stage0EnqueueReady verification.probeWire_laneProbes_6_slots_3_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_6_slots_3_stage0EnqueueValid verification.probeWire_laneProbes_6_slots_3_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_6_slots_3_changingMaskSet verification.probeWire_laneProbes_6_slots_3_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_6_slots_3_slotActive verification.probeWire_laneProbes_6_slots_3_slotActive_probe
`define ref_T1_t1Probe_laneProbes_6_slots_3_slotOccupied verification.probeWire_laneProbes_6_slots_3_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_6_slots_3_pipeFinish verification.probeWire_laneProbes_6_slots_3_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_6_slots_3_slotShiftValid verification.probeWire_laneProbes_6_slots_3_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_6_slots_3_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_6_slots_3_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_6_slots_3_decodeResultIsScheduler verification.probeWire_laneProbes_6_slots_3_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_6_slots_3_executionUnitVfuRequestReady verification.probeWire_laneProbes_6_slots_3_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_6_slots_3_executionUnitVfuRequestValid verification.probeWire_laneProbes_6_slots_3_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_6_slots_3_stage3VrfWriteReady verification.probeWire_laneProbes_6_slots_3_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_6_slots_3_stage3VrfWriteValid verification.probeWire_laneProbes_6_slots_3_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_6_slots_3_writeQueueEnq verification.probeWire_laneProbes_6_slots_3_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_6_slots_3_writeTag verification.probeWire_laneProbes_6_slots_3_writeTag_probe
`define ref_T1_t1Probe_laneProbes_6_slots_3_writeMask verification.probeWire_laneProbes_6_slots_3_writeMask_probe
`define ref_T1_t1Probe_laneProbes_6_laneRequestStall verification.probeWire_laneProbes_6_laneRequestStall_probe
`define ref_T1_t1Probe_laneProbes_6_lastSlotOccupied verification.probeWire_laneProbes_6_lastSlotOccupied_probe
`define ref_T1_t1Probe_laneProbes_6_instructionFinished verification.probeWire_laneProbes_6_instructionFinished_probe
`define ref_T1_t1Probe_laneProbes_6_instructionValid verification.probeWire_laneProbes_6_instructionValid_probe
`define ref_T1_t1Probe_laneProbes_6_crossWriteProbe_0_valid verification.probeWire_laneProbes_6_crossWriteProbe_0_valid_probe
`define ref_T1_t1Probe_laneProbes_6_crossWriteProbe_0_bits_writeTag verification.probeWire_laneProbes_6_crossWriteProbe_0_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_6_crossWriteProbe_0_bits_writeMask verification.probeWire_laneProbes_6_crossWriteProbe_0_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_6_crossWriteProbe_1_valid verification.probeWire_laneProbes_6_crossWriteProbe_1_valid_probe
`define ref_T1_t1Probe_laneProbes_6_crossWriteProbe_1_bits_writeTag verification.probeWire_laneProbes_6_crossWriteProbe_1_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_6_crossWriteProbe_1_bits_writeMask verification.probeWire_laneProbes_6_crossWriteProbe_1_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_6_vrfProbe_valid verification.probeWire_laneProbes_6_vrfProbe_valid_probe
`define ref_T1_t1Probe_laneProbes_6_vrfProbe_requestVd verification.probeWire_laneProbes_6_vrfProbe_requestVd_probe
`define ref_T1_t1Probe_laneProbes_6_vrfProbe_requestOffset verification.probeWire_laneProbes_6_vrfProbe_requestOffset_probe
`define ref_T1_t1Probe_laneProbes_6_vrfProbe_requestMask verification.probeWire_laneProbes_6_vrfProbe_requestMask_probe
`define ref_T1_t1Probe_laneProbes_6_vrfProbe_requestData verification.probeWire_laneProbes_6_vrfProbe_requestData_probe
`define ref_T1_t1Probe_laneProbes_6_vrfProbe_requestInstruction verification.probeWire_laneProbes_6_vrfProbe_requestInstruction_probe
`define ref_T1_t1Probe_laneProbes_7_slots_0_stage0EnqueueReady verification.probeWire_laneProbes_7_slots_0_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_7_slots_0_stage0EnqueueValid verification.probeWire_laneProbes_7_slots_0_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_7_slots_0_changingMaskSet verification.probeWire_laneProbes_7_slots_0_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_7_slots_0_slotActive verification.probeWire_laneProbes_7_slots_0_slotActive_probe
`define ref_T1_t1Probe_laneProbes_7_slots_0_slotOccupied verification.probeWire_laneProbes_7_slots_0_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_7_slots_0_pipeFinish verification.probeWire_laneProbes_7_slots_0_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_7_slots_0_slotShiftValid verification.probeWire_laneProbes_7_slots_0_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_7_slots_0_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_7_slots_0_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_7_slots_0_decodeResultIsScheduler verification.probeWire_laneProbes_7_slots_0_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_7_slots_0_executionUnitVfuRequestReady verification.probeWire_laneProbes_7_slots_0_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_7_slots_0_executionUnitVfuRequestValid verification.probeWire_laneProbes_7_slots_0_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_7_slots_0_stage3VrfWriteReady verification.probeWire_laneProbes_7_slots_0_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_7_slots_0_stage3VrfWriteValid verification.probeWire_laneProbes_7_slots_0_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_7_slots_0_writeQueueEnq verification.probeWire_laneProbes_7_slots_0_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_7_slots_0_writeTag verification.probeWire_laneProbes_7_slots_0_writeTag_probe
`define ref_T1_t1Probe_laneProbes_7_slots_0_writeMask verification.probeWire_laneProbes_7_slots_0_writeMask_probe
`define ref_T1_t1Probe_laneProbes_7_slots_1_stage0EnqueueReady verification.probeWire_laneProbes_7_slots_1_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_7_slots_1_stage0EnqueueValid verification.probeWire_laneProbes_7_slots_1_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_7_slots_1_changingMaskSet verification.probeWire_laneProbes_7_slots_1_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_7_slots_1_slotActive verification.probeWire_laneProbes_7_slots_1_slotActive_probe
`define ref_T1_t1Probe_laneProbes_7_slots_1_slotOccupied verification.probeWire_laneProbes_7_slots_1_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_7_slots_1_pipeFinish verification.probeWire_laneProbes_7_slots_1_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_7_slots_1_slotShiftValid verification.probeWire_laneProbes_7_slots_1_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_7_slots_1_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_7_slots_1_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_7_slots_1_decodeResultIsScheduler verification.probeWire_laneProbes_7_slots_1_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_7_slots_1_executionUnitVfuRequestReady verification.probeWire_laneProbes_7_slots_1_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_7_slots_1_executionUnitVfuRequestValid verification.probeWire_laneProbes_7_slots_1_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_7_slots_1_stage3VrfWriteReady verification.probeWire_laneProbes_7_slots_1_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_7_slots_1_stage3VrfWriteValid verification.probeWire_laneProbes_7_slots_1_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_7_slots_1_writeQueueEnq verification.probeWire_laneProbes_7_slots_1_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_7_slots_1_writeTag verification.probeWire_laneProbes_7_slots_1_writeTag_probe
`define ref_T1_t1Probe_laneProbes_7_slots_1_writeMask verification.probeWire_laneProbes_7_slots_1_writeMask_probe
`define ref_T1_t1Probe_laneProbes_7_slots_2_stage0EnqueueReady verification.probeWire_laneProbes_7_slots_2_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_7_slots_2_stage0EnqueueValid verification.probeWire_laneProbes_7_slots_2_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_7_slots_2_changingMaskSet verification.probeWire_laneProbes_7_slots_2_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_7_slots_2_slotActive verification.probeWire_laneProbes_7_slots_2_slotActive_probe
`define ref_T1_t1Probe_laneProbes_7_slots_2_slotOccupied verification.probeWire_laneProbes_7_slots_2_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_7_slots_2_pipeFinish verification.probeWire_laneProbes_7_slots_2_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_7_slots_2_slotShiftValid verification.probeWire_laneProbes_7_slots_2_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_7_slots_2_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_7_slots_2_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_7_slots_2_decodeResultIsScheduler verification.probeWire_laneProbes_7_slots_2_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_7_slots_2_executionUnitVfuRequestReady verification.probeWire_laneProbes_7_slots_2_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_7_slots_2_executionUnitVfuRequestValid verification.probeWire_laneProbes_7_slots_2_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_7_slots_2_stage3VrfWriteReady verification.probeWire_laneProbes_7_slots_2_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_7_slots_2_stage3VrfWriteValid verification.probeWire_laneProbes_7_slots_2_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_7_slots_2_writeQueueEnq verification.probeWire_laneProbes_7_slots_2_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_7_slots_2_writeTag verification.probeWire_laneProbes_7_slots_2_writeTag_probe
`define ref_T1_t1Probe_laneProbes_7_slots_2_writeMask verification.probeWire_laneProbes_7_slots_2_writeMask_probe
`define ref_T1_t1Probe_laneProbes_7_slots_3_stage0EnqueueReady verification.probeWire_laneProbes_7_slots_3_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_7_slots_3_stage0EnqueueValid verification.probeWire_laneProbes_7_slots_3_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_7_slots_3_changingMaskSet verification.probeWire_laneProbes_7_slots_3_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_7_slots_3_slotActive verification.probeWire_laneProbes_7_slots_3_slotActive_probe
`define ref_T1_t1Probe_laneProbes_7_slots_3_slotOccupied verification.probeWire_laneProbes_7_slots_3_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_7_slots_3_pipeFinish verification.probeWire_laneProbes_7_slots_3_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_7_slots_3_slotShiftValid verification.probeWire_laneProbes_7_slots_3_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_7_slots_3_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_7_slots_3_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_7_slots_3_decodeResultIsScheduler verification.probeWire_laneProbes_7_slots_3_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_7_slots_3_executionUnitVfuRequestReady verification.probeWire_laneProbes_7_slots_3_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_7_slots_3_executionUnitVfuRequestValid verification.probeWire_laneProbes_7_slots_3_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_7_slots_3_stage3VrfWriteReady verification.probeWire_laneProbes_7_slots_3_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_7_slots_3_stage3VrfWriteValid verification.probeWire_laneProbes_7_slots_3_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_7_slots_3_writeQueueEnq verification.probeWire_laneProbes_7_slots_3_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_7_slots_3_writeTag verification.probeWire_laneProbes_7_slots_3_writeTag_probe
`define ref_T1_t1Probe_laneProbes_7_slots_3_writeMask verification.probeWire_laneProbes_7_slots_3_writeMask_probe
`define ref_T1_t1Probe_laneProbes_7_laneRequestStall verification.probeWire_laneProbes_7_laneRequestStall_probe
`define ref_T1_t1Probe_laneProbes_7_lastSlotOccupied verification.probeWire_laneProbes_7_lastSlotOccupied_probe
`define ref_T1_t1Probe_laneProbes_7_instructionFinished verification.probeWire_laneProbes_7_instructionFinished_probe
`define ref_T1_t1Probe_laneProbes_7_instructionValid verification.probeWire_laneProbes_7_instructionValid_probe
`define ref_T1_t1Probe_laneProbes_7_crossWriteProbe_0_valid verification.probeWire_laneProbes_7_crossWriteProbe_0_valid_probe
`define ref_T1_t1Probe_laneProbes_7_crossWriteProbe_0_bits_writeTag verification.probeWire_laneProbes_7_crossWriteProbe_0_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_7_crossWriteProbe_0_bits_writeMask verification.probeWire_laneProbes_7_crossWriteProbe_0_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_7_crossWriteProbe_1_valid verification.probeWire_laneProbes_7_crossWriteProbe_1_valid_probe
`define ref_T1_t1Probe_laneProbes_7_crossWriteProbe_1_bits_writeTag verification.probeWire_laneProbes_7_crossWriteProbe_1_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_7_crossWriteProbe_1_bits_writeMask verification.probeWire_laneProbes_7_crossWriteProbe_1_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_7_vrfProbe_valid verification.probeWire_laneProbes_7_vrfProbe_valid_probe
`define ref_T1_t1Probe_laneProbes_7_vrfProbe_requestVd verification.probeWire_laneProbes_7_vrfProbe_requestVd_probe
`define ref_T1_t1Probe_laneProbes_7_vrfProbe_requestOffset verification.probeWire_laneProbes_7_vrfProbe_requestOffset_probe
`define ref_T1_t1Probe_laneProbes_7_vrfProbe_requestMask verification.probeWire_laneProbes_7_vrfProbe_requestMask_probe
`define ref_T1_t1Probe_laneProbes_7_vrfProbe_requestData verification.probeWire_laneProbes_7_vrfProbe_requestData_probe
`define ref_T1_t1Probe_laneProbes_7_vrfProbe_requestInstruction verification.probeWire_laneProbes_7_vrfProbe_requestInstruction_probe
`define ref_T1_t1Probe_laneProbes_8_slots_0_stage0EnqueueReady verification.probeWire_laneProbes_8_slots_0_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_8_slots_0_stage0EnqueueValid verification.probeWire_laneProbes_8_slots_0_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_8_slots_0_changingMaskSet verification.probeWire_laneProbes_8_slots_0_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_8_slots_0_slotActive verification.probeWire_laneProbes_8_slots_0_slotActive_probe
`define ref_T1_t1Probe_laneProbes_8_slots_0_slotOccupied verification.probeWire_laneProbes_8_slots_0_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_8_slots_0_pipeFinish verification.probeWire_laneProbes_8_slots_0_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_8_slots_0_slotShiftValid verification.probeWire_laneProbes_8_slots_0_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_8_slots_0_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_8_slots_0_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_8_slots_0_decodeResultIsScheduler verification.probeWire_laneProbes_8_slots_0_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_8_slots_0_executionUnitVfuRequestReady verification.probeWire_laneProbes_8_slots_0_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_8_slots_0_executionUnitVfuRequestValid verification.probeWire_laneProbes_8_slots_0_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_8_slots_0_stage3VrfWriteReady verification.probeWire_laneProbes_8_slots_0_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_8_slots_0_stage3VrfWriteValid verification.probeWire_laneProbes_8_slots_0_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_8_slots_0_writeQueueEnq verification.probeWire_laneProbes_8_slots_0_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_8_slots_0_writeTag verification.probeWire_laneProbes_8_slots_0_writeTag_probe
`define ref_T1_t1Probe_laneProbes_8_slots_0_writeMask verification.probeWire_laneProbes_8_slots_0_writeMask_probe
`define ref_T1_t1Probe_laneProbes_8_slots_1_stage0EnqueueReady verification.probeWire_laneProbes_8_slots_1_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_8_slots_1_stage0EnqueueValid verification.probeWire_laneProbes_8_slots_1_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_8_slots_1_changingMaskSet verification.probeWire_laneProbes_8_slots_1_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_8_slots_1_slotActive verification.probeWire_laneProbes_8_slots_1_slotActive_probe
`define ref_T1_t1Probe_laneProbes_8_slots_1_slotOccupied verification.probeWire_laneProbes_8_slots_1_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_8_slots_1_pipeFinish verification.probeWire_laneProbes_8_slots_1_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_8_slots_1_slotShiftValid verification.probeWire_laneProbes_8_slots_1_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_8_slots_1_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_8_slots_1_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_8_slots_1_decodeResultIsScheduler verification.probeWire_laneProbes_8_slots_1_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_8_slots_1_executionUnitVfuRequestReady verification.probeWire_laneProbes_8_slots_1_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_8_slots_1_executionUnitVfuRequestValid verification.probeWire_laneProbes_8_slots_1_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_8_slots_1_stage3VrfWriteReady verification.probeWire_laneProbes_8_slots_1_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_8_slots_1_stage3VrfWriteValid verification.probeWire_laneProbes_8_slots_1_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_8_slots_1_writeQueueEnq verification.probeWire_laneProbes_8_slots_1_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_8_slots_1_writeTag verification.probeWire_laneProbes_8_slots_1_writeTag_probe
`define ref_T1_t1Probe_laneProbes_8_slots_1_writeMask verification.probeWire_laneProbes_8_slots_1_writeMask_probe
`define ref_T1_t1Probe_laneProbes_8_slots_2_stage0EnqueueReady verification.probeWire_laneProbes_8_slots_2_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_8_slots_2_stage0EnqueueValid verification.probeWire_laneProbes_8_slots_2_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_8_slots_2_changingMaskSet verification.probeWire_laneProbes_8_slots_2_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_8_slots_2_slotActive verification.probeWire_laneProbes_8_slots_2_slotActive_probe
`define ref_T1_t1Probe_laneProbes_8_slots_2_slotOccupied verification.probeWire_laneProbes_8_slots_2_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_8_slots_2_pipeFinish verification.probeWire_laneProbes_8_slots_2_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_8_slots_2_slotShiftValid verification.probeWire_laneProbes_8_slots_2_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_8_slots_2_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_8_slots_2_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_8_slots_2_decodeResultIsScheduler verification.probeWire_laneProbes_8_slots_2_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_8_slots_2_executionUnitVfuRequestReady verification.probeWire_laneProbes_8_slots_2_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_8_slots_2_executionUnitVfuRequestValid verification.probeWire_laneProbes_8_slots_2_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_8_slots_2_stage3VrfWriteReady verification.probeWire_laneProbes_8_slots_2_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_8_slots_2_stage3VrfWriteValid verification.probeWire_laneProbes_8_slots_2_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_8_slots_2_writeQueueEnq verification.probeWire_laneProbes_8_slots_2_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_8_slots_2_writeTag verification.probeWire_laneProbes_8_slots_2_writeTag_probe
`define ref_T1_t1Probe_laneProbes_8_slots_2_writeMask verification.probeWire_laneProbes_8_slots_2_writeMask_probe
`define ref_T1_t1Probe_laneProbes_8_slots_3_stage0EnqueueReady verification.probeWire_laneProbes_8_slots_3_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_8_slots_3_stage0EnqueueValid verification.probeWire_laneProbes_8_slots_3_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_8_slots_3_changingMaskSet verification.probeWire_laneProbes_8_slots_3_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_8_slots_3_slotActive verification.probeWire_laneProbes_8_slots_3_slotActive_probe
`define ref_T1_t1Probe_laneProbes_8_slots_3_slotOccupied verification.probeWire_laneProbes_8_slots_3_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_8_slots_3_pipeFinish verification.probeWire_laneProbes_8_slots_3_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_8_slots_3_slotShiftValid verification.probeWire_laneProbes_8_slots_3_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_8_slots_3_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_8_slots_3_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_8_slots_3_decodeResultIsScheduler verification.probeWire_laneProbes_8_slots_3_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_8_slots_3_executionUnitVfuRequestReady verification.probeWire_laneProbes_8_slots_3_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_8_slots_3_executionUnitVfuRequestValid verification.probeWire_laneProbes_8_slots_3_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_8_slots_3_stage3VrfWriteReady verification.probeWire_laneProbes_8_slots_3_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_8_slots_3_stage3VrfWriteValid verification.probeWire_laneProbes_8_slots_3_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_8_slots_3_writeQueueEnq verification.probeWire_laneProbes_8_slots_3_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_8_slots_3_writeTag verification.probeWire_laneProbes_8_slots_3_writeTag_probe
`define ref_T1_t1Probe_laneProbes_8_slots_3_writeMask verification.probeWire_laneProbes_8_slots_3_writeMask_probe
`define ref_T1_t1Probe_laneProbes_8_laneRequestStall verification.probeWire_laneProbes_8_laneRequestStall_probe
`define ref_T1_t1Probe_laneProbes_8_lastSlotOccupied verification.probeWire_laneProbes_8_lastSlotOccupied_probe
`define ref_T1_t1Probe_laneProbes_8_instructionFinished verification.probeWire_laneProbes_8_instructionFinished_probe
`define ref_T1_t1Probe_laneProbes_8_instructionValid verification.probeWire_laneProbes_8_instructionValid_probe
`define ref_T1_t1Probe_laneProbes_8_crossWriteProbe_0_valid verification.probeWire_laneProbes_8_crossWriteProbe_0_valid_probe
`define ref_T1_t1Probe_laneProbes_8_crossWriteProbe_0_bits_writeTag verification.probeWire_laneProbes_8_crossWriteProbe_0_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_8_crossWriteProbe_0_bits_writeMask verification.probeWire_laneProbes_8_crossWriteProbe_0_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_8_crossWriteProbe_1_valid verification.probeWire_laneProbes_8_crossWriteProbe_1_valid_probe
`define ref_T1_t1Probe_laneProbes_8_crossWriteProbe_1_bits_writeTag verification.probeWire_laneProbes_8_crossWriteProbe_1_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_8_crossWriteProbe_1_bits_writeMask verification.probeWire_laneProbes_8_crossWriteProbe_1_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_8_vrfProbe_valid verification.probeWire_laneProbes_8_vrfProbe_valid_probe
`define ref_T1_t1Probe_laneProbes_8_vrfProbe_requestVd verification.probeWire_laneProbes_8_vrfProbe_requestVd_probe
`define ref_T1_t1Probe_laneProbes_8_vrfProbe_requestOffset verification.probeWire_laneProbes_8_vrfProbe_requestOffset_probe
`define ref_T1_t1Probe_laneProbes_8_vrfProbe_requestMask verification.probeWire_laneProbes_8_vrfProbe_requestMask_probe
`define ref_T1_t1Probe_laneProbes_8_vrfProbe_requestData verification.probeWire_laneProbes_8_vrfProbe_requestData_probe
`define ref_T1_t1Probe_laneProbes_8_vrfProbe_requestInstruction verification.probeWire_laneProbes_8_vrfProbe_requestInstruction_probe
`define ref_T1_t1Probe_laneProbes_9_slots_0_stage0EnqueueReady verification.probeWire_laneProbes_9_slots_0_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_9_slots_0_stage0EnqueueValid verification.probeWire_laneProbes_9_slots_0_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_9_slots_0_changingMaskSet verification.probeWire_laneProbes_9_slots_0_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_9_slots_0_slotActive verification.probeWire_laneProbes_9_slots_0_slotActive_probe
`define ref_T1_t1Probe_laneProbes_9_slots_0_slotOccupied verification.probeWire_laneProbes_9_slots_0_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_9_slots_0_pipeFinish verification.probeWire_laneProbes_9_slots_0_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_9_slots_0_slotShiftValid verification.probeWire_laneProbes_9_slots_0_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_9_slots_0_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_9_slots_0_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_9_slots_0_decodeResultIsScheduler verification.probeWire_laneProbes_9_slots_0_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_9_slots_0_executionUnitVfuRequestReady verification.probeWire_laneProbes_9_slots_0_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_9_slots_0_executionUnitVfuRequestValid verification.probeWire_laneProbes_9_slots_0_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_9_slots_0_stage3VrfWriteReady verification.probeWire_laneProbes_9_slots_0_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_9_slots_0_stage3VrfWriteValid verification.probeWire_laneProbes_9_slots_0_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_9_slots_0_writeQueueEnq verification.probeWire_laneProbes_9_slots_0_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_9_slots_0_writeTag verification.probeWire_laneProbes_9_slots_0_writeTag_probe
`define ref_T1_t1Probe_laneProbes_9_slots_0_writeMask verification.probeWire_laneProbes_9_slots_0_writeMask_probe
`define ref_T1_t1Probe_laneProbes_9_slots_1_stage0EnqueueReady verification.probeWire_laneProbes_9_slots_1_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_9_slots_1_stage0EnqueueValid verification.probeWire_laneProbes_9_slots_1_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_9_slots_1_changingMaskSet verification.probeWire_laneProbes_9_slots_1_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_9_slots_1_slotActive verification.probeWire_laneProbes_9_slots_1_slotActive_probe
`define ref_T1_t1Probe_laneProbes_9_slots_1_slotOccupied verification.probeWire_laneProbes_9_slots_1_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_9_slots_1_pipeFinish verification.probeWire_laneProbes_9_slots_1_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_9_slots_1_slotShiftValid verification.probeWire_laneProbes_9_slots_1_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_9_slots_1_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_9_slots_1_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_9_slots_1_decodeResultIsScheduler verification.probeWire_laneProbes_9_slots_1_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_9_slots_1_executionUnitVfuRequestReady verification.probeWire_laneProbes_9_slots_1_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_9_slots_1_executionUnitVfuRequestValid verification.probeWire_laneProbes_9_slots_1_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_9_slots_1_stage3VrfWriteReady verification.probeWire_laneProbes_9_slots_1_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_9_slots_1_stage3VrfWriteValid verification.probeWire_laneProbes_9_slots_1_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_9_slots_1_writeQueueEnq verification.probeWire_laneProbes_9_slots_1_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_9_slots_1_writeTag verification.probeWire_laneProbes_9_slots_1_writeTag_probe
`define ref_T1_t1Probe_laneProbes_9_slots_1_writeMask verification.probeWire_laneProbes_9_slots_1_writeMask_probe
`define ref_T1_t1Probe_laneProbes_9_slots_2_stage0EnqueueReady verification.probeWire_laneProbes_9_slots_2_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_9_slots_2_stage0EnqueueValid verification.probeWire_laneProbes_9_slots_2_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_9_slots_2_changingMaskSet verification.probeWire_laneProbes_9_slots_2_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_9_slots_2_slotActive verification.probeWire_laneProbes_9_slots_2_slotActive_probe
`define ref_T1_t1Probe_laneProbes_9_slots_2_slotOccupied verification.probeWire_laneProbes_9_slots_2_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_9_slots_2_pipeFinish verification.probeWire_laneProbes_9_slots_2_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_9_slots_2_slotShiftValid verification.probeWire_laneProbes_9_slots_2_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_9_slots_2_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_9_slots_2_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_9_slots_2_decodeResultIsScheduler verification.probeWire_laneProbes_9_slots_2_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_9_slots_2_executionUnitVfuRequestReady verification.probeWire_laneProbes_9_slots_2_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_9_slots_2_executionUnitVfuRequestValid verification.probeWire_laneProbes_9_slots_2_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_9_slots_2_stage3VrfWriteReady verification.probeWire_laneProbes_9_slots_2_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_9_slots_2_stage3VrfWriteValid verification.probeWire_laneProbes_9_slots_2_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_9_slots_2_writeQueueEnq verification.probeWire_laneProbes_9_slots_2_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_9_slots_2_writeTag verification.probeWire_laneProbes_9_slots_2_writeTag_probe
`define ref_T1_t1Probe_laneProbes_9_slots_2_writeMask verification.probeWire_laneProbes_9_slots_2_writeMask_probe
`define ref_T1_t1Probe_laneProbes_9_slots_3_stage0EnqueueReady verification.probeWire_laneProbes_9_slots_3_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_9_slots_3_stage0EnqueueValid verification.probeWire_laneProbes_9_slots_3_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_9_slots_3_changingMaskSet verification.probeWire_laneProbes_9_slots_3_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_9_slots_3_slotActive verification.probeWire_laneProbes_9_slots_3_slotActive_probe
`define ref_T1_t1Probe_laneProbes_9_slots_3_slotOccupied verification.probeWire_laneProbes_9_slots_3_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_9_slots_3_pipeFinish verification.probeWire_laneProbes_9_slots_3_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_9_slots_3_slotShiftValid verification.probeWire_laneProbes_9_slots_3_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_9_slots_3_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_9_slots_3_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_9_slots_3_decodeResultIsScheduler verification.probeWire_laneProbes_9_slots_3_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_9_slots_3_executionUnitVfuRequestReady verification.probeWire_laneProbes_9_slots_3_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_9_slots_3_executionUnitVfuRequestValid verification.probeWire_laneProbes_9_slots_3_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_9_slots_3_stage3VrfWriteReady verification.probeWire_laneProbes_9_slots_3_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_9_slots_3_stage3VrfWriteValid verification.probeWire_laneProbes_9_slots_3_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_9_slots_3_writeQueueEnq verification.probeWire_laneProbes_9_slots_3_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_9_slots_3_writeTag verification.probeWire_laneProbes_9_slots_3_writeTag_probe
`define ref_T1_t1Probe_laneProbes_9_slots_3_writeMask verification.probeWire_laneProbes_9_slots_3_writeMask_probe
`define ref_T1_t1Probe_laneProbes_9_laneRequestStall verification.probeWire_laneProbes_9_laneRequestStall_probe
`define ref_T1_t1Probe_laneProbes_9_lastSlotOccupied verification.probeWire_laneProbes_9_lastSlotOccupied_probe
`define ref_T1_t1Probe_laneProbes_9_instructionFinished verification.probeWire_laneProbes_9_instructionFinished_probe
`define ref_T1_t1Probe_laneProbes_9_instructionValid verification.probeWire_laneProbes_9_instructionValid_probe
`define ref_T1_t1Probe_laneProbes_9_crossWriteProbe_0_valid verification.probeWire_laneProbes_9_crossWriteProbe_0_valid_probe
`define ref_T1_t1Probe_laneProbes_9_crossWriteProbe_0_bits_writeTag verification.probeWire_laneProbes_9_crossWriteProbe_0_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_9_crossWriteProbe_0_bits_writeMask verification.probeWire_laneProbes_9_crossWriteProbe_0_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_9_crossWriteProbe_1_valid verification.probeWire_laneProbes_9_crossWriteProbe_1_valid_probe
`define ref_T1_t1Probe_laneProbes_9_crossWriteProbe_1_bits_writeTag verification.probeWire_laneProbes_9_crossWriteProbe_1_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_9_crossWriteProbe_1_bits_writeMask verification.probeWire_laneProbes_9_crossWriteProbe_1_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_9_vrfProbe_valid verification.probeWire_laneProbes_9_vrfProbe_valid_probe
`define ref_T1_t1Probe_laneProbes_9_vrfProbe_requestVd verification.probeWire_laneProbes_9_vrfProbe_requestVd_probe
`define ref_T1_t1Probe_laneProbes_9_vrfProbe_requestOffset verification.probeWire_laneProbes_9_vrfProbe_requestOffset_probe
`define ref_T1_t1Probe_laneProbes_9_vrfProbe_requestMask verification.probeWire_laneProbes_9_vrfProbe_requestMask_probe
`define ref_T1_t1Probe_laneProbes_9_vrfProbe_requestData verification.probeWire_laneProbes_9_vrfProbe_requestData_probe
`define ref_T1_t1Probe_laneProbes_9_vrfProbe_requestInstruction verification.probeWire_laneProbes_9_vrfProbe_requestInstruction_probe
`define ref_T1_t1Probe_laneProbes_10_slots_0_stage0EnqueueReady verification.probeWire_laneProbes_10_slots_0_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_10_slots_0_stage0EnqueueValid verification.probeWire_laneProbes_10_slots_0_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_10_slots_0_changingMaskSet verification.probeWire_laneProbes_10_slots_0_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_10_slots_0_slotActive verification.probeWire_laneProbes_10_slots_0_slotActive_probe
`define ref_T1_t1Probe_laneProbes_10_slots_0_slotOccupied verification.probeWire_laneProbes_10_slots_0_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_10_slots_0_pipeFinish verification.probeWire_laneProbes_10_slots_0_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_10_slots_0_slotShiftValid verification.probeWire_laneProbes_10_slots_0_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_10_slots_0_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_10_slots_0_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_10_slots_0_decodeResultIsScheduler verification.probeWire_laneProbes_10_slots_0_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_10_slots_0_executionUnitVfuRequestReady verification.probeWire_laneProbes_10_slots_0_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_10_slots_0_executionUnitVfuRequestValid verification.probeWire_laneProbes_10_slots_0_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_10_slots_0_stage3VrfWriteReady verification.probeWire_laneProbes_10_slots_0_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_10_slots_0_stage3VrfWriteValid verification.probeWire_laneProbes_10_slots_0_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_10_slots_0_writeQueueEnq verification.probeWire_laneProbes_10_slots_0_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_10_slots_0_writeTag verification.probeWire_laneProbes_10_slots_0_writeTag_probe
`define ref_T1_t1Probe_laneProbes_10_slots_0_writeMask verification.probeWire_laneProbes_10_slots_0_writeMask_probe
`define ref_T1_t1Probe_laneProbes_10_slots_1_stage0EnqueueReady verification.probeWire_laneProbes_10_slots_1_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_10_slots_1_stage0EnqueueValid verification.probeWire_laneProbes_10_slots_1_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_10_slots_1_changingMaskSet verification.probeWire_laneProbes_10_slots_1_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_10_slots_1_slotActive verification.probeWire_laneProbes_10_slots_1_slotActive_probe
`define ref_T1_t1Probe_laneProbes_10_slots_1_slotOccupied verification.probeWire_laneProbes_10_slots_1_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_10_slots_1_pipeFinish verification.probeWire_laneProbes_10_slots_1_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_10_slots_1_slotShiftValid verification.probeWire_laneProbes_10_slots_1_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_10_slots_1_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_10_slots_1_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_10_slots_1_decodeResultIsScheduler verification.probeWire_laneProbes_10_slots_1_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_10_slots_1_executionUnitVfuRequestReady verification.probeWire_laneProbes_10_slots_1_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_10_slots_1_executionUnitVfuRequestValid verification.probeWire_laneProbes_10_slots_1_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_10_slots_1_stage3VrfWriteReady verification.probeWire_laneProbes_10_slots_1_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_10_slots_1_stage3VrfWriteValid verification.probeWire_laneProbes_10_slots_1_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_10_slots_1_writeQueueEnq verification.probeWire_laneProbes_10_slots_1_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_10_slots_1_writeTag verification.probeWire_laneProbes_10_slots_1_writeTag_probe
`define ref_T1_t1Probe_laneProbes_10_slots_1_writeMask verification.probeWire_laneProbes_10_slots_1_writeMask_probe
`define ref_T1_t1Probe_laneProbes_10_slots_2_stage0EnqueueReady verification.probeWire_laneProbes_10_slots_2_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_10_slots_2_stage0EnqueueValid verification.probeWire_laneProbes_10_slots_2_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_10_slots_2_changingMaskSet verification.probeWire_laneProbes_10_slots_2_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_10_slots_2_slotActive verification.probeWire_laneProbes_10_slots_2_slotActive_probe
`define ref_T1_t1Probe_laneProbes_10_slots_2_slotOccupied verification.probeWire_laneProbes_10_slots_2_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_10_slots_2_pipeFinish verification.probeWire_laneProbes_10_slots_2_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_10_slots_2_slotShiftValid verification.probeWire_laneProbes_10_slots_2_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_10_slots_2_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_10_slots_2_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_10_slots_2_decodeResultIsScheduler verification.probeWire_laneProbes_10_slots_2_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_10_slots_2_executionUnitVfuRequestReady verification.probeWire_laneProbes_10_slots_2_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_10_slots_2_executionUnitVfuRequestValid verification.probeWire_laneProbes_10_slots_2_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_10_slots_2_stage3VrfWriteReady verification.probeWire_laneProbes_10_slots_2_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_10_slots_2_stage3VrfWriteValid verification.probeWire_laneProbes_10_slots_2_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_10_slots_2_writeQueueEnq verification.probeWire_laneProbes_10_slots_2_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_10_slots_2_writeTag verification.probeWire_laneProbes_10_slots_2_writeTag_probe
`define ref_T1_t1Probe_laneProbes_10_slots_2_writeMask verification.probeWire_laneProbes_10_slots_2_writeMask_probe
`define ref_T1_t1Probe_laneProbes_10_slots_3_stage0EnqueueReady verification.probeWire_laneProbes_10_slots_3_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_10_slots_3_stage0EnqueueValid verification.probeWire_laneProbes_10_slots_3_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_10_slots_3_changingMaskSet verification.probeWire_laneProbes_10_slots_3_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_10_slots_3_slotActive verification.probeWire_laneProbes_10_slots_3_slotActive_probe
`define ref_T1_t1Probe_laneProbes_10_slots_3_slotOccupied verification.probeWire_laneProbes_10_slots_3_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_10_slots_3_pipeFinish verification.probeWire_laneProbes_10_slots_3_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_10_slots_3_slotShiftValid verification.probeWire_laneProbes_10_slots_3_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_10_slots_3_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_10_slots_3_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_10_slots_3_decodeResultIsScheduler verification.probeWire_laneProbes_10_slots_3_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_10_slots_3_executionUnitVfuRequestReady verification.probeWire_laneProbes_10_slots_3_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_10_slots_3_executionUnitVfuRequestValid verification.probeWire_laneProbes_10_slots_3_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_10_slots_3_stage3VrfWriteReady verification.probeWire_laneProbes_10_slots_3_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_10_slots_3_stage3VrfWriteValid verification.probeWire_laneProbes_10_slots_3_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_10_slots_3_writeQueueEnq verification.probeWire_laneProbes_10_slots_3_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_10_slots_3_writeTag verification.probeWire_laneProbes_10_slots_3_writeTag_probe
`define ref_T1_t1Probe_laneProbes_10_slots_3_writeMask verification.probeWire_laneProbes_10_slots_3_writeMask_probe
`define ref_T1_t1Probe_laneProbes_10_laneRequestStall verification.probeWire_laneProbes_10_laneRequestStall_probe
`define ref_T1_t1Probe_laneProbes_10_lastSlotOccupied verification.probeWire_laneProbes_10_lastSlotOccupied_probe
`define ref_T1_t1Probe_laneProbes_10_instructionFinished verification.probeWire_laneProbes_10_instructionFinished_probe
`define ref_T1_t1Probe_laneProbes_10_instructionValid verification.probeWire_laneProbes_10_instructionValid_probe
`define ref_T1_t1Probe_laneProbes_10_crossWriteProbe_0_valid verification.probeWire_laneProbes_10_crossWriteProbe_0_valid_probe
`define ref_T1_t1Probe_laneProbes_10_crossWriteProbe_0_bits_writeTag verification.probeWire_laneProbes_10_crossWriteProbe_0_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_10_crossWriteProbe_0_bits_writeMask verification.probeWire_laneProbes_10_crossWriteProbe_0_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_10_crossWriteProbe_1_valid verification.probeWire_laneProbes_10_crossWriteProbe_1_valid_probe
`define ref_T1_t1Probe_laneProbes_10_crossWriteProbe_1_bits_writeTag verification.probeWire_laneProbes_10_crossWriteProbe_1_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_10_crossWriteProbe_1_bits_writeMask verification.probeWire_laneProbes_10_crossWriteProbe_1_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_10_vrfProbe_valid verification.probeWire_laneProbes_10_vrfProbe_valid_probe
`define ref_T1_t1Probe_laneProbes_10_vrfProbe_requestVd verification.probeWire_laneProbes_10_vrfProbe_requestVd_probe
`define ref_T1_t1Probe_laneProbes_10_vrfProbe_requestOffset verification.probeWire_laneProbes_10_vrfProbe_requestOffset_probe
`define ref_T1_t1Probe_laneProbes_10_vrfProbe_requestMask verification.probeWire_laneProbes_10_vrfProbe_requestMask_probe
`define ref_T1_t1Probe_laneProbes_10_vrfProbe_requestData verification.probeWire_laneProbes_10_vrfProbe_requestData_probe
`define ref_T1_t1Probe_laneProbes_10_vrfProbe_requestInstruction verification.probeWire_laneProbes_10_vrfProbe_requestInstruction_probe
`define ref_T1_t1Probe_laneProbes_11_slots_0_stage0EnqueueReady verification.probeWire_laneProbes_11_slots_0_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_11_slots_0_stage0EnqueueValid verification.probeWire_laneProbes_11_slots_0_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_11_slots_0_changingMaskSet verification.probeWire_laneProbes_11_slots_0_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_11_slots_0_slotActive verification.probeWire_laneProbes_11_slots_0_slotActive_probe
`define ref_T1_t1Probe_laneProbes_11_slots_0_slotOccupied verification.probeWire_laneProbes_11_slots_0_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_11_slots_0_pipeFinish verification.probeWire_laneProbes_11_slots_0_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_11_slots_0_slotShiftValid verification.probeWire_laneProbes_11_slots_0_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_11_slots_0_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_11_slots_0_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_11_slots_0_decodeResultIsScheduler verification.probeWire_laneProbes_11_slots_0_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_11_slots_0_executionUnitVfuRequestReady verification.probeWire_laneProbes_11_slots_0_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_11_slots_0_executionUnitVfuRequestValid verification.probeWire_laneProbes_11_slots_0_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_11_slots_0_stage3VrfWriteReady verification.probeWire_laneProbes_11_slots_0_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_11_slots_0_stage3VrfWriteValid verification.probeWire_laneProbes_11_slots_0_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_11_slots_0_writeQueueEnq verification.probeWire_laneProbes_11_slots_0_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_11_slots_0_writeTag verification.probeWire_laneProbes_11_slots_0_writeTag_probe
`define ref_T1_t1Probe_laneProbes_11_slots_0_writeMask verification.probeWire_laneProbes_11_slots_0_writeMask_probe
`define ref_T1_t1Probe_laneProbes_11_slots_1_stage0EnqueueReady verification.probeWire_laneProbes_11_slots_1_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_11_slots_1_stage0EnqueueValid verification.probeWire_laneProbes_11_slots_1_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_11_slots_1_changingMaskSet verification.probeWire_laneProbes_11_slots_1_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_11_slots_1_slotActive verification.probeWire_laneProbes_11_slots_1_slotActive_probe
`define ref_T1_t1Probe_laneProbes_11_slots_1_slotOccupied verification.probeWire_laneProbes_11_slots_1_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_11_slots_1_pipeFinish verification.probeWire_laneProbes_11_slots_1_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_11_slots_1_slotShiftValid verification.probeWire_laneProbes_11_slots_1_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_11_slots_1_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_11_slots_1_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_11_slots_1_decodeResultIsScheduler verification.probeWire_laneProbes_11_slots_1_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_11_slots_1_executionUnitVfuRequestReady verification.probeWire_laneProbes_11_slots_1_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_11_slots_1_executionUnitVfuRequestValid verification.probeWire_laneProbes_11_slots_1_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_11_slots_1_stage3VrfWriteReady verification.probeWire_laneProbes_11_slots_1_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_11_slots_1_stage3VrfWriteValid verification.probeWire_laneProbes_11_slots_1_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_11_slots_1_writeQueueEnq verification.probeWire_laneProbes_11_slots_1_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_11_slots_1_writeTag verification.probeWire_laneProbes_11_slots_1_writeTag_probe
`define ref_T1_t1Probe_laneProbes_11_slots_1_writeMask verification.probeWire_laneProbes_11_slots_1_writeMask_probe
`define ref_T1_t1Probe_laneProbes_11_slots_2_stage0EnqueueReady verification.probeWire_laneProbes_11_slots_2_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_11_slots_2_stage0EnqueueValid verification.probeWire_laneProbes_11_slots_2_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_11_slots_2_changingMaskSet verification.probeWire_laneProbes_11_slots_2_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_11_slots_2_slotActive verification.probeWire_laneProbes_11_slots_2_slotActive_probe
`define ref_T1_t1Probe_laneProbes_11_slots_2_slotOccupied verification.probeWire_laneProbes_11_slots_2_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_11_slots_2_pipeFinish verification.probeWire_laneProbes_11_slots_2_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_11_slots_2_slotShiftValid verification.probeWire_laneProbes_11_slots_2_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_11_slots_2_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_11_slots_2_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_11_slots_2_decodeResultIsScheduler verification.probeWire_laneProbes_11_slots_2_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_11_slots_2_executionUnitVfuRequestReady verification.probeWire_laneProbes_11_slots_2_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_11_slots_2_executionUnitVfuRequestValid verification.probeWire_laneProbes_11_slots_2_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_11_slots_2_stage3VrfWriteReady verification.probeWire_laneProbes_11_slots_2_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_11_slots_2_stage3VrfWriteValid verification.probeWire_laneProbes_11_slots_2_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_11_slots_2_writeQueueEnq verification.probeWire_laneProbes_11_slots_2_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_11_slots_2_writeTag verification.probeWire_laneProbes_11_slots_2_writeTag_probe
`define ref_T1_t1Probe_laneProbes_11_slots_2_writeMask verification.probeWire_laneProbes_11_slots_2_writeMask_probe
`define ref_T1_t1Probe_laneProbes_11_slots_3_stage0EnqueueReady verification.probeWire_laneProbes_11_slots_3_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_11_slots_3_stage0EnqueueValid verification.probeWire_laneProbes_11_slots_3_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_11_slots_3_changingMaskSet verification.probeWire_laneProbes_11_slots_3_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_11_slots_3_slotActive verification.probeWire_laneProbes_11_slots_3_slotActive_probe
`define ref_T1_t1Probe_laneProbes_11_slots_3_slotOccupied verification.probeWire_laneProbes_11_slots_3_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_11_slots_3_pipeFinish verification.probeWire_laneProbes_11_slots_3_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_11_slots_3_slotShiftValid verification.probeWire_laneProbes_11_slots_3_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_11_slots_3_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_11_slots_3_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_11_slots_3_decodeResultIsScheduler verification.probeWire_laneProbes_11_slots_3_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_11_slots_3_executionUnitVfuRequestReady verification.probeWire_laneProbes_11_slots_3_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_11_slots_3_executionUnitVfuRequestValid verification.probeWire_laneProbes_11_slots_3_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_11_slots_3_stage3VrfWriteReady verification.probeWire_laneProbes_11_slots_3_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_11_slots_3_stage3VrfWriteValid verification.probeWire_laneProbes_11_slots_3_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_11_slots_3_writeQueueEnq verification.probeWire_laneProbes_11_slots_3_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_11_slots_3_writeTag verification.probeWire_laneProbes_11_slots_3_writeTag_probe
`define ref_T1_t1Probe_laneProbes_11_slots_3_writeMask verification.probeWire_laneProbes_11_slots_3_writeMask_probe
`define ref_T1_t1Probe_laneProbes_11_laneRequestStall verification.probeWire_laneProbes_11_laneRequestStall_probe
`define ref_T1_t1Probe_laneProbes_11_lastSlotOccupied verification.probeWire_laneProbes_11_lastSlotOccupied_probe
`define ref_T1_t1Probe_laneProbes_11_instructionFinished verification.probeWire_laneProbes_11_instructionFinished_probe
`define ref_T1_t1Probe_laneProbes_11_instructionValid verification.probeWire_laneProbes_11_instructionValid_probe
`define ref_T1_t1Probe_laneProbes_11_crossWriteProbe_0_valid verification.probeWire_laneProbes_11_crossWriteProbe_0_valid_probe
`define ref_T1_t1Probe_laneProbes_11_crossWriteProbe_0_bits_writeTag verification.probeWire_laneProbes_11_crossWriteProbe_0_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_11_crossWriteProbe_0_bits_writeMask verification.probeWire_laneProbes_11_crossWriteProbe_0_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_11_crossWriteProbe_1_valid verification.probeWire_laneProbes_11_crossWriteProbe_1_valid_probe
`define ref_T1_t1Probe_laneProbes_11_crossWriteProbe_1_bits_writeTag verification.probeWire_laneProbes_11_crossWriteProbe_1_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_11_crossWriteProbe_1_bits_writeMask verification.probeWire_laneProbes_11_crossWriteProbe_1_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_11_vrfProbe_valid verification.probeWire_laneProbes_11_vrfProbe_valid_probe
`define ref_T1_t1Probe_laneProbes_11_vrfProbe_requestVd verification.probeWire_laneProbes_11_vrfProbe_requestVd_probe
`define ref_T1_t1Probe_laneProbes_11_vrfProbe_requestOffset verification.probeWire_laneProbes_11_vrfProbe_requestOffset_probe
`define ref_T1_t1Probe_laneProbes_11_vrfProbe_requestMask verification.probeWire_laneProbes_11_vrfProbe_requestMask_probe
`define ref_T1_t1Probe_laneProbes_11_vrfProbe_requestData verification.probeWire_laneProbes_11_vrfProbe_requestData_probe
`define ref_T1_t1Probe_laneProbes_11_vrfProbe_requestInstruction verification.probeWire_laneProbes_11_vrfProbe_requestInstruction_probe
`define ref_T1_t1Probe_laneProbes_12_slots_0_stage0EnqueueReady verification.probeWire_laneProbes_12_slots_0_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_12_slots_0_stage0EnqueueValid verification.probeWire_laneProbes_12_slots_0_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_12_slots_0_changingMaskSet verification.probeWire_laneProbes_12_slots_0_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_12_slots_0_slotActive verification.probeWire_laneProbes_12_slots_0_slotActive_probe
`define ref_T1_t1Probe_laneProbes_12_slots_0_slotOccupied verification.probeWire_laneProbes_12_slots_0_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_12_slots_0_pipeFinish verification.probeWire_laneProbes_12_slots_0_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_12_slots_0_slotShiftValid verification.probeWire_laneProbes_12_slots_0_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_12_slots_0_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_12_slots_0_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_12_slots_0_decodeResultIsScheduler verification.probeWire_laneProbes_12_slots_0_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_12_slots_0_executionUnitVfuRequestReady verification.probeWire_laneProbes_12_slots_0_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_12_slots_0_executionUnitVfuRequestValid verification.probeWire_laneProbes_12_slots_0_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_12_slots_0_stage3VrfWriteReady verification.probeWire_laneProbes_12_slots_0_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_12_slots_0_stage3VrfWriteValid verification.probeWire_laneProbes_12_slots_0_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_12_slots_0_writeQueueEnq verification.probeWire_laneProbes_12_slots_0_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_12_slots_0_writeTag verification.probeWire_laneProbes_12_slots_0_writeTag_probe
`define ref_T1_t1Probe_laneProbes_12_slots_0_writeMask verification.probeWire_laneProbes_12_slots_0_writeMask_probe
`define ref_T1_t1Probe_laneProbes_12_slots_1_stage0EnqueueReady verification.probeWire_laneProbes_12_slots_1_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_12_slots_1_stage0EnqueueValid verification.probeWire_laneProbes_12_slots_1_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_12_slots_1_changingMaskSet verification.probeWire_laneProbes_12_slots_1_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_12_slots_1_slotActive verification.probeWire_laneProbes_12_slots_1_slotActive_probe
`define ref_T1_t1Probe_laneProbes_12_slots_1_slotOccupied verification.probeWire_laneProbes_12_slots_1_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_12_slots_1_pipeFinish verification.probeWire_laneProbes_12_slots_1_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_12_slots_1_slotShiftValid verification.probeWire_laneProbes_12_slots_1_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_12_slots_1_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_12_slots_1_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_12_slots_1_decodeResultIsScheduler verification.probeWire_laneProbes_12_slots_1_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_12_slots_1_executionUnitVfuRequestReady verification.probeWire_laneProbes_12_slots_1_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_12_slots_1_executionUnitVfuRequestValid verification.probeWire_laneProbes_12_slots_1_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_12_slots_1_stage3VrfWriteReady verification.probeWire_laneProbes_12_slots_1_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_12_slots_1_stage3VrfWriteValid verification.probeWire_laneProbes_12_slots_1_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_12_slots_1_writeQueueEnq verification.probeWire_laneProbes_12_slots_1_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_12_slots_1_writeTag verification.probeWire_laneProbes_12_slots_1_writeTag_probe
`define ref_T1_t1Probe_laneProbes_12_slots_1_writeMask verification.probeWire_laneProbes_12_slots_1_writeMask_probe
`define ref_T1_t1Probe_laneProbes_12_slots_2_stage0EnqueueReady verification.probeWire_laneProbes_12_slots_2_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_12_slots_2_stage0EnqueueValid verification.probeWire_laneProbes_12_slots_2_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_12_slots_2_changingMaskSet verification.probeWire_laneProbes_12_slots_2_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_12_slots_2_slotActive verification.probeWire_laneProbes_12_slots_2_slotActive_probe
`define ref_T1_t1Probe_laneProbes_12_slots_2_slotOccupied verification.probeWire_laneProbes_12_slots_2_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_12_slots_2_pipeFinish verification.probeWire_laneProbes_12_slots_2_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_12_slots_2_slotShiftValid verification.probeWire_laneProbes_12_slots_2_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_12_slots_2_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_12_slots_2_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_12_slots_2_decodeResultIsScheduler verification.probeWire_laneProbes_12_slots_2_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_12_slots_2_executionUnitVfuRequestReady verification.probeWire_laneProbes_12_slots_2_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_12_slots_2_executionUnitVfuRequestValid verification.probeWire_laneProbes_12_slots_2_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_12_slots_2_stage3VrfWriteReady verification.probeWire_laneProbes_12_slots_2_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_12_slots_2_stage3VrfWriteValid verification.probeWire_laneProbes_12_slots_2_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_12_slots_2_writeQueueEnq verification.probeWire_laneProbes_12_slots_2_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_12_slots_2_writeTag verification.probeWire_laneProbes_12_slots_2_writeTag_probe
`define ref_T1_t1Probe_laneProbes_12_slots_2_writeMask verification.probeWire_laneProbes_12_slots_2_writeMask_probe
`define ref_T1_t1Probe_laneProbes_12_slots_3_stage0EnqueueReady verification.probeWire_laneProbes_12_slots_3_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_12_slots_3_stage0EnqueueValid verification.probeWire_laneProbes_12_slots_3_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_12_slots_3_changingMaskSet verification.probeWire_laneProbes_12_slots_3_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_12_slots_3_slotActive verification.probeWire_laneProbes_12_slots_3_slotActive_probe
`define ref_T1_t1Probe_laneProbes_12_slots_3_slotOccupied verification.probeWire_laneProbes_12_slots_3_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_12_slots_3_pipeFinish verification.probeWire_laneProbes_12_slots_3_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_12_slots_3_slotShiftValid verification.probeWire_laneProbes_12_slots_3_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_12_slots_3_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_12_slots_3_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_12_slots_3_decodeResultIsScheduler verification.probeWire_laneProbes_12_slots_3_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_12_slots_3_executionUnitVfuRequestReady verification.probeWire_laneProbes_12_slots_3_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_12_slots_3_executionUnitVfuRequestValid verification.probeWire_laneProbes_12_slots_3_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_12_slots_3_stage3VrfWriteReady verification.probeWire_laneProbes_12_slots_3_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_12_slots_3_stage3VrfWriteValid verification.probeWire_laneProbes_12_slots_3_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_12_slots_3_writeQueueEnq verification.probeWire_laneProbes_12_slots_3_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_12_slots_3_writeTag verification.probeWire_laneProbes_12_slots_3_writeTag_probe
`define ref_T1_t1Probe_laneProbes_12_slots_3_writeMask verification.probeWire_laneProbes_12_slots_3_writeMask_probe
`define ref_T1_t1Probe_laneProbes_12_laneRequestStall verification.probeWire_laneProbes_12_laneRequestStall_probe
`define ref_T1_t1Probe_laneProbes_12_lastSlotOccupied verification.probeWire_laneProbes_12_lastSlotOccupied_probe
`define ref_T1_t1Probe_laneProbes_12_instructionFinished verification.probeWire_laneProbes_12_instructionFinished_probe
`define ref_T1_t1Probe_laneProbes_12_instructionValid verification.probeWire_laneProbes_12_instructionValid_probe
`define ref_T1_t1Probe_laneProbes_12_crossWriteProbe_0_valid verification.probeWire_laneProbes_12_crossWriteProbe_0_valid_probe
`define ref_T1_t1Probe_laneProbes_12_crossWriteProbe_0_bits_writeTag verification.probeWire_laneProbes_12_crossWriteProbe_0_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_12_crossWriteProbe_0_bits_writeMask verification.probeWire_laneProbes_12_crossWriteProbe_0_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_12_crossWriteProbe_1_valid verification.probeWire_laneProbes_12_crossWriteProbe_1_valid_probe
`define ref_T1_t1Probe_laneProbes_12_crossWriteProbe_1_bits_writeTag verification.probeWire_laneProbes_12_crossWriteProbe_1_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_12_crossWriteProbe_1_bits_writeMask verification.probeWire_laneProbes_12_crossWriteProbe_1_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_12_vrfProbe_valid verification.probeWire_laneProbes_12_vrfProbe_valid_probe
`define ref_T1_t1Probe_laneProbes_12_vrfProbe_requestVd verification.probeWire_laneProbes_12_vrfProbe_requestVd_probe
`define ref_T1_t1Probe_laneProbes_12_vrfProbe_requestOffset verification.probeWire_laneProbes_12_vrfProbe_requestOffset_probe
`define ref_T1_t1Probe_laneProbes_12_vrfProbe_requestMask verification.probeWire_laneProbes_12_vrfProbe_requestMask_probe
`define ref_T1_t1Probe_laneProbes_12_vrfProbe_requestData verification.probeWire_laneProbes_12_vrfProbe_requestData_probe
`define ref_T1_t1Probe_laneProbes_12_vrfProbe_requestInstruction verification.probeWire_laneProbes_12_vrfProbe_requestInstruction_probe
`define ref_T1_t1Probe_laneProbes_13_slots_0_stage0EnqueueReady verification.probeWire_laneProbes_13_slots_0_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_13_slots_0_stage0EnqueueValid verification.probeWire_laneProbes_13_slots_0_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_13_slots_0_changingMaskSet verification.probeWire_laneProbes_13_slots_0_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_13_slots_0_slotActive verification.probeWire_laneProbes_13_slots_0_slotActive_probe
`define ref_T1_t1Probe_laneProbes_13_slots_0_slotOccupied verification.probeWire_laneProbes_13_slots_0_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_13_slots_0_pipeFinish verification.probeWire_laneProbes_13_slots_0_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_13_slots_0_slotShiftValid verification.probeWire_laneProbes_13_slots_0_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_13_slots_0_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_13_slots_0_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_13_slots_0_decodeResultIsScheduler verification.probeWire_laneProbes_13_slots_0_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_13_slots_0_executionUnitVfuRequestReady verification.probeWire_laneProbes_13_slots_0_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_13_slots_0_executionUnitVfuRequestValid verification.probeWire_laneProbes_13_slots_0_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_13_slots_0_stage3VrfWriteReady verification.probeWire_laneProbes_13_slots_0_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_13_slots_0_stage3VrfWriteValid verification.probeWire_laneProbes_13_slots_0_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_13_slots_0_writeQueueEnq verification.probeWire_laneProbes_13_slots_0_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_13_slots_0_writeTag verification.probeWire_laneProbes_13_slots_0_writeTag_probe
`define ref_T1_t1Probe_laneProbes_13_slots_0_writeMask verification.probeWire_laneProbes_13_slots_0_writeMask_probe
`define ref_T1_t1Probe_laneProbes_13_slots_1_stage0EnqueueReady verification.probeWire_laneProbes_13_slots_1_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_13_slots_1_stage0EnqueueValid verification.probeWire_laneProbes_13_slots_1_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_13_slots_1_changingMaskSet verification.probeWire_laneProbes_13_slots_1_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_13_slots_1_slotActive verification.probeWire_laneProbes_13_slots_1_slotActive_probe
`define ref_T1_t1Probe_laneProbes_13_slots_1_slotOccupied verification.probeWire_laneProbes_13_slots_1_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_13_slots_1_pipeFinish verification.probeWire_laneProbes_13_slots_1_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_13_slots_1_slotShiftValid verification.probeWire_laneProbes_13_slots_1_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_13_slots_1_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_13_slots_1_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_13_slots_1_decodeResultIsScheduler verification.probeWire_laneProbes_13_slots_1_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_13_slots_1_executionUnitVfuRequestReady verification.probeWire_laneProbes_13_slots_1_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_13_slots_1_executionUnitVfuRequestValid verification.probeWire_laneProbes_13_slots_1_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_13_slots_1_stage3VrfWriteReady verification.probeWire_laneProbes_13_slots_1_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_13_slots_1_stage3VrfWriteValid verification.probeWire_laneProbes_13_slots_1_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_13_slots_1_writeQueueEnq verification.probeWire_laneProbes_13_slots_1_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_13_slots_1_writeTag verification.probeWire_laneProbes_13_slots_1_writeTag_probe
`define ref_T1_t1Probe_laneProbes_13_slots_1_writeMask verification.probeWire_laneProbes_13_slots_1_writeMask_probe
`define ref_T1_t1Probe_laneProbes_13_slots_2_stage0EnqueueReady verification.probeWire_laneProbes_13_slots_2_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_13_slots_2_stage0EnqueueValid verification.probeWire_laneProbes_13_slots_2_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_13_slots_2_changingMaskSet verification.probeWire_laneProbes_13_slots_2_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_13_slots_2_slotActive verification.probeWire_laneProbes_13_slots_2_slotActive_probe
`define ref_T1_t1Probe_laneProbes_13_slots_2_slotOccupied verification.probeWire_laneProbes_13_slots_2_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_13_slots_2_pipeFinish verification.probeWire_laneProbes_13_slots_2_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_13_slots_2_slotShiftValid verification.probeWire_laneProbes_13_slots_2_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_13_slots_2_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_13_slots_2_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_13_slots_2_decodeResultIsScheduler verification.probeWire_laneProbes_13_slots_2_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_13_slots_2_executionUnitVfuRequestReady verification.probeWire_laneProbes_13_slots_2_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_13_slots_2_executionUnitVfuRequestValid verification.probeWire_laneProbes_13_slots_2_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_13_slots_2_stage3VrfWriteReady verification.probeWire_laneProbes_13_slots_2_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_13_slots_2_stage3VrfWriteValid verification.probeWire_laneProbes_13_slots_2_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_13_slots_2_writeQueueEnq verification.probeWire_laneProbes_13_slots_2_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_13_slots_2_writeTag verification.probeWire_laneProbes_13_slots_2_writeTag_probe
`define ref_T1_t1Probe_laneProbes_13_slots_2_writeMask verification.probeWire_laneProbes_13_slots_2_writeMask_probe
`define ref_T1_t1Probe_laneProbes_13_slots_3_stage0EnqueueReady verification.probeWire_laneProbes_13_slots_3_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_13_slots_3_stage0EnqueueValid verification.probeWire_laneProbes_13_slots_3_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_13_slots_3_changingMaskSet verification.probeWire_laneProbes_13_slots_3_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_13_slots_3_slotActive verification.probeWire_laneProbes_13_slots_3_slotActive_probe
`define ref_T1_t1Probe_laneProbes_13_slots_3_slotOccupied verification.probeWire_laneProbes_13_slots_3_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_13_slots_3_pipeFinish verification.probeWire_laneProbes_13_slots_3_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_13_slots_3_slotShiftValid verification.probeWire_laneProbes_13_slots_3_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_13_slots_3_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_13_slots_3_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_13_slots_3_decodeResultIsScheduler verification.probeWire_laneProbes_13_slots_3_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_13_slots_3_executionUnitVfuRequestReady verification.probeWire_laneProbes_13_slots_3_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_13_slots_3_executionUnitVfuRequestValid verification.probeWire_laneProbes_13_slots_3_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_13_slots_3_stage3VrfWriteReady verification.probeWire_laneProbes_13_slots_3_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_13_slots_3_stage3VrfWriteValid verification.probeWire_laneProbes_13_slots_3_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_13_slots_3_writeQueueEnq verification.probeWire_laneProbes_13_slots_3_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_13_slots_3_writeTag verification.probeWire_laneProbes_13_slots_3_writeTag_probe
`define ref_T1_t1Probe_laneProbes_13_slots_3_writeMask verification.probeWire_laneProbes_13_slots_3_writeMask_probe
`define ref_T1_t1Probe_laneProbes_13_laneRequestStall verification.probeWire_laneProbes_13_laneRequestStall_probe
`define ref_T1_t1Probe_laneProbes_13_lastSlotOccupied verification.probeWire_laneProbes_13_lastSlotOccupied_probe
`define ref_T1_t1Probe_laneProbes_13_instructionFinished verification.probeWire_laneProbes_13_instructionFinished_probe
`define ref_T1_t1Probe_laneProbes_13_instructionValid verification.probeWire_laneProbes_13_instructionValid_probe
`define ref_T1_t1Probe_laneProbes_13_crossWriteProbe_0_valid verification.probeWire_laneProbes_13_crossWriteProbe_0_valid_probe
`define ref_T1_t1Probe_laneProbes_13_crossWriteProbe_0_bits_writeTag verification.probeWire_laneProbes_13_crossWriteProbe_0_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_13_crossWriteProbe_0_bits_writeMask verification.probeWire_laneProbes_13_crossWriteProbe_0_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_13_crossWriteProbe_1_valid verification.probeWire_laneProbes_13_crossWriteProbe_1_valid_probe
`define ref_T1_t1Probe_laneProbes_13_crossWriteProbe_1_bits_writeTag verification.probeWire_laneProbes_13_crossWriteProbe_1_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_13_crossWriteProbe_1_bits_writeMask verification.probeWire_laneProbes_13_crossWriteProbe_1_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_13_vrfProbe_valid verification.probeWire_laneProbes_13_vrfProbe_valid_probe
`define ref_T1_t1Probe_laneProbes_13_vrfProbe_requestVd verification.probeWire_laneProbes_13_vrfProbe_requestVd_probe
`define ref_T1_t1Probe_laneProbes_13_vrfProbe_requestOffset verification.probeWire_laneProbes_13_vrfProbe_requestOffset_probe
`define ref_T1_t1Probe_laneProbes_13_vrfProbe_requestMask verification.probeWire_laneProbes_13_vrfProbe_requestMask_probe
`define ref_T1_t1Probe_laneProbes_13_vrfProbe_requestData verification.probeWire_laneProbes_13_vrfProbe_requestData_probe
`define ref_T1_t1Probe_laneProbes_13_vrfProbe_requestInstruction verification.probeWire_laneProbes_13_vrfProbe_requestInstruction_probe
`define ref_T1_t1Probe_laneProbes_14_slots_0_stage0EnqueueReady verification.probeWire_laneProbes_14_slots_0_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_14_slots_0_stage0EnqueueValid verification.probeWire_laneProbes_14_slots_0_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_14_slots_0_changingMaskSet verification.probeWire_laneProbes_14_slots_0_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_14_slots_0_slotActive verification.probeWire_laneProbes_14_slots_0_slotActive_probe
`define ref_T1_t1Probe_laneProbes_14_slots_0_slotOccupied verification.probeWire_laneProbes_14_slots_0_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_14_slots_0_pipeFinish verification.probeWire_laneProbes_14_slots_0_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_14_slots_0_slotShiftValid verification.probeWire_laneProbes_14_slots_0_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_14_slots_0_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_14_slots_0_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_14_slots_0_decodeResultIsScheduler verification.probeWire_laneProbes_14_slots_0_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_14_slots_0_executionUnitVfuRequestReady verification.probeWire_laneProbes_14_slots_0_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_14_slots_0_executionUnitVfuRequestValid verification.probeWire_laneProbes_14_slots_0_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_14_slots_0_stage3VrfWriteReady verification.probeWire_laneProbes_14_slots_0_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_14_slots_0_stage3VrfWriteValid verification.probeWire_laneProbes_14_slots_0_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_14_slots_0_writeQueueEnq verification.probeWire_laneProbes_14_slots_0_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_14_slots_0_writeTag verification.probeWire_laneProbes_14_slots_0_writeTag_probe
`define ref_T1_t1Probe_laneProbes_14_slots_0_writeMask verification.probeWire_laneProbes_14_slots_0_writeMask_probe
`define ref_T1_t1Probe_laneProbes_14_slots_1_stage0EnqueueReady verification.probeWire_laneProbes_14_slots_1_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_14_slots_1_stage0EnqueueValid verification.probeWire_laneProbes_14_slots_1_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_14_slots_1_changingMaskSet verification.probeWire_laneProbes_14_slots_1_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_14_slots_1_slotActive verification.probeWire_laneProbes_14_slots_1_slotActive_probe
`define ref_T1_t1Probe_laneProbes_14_slots_1_slotOccupied verification.probeWire_laneProbes_14_slots_1_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_14_slots_1_pipeFinish verification.probeWire_laneProbes_14_slots_1_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_14_slots_1_slotShiftValid verification.probeWire_laneProbes_14_slots_1_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_14_slots_1_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_14_slots_1_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_14_slots_1_decodeResultIsScheduler verification.probeWire_laneProbes_14_slots_1_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_14_slots_1_executionUnitVfuRequestReady verification.probeWire_laneProbes_14_slots_1_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_14_slots_1_executionUnitVfuRequestValid verification.probeWire_laneProbes_14_slots_1_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_14_slots_1_stage3VrfWriteReady verification.probeWire_laneProbes_14_slots_1_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_14_slots_1_stage3VrfWriteValid verification.probeWire_laneProbes_14_slots_1_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_14_slots_1_writeQueueEnq verification.probeWire_laneProbes_14_slots_1_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_14_slots_1_writeTag verification.probeWire_laneProbes_14_slots_1_writeTag_probe
`define ref_T1_t1Probe_laneProbes_14_slots_1_writeMask verification.probeWire_laneProbes_14_slots_1_writeMask_probe
`define ref_T1_t1Probe_laneProbes_14_slots_2_stage0EnqueueReady verification.probeWire_laneProbes_14_slots_2_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_14_slots_2_stage0EnqueueValid verification.probeWire_laneProbes_14_slots_2_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_14_slots_2_changingMaskSet verification.probeWire_laneProbes_14_slots_2_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_14_slots_2_slotActive verification.probeWire_laneProbes_14_slots_2_slotActive_probe
`define ref_T1_t1Probe_laneProbes_14_slots_2_slotOccupied verification.probeWire_laneProbes_14_slots_2_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_14_slots_2_pipeFinish verification.probeWire_laneProbes_14_slots_2_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_14_slots_2_slotShiftValid verification.probeWire_laneProbes_14_slots_2_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_14_slots_2_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_14_slots_2_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_14_slots_2_decodeResultIsScheduler verification.probeWire_laneProbes_14_slots_2_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_14_slots_2_executionUnitVfuRequestReady verification.probeWire_laneProbes_14_slots_2_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_14_slots_2_executionUnitVfuRequestValid verification.probeWire_laneProbes_14_slots_2_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_14_slots_2_stage3VrfWriteReady verification.probeWire_laneProbes_14_slots_2_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_14_slots_2_stage3VrfWriteValid verification.probeWire_laneProbes_14_slots_2_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_14_slots_2_writeQueueEnq verification.probeWire_laneProbes_14_slots_2_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_14_slots_2_writeTag verification.probeWire_laneProbes_14_slots_2_writeTag_probe
`define ref_T1_t1Probe_laneProbes_14_slots_2_writeMask verification.probeWire_laneProbes_14_slots_2_writeMask_probe
`define ref_T1_t1Probe_laneProbes_14_slots_3_stage0EnqueueReady verification.probeWire_laneProbes_14_slots_3_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_14_slots_3_stage0EnqueueValid verification.probeWire_laneProbes_14_slots_3_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_14_slots_3_changingMaskSet verification.probeWire_laneProbes_14_slots_3_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_14_slots_3_slotActive verification.probeWire_laneProbes_14_slots_3_slotActive_probe
`define ref_T1_t1Probe_laneProbes_14_slots_3_slotOccupied verification.probeWire_laneProbes_14_slots_3_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_14_slots_3_pipeFinish verification.probeWire_laneProbes_14_slots_3_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_14_slots_3_slotShiftValid verification.probeWire_laneProbes_14_slots_3_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_14_slots_3_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_14_slots_3_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_14_slots_3_decodeResultIsScheduler verification.probeWire_laneProbes_14_slots_3_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_14_slots_3_executionUnitVfuRequestReady verification.probeWire_laneProbes_14_slots_3_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_14_slots_3_executionUnitVfuRequestValid verification.probeWire_laneProbes_14_slots_3_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_14_slots_3_stage3VrfWriteReady verification.probeWire_laneProbes_14_slots_3_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_14_slots_3_stage3VrfWriteValid verification.probeWire_laneProbes_14_slots_3_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_14_slots_3_writeQueueEnq verification.probeWire_laneProbes_14_slots_3_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_14_slots_3_writeTag verification.probeWire_laneProbes_14_slots_3_writeTag_probe
`define ref_T1_t1Probe_laneProbes_14_slots_3_writeMask verification.probeWire_laneProbes_14_slots_3_writeMask_probe
`define ref_T1_t1Probe_laneProbes_14_laneRequestStall verification.probeWire_laneProbes_14_laneRequestStall_probe
`define ref_T1_t1Probe_laneProbes_14_lastSlotOccupied verification.probeWire_laneProbes_14_lastSlotOccupied_probe
`define ref_T1_t1Probe_laneProbes_14_instructionFinished verification.probeWire_laneProbes_14_instructionFinished_probe
`define ref_T1_t1Probe_laneProbes_14_instructionValid verification.probeWire_laneProbes_14_instructionValid_probe
`define ref_T1_t1Probe_laneProbes_14_crossWriteProbe_0_valid verification.probeWire_laneProbes_14_crossWriteProbe_0_valid_probe
`define ref_T1_t1Probe_laneProbes_14_crossWriteProbe_0_bits_writeTag verification.probeWire_laneProbes_14_crossWriteProbe_0_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_14_crossWriteProbe_0_bits_writeMask verification.probeWire_laneProbes_14_crossWriteProbe_0_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_14_crossWriteProbe_1_valid verification.probeWire_laneProbes_14_crossWriteProbe_1_valid_probe
`define ref_T1_t1Probe_laneProbes_14_crossWriteProbe_1_bits_writeTag verification.probeWire_laneProbes_14_crossWriteProbe_1_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_14_crossWriteProbe_1_bits_writeMask verification.probeWire_laneProbes_14_crossWriteProbe_1_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_14_vrfProbe_valid verification.probeWire_laneProbes_14_vrfProbe_valid_probe
`define ref_T1_t1Probe_laneProbes_14_vrfProbe_requestVd verification.probeWire_laneProbes_14_vrfProbe_requestVd_probe
`define ref_T1_t1Probe_laneProbes_14_vrfProbe_requestOffset verification.probeWire_laneProbes_14_vrfProbe_requestOffset_probe
`define ref_T1_t1Probe_laneProbes_14_vrfProbe_requestMask verification.probeWire_laneProbes_14_vrfProbe_requestMask_probe
`define ref_T1_t1Probe_laneProbes_14_vrfProbe_requestData verification.probeWire_laneProbes_14_vrfProbe_requestData_probe
`define ref_T1_t1Probe_laneProbes_14_vrfProbe_requestInstruction verification.probeWire_laneProbes_14_vrfProbe_requestInstruction_probe
`define ref_T1_t1Probe_laneProbes_15_slots_0_stage0EnqueueReady verification.probeWire_laneProbes_15_slots_0_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_15_slots_0_stage0EnqueueValid verification.probeWire_laneProbes_15_slots_0_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_15_slots_0_changingMaskSet verification.probeWire_laneProbes_15_slots_0_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_15_slots_0_slotActive verification.probeWire_laneProbes_15_slots_0_slotActive_probe
`define ref_T1_t1Probe_laneProbes_15_slots_0_slotOccupied verification.probeWire_laneProbes_15_slots_0_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_15_slots_0_pipeFinish verification.probeWire_laneProbes_15_slots_0_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_15_slots_0_slotShiftValid verification.probeWire_laneProbes_15_slots_0_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_15_slots_0_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_15_slots_0_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_15_slots_0_decodeResultIsScheduler verification.probeWire_laneProbes_15_slots_0_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_15_slots_0_executionUnitVfuRequestReady verification.probeWire_laneProbes_15_slots_0_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_15_slots_0_executionUnitVfuRequestValid verification.probeWire_laneProbes_15_slots_0_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_15_slots_0_stage3VrfWriteReady verification.probeWire_laneProbes_15_slots_0_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_15_slots_0_stage3VrfWriteValid verification.probeWire_laneProbes_15_slots_0_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_15_slots_0_writeQueueEnq verification.probeWire_laneProbes_15_slots_0_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_15_slots_0_writeTag verification.probeWire_laneProbes_15_slots_0_writeTag_probe
`define ref_T1_t1Probe_laneProbes_15_slots_0_writeMask verification.probeWire_laneProbes_15_slots_0_writeMask_probe
`define ref_T1_t1Probe_laneProbes_15_slots_1_stage0EnqueueReady verification.probeWire_laneProbes_15_slots_1_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_15_slots_1_stage0EnqueueValid verification.probeWire_laneProbes_15_slots_1_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_15_slots_1_changingMaskSet verification.probeWire_laneProbes_15_slots_1_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_15_slots_1_slotActive verification.probeWire_laneProbes_15_slots_1_slotActive_probe
`define ref_T1_t1Probe_laneProbes_15_slots_1_slotOccupied verification.probeWire_laneProbes_15_slots_1_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_15_slots_1_pipeFinish verification.probeWire_laneProbes_15_slots_1_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_15_slots_1_slotShiftValid verification.probeWire_laneProbes_15_slots_1_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_15_slots_1_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_15_slots_1_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_15_slots_1_decodeResultIsScheduler verification.probeWire_laneProbes_15_slots_1_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_15_slots_1_executionUnitVfuRequestReady verification.probeWire_laneProbes_15_slots_1_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_15_slots_1_executionUnitVfuRequestValid verification.probeWire_laneProbes_15_slots_1_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_15_slots_1_stage3VrfWriteReady verification.probeWire_laneProbes_15_slots_1_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_15_slots_1_stage3VrfWriteValid verification.probeWire_laneProbes_15_slots_1_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_15_slots_1_writeQueueEnq verification.probeWire_laneProbes_15_slots_1_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_15_slots_1_writeTag verification.probeWire_laneProbes_15_slots_1_writeTag_probe
`define ref_T1_t1Probe_laneProbes_15_slots_1_writeMask verification.probeWire_laneProbes_15_slots_1_writeMask_probe
`define ref_T1_t1Probe_laneProbes_15_slots_2_stage0EnqueueReady verification.probeWire_laneProbes_15_slots_2_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_15_slots_2_stage0EnqueueValid verification.probeWire_laneProbes_15_slots_2_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_15_slots_2_changingMaskSet verification.probeWire_laneProbes_15_slots_2_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_15_slots_2_slotActive verification.probeWire_laneProbes_15_slots_2_slotActive_probe
`define ref_T1_t1Probe_laneProbes_15_slots_2_slotOccupied verification.probeWire_laneProbes_15_slots_2_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_15_slots_2_pipeFinish verification.probeWire_laneProbes_15_slots_2_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_15_slots_2_slotShiftValid verification.probeWire_laneProbes_15_slots_2_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_15_slots_2_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_15_slots_2_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_15_slots_2_decodeResultIsScheduler verification.probeWire_laneProbes_15_slots_2_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_15_slots_2_executionUnitVfuRequestReady verification.probeWire_laneProbes_15_slots_2_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_15_slots_2_executionUnitVfuRequestValid verification.probeWire_laneProbes_15_slots_2_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_15_slots_2_stage3VrfWriteReady verification.probeWire_laneProbes_15_slots_2_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_15_slots_2_stage3VrfWriteValid verification.probeWire_laneProbes_15_slots_2_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_15_slots_2_writeQueueEnq verification.probeWire_laneProbes_15_slots_2_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_15_slots_2_writeTag verification.probeWire_laneProbes_15_slots_2_writeTag_probe
`define ref_T1_t1Probe_laneProbes_15_slots_2_writeMask verification.probeWire_laneProbes_15_slots_2_writeMask_probe
`define ref_T1_t1Probe_laneProbes_15_slots_3_stage0EnqueueReady verification.probeWire_laneProbes_15_slots_3_stage0EnqueueReady_probe
`define ref_T1_t1Probe_laneProbes_15_slots_3_stage0EnqueueValid verification.probeWire_laneProbes_15_slots_3_stage0EnqueueValid_probe
`define ref_T1_t1Probe_laneProbes_15_slots_3_changingMaskSet verification.probeWire_laneProbes_15_slots_3_changingMaskSet_probe
`define ref_T1_t1Probe_laneProbes_15_slots_3_slotActive verification.probeWire_laneProbes_15_slots_3_slotActive_probe
`define ref_T1_t1Probe_laneProbes_15_slots_3_slotOccupied verification.probeWire_laneProbes_15_slots_3_slotOccupied_probe
`define ref_T1_t1Probe_laneProbes_15_slots_3_pipeFinish verification.probeWire_laneProbes_15_slots_3_pipeFinish_probe
`define ref_T1_t1Probe_laneProbes_15_slots_3_slotShiftValid verification.probeWire_laneProbes_15_slots_3_slotShiftValid_probe
`define ref_T1_t1Probe_laneProbes_15_slots_3_decodeResultIsCrossReadOrWrite verification.probeWire_laneProbes_15_slots_3_decodeResultIsCrossReadOrWrite_probe
`define ref_T1_t1Probe_laneProbes_15_slots_3_decodeResultIsScheduler verification.probeWire_laneProbes_15_slots_3_decodeResultIsScheduler_probe
`define ref_T1_t1Probe_laneProbes_15_slots_3_executionUnitVfuRequestReady verification.probeWire_laneProbes_15_slots_3_executionUnitVfuRequestReady_probe
`define ref_T1_t1Probe_laneProbes_15_slots_3_executionUnitVfuRequestValid verification.probeWire_laneProbes_15_slots_3_executionUnitVfuRequestValid_probe
`define ref_T1_t1Probe_laneProbes_15_slots_3_stage3VrfWriteReady verification.probeWire_laneProbes_15_slots_3_stage3VrfWriteReady_probe
`define ref_T1_t1Probe_laneProbes_15_slots_3_stage3VrfWriteValid verification.probeWire_laneProbes_15_slots_3_stage3VrfWriteValid_probe
`define ref_T1_t1Probe_laneProbes_15_slots_3_writeQueueEnq verification.probeWire_laneProbes_15_slots_3_writeQueueEnq_probe
`define ref_T1_t1Probe_laneProbes_15_slots_3_writeTag verification.probeWire_laneProbes_15_slots_3_writeTag_probe
`define ref_T1_t1Probe_laneProbes_15_slots_3_writeMask verification.probeWire_laneProbes_15_slots_3_writeMask_probe
`define ref_T1_t1Probe_laneProbes_15_laneRequestStall verification.probeWire_laneProbes_15_laneRequestStall_probe
`define ref_T1_t1Probe_laneProbes_15_lastSlotOccupied verification.probeWire_laneProbes_15_lastSlotOccupied_probe
`define ref_T1_t1Probe_laneProbes_15_instructionFinished verification.probeWire_laneProbes_15_instructionFinished_probe
`define ref_T1_t1Probe_laneProbes_15_instructionValid verification.probeWire_laneProbes_15_instructionValid_probe
`define ref_T1_t1Probe_laneProbes_15_crossWriteProbe_0_valid verification.probeWire_laneProbes_15_crossWriteProbe_0_valid_probe
`define ref_T1_t1Probe_laneProbes_15_crossWriteProbe_0_bits_writeTag verification.probeWire_laneProbes_15_crossWriteProbe_0_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_15_crossWriteProbe_0_bits_writeMask verification.probeWire_laneProbes_15_crossWriteProbe_0_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_15_crossWriteProbe_1_valid verification.probeWire_laneProbes_15_crossWriteProbe_1_valid_probe
`define ref_T1_t1Probe_laneProbes_15_crossWriteProbe_1_bits_writeTag verification.probeWire_laneProbes_15_crossWriteProbe_1_bits_writeTag_probe
`define ref_T1_t1Probe_laneProbes_15_crossWriteProbe_1_bits_writeMask verification.probeWire_laneProbes_15_crossWriteProbe_1_bits_writeMask_probe
`define ref_T1_t1Probe_laneProbes_15_vrfProbe_valid verification.probeWire_laneProbes_15_vrfProbe_valid_probe
`define ref_T1_t1Probe_laneProbes_15_vrfProbe_requestVd verification.probeWire_laneProbes_15_vrfProbe_requestVd_probe
`define ref_T1_t1Probe_laneProbes_15_vrfProbe_requestOffset verification.probeWire_laneProbes_15_vrfProbe_requestOffset_probe
`define ref_T1_t1Probe_laneProbes_15_vrfProbe_requestMask verification.probeWire_laneProbes_15_vrfProbe_requestMask_probe
`define ref_T1_t1Probe_laneProbes_15_vrfProbe_requestData verification.probeWire_laneProbes_15_vrfProbe_requestData_probe
`define ref_T1_t1Probe_laneProbes_15_vrfProbe_requestInstruction verification.probeWire_laneProbes_15_vrfProbe_requestInstruction_probe
`define ref_T1_t1Probe_issue_valid verification.probeWire_issue_valid_probe
`define ref_T1_t1Probe_issue_bits verification.probeWire_issue_bits_probe
`define ref_T1_t1Probe_retire_valid verification.probeWire_retire_valid_probe
`define ref_T1_t1Probe_retire_bits verification.probeWire_retire_bits_probe
`define ref_T1_t1Probe_idle verification.probeWire_idle_probe
