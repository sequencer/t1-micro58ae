module Rec7Fn(
  input  [31:0] in_data,
  input  [9:0]  in_classifyIn,
  input  [2:0]  in_roundingMode,
  output [31:0] out_data,
  output [4:0]  out_exceptionFlags
);

  wire         sign = in_data[31];
  wire [7:0]   expIn = in_data[30:23];
  wire [22:0]  fractIn = in_data[22:0];
  wire         inIsPositiveInf = in_classifyIn[7];
  wire         inIsNegativeInf = in_classifyIn[0];
  wire         inIsNegativeZero = in_classifyIn[3];
  wire         inIsPositveZero = in_classifyIn[4];
  wire         inIsSNaN = in_classifyIn[8];
  wire         inIsQNaN = in_classifyIn[9];
  wire         inIsSub = in_classifyIn[2] | in_classifyIn[5];
  wire         inIsSubMayberound = inIsSub & in_data[22:21] == 2'h0;
  wire         _maybyRoundToNegaInf_T_3 = in_roundingMode == 3'h2;
  wire         _maybyRoundToPosInf_T_4 = in_roundingMode == 3'h3;
  wire         maybeRoundToMax = in_roundingMode == 3'h1 | _maybyRoundToNegaInf_T_3 & ~sign | _maybyRoundToPosInf_T_4 & sign;
  wire         _maybyRoundToPosInf_T_1 = in_roundingMode == 3'h0;
  wire         _maybyRoundToPosInf_T_2 = in_roundingMode == 3'h4;
  wire         maybyRoundToNegaInf = sign & (_maybyRoundToPosInf_T_1 | _maybyRoundToPosInf_T_2 | _maybyRoundToNegaInf_T_3);
  wire         maybyRoundToPosInf = ~sign & (_maybyRoundToPosInf_T_1 | _maybyRoundToPosInf_T_2 | _maybyRoundToPosInf_T_4);
  wire         roundAbnormalToMax = inIsSubMayberound & maybeRoundToMax;
  wire         roundAbnormalToNegaInf = inIsSubMayberound & maybyRoundToNegaInf;
  wire         roundAbnormalToPosInf = inIsSubMayberound & maybyRoundToPosInf;
  wire         roundAbnormal = roundAbnormalToPosInf | roundAbnormalToNegaInf | roundAbnormalToMax;
  wire [7:0]   normDist =
    {3'h0,
     fractIn[22]
       ? 5'h0
       : fractIn[21]
           ? 5'h1
           : fractIn[20]
               ? 5'h2
               : fractIn[19]
                   ? 5'h3
                   : fractIn[18]
                       ? 5'h4
                       : fractIn[17]
                           ? 5'h5
                           : fractIn[16]
                               ? 5'h6
                               : fractIn[15]
                                   ? 5'h7
                                   : fractIn[14]
                                       ? 5'h8
                                       : fractIn[13]
                                           ? 5'h9
                                           : fractIn[12]
                                               ? 5'hA
                                               : fractIn[11]
                                                   ? 5'hB
                                                   : fractIn[10]
                                                       ? 5'hC
                                                       : fractIn[9]
                                                           ? 5'hD
                                                           : fractIn[8] ? 5'hE : fractIn[7] ? 5'hF : fractIn[6] ? 5'h10 : fractIn[5] ? 5'h11 : fractIn[4] ? 5'h12 : fractIn[3] ? 5'h13 : fractIn[2] ? 5'h14 : fractIn[1] ? 5'h15 : 5'h16};
  wire [7:0]   normExpIn = inIsSub ? 8'h0 - normDist : expIn;
  wire [278:0] _normSigIn_T_1 = {255'h0, fractIn, 1'h0} << normDist;
  wire [22:0]  normSigIn = inIsSub ? _normSigIn_T_1[22:0] : fractIn;
  wire [6:0]   normSigOut_plaInput = normSigIn[22:16];
  wire [6:0]   normSigOut_invInputs = ~normSigOut_plaInput;
  wire [6:0]   normSigOut_invMatrixOutputs;
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_2 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_4 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_5 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_7 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_10 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_14 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_16 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_17 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_18 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_19 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_22 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_25 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_27 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_28 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_34 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_39 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_42 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_43 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_46 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_47 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_52 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_56 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_62 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_63 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_66 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_67 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_75 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_79 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_80 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_84 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_87 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_88 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_91 = normSigOut_invInputs[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_2 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_5 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_8 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_10 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_12 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_13 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_17 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_18 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_19 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_21 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_24 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_27 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_28 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_30 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_32 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_33 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_35 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_40 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_41 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_42 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_44 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_47 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_54 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_55 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_58 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_61 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_62 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_63 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_64 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_68 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_70 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_71 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_72 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_76 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_79 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_80 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_82 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_86 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_87 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_89 = normSigOut_invInputs[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_1 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_1 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_3 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_4 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_4 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_6 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_9 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_8 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_11 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_12 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_6 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_7 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_15 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_14 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_9 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_12 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_13 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_22 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_38 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_39 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_45 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_44 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_37 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_49 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_53 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_60 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_62 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_65 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_68 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_59 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_72 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_83 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_85 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_84 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_85 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_86 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_87 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_88 = normSigOut_invInputs[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_1 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_2 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_6 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_7 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_9 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_4 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_11 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_10 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_13 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_17 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_2 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_3 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_20 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_17 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_24 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_19 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_4 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_28 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_29 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_5 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_26 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_27 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_34 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_29 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_30 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_63 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_64 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_65 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_66 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_67 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_58 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_60 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_71 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_62 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_73 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_74 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_77 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_67 = normSigOut_invInputs[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_79 = normSigOut_invInputs[5];
  wire [1:0]   normSigOut_andMatrixOutputs_lo = {normSigOut_andMatrixOutputs_andMatrixInput_2, normSigOut_andMatrixOutputs_andMatrixInput_3};
  wire [1:0]   normSigOut_andMatrixOutputs_hi = {normSigOut_andMatrixOutputs_andMatrixInput_0, normSigOut_andMatrixOutputs_andMatrixInput_1};
  wire         normSigOut_andMatrixOutputs_37_2 = &{normSigOut_andMatrixOutputs_hi, normSigOut_andMatrixOutputs_lo};
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_1 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_3 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_4 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_6 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_7 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_8 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_10 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_13 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_14 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_15 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_21 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_23 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_27 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_28 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_29 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_35 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_36 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_39 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_40 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_47 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_48 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_50 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_55 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_56 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_58 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_59 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_67 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_68 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_69 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_75 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_76 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_78 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_79 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_81 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_82 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_83 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_84 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_88 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_89 = normSigOut_invInputs[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_92 = normSigOut_invInputs[2];
  wire [1:0]   normSigOut_andMatrixOutputs_hi_1 = {normSigOut_andMatrixOutputs_andMatrixInput_0_1, normSigOut_andMatrixOutputs_andMatrixInput_1_1};
  wire         normSigOut_andMatrixOutputs_62_2 = &{normSigOut_andMatrixOutputs_hi_1, normSigOut_andMatrixOutputs_andMatrixInput_2_1};
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_2 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_3 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_5 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_6 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_7 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_8 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_11 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_12 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_11 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_12 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_16 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_15 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_16 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_18 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_27 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_31 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_30 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_31 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_39 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_41 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_43 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_44 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_45 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_46 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_55 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_57 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_57 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_62 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_61 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_64 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_65 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_77 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_76 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_83 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_82 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_85 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_86 = normSigOut_invInputs[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_93 = normSigOut_invInputs[3];
  wire [1:0]   normSigOut_andMatrixOutputs_lo_1 = {normSigOut_andMatrixOutputs_andMatrixInput_3_1, normSigOut_andMatrixOutputs_andMatrixInput_4};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi = {normSigOut_andMatrixOutputs_andMatrixInput_0_2, normSigOut_andMatrixOutputs_andMatrixInput_1_2};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_2 = {normSigOut_andMatrixOutputs_hi_hi, normSigOut_andMatrixOutputs_andMatrixInput_2_2};
  wire         normSigOut_andMatrixOutputs_61_2 = &{normSigOut_andMatrixOutputs_hi_2, normSigOut_andMatrixOutputs_lo_1};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_2 = {normSigOut_andMatrixOutputs_andMatrixInput_2_3, normSigOut_andMatrixOutputs_andMatrixInput_3_2};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_3 = {normSigOut_andMatrixOutputs_andMatrixInput_0_3, normSigOut_andMatrixOutputs_andMatrixInput_1_3};
  wire         normSigOut_andMatrixOutputs_41_2 = &{normSigOut_andMatrixOutputs_hi_3, normSigOut_andMatrixOutputs_lo_2};
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_3 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_1 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_5 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_2 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_3 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_9 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_9 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_5 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_1 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_8 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_10 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_11 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_6 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_6_1 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_14 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_15 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_16 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_18 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_20 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_6_2 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_22 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_23 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_6_3 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_6 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_28 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_7 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_31 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_8 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_9 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_34 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_10 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_11 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_38 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_13 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_14 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_41 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_42 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_15 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_45 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_55 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_16 = normSigOut_invInputs[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_48 = normSigOut_invInputs[6];
  wire [1:0]   normSigOut_andMatrixOutputs_lo_3 = {normSigOut_andMatrixOutputs_andMatrixInput_2_4, normSigOut_andMatrixOutputs_andMatrixInput_3_3};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_4 = {normSigOut_andMatrixOutputs_andMatrixInput_0_4, normSigOut_andMatrixOutputs_andMatrixInput_1_4};
  wire         normSigOut_andMatrixOutputs_13_2 = &{normSigOut_andMatrixOutputs_hi_4, normSigOut_andMatrixOutputs_lo_3};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_4 = {normSigOut_andMatrixOutputs_andMatrixInput_3_4, normSigOut_andMatrixOutputs_andMatrixInput_4_1};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_1 = {normSigOut_andMatrixOutputs_andMatrixInput_0_5, normSigOut_andMatrixOutputs_andMatrixInput_1_5};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_5 = {normSigOut_andMatrixOutputs_hi_hi_1, normSigOut_andMatrixOutputs_andMatrixInput_2_5};
  wire         normSigOut_andMatrixOutputs_65_2 = &{normSigOut_andMatrixOutputs_hi_5, normSigOut_andMatrixOutputs_lo_4};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_5 = {normSigOut_andMatrixOutputs_andMatrixInput_2_6, normSigOut_andMatrixOutputs_andMatrixInput_3_5};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_6 = {normSigOut_andMatrixOutputs_andMatrixInput_0_6, normSigOut_andMatrixOutputs_andMatrixInput_1_6};
  wire         normSigOut_andMatrixOutputs_83_2 = &{normSigOut_andMatrixOutputs_hi_6, normSigOut_andMatrixOutputs_lo_5};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_6 = {normSigOut_andMatrixOutputs_andMatrixInput_3_6, normSigOut_andMatrixOutputs_andMatrixInput_4_2};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_2 = {normSigOut_andMatrixOutputs_andMatrixInput_0_7, normSigOut_andMatrixOutputs_andMatrixInput_1_7};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_7 = {normSigOut_andMatrixOutputs_hi_hi_2, normSigOut_andMatrixOutputs_andMatrixInput_2_7};
  wire         normSigOut_andMatrixOutputs_35_2 = &{normSigOut_andMatrixOutputs_hi_7, normSigOut_andMatrixOutputs_lo_6};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_7 = {normSigOut_andMatrixOutputs_andMatrixInput_3_7, normSigOut_andMatrixOutputs_andMatrixInput_4_3};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_3 = {normSigOut_andMatrixOutputs_andMatrixInput_0_8, normSigOut_andMatrixOutputs_andMatrixInput_1_8};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_8 = {normSigOut_andMatrixOutputs_hi_hi_3, normSigOut_andMatrixOutputs_andMatrixInput_2_8};
  wire         normSigOut_andMatrixOutputs_47_2 = &{normSigOut_andMatrixOutputs_hi_8, normSigOut_andMatrixOutputs_lo_7};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_9 = {normSigOut_andMatrixOutputs_andMatrixInput_0_9, normSigOut_andMatrixOutputs_andMatrixInput_1_9};
  wire         normSigOut_andMatrixOutputs_39_2 = &{normSigOut_andMatrixOutputs_hi_9, normSigOut_andMatrixOutputs_andMatrixInput_2_9};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi = {normSigOut_andMatrixOutputs_andMatrixInput_3_8, normSigOut_andMatrixOutputs_andMatrixInput_4_4};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_8 = {normSigOut_andMatrixOutputs_lo_hi, normSigOut_andMatrixOutputs_andMatrixInput_5};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_4 = {normSigOut_andMatrixOutputs_andMatrixInput_0_10, normSigOut_andMatrixOutputs_andMatrixInput_1_10};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_10 = {normSigOut_andMatrixOutputs_hi_hi_4, normSigOut_andMatrixOutputs_andMatrixInput_2_10};
  wire         normSigOut_andMatrixOutputs_11_2 = &{normSigOut_andMatrixOutputs_hi_10, normSigOut_andMatrixOutputs_lo_8};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_9 = {normSigOut_andMatrixOutputs_andMatrixInput_2_11, normSigOut_andMatrixOutputs_andMatrixInput_3_9};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_11 = {normSigOut_andMatrixOutputs_andMatrixInput_0_11, normSigOut_andMatrixOutputs_andMatrixInput_1_11};
  wire         normSigOut_andMatrixOutputs_78_2 = &{normSigOut_andMatrixOutputs_hi_11, normSigOut_andMatrixOutputs_lo_9};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_10 = {normSigOut_andMatrixOutputs_andMatrixInput_3_10, normSigOut_andMatrixOutputs_andMatrixInput_4_5};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_5 = {normSigOut_andMatrixOutputs_andMatrixInput_0_12, normSigOut_andMatrixOutputs_andMatrixInput_1_12};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_12 = {normSigOut_andMatrixOutputs_hi_hi_5, normSigOut_andMatrixOutputs_andMatrixInput_2_12};
  wire         normSigOut_andMatrixOutputs_7_2 = &{normSigOut_andMatrixOutputs_hi_12, normSigOut_andMatrixOutputs_lo_10};
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_13 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_20 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_21 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_23 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_29 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_32 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_33 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_37 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_40 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_41 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_48 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_49 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_50 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_51 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_54 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_58 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_59 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_60 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_61 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_69 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_70 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_71 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_72 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_78 = normSigOut_plaInput[0];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_82 = normSigOut_plaInput[0];
  wire [1:0]   normSigOut_andMatrixOutputs_lo_11 = {normSigOut_andMatrixOutputs_andMatrixInput_3_11, normSigOut_andMatrixOutputs_andMatrixInput_4_6};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_6 = {normSigOut_andMatrixOutputs_andMatrixInput_0_13, normSigOut_andMatrixOutputs_andMatrixInput_1_13};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_13 = {normSigOut_andMatrixOutputs_hi_hi_6, normSigOut_andMatrixOutputs_andMatrixInput_2_13};
  wire         normSigOut_andMatrixOutputs_52_2 = &{normSigOut_andMatrixOutputs_hi_13, normSigOut_andMatrixOutputs_lo_11};
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_14 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_15 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_20 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_22 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_23 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_25 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_26 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_29 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_34 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_37 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_38 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_48 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_49 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_50 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_51 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_59 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_60 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_66 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_73 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_74 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_78 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_84 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_90 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_91 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_92 = normSigOut_plaInput[1];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_93 = normSigOut_plaInput[1];
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_1 = {normSigOut_andMatrixOutputs_andMatrixInput_3_12, normSigOut_andMatrixOutputs_andMatrixInput_4_7};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_12 = {normSigOut_andMatrixOutputs_lo_hi_1, normSigOut_andMatrixOutputs_andMatrixInput_5_1};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_7 = {normSigOut_andMatrixOutputs_andMatrixInput_0_14, normSigOut_andMatrixOutputs_andMatrixInput_1_14};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_14 = {normSigOut_andMatrixOutputs_hi_hi_7, normSigOut_andMatrixOutputs_andMatrixInput_2_14};
  wire         normSigOut_andMatrixOutputs_67_2 = &{normSigOut_andMatrixOutputs_hi_14, normSigOut_andMatrixOutputs_lo_12};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_13 = {normSigOut_andMatrixOutputs_andMatrixInput_3_13, normSigOut_andMatrixOutputs_andMatrixInput_4_8};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_8 = {normSigOut_andMatrixOutputs_andMatrixInput_0_15, normSigOut_andMatrixOutputs_andMatrixInput_1_15};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_15 = {normSigOut_andMatrixOutputs_hi_hi_8, normSigOut_andMatrixOutputs_andMatrixInput_2_15};
  wire         normSigOut_andMatrixOutputs_64_2 = &{normSigOut_andMatrixOutputs_hi_15, normSigOut_andMatrixOutputs_lo_13};
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_16 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_17 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_18 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_19 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_20 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_24 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_25 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_26 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_30 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_31 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_32 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_33 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_34 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_38 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_42 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_43 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_44 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_45 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_46 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_52 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_53 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_54 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_61 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_63 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_64 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_65 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_66 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_71 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_72 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_73 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_74 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_0_85 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_86 = normSigOut_plaInput[2];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_90 = normSigOut_plaInput[2];
  wire [1:0]   normSigOut_andMatrixOutputs_lo_14 = {normSigOut_andMatrixOutputs_andMatrixInput_2_16, normSigOut_andMatrixOutputs_andMatrixInput_3_14};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_16 = {normSigOut_andMatrixOutputs_andMatrixInput_0_16, normSigOut_andMatrixOutputs_andMatrixInput_1_16};
  wire         normSigOut_andMatrixOutputs_51_2 = &{normSigOut_andMatrixOutputs_hi_16, normSigOut_andMatrixOutputs_lo_14};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_15 = {normSigOut_andMatrixOutputs_andMatrixInput_3_15, normSigOut_andMatrixOutputs_andMatrixInput_4_9};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_9 = {normSigOut_andMatrixOutputs_andMatrixInput_0_17, normSigOut_andMatrixOutputs_andMatrixInput_1_17};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_17 = {normSigOut_andMatrixOutputs_hi_hi_9, normSigOut_andMatrixOutputs_andMatrixInput_2_17};
  wire         normSigOut_andMatrixOutputs_90_2 = &{normSigOut_andMatrixOutputs_hi_17, normSigOut_andMatrixOutputs_lo_15};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_16 = {normSigOut_andMatrixOutputs_andMatrixInput_3_16, normSigOut_andMatrixOutputs_andMatrixInput_4_10};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_10 = {normSigOut_andMatrixOutputs_andMatrixInput_0_18, normSigOut_andMatrixOutputs_andMatrixInput_1_18};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_18 = {normSigOut_andMatrixOutputs_hi_hi_10, normSigOut_andMatrixOutputs_andMatrixInput_2_18};
  wire         normSigOut_andMatrixOutputs_63_2 = &{normSigOut_andMatrixOutputs_hi_18, normSigOut_andMatrixOutputs_lo_16};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_17 = {normSigOut_andMatrixOutputs_andMatrixInput_3_17, normSigOut_andMatrixOutputs_andMatrixInput_4_11};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_11 = {normSigOut_andMatrixOutputs_andMatrixInput_0_19, normSigOut_andMatrixOutputs_andMatrixInput_1_19};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_19 = {normSigOut_andMatrixOutputs_hi_hi_11, normSigOut_andMatrixOutputs_andMatrixInput_2_19};
  wire         normSigOut_andMatrixOutputs_71_2 = &{normSigOut_andMatrixOutputs_hi_19, normSigOut_andMatrixOutputs_lo_17};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_2 = {normSigOut_andMatrixOutputs_andMatrixInput_4_12, normSigOut_andMatrixOutputs_andMatrixInput_5_2};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_18 = {normSigOut_andMatrixOutputs_lo_hi_2, normSigOut_andMatrixOutputs_andMatrixInput_6};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_lo = {normSigOut_andMatrixOutputs_andMatrixInput_2_20, normSigOut_andMatrixOutputs_andMatrixInput_3_18};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_12 = {normSigOut_andMatrixOutputs_andMatrixInput_0_20, normSigOut_andMatrixOutputs_andMatrixInput_1_20};
  wire [3:0]   normSigOut_andMatrixOutputs_hi_20 = {normSigOut_andMatrixOutputs_hi_hi_12, normSigOut_andMatrixOutputs_hi_lo};
  wire         normSigOut_andMatrixOutputs_92_2 = &{normSigOut_andMatrixOutputs_hi_20, normSigOut_andMatrixOutputs_lo_18};
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_19 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_22 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_21 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_24 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_23 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_26 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_35 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_36 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_37 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_38 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_45 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_46 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_49 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_48 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_51 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_52 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_53 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_52 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_67 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_68 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_69 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_70 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_69 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_70 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_73 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_74 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_77 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_80 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_81 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_80 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_87 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_88 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_89 = normSigOut_plaInput[3];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_90 = normSigOut_plaInput[3];
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_3 = {normSigOut_andMatrixOutputs_andMatrixInput_4_13, normSigOut_andMatrixOutputs_andMatrixInput_5_3};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_19 = {normSigOut_andMatrixOutputs_lo_hi_3, normSigOut_andMatrixOutputs_andMatrixInput_6_1};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_lo_1 = {normSigOut_andMatrixOutputs_andMatrixInput_2_21, normSigOut_andMatrixOutputs_andMatrixInput_3_19};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_13 = {normSigOut_andMatrixOutputs_andMatrixInput_0_21, normSigOut_andMatrixOutputs_andMatrixInput_1_21};
  wire [3:0]   normSigOut_andMatrixOutputs_hi_21 = {normSigOut_andMatrixOutputs_hi_hi_13, normSigOut_andMatrixOutputs_hi_lo_1};
  wire         normSigOut_andMatrixOutputs_86_2 = &{normSigOut_andMatrixOutputs_hi_21, normSigOut_andMatrixOutputs_lo_19};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_20 = {normSigOut_andMatrixOutputs_andMatrixInput_3_20, normSigOut_andMatrixOutputs_andMatrixInput_4_14};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_14 = {normSigOut_andMatrixOutputs_andMatrixInput_0_22, normSigOut_andMatrixOutputs_andMatrixInput_1_22};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_22 = {normSigOut_andMatrixOutputs_hi_hi_14, normSigOut_andMatrixOutputs_andMatrixInput_2_22};
  wire         normSigOut_andMatrixOutputs_81_2 = &{normSigOut_andMatrixOutputs_hi_22, normSigOut_andMatrixOutputs_lo_20};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_21 = {normSigOut_andMatrixOutputs_andMatrixInput_3_21, normSigOut_andMatrixOutputs_andMatrixInput_4_15};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_15 = {normSigOut_andMatrixOutputs_andMatrixInput_0_23, normSigOut_andMatrixOutputs_andMatrixInput_1_23};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_23 = {normSigOut_andMatrixOutputs_hi_hi_15, normSigOut_andMatrixOutputs_andMatrixInput_2_23};
  wire         normSigOut_andMatrixOutputs_87_2 = &{normSigOut_andMatrixOutputs_hi_23, normSigOut_andMatrixOutputs_lo_21};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_22 = {normSigOut_andMatrixOutputs_andMatrixInput_3_22, normSigOut_andMatrixOutputs_andMatrixInput_4_16};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_16 = {normSigOut_andMatrixOutputs_andMatrixInput_0_24, normSigOut_andMatrixOutputs_andMatrixInput_1_24};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_24 = {normSigOut_andMatrixOutputs_hi_hi_16, normSigOut_andMatrixOutputs_andMatrixInput_2_24};
  wire         normSigOut_andMatrixOutputs_27_2 = &{normSigOut_andMatrixOutputs_hi_24, normSigOut_andMatrixOutputs_lo_22};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_23 = {normSigOut_andMatrixOutputs_andMatrixInput_3_23, normSigOut_andMatrixOutputs_andMatrixInput_4_17};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_17 = {normSigOut_andMatrixOutputs_andMatrixInput_0_25, normSigOut_andMatrixOutputs_andMatrixInput_1_25};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_25 = {normSigOut_andMatrixOutputs_hi_hi_17, normSigOut_andMatrixOutputs_andMatrixInput_2_25};
  wire         normSigOut_andMatrixOutputs_85_2 = &{normSigOut_andMatrixOutputs_hi_25, normSigOut_andMatrixOutputs_lo_23};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_24 = {normSigOut_andMatrixOutputs_andMatrixInput_3_24, normSigOut_andMatrixOutputs_andMatrixInput_4_18};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_18 = {normSigOut_andMatrixOutputs_andMatrixInput_0_26, normSigOut_andMatrixOutputs_andMatrixInput_1_26};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_26 = {normSigOut_andMatrixOutputs_hi_hi_18, normSigOut_andMatrixOutputs_andMatrixInput_2_26};
  wire         normSigOut_andMatrixOutputs_12_2 = &{normSigOut_andMatrixOutputs_hi_26, normSigOut_andMatrixOutputs_lo_24};
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_25 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_26 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_21 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_30 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_31 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_24 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_25 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_32 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_33 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_36 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_35 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_36 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_53 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_56 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_57 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_56 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_47 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_60 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_59 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_75 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_76 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_1_77 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_65 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_66 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_78 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_81 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_69 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_91 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_92 = normSigOut_plaInput[4];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_93 = normSigOut_plaInput[4];
  wire [1:0]   normSigOut_andMatrixOutputs_lo_25 = {normSigOut_andMatrixOutputs_andMatrixInput_3_25, normSigOut_andMatrixOutputs_andMatrixInput_4_19};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_19 = {normSigOut_andMatrixOutputs_andMatrixInput_0_27, normSigOut_andMatrixOutputs_andMatrixInput_1_27};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_27 = {normSigOut_andMatrixOutputs_hi_hi_19, normSigOut_andMatrixOutputs_andMatrixInput_2_27};
  wire         normSigOut_andMatrixOutputs_45_2 = &{normSigOut_andMatrixOutputs_hi_27, normSigOut_andMatrixOutputs_lo_25};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_26 = {normSigOut_andMatrixOutputs_andMatrixInput_3_26, normSigOut_andMatrixOutputs_andMatrixInput_4_20};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_20 = {normSigOut_andMatrixOutputs_andMatrixInput_0_28, normSigOut_andMatrixOutputs_andMatrixInput_1_28};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_28 = {normSigOut_andMatrixOutputs_hi_hi_20, normSigOut_andMatrixOutputs_andMatrixInput_2_28};
  wire         normSigOut_andMatrixOutputs_59_2 = &{normSigOut_andMatrixOutputs_hi_28, normSigOut_andMatrixOutputs_lo_26};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_4 = {normSigOut_andMatrixOutputs_andMatrixInput_4_21, normSigOut_andMatrixOutputs_andMatrixInput_5_4};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_27 = {normSigOut_andMatrixOutputs_lo_hi_4, normSigOut_andMatrixOutputs_andMatrixInput_6_2};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_lo_2 = {normSigOut_andMatrixOutputs_andMatrixInput_2_29, normSigOut_andMatrixOutputs_andMatrixInput_3_27};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_21 = {normSigOut_andMatrixOutputs_andMatrixInput_0_29, normSigOut_andMatrixOutputs_andMatrixInput_1_29};
  wire [3:0]   normSigOut_andMatrixOutputs_hi_29 = {normSigOut_andMatrixOutputs_hi_hi_21, normSigOut_andMatrixOutputs_hi_lo_2};
  wire         normSigOut_andMatrixOutputs_6_2 = &{normSigOut_andMatrixOutputs_hi_29, normSigOut_andMatrixOutputs_lo_27};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_28 = {normSigOut_andMatrixOutputs_andMatrixInput_3_28, normSigOut_andMatrixOutputs_andMatrixInput_4_22};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_22 = {normSigOut_andMatrixOutputs_andMatrixInput_0_30, normSigOut_andMatrixOutputs_andMatrixInput_1_30};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_30 = {normSigOut_andMatrixOutputs_hi_hi_22, normSigOut_andMatrixOutputs_andMatrixInput_2_30};
  wire         normSigOut_andMatrixOutputs_14_2 = &{normSigOut_andMatrixOutputs_hi_30, normSigOut_andMatrixOutputs_lo_28};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_29 = {normSigOut_andMatrixOutputs_andMatrixInput_3_29, normSigOut_andMatrixOutputs_andMatrixInput_4_23};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_23 = {normSigOut_andMatrixOutputs_andMatrixInput_0_31, normSigOut_andMatrixOutputs_andMatrixInput_1_31};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_31 = {normSigOut_andMatrixOutputs_hi_hi_23, normSigOut_andMatrixOutputs_andMatrixInput_2_31};
  wire         normSigOut_andMatrixOutputs_1_2 = &{normSigOut_andMatrixOutputs_hi_31, normSigOut_andMatrixOutputs_lo_29};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_30 = {normSigOut_andMatrixOutputs_andMatrixInput_3_30, normSigOut_andMatrixOutputs_andMatrixInput_4_24};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_24 = {normSigOut_andMatrixOutputs_andMatrixInput_0_32, normSigOut_andMatrixOutputs_andMatrixInput_1_32};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_32 = {normSigOut_andMatrixOutputs_hi_hi_24, normSigOut_andMatrixOutputs_andMatrixInput_2_32};
  wire         normSigOut_andMatrixOutputs_80_2 = &{normSigOut_andMatrixOutputs_hi_32, normSigOut_andMatrixOutputs_lo_30};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_5 = {normSigOut_andMatrixOutputs_andMatrixInput_4_25, normSigOut_andMatrixOutputs_andMatrixInput_5_5};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_31 = {normSigOut_andMatrixOutputs_lo_hi_5, normSigOut_andMatrixOutputs_andMatrixInput_6_3};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_lo_3 = {normSigOut_andMatrixOutputs_andMatrixInput_2_33, normSigOut_andMatrixOutputs_andMatrixInput_3_31};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_25 = {normSigOut_andMatrixOutputs_andMatrixInput_0_33, normSigOut_andMatrixOutputs_andMatrixInput_1_33};
  wire [3:0]   normSigOut_andMatrixOutputs_hi_33 = {normSigOut_andMatrixOutputs_hi_hi_25, normSigOut_andMatrixOutputs_hi_lo_3};
  wire         normSigOut_andMatrixOutputs_70_2 = &{normSigOut_andMatrixOutputs_hi_33, normSigOut_andMatrixOutputs_lo_31};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_6 = {normSigOut_andMatrixOutputs_andMatrixInput_3_32, normSigOut_andMatrixOutputs_andMatrixInput_4_26};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_32 = {normSigOut_andMatrixOutputs_lo_hi_6, normSigOut_andMatrixOutputs_andMatrixInput_5_6};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_26 = {normSigOut_andMatrixOutputs_andMatrixInput_0_34, normSigOut_andMatrixOutputs_andMatrixInput_1_34};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_34 = {normSigOut_andMatrixOutputs_hi_hi_26, normSigOut_andMatrixOutputs_andMatrixInput_2_34};
  wire         normSigOut_andMatrixOutputs_23_2 = &{normSigOut_andMatrixOutputs_hi_34, normSigOut_andMatrixOutputs_lo_32};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_33 = {normSigOut_andMatrixOutputs_andMatrixInput_3_33, normSigOut_andMatrixOutputs_andMatrixInput_4_27};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_27 = {normSigOut_andMatrixOutputs_andMatrixInput_0_35, normSigOut_andMatrixOutputs_andMatrixInput_1_35};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_35 = {normSigOut_andMatrixOutputs_hi_hi_27, normSigOut_andMatrixOutputs_andMatrixInput_2_35};
  wire         normSigOut_andMatrixOutputs_88_2 = &{normSigOut_andMatrixOutputs_hi_35, normSigOut_andMatrixOutputs_lo_33};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_34 = {normSigOut_andMatrixOutputs_andMatrixInput_3_34, normSigOut_andMatrixOutputs_andMatrixInput_4_28};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_28 = {normSigOut_andMatrixOutputs_andMatrixInput_0_36, normSigOut_andMatrixOutputs_andMatrixInput_1_36};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_36 = {normSigOut_andMatrixOutputs_hi_hi_28, normSigOut_andMatrixOutputs_andMatrixInput_2_36};
  wire         normSigOut_andMatrixOutputs_34_2 = &{normSigOut_andMatrixOutputs_hi_36, normSigOut_andMatrixOutputs_lo_34};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_35 = {normSigOut_andMatrixOutputs_andMatrixInput_3_35, normSigOut_andMatrixOutputs_andMatrixInput_4_29};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_29 = {normSigOut_andMatrixOutputs_andMatrixInput_0_37, normSigOut_andMatrixOutputs_andMatrixInput_1_37};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_37 = {normSigOut_andMatrixOutputs_hi_hi_29, normSigOut_andMatrixOutputs_andMatrixInput_2_37};
  wire         normSigOut_andMatrixOutputs_75_2 = &{normSigOut_andMatrixOutputs_hi_37, normSigOut_andMatrixOutputs_lo_35};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_7 = {normSigOut_andMatrixOutputs_andMatrixInput_3_36, normSigOut_andMatrixOutputs_andMatrixInput_4_30};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_36 = {normSigOut_andMatrixOutputs_lo_hi_7, normSigOut_andMatrixOutputs_andMatrixInput_5_7};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_30 = {normSigOut_andMatrixOutputs_andMatrixInput_0_38, normSigOut_andMatrixOutputs_andMatrixInput_1_38};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_38 = {normSigOut_andMatrixOutputs_hi_hi_30, normSigOut_andMatrixOutputs_andMatrixInput_2_38};
  wire         normSigOut_andMatrixOutputs_3_2 = &{normSigOut_andMatrixOutputs_hi_38, normSigOut_andMatrixOutputs_lo_36};
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_37 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_32 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_33 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_40 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_41 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_42 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_43 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_35 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_36 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_12 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_47 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_39 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_40 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_50 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_51 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_43 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_44 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_54 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_2_57 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_46 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_17 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_58 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_49 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_81 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_71 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_83 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_73 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_74 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_75 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_76 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_77 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_89 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_90 = normSigOut_plaInput[5];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_91 = normSigOut_plaInput[5];
  wire [1:0]   normSigOut_andMatrixOutputs_lo_37 = {normSigOut_andMatrixOutputs_andMatrixInput_3_37, normSigOut_andMatrixOutputs_andMatrixInput_4_31};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_31 = {normSigOut_andMatrixOutputs_andMatrixInput_0_39, normSigOut_andMatrixOutputs_andMatrixInput_1_39};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_39 = {normSigOut_andMatrixOutputs_hi_hi_31, normSigOut_andMatrixOutputs_andMatrixInput_2_39};
  wire         normSigOut_andMatrixOutputs_93_2 = &{normSigOut_andMatrixOutputs_hi_39, normSigOut_andMatrixOutputs_lo_37};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_8 = {normSigOut_andMatrixOutputs_andMatrixInput_3_38, normSigOut_andMatrixOutputs_andMatrixInput_4_32};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_38 = {normSigOut_andMatrixOutputs_lo_hi_8, normSigOut_andMatrixOutputs_andMatrixInput_5_8};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_32 = {normSigOut_andMatrixOutputs_andMatrixInput_0_40, normSigOut_andMatrixOutputs_andMatrixInput_1_40};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_40 = {normSigOut_andMatrixOutputs_hi_hi_32, normSigOut_andMatrixOutputs_andMatrixInput_2_40};
  wire         normSigOut_andMatrixOutputs_8_2 = &{normSigOut_andMatrixOutputs_hi_40, normSigOut_andMatrixOutputs_lo_38};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_9 = {normSigOut_andMatrixOutputs_andMatrixInput_3_39, normSigOut_andMatrixOutputs_andMatrixInput_4_33};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_39 = {normSigOut_andMatrixOutputs_lo_hi_9, normSigOut_andMatrixOutputs_andMatrixInput_5_9};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_33 = {normSigOut_andMatrixOutputs_andMatrixInput_0_41, normSigOut_andMatrixOutputs_andMatrixInput_1_41};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_41 = {normSigOut_andMatrixOutputs_hi_hi_33, normSigOut_andMatrixOutputs_andMatrixInput_2_41};
  wire         normSigOut_andMatrixOutputs_10_2 = &{normSigOut_andMatrixOutputs_hi_41, normSigOut_andMatrixOutputs_lo_39};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_40 = {normSigOut_andMatrixOutputs_andMatrixInput_2_42, normSigOut_andMatrixOutputs_andMatrixInput_3_40};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_42 = {normSigOut_andMatrixOutputs_andMatrixInput_0_42, normSigOut_andMatrixOutputs_andMatrixInput_1_42};
  wire         normSigOut_andMatrixOutputs_79_2 = &{normSigOut_andMatrixOutputs_hi_42, normSigOut_andMatrixOutputs_lo_40};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_41 = {normSigOut_andMatrixOutputs_andMatrixInput_2_43, normSigOut_andMatrixOutputs_andMatrixInput_3_41};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_43 = {normSigOut_andMatrixOutputs_andMatrixInput_0_43, normSigOut_andMatrixOutputs_andMatrixInput_1_43};
  wire         normSigOut_andMatrixOutputs_2_2 = &{normSigOut_andMatrixOutputs_hi_43, normSigOut_andMatrixOutputs_lo_41};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_42 = {normSigOut_andMatrixOutputs_andMatrixInput_2_44, normSigOut_andMatrixOutputs_andMatrixInput_3_42};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_44 = {normSigOut_andMatrixOutputs_andMatrixInput_0_44, normSigOut_andMatrixOutputs_andMatrixInput_1_44};
  wire         normSigOut_andMatrixOutputs_17_2 = &{normSigOut_andMatrixOutputs_hi_44, normSigOut_andMatrixOutputs_lo_42};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_43 = {normSigOut_andMatrixOutputs_andMatrixInput_3_43, normSigOut_andMatrixOutputs_andMatrixInput_4_34};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_34 = {normSigOut_andMatrixOutputs_andMatrixInput_0_45, normSigOut_andMatrixOutputs_andMatrixInput_1_45};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_45 = {normSigOut_andMatrixOutputs_hi_hi_34, normSigOut_andMatrixOutputs_andMatrixInput_2_45};
  wire         normSigOut_andMatrixOutputs_43_2 = &{normSigOut_andMatrixOutputs_hi_45, normSigOut_andMatrixOutputs_lo_43};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_10 = {normSigOut_andMatrixOutputs_andMatrixInput_3_44, normSigOut_andMatrixOutputs_andMatrixInput_4_35};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_44 = {normSigOut_andMatrixOutputs_lo_hi_10, normSigOut_andMatrixOutputs_andMatrixInput_5_10};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_35 = {normSigOut_andMatrixOutputs_andMatrixInput_0_46, normSigOut_andMatrixOutputs_andMatrixInput_1_46};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_46 = {normSigOut_andMatrixOutputs_hi_hi_35, normSigOut_andMatrixOutputs_andMatrixInput_2_46};
  wire         normSigOut_andMatrixOutputs_48_2 = &{normSigOut_andMatrixOutputs_hi_46, normSigOut_andMatrixOutputs_lo_44};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_11 = {normSigOut_andMatrixOutputs_andMatrixInput_3_45, normSigOut_andMatrixOutputs_andMatrixInput_4_36};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_45 = {normSigOut_andMatrixOutputs_lo_hi_11, normSigOut_andMatrixOutputs_andMatrixInput_5_11};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_36 = {normSigOut_andMatrixOutputs_andMatrixInput_0_47, normSigOut_andMatrixOutputs_andMatrixInput_1_47};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_47 = {normSigOut_andMatrixOutputs_hi_hi_36, normSigOut_andMatrixOutputs_andMatrixInput_2_47};
  wire         normSigOut_andMatrixOutputs_74_2 = &{normSigOut_andMatrixOutputs_hi_47, normSigOut_andMatrixOutputs_lo_45};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_12 = {normSigOut_andMatrixOutputs_andMatrixInput_3_46, normSigOut_andMatrixOutputs_andMatrixInput_4_37};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_46 = {normSigOut_andMatrixOutputs_lo_hi_12, normSigOut_andMatrixOutputs_andMatrixInput_5_12};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_37 = {normSigOut_andMatrixOutputs_andMatrixInput_0_48, normSigOut_andMatrixOutputs_andMatrixInput_1_48};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_48 = {normSigOut_andMatrixOutputs_hi_hi_37, normSigOut_andMatrixOutputs_andMatrixInput_2_48};
  wire         normSigOut_andMatrixOutputs_60_2 = &{normSigOut_andMatrixOutputs_hi_48, normSigOut_andMatrixOutputs_lo_46};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_47 = {normSigOut_andMatrixOutputs_andMatrixInput_3_47, normSigOut_andMatrixOutputs_andMatrixInput_4_38};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_38 = {normSigOut_andMatrixOutputs_andMatrixInput_0_49, normSigOut_andMatrixOutputs_andMatrixInput_1_49};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_49 = {normSigOut_andMatrixOutputs_hi_hi_38, normSigOut_andMatrixOutputs_andMatrixInput_2_49};
  wire         normSigOut_andMatrixOutputs_4_2 = &{normSigOut_andMatrixOutputs_hi_49, normSigOut_andMatrixOutputs_lo_47};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_13 = {normSigOut_andMatrixOutputs_andMatrixInput_3_48, normSigOut_andMatrixOutputs_andMatrixInput_4_39};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_48 = {normSigOut_andMatrixOutputs_lo_hi_13, normSigOut_andMatrixOutputs_andMatrixInput_5_13};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_39 = {normSigOut_andMatrixOutputs_andMatrixInput_0_50, normSigOut_andMatrixOutputs_andMatrixInput_1_50};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_50 = {normSigOut_andMatrixOutputs_hi_hi_39, normSigOut_andMatrixOutputs_andMatrixInput_2_50};
  wire         normSigOut_andMatrixOutputs_30_2 = &{normSigOut_andMatrixOutputs_hi_50, normSigOut_andMatrixOutputs_lo_48};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_14 = {normSigOut_andMatrixOutputs_andMatrixInput_3_49, normSigOut_andMatrixOutputs_andMatrixInput_4_40};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_49 = {normSigOut_andMatrixOutputs_lo_hi_14, normSigOut_andMatrixOutputs_andMatrixInput_5_14};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_40 = {normSigOut_andMatrixOutputs_andMatrixInput_0_51, normSigOut_andMatrixOutputs_andMatrixInput_1_51};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_51 = {normSigOut_andMatrixOutputs_hi_hi_40, normSigOut_andMatrixOutputs_andMatrixInput_2_51};
  wire         normSigOut_andMatrixOutputs_56_2 = &{normSigOut_andMatrixOutputs_hi_51, normSigOut_andMatrixOutputs_lo_49};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_50 = {normSigOut_andMatrixOutputs_andMatrixInput_3_50, normSigOut_andMatrixOutputs_andMatrixInput_4_41};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_41 = {normSigOut_andMatrixOutputs_andMatrixInput_0_52, normSigOut_andMatrixOutputs_andMatrixInput_1_52};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_52 = {normSigOut_andMatrixOutputs_hi_hi_41, normSigOut_andMatrixOutputs_andMatrixInput_2_52};
  wire         normSigOut_andMatrixOutputs_66_2 = &{normSigOut_andMatrixOutputs_hi_52, normSigOut_andMatrixOutputs_lo_50};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_51 = {normSigOut_andMatrixOutputs_andMatrixInput_3_51, normSigOut_andMatrixOutputs_andMatrixInput_4_42};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_42 = {normSigOut_andMatrixOutputs_andMatrixInput_0_53, normSigOut_andMatrixOutputs_andMatrixInput_1_53};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_53 = {normSigOut_andMatrixOutputs_hi_hi_42, normSigOut_andMatrixOutputs_andMatrixInput_2_53};
  wire         normSigOut_andMatrixOutputs_9_2 = &{normSigOut_andMatrixOutputs_hi_53, normSigOut_andMatrixOutputs_lo_51};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_15 = {normSigOut_andMatrixOutputs_andMatrixInput_3_52, normSigOut_andMatrixOutputs_andMatrixInput_4_43};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_52 = {normSigOut_andMatrixOutputs_lo_hi_15, normSigOut_andMatrixOutputs_andMatrixInput_5_15};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_43 = {normSigOut_andMatrixOutputs_andMatrixInput_0_54, normSigOut_andMatrixOutputs_andMatrixInput_1_54};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_54 = {normSigOut_andMatrixOutputs_hi_hi_43, normSigOut_andMatrixOutputs_andMatrixInput_2_54};
  wire         normSigOut_andMatrixOutputs_57_2 = &{normSigOut_andMatrixOutputs_hi_54, normSigOut_andMatrixOutputs_lo_52};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_53 = {normSigOut_andMatrixOutputs_andMatrixInput_3_53, normSigOut_andMatrixOutputs_andMatrixInput_4_44};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_44 = {normSigOut_andMatrixOutputs_andMatrixInput_0_55, normSigOut_andMatrixOutputs_andMatrixInput_1_55};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_55 = {normSigOut_andMatrixOutputs_hi_hi_44, normSigOut_andMatrixOutputs_andMatrixInput_2_55};
  wire         normSigOut_andMatrixOutputs_18_2 = &{normSigOut_andMatrixOutputs_hi_55, normSigOut_andMatrixOutputs_lo_53};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_54 = {normSigOut_andMatrixOutputs_andMatrixInput_3_54, normSigOut_andMatrixOutputs_andMatrixInput_4_45};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_45 = {normSigOut_andMatrixOutputs_andMatrixInput_0_56, normSigOut_andMatrixOutputs_andMatrixInput_1_56};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_56 = {normSigOut_andMatrixOutputs_hi_hi_45, normSigOut_andMatrixOutputs_andMatrixInput_2_56};
  wire         normSigOut_andMatrixOutputs_16_2 = &{normSigOut_andMatrixOutputs_hi_56, normSigOut_andMatrixOutputs_lo_54};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_55 = {normSigOut_andMatrixOutputs_andMatrixInput_2_57, normSigOut_andMatrixOutputs_andMatrixInput_3_55};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_57 = {normSigOut_andMatrixOutputs_andMatrixInput_0_57, normSigOut_andMatrixOutputs_andMatrixInput_1_57};
  wire         normSigOut_andMatrixOutputs_82_2 = &{normSigOut_andMatrixOutputs_hi_57, normSigOut_andMatrixOutputs_lo_55};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_16 = {normSigOut_andMatrixOutputs_andMatrixInput_3_56, normSigOut_andMatrixOutputs_andMatrixInput_4_46};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_56 = {normSigOut_andMatrixOutputs_lo_hi_16, normSigOut_andMatrixOutputs_andMatrixInput_5_16};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_46 = {normSigOut_andMatrixOutputs_andMatrixInput_0_58, normSigOut_andMatrixOutputs_andMatrixInput_1_58};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_58 = {normSigOut_andMatrixOutputs_hi_hi_46, normSigOut_andMatrixOutputs_andMatrixInput_2_58};
  wire         normSigOut_andMatrixOutputs_50_2 = &{normSigOut_andMatrixOutputs_hi_58, normSigOut_andMatrixOutputs_lo_56};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_17 = {normSigOut_andMatrixOutputs_andMatrixInput_3_57, normSigOut_andMatrixOutputs_andMatrixInput_4_47};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_57 = {normSigOut_andMatrixOutputs_lo_hi_17, normSigOut_andMatrixOutputs_andMatrixInput_5_17};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_47 = {normSigOut_andMatrixOutputs_andMatrixInput_0_59, normSigOut_andMatrixOutputs_andMatrixInput_1_59};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_59 = {normSigOut_andMatrixOutputs_hi_hi_47, normSigOut_andMatrixOutputs_andMatrixInput_2_59};
  wire         normSigOut_andMatrixOutputs_77_2 = &{normSigOut_andMatrixOutputs_hi_59, normSigOut_andMatrixOutputs_lo_57};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_58 = {normSigOut_andMatrixOutputs_andMatrixInput_3_58, normSigOut_andMatrixOutputs_andMatrixInput_4_48};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_48 = {normSigOut_andMatrixOutputs_andMatrixInput_0_60, normSigOut_andMatrixOutputs_andMatrixInput_1_60};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_60 = {normSigOut_andMatrixOutputs_hi_hi_48, normSigOut_andMatrixOutputs_andMatrixInput_2_60};
  wire         normSigOut_andMatrixOutputs_22_2 = &{normSigOut_andMatrixOutputs_hi_60, normSigOut_andMatrixOutputs_lo_58};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_59 = {normSigOut_andMatrixOutputs_andMatrixInput_3_59, normSigOut_andMatrixOutputs_andMatrixInput_4_49};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_49 = {normSigOut_andMatrixOutputs_andMatrixInput_0_61, normSigOut_andMatrixOutputs_andMatrixInput_1_61};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_61 = {normSigOut_andMatrixOutputs_hi_hi_49, normSigOut_andMatrixOutputs_andMatrixInput_2_61};
  wire         normSigOut_andMatrixOutputs_91_2 = &{normSigOut_andMatrixOutputs_hi_61, normSigOut_andMatrixOutputs_lo_59};
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_50 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_51 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_52 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_53 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_54 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_55 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_56 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_57 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_18 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_19 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_20 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_61 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_21 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_63 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_64 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_3_75 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_22 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_23 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_24 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_68 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_25 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_70 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_26 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_72 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_27 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_28 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_29 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_30 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_5_31 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_78 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_79 = normSigOut_plaInput[6];
  wire         normSigOut_andMatrixOutputs_andMatrixInput_4_80 = normSigOut_plaInput[6];
  wire [1:0]   normSigOut_andMatrixOutputs_lo_60 = {normSigOut_andMatrixOutputs_andMatrixInput_3_60, normSigOut_andMatrixOutputs_andMatrixInput_4_50};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_50 = {normSigOut_andMatrixOutputs_andMatrixInput_0_62, normSigOut_andMatrixOutputs_andMatrixInput_1_62};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_62 = {normSigOut_andMatrixOutputs_hi_hi_50, normSigOut_andMatrixOutputs_andMatrixInput_2_62};
  wire         normSigOut_andMatrixOutputs_32_2 = &{normSigOut_andMatrixOutputs_hi_62, normSigOut_andMatrixOutputs_lo_60};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_61 = {normSigOut_andMatrixOutputs_andMatrixInput_3_61, normSigOut_andMatrixOutputs_andMatrixInput_4_51};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_51 = {normSigOut_andMatrixOutputs_andMatrixInput_0_63, normSigOut_andMatrixOutputs_andMatrixInput_1_63};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_63 = {normSigOut_andMatrixOutputs_hi_hi_51, normSigOut_andMatrixOutputs_andMatrixInput_2_63};
  wire         normSigOut_andMatrixOutputs_25_2 = &{normSigOut_andMatrixOutputs_hi_63, normSigOut_andMatrixOutputs_lo_61};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_62 = {normSigOut_andMatrixOutputs_andMatrixInput_3_62, normSigOut_andMatrixOutputs_andMatrixInput_4_52};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_52 = {normSigOut_andMatrixOutputs_andMatrixInput_0_64, normSigOut_andMatrixOutputs_andMatrixInput_1_64};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_64 = {normSigOut_andMatrixOutputs_hi_hi_52, normSigOut_andMatrixOutputs_andMatrixInput_2_64};
  wire         normSigOut_andMatrixOutputs_40_2 = &{normSigOut_andMatrixOutputs_hi_64, normSigOut_andMatrixOutputs_lo_62};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_63 = {normSigOut_andMatrixOutputs_andMatrixInput_3_63, normSigOut_andMatrixOutputs_andMatrixInput_4_53};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_53 = {normSigOut_andMatrixOutputs_andMatrixInput_0_65, normSigOut_andMatrixOutputs_andMatrixInput_1_65};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_65 = {normSigOut_andMatrixOutputs_hi_hi_53, normSigOut_andMatrixOutputs_andMatrixInput_2_65};
  wire         normSigOut_andMatrixOutputs_31_2 = &{normSigOut_andMatrixOutputs_hi_65, normSigOut_andMatrixOutputs_lo_63};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_64 = {normSigOut_andMatrixOutputs_andMatrixInput_3_64, normSigOut_andMatrixOutputs_andMatrixInput_4_54};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_54 = {normSigOut_andMatrixOutputs_andMatrixInput_0_66, normSigOut_andMatrixOutputs_andMatrixInput_1_66};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_66 = {normSigOut_andMatrixOutputs_hi_hi_54, normSigOut_andMatrixOutputs_andMatrixInput_2_66};
  wire         normSigOut_andMatrixOutputs_58_2 = &{normSigOut_andMatrixOutputs_hi_66, normSigOut_andMatrixOutputs_lo_64};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_65 = {normSigOut_andMatrixOutputs_andMatrixInput_3_65, normSigOut_andMatrixOutputs_andMatrixInput_4_55};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_55 = {normSigOut_andMatrixOutputs_andMatrixInput_0_67, normSigOut_andMatrixOutputs_andMatrixInput_1_67};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_67 = {normSigOut_andMatrixOutputs_hi_hi_55, normSigOut_andMatrixOutputs_andMatrixInput_2_67};
  wire         normSigOut_andMatrixOutputs_29_2 = &{normSigOut_andMatrixOutputs_hi_67, normSigOut_andMatrixOutputs_lo_65};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_66 = {normSigOut_andMatrixOutputs_andMatrixInput_3_66, normSigOut_andMatrixOutputs_andMatrixInput_4_56};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_56 = {normSigOut_andMatrixOutputs_andMatrixInput_0_68, normSigOut_andMatrixOutputs_andMatrixInput_1_68};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_68 = {normSigOut_andMatrixOutputs_hi_hi_56, normSigOut_andMatrixOutputs_andMatrixInput_2_68};
  wire         normSigOut_andMatrixOutputs_20_2 = &{normSigOut_andMatrixOutputs_hi_68, normSigOut_andMatrixOutputs_lo_66};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_67 = {normSigOut_andMatrixOutputs_andMatrixInput_3_67, normSigOut_andMatrixOutputs_andMatrixInput_4_57};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_57 = {normSigOut_andMatrixOutputs_andMatrixInput_0_69, normSigOut_andMatrixOutputs_andMatrixInput_1_69};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_69 = {normSigOut_andMatrixOutputs_hi_hi_57, normSigOut_andMatrixOutputs_andMatrixInput_2_69};
  wire         normSigOut_andMatrixOutputs_54_2 = &{normSigOut_andMatrixOutputs_hi_69, normSigOut_andMatrixOutputs_lo_67};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_18 = {normSigOut_andMatrixOutputs_andMatrixInput_3_68, normSigOut_andMatrixOutputs_andMatrixInput_4_58};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_68 = {normSigOut_andMatrixOutputs_lo_hi_18, normSigOut_andMatrixOutputs_andMatrixInput_5_18};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_58 = {normSigOut_andMatrixOutputs_andMatrixInput_0_70, normSigOut_andMatrixOutputs_andMatrixInput_1_70};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_70 = {normSigOut_andMatrixOutputs_hi_hi_58, normSigOut_andMatrixOutputs_andMatrixInput_2_70};
  wire         normSigOut_andMatrixOutputs_38_2 = &{normSigOut_andMatrixOutputs_hi_70, normSigOut_andMatrixOutputs_lo_68};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_19 = {normSigOut_andMatrixOutputs_andMatrixInput_3_69, normSigOut_andMatrixOutputs_andMatrixInput_4_59};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_69 = {normSigOut_andMatrixOutputs_lo_hi_19, normSigOut_andMatrixOutputs_andMatrixInput_5_19};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_59 = {normSigOut_andMatrixOutputs_andMatrixInput_0_71, normSigOut_andMatrixOutputs_andMatrixInput_1_71};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_71 = {normSigOut_andMatrixOutputs_hi_hi_59, normSigOut_andMatrixOutputs_andMatrixInput_2_71};
  wire         normSigOut_andMatrixOutputs_44_2 = &{normSigOut_andMatrixOutputs_hi_71, normSigOut_andMatrixOutputs_lo_69};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_20 = {normSigOut_andMatrixOutputs_andMatrixInput_3_70, normSigOut_andMatrixOutputs_andMatrixInput_4_60};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_70 = {normSigOut_andMatrixOutputs_lo_hi_20, normSigOut_andMatrixOutputs_andMatrixInput_5_20};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_60 = {normSigOut_andMatrixOutputs_andMatrixInput_0_72, normSigOut_andMatrixOutputs_andMatrixInput_1_72};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_72 = {normSigOut_andMatrixOutputs_hi_hi_60, normSigOut_andMatrixOutputs_andMatrixInput_2_72};
  wire         normSigOut_andMatrixOutputs_46_2 = &{normSigOut_andMatrixOutputs_hi_72, normSigOut_andMatrixOutputs_lo_70};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_71 = {normSigOut_andMatrixOutputs_andMatrixInput_3_71, normSigOut_andMatrixOutputs_andMatrixInput_4_61};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_61 = {normSigOut_andMatrixOutputs_andMatrixInput_0_73, normSigOut_andMatrixOutputs_andMatrixInput_1_73};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_73 = {normSigOut_andMatrixOutputs_hi_hi_61, normSigOut_andMatrixOutputs_andMatrixInput_2_73};
  wire         normSigOut_andMatrixOutputs_26_2 = &{normSigOut_andMatrixOutputs_hi_73, normSigOut_andMatrixOutputs_lo_71};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_21 = {normSigOut_andMatrixOutputs_andMatrixInput_3_72, normSigOut_andMatrixOutputs_andMatrixInput_4_62};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_72 = {normSigOut_andMatrixOutputs_lo_hi_21, normSigOut_andMatrixOutputs_andMatrixInput_5_21};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_62 = {normSigOut_andMatrixOutputs_andMatrixInput_0_74, normSigOut_andMatrixOutputs_andMatrixInput_1_74};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_74 = {normSigOut_andMatrixOutputs_hi_hi_62, normSigOut_andMatrixOutputs_andMatrixInput_2_74};
  wire         normSigOut_andMatrixOutputs_49_2 = &{normSigOut_andMatrixOutputs_hi_74, normSigOut_andMatrixOutputs_lo_72};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_73 = {normSigOut_andMatrixOutputs_andMatrixInput_3_73, normSigOut_andMatrixOutputs_andMatrixInput_4_63};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_63 = {normSigOut_andMatrixOutputs_andMatrixInput_0_75, normSigOut_andMatrixOutputs_andMatrixInput_1_75};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_75 = {normSigOut_andMatrixOutputs_hi_hi_63, normSigOut_andMatrixOutputs_andMatrixInput_2_75};
  wire         normSigOut_andMatrixOutputs_42_2 = &{normSigOut_andMatrixOutputs_hi_75, normSigOut_andMatrixOutputs_lo_73};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_74 = {normSigOut_andMatrixOutputs_andMatrixInput_3_74, normSigOut_andMatrixOutputs_andMatrixInput_4_64};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_64 = {normSigOut_andMatrixOutputs_andMatrixInput_0_76, normSigOut_andMatrixOutputs_andMatrixInput_1_76};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_76 = {normSigOut_andMatrixOutputs_hi_hi_64, normSigOut_andMatrixOutputs_andMatrixInput_2_76};
  wire         normSigOut_andMatrixOutputs_55_2 = &{normSigOut_andMatrixOutputs_hi_76, normSigOut_andMatrixOutputs_lo_74};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_75 = {normSigOut_andMatrixOutputs_andMatrixInput_2_77, normSigOut_andMatrixOutputs_andMatrixInput_3_75};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_77 = {normSigOut_andMatrixOutputs_andMatrixInput_0_77, normSigOut_andMatrixOutputs_andMatrixInput_1_77};
  wire         normSigOut_andMatrixOutputs_69_2 = &{normSigOut_andMatrixOutputs_hi_77, normSigOut_andMatrixOutputs_lo_75};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_22 = {normSigOut_andMatrixOutputs_andMatrixInput_3_76, normSigOut_andMatrixOutputs_andMatrixInput_4_65};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_76 = {normSigOut_andMatrixOutputs_lo_hi_22, normSigOut_andMatrixOutputs_andMatrixInput_5_22};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_65 = {normSigOut_andMatrixOutputs_andMatrixInput_0_78, normSigOut_andMatrixOutputs_andMatrixInput_1_78};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_78 = {normSigOut_andMatrixOutputs_hi_hi_65, normSigOut_andMatrixOutputs_andMatrixInput_2_78};
  wire         normSigOut_andMatrixOutputs_68_2 = &{normSigOut_andMatrixOutputs_hi_78, normSigOut_andMatrixOutputs_lo_76};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_23 = {normSigOut_andMatrixOutputs_andMatrixInput_3_77, normSigOut_andMatrixOutputs_andMatrixInput_4_66};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_77 = {normSigOut_andMatrixOutputs_lo_hi_23, normSigOut_andMatrixOutputs_andMatrixInput_5_23};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_66 = {normSigOut_andMatrixOutputs_andMatrixInput_0_79, normSigOut_andMatrixOutputs_andMatrixInput_1_79};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_79 = {normSigOut_andMatrixOutputs_hi_hi_66, normSigOut_andMatrixOutputs_andMatrixInput_2_79};
  wire         normSigOut_andMatrixOutputs_19_2 = &{normSigOut_andMatrixOutputs_hi_79, normSigOut_andMatrixOutputs_lo_77};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_24 = {normSigOut_andMatrixOutputs_andMatrixInput_3_78, normSigOut_andMatrixOutputs_andMatrixInput_4_67};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_78 = {normSigOut_andMatrixOutputs_lo_hi_24, normSigOut_andMatrixOutputs_andMatrixInput_5_24};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_67 = {normSigOut_andMatrixOutputs_andMatrixInput_0_80, normSigOut_andMatrixOutputs_andMatrixInput_1_80};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_80 = {normSigOut_andMatrixOutputs_hi_hi_67, normSigOut_andMatrixOutputs_andMatrixInput_2_80};
  wire         normSigOut_andMatrixOutputs_5_2 = &{normSigOut_andMatrixOutputs_hi_80, normSigOut_andMatrixOutputs_lo_78};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_79 = {normSigOut_andMatrixOutputs_andMatrixInput_3_79, normSigOut_andMatrixOutputs_andMatrixInput_4_68};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_68 = {normSigOut_andMatrixOutputs_andMatrixInput_0_81, normSigOut_andMatrixOutputs_andMatrixInput_1_81};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_81 = {normSigOut_andMatrixOutputs_hi_hi_68, normSigOut_andMatrixOutputs_andMatrixInput_2_81};
  wire         normSigOut_andMatrixOutputs_21_2 = &{normSigOut_andMatrixOutputs_hi_81, normSigOut_andMatrixOutputs_lo_79};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_25 = {normSigOut_andMatrixOutputs_andMatrixInput_3_80, normSigOut_andMatrixOutputs_andMatrixInput_4_69};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_80 = {normSigOut_andMatrixOutputs_lo_hi_25, normSigOut_andMatrixOutputs_andMatrixInput_5_25};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_69 = {normSigOut_andMatrixOutputs_andMatrixInput_0_82, normSigOut_andMatrixOutputs_andMatrixInput_1_82};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_82 = {normSigOut_andMatrixOutputs_hi_hi_69, normSigOut_andMatrixOutputs_andMatrixInput_2_82};
  wire         normSigOut_andMatrixOutputs_53_2 = &{normSigOut_andMatrixOutputs_hi_82, normSigOut_andMatrixOutputs_lo_80};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_81 = {normSigOut_andMatrixOutputs_andMatrixInput_3_81, normSigOut_andMatrixOutputs_andMatrixInput_4_70};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_70 = {normSigOut_andMatrixOutputs_andMatrixInput_0_83, normSigOut_andMatrixOutputs_andMatrixInput_1_83};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_83 = {normSigOut_andMatrixOutputs_hi_hi_70, normSigOut_andMatrixOutputs_andMatrixInput_2_83};
  wire         normSigOut_andMatrixOutputs_36_2 = &{normSigOut_andMatrixOutputs_hi_83, normSigOut_andMatrixOutputs_lo_81};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_26 = {normSigOut_andMatrixOutputs_andMatrixInput_3_82, normSigOut_andMatrixOutputs_andMatrixInput_4_71};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_82 = {normSigOut_andMatrixOutputs_lo_hi_26, normSigOut_andMatrixOutputs_andMatrixInput_5_26};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_71 = {normSigOut_andMatrixOutputs_andMatrixInput_0_84, normSigOut_andMatrixOutputs_andMatrixInput_1_84};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_84 = {normSigOut_andMatrixOutputs_hi_hi_71, normSigOut_andMatrixOutputs_andMatrixInput_2_84};
  wire         normSigOut_andMatrixOutputs_15_2 = &{normSigOut_andMatrixOutputs_hi_84, normSigOut_andMatrixOutputs_lo_82};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_83 = {normSigOut_andMatrixOutputs_andMatrixInput_3_83, normSigOut_andMatrixOutputs_andMatrixInput_4_72};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_72 = {normSigOut_andMatrixOutputs_andMatrixInput_0_85, normSigOut_andMatrixOutputs_andMatrixInput_1_85};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_85 = {normSigOut_andMatrixOutputs_hi_hi_72, normSigOut_andMatrixOutputs_andMatrixInput_2_85};
  wire         normSigOut_andMatrixOutputs_73_2 = &{normSigOut_andMatrixOutputs_hi_85, normSigOut_andMatrixOutputs_lo_83};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_27 = {normSigOut_andMatrixOutputs_andMatrixInput_3_84, normSigOut_andMatrixOutputs_andMatrixInput_4_73};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_84 = {normSigOut_andMatrixOutputs_lo_hi_27, normSigOut_andMatrixOutputs_andMatrixInput_5_27};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_73 = {normSigOut_andMatrixOutputs_andMatrixInput_0_86, normSigOut_andMatrixOutputs_andMatrixInput_1_86};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_86 = {normSigOut_andMatrixOutputs_hi_hi_73, normSigOut_andMatrixOutputs_andMatrixInput_2_86};
  wire         normSigOut_andMatrixOutputs_89_2 = &{normSigOut_andMatrixOutputs_hi_86, normSigOut_andMatrixOutputs_lo_84};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_28 = {normSigOut_andMatrixOutputs_andMatrixInput_3_85, normSigOut_andMatrixOutputs_andMatrixInput_4_74};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_85 = {normSigOut_andMatrixOutputs_lo_hi_28, normSigOut_andMatrixOutputs_andMatrixInput_5_28};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_74 = {normSigOut_andMatrixOutputs_andMatrixInput_0_87, normSigOut_andMatrixOutputs_andMatrixInput_1_87};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_87 = {normSigOut_andMatrixOutputs_hi_hi_74, normSigOut_andMatrixOutputs_andMatrixInput_2_87};
  wire         normSigOut_andMatrixOutputs_72_2 = &{normSigOut_andMatrixOutputs_hi_87, normSigOut_andMatrixOutputs_lo_85};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_29 = {normSigOut_andMatrixOutputs_andMatrixInput_3_86, normSigOut_andMatrixOutputs_andMatrixInput_4_75};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_86 = {normSigOut_andMatrixOutputs_lo_hi_29, normSigOut_andMatrixOutputs_andMatrixInput_5_29};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_75 = {normSigOut_andMatrixOutputs_andMatrixInput_0_88, normSigOut_andMatrixOutputs_andMatrixInput_1_88};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_88 = {normSigOut_andMatrixOutputs_hi_hi_75, normSigOut_andMatrixOutputs_andMatrixInput_2_88};
  wire         normSigOut_andMatrixOutputs_84_2 = &{normSigOut_andMatrixOutputs_hi_88, normSigOut_andMatrixOutputs_lo_86};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_30 = {normSigOut_andMatrixOutputs_andMatrixInput_3_87, normSigOut_andMatrixOutputs_andMatrixInput_4_76};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_87 = {normSigOut_andMatrixOutputs_lo_hi_30, normSigOut_andMatrixOutputs_andMatrixInput_5_30};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_76 = {normSigOut_andMatrixOutputs_andMatrixInput_0_89, normSigOut_andMatrixOutputs_andMatrixInput_1_89};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_89 = {normSigOut_andMatrixOutputs_hi_hi_76, normSigOut_andMatrixOutputs_andMatrixInput_2_89};
  wire         normSigOut_andMatrixOutputs_76_2 = &{normSigOut_andMatrixOutputs_hi_89, normSigOut_andMatrixOutputs_lo_87};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_hi_31 = {normSigOut_andMatrixOutputs_andMatrixInput_3_88, normSigOut_andMatrixOutputs_andMatrixInput_4_77};
  wire [2:0]   normSigOut_andMatrixOutputs_lo_88 = {normSigOut_andMatrixOutputs_lo_hi_31, normSigOut_andMatrixOutputs_andMatrixInput_5_31};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_77 = {normSigOut_andMatrixOutputs_andMatrixInput_0_90, normSigOut_andMatrixOutputs_andMatrixInput_1_90};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_90 = {normSigOut_andMatrixOutputs_hi_hi_77, normSigOut_andMatrixOutputs_andMatrixInput_2_90};
  wire         normSigOut_andMatrixOutputs_28_2 = &{normSigOut_andMatrixOutputs_hi_90, normSigOut_andMatrixOutputs_lo_88};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_89 = {normSigOut_andMatrixOutputs_andMatrixInput_3_89, normSigOut_andMatrixOutputs_andMatrixInput_4_78};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_78 = {normSigOut_andMatrixOutputs_andMatrixInput_0_91, normSigOut_andMatrixOutputs_andMatrixInput_1_91};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_91 = {normSigOut_andMatrixOutputs_hi_hi_78, normSigOut_andMatrixOutputs_andMatrixInput_2_91};
  wire         normSigOut_andMatrixOutputs_33_2 = &{normSigOut_andMatrixOutputs_hi_91, normSigOut_andMatrixOutputs_lo_89};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_90 = {normSigOut_andMatrixOutputs_andMatrixInput_3_90, normSigOut_andMatrixOutputs_andMatrixInput_4_79};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_79 = {normSigOut_andMatrixOutputs_andMatrixInput_0_92, normSigOut_andMatrixOutputs_andMatrixInput_1_92};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_92 = {normSigOut_andMatrixOutputs_hi_hi_79, normSigOut_andMatrixOutputs_andMatrixInput_2_92};
  wire         normSigOut_andMatrixOutputs_0_2 = &{normSigOut_andMatrixOutputs_hi_92, normSigOut_andMatrixOutputs_lo_90};
  wire [1:0]   normSigOut_andMatrixOutputs_lo_91 = {normSigOut_andMatrixOutputs_andMatrixInput_3_91, normSigOut_andMatrixOutputs_andMatrixInput_4_80};
  wire [1:0]   normSigOut_andMatrixOutputs_hi_hi_80 = {normSigOut_andMatrixOutputs_andMatrixInput_0_93, normSigOut_andMatrixOutputs_andMatrixInput_1_93};
  wire [2:0]   normSigOut_andMatrixOutputs_hi_93 = {normSigOut_andMatrixOutputs_hi_hi_80, normSigOut_andMatrixOutputs_andMatrixInput_2_93};
  wire         normSigOut_andMatrixOutputs_24_2 = &{normSigOut_andMatrixOutputs_hi_93, normSigOut_andMatrixOutputs_lo_91};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_lo_lo_hi = {normSigOut_andMatrixOutputs_72_2, normSigOut_andMatrixOutputs_28_2};
  wire [2:0]   normSigOut_orMatrixOutputs_lo_lo_lo = {normSigOut_orMatrixOutputs_lo_lo_lo_hi, normSigOut_andMatrixOutputs_33_2};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_lo_hi_lo = {normSigOut_andMatrixOutputs_15_2, normSigOut_andMatrixOutputs_89_2};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_lo_hi_hi = {normSigOut_andMatrixOutputs_5_2, normSigOut_andMatrixOutputs_53_2};
  wire [3:0]   normSigOut_orMatrixOutputs_lo_lo_hi = {normSigOut_orMatrixOutputs_lo_lo_hi_hi, normSigOut_orMatrixOutputs_lo_lo_hi_lo};
  wire [6:0]   normSigOut_orMatrixOutputs_lo_lo = {normSigOut_orMatrixOutputs_lo_lo_hi, normSigOut_orMatrixOutputs_lo_lo_lo};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_hi_lo_lo = {normSigOut_andMatrixOutputs_38_2, normSigOut_andMatrixOutputs_68_2};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_hi_lo_hi = {normSigOut_andMatrixOutputs_20_2, normSigOut_andMatrixOutputs_54_2};
  wire [3:0]   normSigOut_orMatrixOutputs_lo_hi_lo = {normSigOut_orMatrixOutputs_lo_hi_lo_hi, normSigOut_orMatrixOutputs_lo_hi_lo_lo};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_hi_hi_lo = {normSigOut_andMatrixOutputs_91_2, normSigOut_andMatrixOutputs_58_2};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_hi_hi_hi = {normSigOut_andMatrixOutputs_50_2, normSigOut_andMatrixOutputs_22_2};
  wire [3:0]   normSigOut_orMatrixOutputs_lo_hi_hi = {normSigOut_orMatrixOutputs_lo_hi_hi_hi, normSigOut_orMatrixOutputs_lo_hi_hi_lo};
  wire [7:0]   normSigOut_orMatrixOutputs_lo_hi = {normSigOut_orMatrixOutputs_lo_hi_hi, normSigOut_orMatrixOutputs_lo_hi_lo};
  wire [14:0]  normSigOut_orMatrixOutputs_lo = {normSigOut_orMatrixOutputs_lo_hi, normSigOut_orMatrixOutputs_lo_lo};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_lo_lo_lo = {normSigOut_andMatrixOutputs_4_2, normSigOut_andMatrixOutputs_57_2};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_lo_lo_hi = {normSigOut_andMatrixOutputs_48_2, normSigOut_andMatrixOutputs_60_2};
  wire [3:0]   normSigOut_orMatrixOutputs_hi_lo_lo = {normSigOut_orMatrixOutputs_hi_lo_lo_hi, normSigOut_orMatrixOutputs_hi_lo_lo_lo};
  wire [1:0]   _GEN = {normSigOut_andMatrixOutputs_3_2, normSigOut_andMatrixOutputs_8_2};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_lo_hi_lo;
  assign normSigOut_orMatrixOutputs_hi_lo_hi_lo = _GEN;
  wire [1:0]   normSigOut_orMatrixOutputs_lo_lo_hi_6;
  assign normSigOut_orMatrixOutputs_lo_lo_hi_6 = _GEN;
  wire [1:0]   normSigOut_orMatrixOutputs_hi_lo_hi_hi = {normSigOut_andMatrixOutputs_88_2, normSigOut_andMatrixOutputs_75_2};
  wire [3:0]   normSigOut_orMatrixOutputs_hi_lo_hi = {normSigOut_orMatrixOutputs_hi_lo_hi_hi, normSigOut_orMatrixOutputs_hi_lo_hi_lo};
  wire [7:0]   normSigOut_orMatrixOutputs_hi_lo = {normSigOut_orMatrixOutputs_hi_lo_hi, normSigOut_orMatrixOutputs_hi_lo_lo};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_hi_lo_lo = {normSigOut_andMatrixOutputs_45_2, normSigOut_andMatrixOutputs_80_2};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_hi_lo_hi = {normSigOut_andMatrixOutputs_90_2, normSigOut_andMatrixOutputs_71_2};
  wire [3:0]   normSigOut_orMatrixOutputs_hi_hi_lo = {normSigOut_orMatrixOutputs_hi_hi_lo_hi, normSigOut_orMatrixOutputs_hi_hi_lo_lo};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_hi_hi_lo = {normSigOut_andMatrixOutputs_52_2, normSigOut_andMatrixOutputs_64_2};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_hi_hi_hi = {normSigOut_andMatrixOutputs_47_2, normSigOut_andMatrixOutputs_7_2};
  wire [3:0]   normSigOut_orMatrixOutputs_hi_hi_hi = {normSigOut_orMatrixOutputs_hi_hi_hi_hi, normSigOut_orMatrixOutputs_hi_hi_hi_lo};
  wire [7:0]   normSigOut_orMatrixOutputs_hi_hi = {normSigOut_orMatrixOutputs_hi_hi_hi, normSigOut_orMatrixOutputs_hi_hi_lo};
  wire [15:0]  normSigOut_orMatrixOutputs_hi = {normSigOut_orMatrixOutputs_hi_hi, normSigOut_orMatrixOutputs_hi_lo};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_lo_lo_hi_1 = {normSigOut_andMatrixOutputs_53_2, normSigOut_andMatrixOutputs_73_2};
  wire [2:0]   normSigOut_orMatrixOutputs_lo_lo_lo_1 = {normSigOut_orMatrixOutputs_lo_lo_lo_hi_1, normSigOut_andMatrixOutputs_0_2};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_lo_hi_hi_1 = {normSigOut_andMatrixOutputs_44_2, normSigOut_andMatrixOutputs_26_2};
  wire [2:0]   normSigOut_orMatrixOutputs_lo_lo_hi_1 = {normSigOut_orMatrixOutputs_lo_lo_hi_hi_1, normSigOut_andMatrixOutputs_68_2};
  wire [5:0]   normSigOut_orMatrixOutputs_lo_lo_1 = {normSigOut_orMatrixOutputs_lo_lo_hi_1, normSigOut_orMatrixOutputs_lo_lo_lo_1};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_hi_lo_hi_1 = {normSigOut_andMatrixOutputs_40_2, normSigOut_andMatrixOutputs_29_2};
  wire [2:0]   normSigOut_orMatrixOutputs_lo_hi_lo_1 = {normSigOut_orMatrixOutputs_lo_hi_lo_hi_1, normSigOut_andMatrixOutputs_20_2};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_hi_hi_lo_1 = {normSigOut_andMatrixOutputs_32_2, normSigOut_andMatrixOutputs_25_2};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_hi_hi_hi_1 = {normSigOut_andMatrixOutputs_4_2, normSigOut_andMatrixOutputs_22_2};
  wire [3:0]   normSigOut_orMatrixOutputs_lo_hi_hi_1 = {normSigOut_orMatrixOutputs_lo_hi_hi_hi_1, normSigOut_orMatrixOutputs_lo_hi_hi_lo_1};
  wire [6:0]   normSigOut_orMatrixOutputs_lo_hi_1 = {normSigOut_orMatrixOutputs_lo_hi_hi_1, normSigOut_orMatrixOutputs_lo_hi_lo_1};
  wire [12:0]  normSigOut_orMatrixOutputs_lo_1 = {normSigOut_orMatrixOutputs_lo_hi_1, normSigOut_orMatrixOutputs_lo_lo_1};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_lo_lo_hi_1 = {normSigOut_andMatrixOutputs_79_2, normSigOut_andMatrixOutputs_74_2};
  wire [2:0]   normSigOut_orMatrixOutputs_hi_lo_lo_1 = {normSigOut_orMatrixOutputs_hi_lo_lo_hi_1, normSigOut_andMatrixOutputs_60_2};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_lo_hi_lo_1 = {normSigOut_andMatrixOutputs_23_2, normSigOut_andMatrixOutputs_10_2};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_lo_hi_hi_1 = {normSigOut_andMatrixOutputs_6_2, normSigOut_andMatrixOutputs_70_2};
  wire [3:0]   normSigOut_orMatrixOutputs_hi_lo_hi_1 = {normSigOut_orMatrixOutputs_hi_lo_hi_hi_1, normSigOut_orMatrixOutputs_hi_lo_hi_lo_1};
  wire [6:0]   normSigOut_orMatrixOutputs_hi_lo_1 = {normSigOut_orMatrixOutputs_hi_lo_hi_1, normSigOut_orMatrixOutputs_hi_lo_lo_1};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_hi_lo_hi_1 = {normSigOut_andMatrixOutputs_87_2, normSigOut_andMatrixOutputs_85_2};
  wire [2:0]   normSigOut_orMatrixOutputs_hi_hi_lo_1 = {normSigOut_orMatrixOutputs_hi_hi_lo_hi_1, normSigOut_andMatrixOutputs_59_2};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_hi_hi_lo_1 = {normSigOut_andMatrixOutputs_92_2, normSigOut_andMatrixOutputs_86_2};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_hi_hi_hi_1 = {normSigOut_andMatrixOutputs_61_2, normSigOut_andMatrixOutputs_67_2};
  wire [3:0]   normSigOut_orMatrixOutputs_hi_hi_hi_1 = {normSigOut_orMatrixOutputs_hi_hi_hi_hi_1, normSigOut_orMatrixOutputs_hi_hi_hi_lo_1};
  wire [6:0]   normSigOut_orMatrixOutputs_hi_hi_1 = {normSigOut_orMatrixOutputs_hi_hi_hi_1, normSigOut_orMatrixOutputs_hi_hi_lo_1};
  wire [13:0]  normSigOut_orMatrixOutputs_hi_1 = {normSigOut_orMatrixOutputs_hi_hi_1, normSigOut_orMatrixOutputs_hi_lo_1};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_lo_lo_hi_2 = {normSigOut_andMatrixOutputs_84_2, normSigOut_andMatrixOutputs_76_2};
  wire [2:0]   normSigOut_orMatrixOutputs_lo_lo_lo_2 = {normSigOut_orMatrixOutputs_lo_lo_lo_hi_2, normSigOut_andMatrixOutputs_24_2};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_lo_hi_lo_1 = {normSigOut_andMatrixOutputs_21_2, normSigOut_andMatrixOutputs_73_2};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_lo_hi_hi_2 = {normSigOut_andMatrixOutputs_19_2, normSigOut_andMatrixOutputs_5_2};
  wire [3:0]   normSigOut_orMatrixOutputs_lo_lo_hi_2 = {normSigOut_orMatrixOutputs_lo_lo_hi_hi_2, normSigOut_orMatrixOutputs_lo_lo_hi_lo_1};
  wire [6:0]   normSigOut_orMatrixOutputs_lo_lo_2 = {normSigOut_orMatrixOutputs_lo_lo_hi_2, normSigOut_orMatrixOutputs_lo_lo_lo_2};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_hi_lo_hi_2 = {normSigOut_andMatrixOutputs_49_2, normSigOut_andMatrixOutputs_42_2};
  wire [2:0]   normSigOut_orMatrixOutputs_lo_hi_lo_2 = {normSigOut_orMatrixOutputs_lo_hi_lo_hi_2, normSigOut_andMatrixOutputs_55_2};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_hi_hi_lo_2 = {normSigOut_andMatrixOutputs_31_2, normSigOut_andMatrixOutputs_46_2};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_hi_hi_hi_2 = {normSigOut_andMatrixOutputs_57_2, normSigOut_andMatrixOutputs_77_2};
  wire [3:0]   normSigOut_orMatrixOutputs_lo_hi_hi_2 = {normSigOut_orMatrixOutputs_lo_hi_hi_hi_2, normSigOut_orMatrixOutputs_lo_hi_hi_lo_2};
  wire [6:0]   normSigOut_orMatrixOutputs_lo_hi_2 = {normSigOut_orMatrixOutputs_lo_hi_hi_2, normSigOut_orMatrixOutputs_lo_hi_lo_2};
  wire [13:0]  normSigOut_orMatrixOutputs_lo_2 = {normSigOut_orMatrixOutputs_lo_hi_2, normSigOut_orMatrixOutputs_lo_lo_2};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_lo_lo_hi_2 = {normSigOut_andMatrixOutputs_43_2, normSigOut_andMatrixOutputs_30_2};
  wire [2:0]   normSigOut_orMatrixOutputs_hi_lo_lo_2 = {normSigOut_orMatrixOutputs_hi_lo_lo_hi_2, normSigOut_andMatrixOutputs_66_2};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_lo_hi_lo_2 = {normSigOut_andMatrixOutputs_2_2, normSigOut_andMatrixOutputs_17_2};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_lo_hi_hi_2 = {normSigOut_andMatrixOutputs_6_2, normSigOut_andMatrixOutputs_88_2};
  wire [3:0]   normSigOut_orMatrixOutputs_hi_lo_hi_2 = {normSigOut_orMatrixOutputs_hi_lo_hi_hi_2, normSigOut_orMatrixOutputs_hi_lo_hi_lo_2};
  wire [6:0]   normSigOut_orMatrixOutputs_hi_lo_2 = {normSigOut_orMatrixOutputs_hi_lo_hi_2, normSigOut_orMatrixOutputs_hi_lo_lo_2};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_hi_lo_hi_2 = {normSigOut_andMatrixOutputs_86_2, normSigOut_andMatrixOutputs_81_2};
  wire [2:0]   normSigOut_orMatrixOutputs_hi_hi_lo_2 = {normSigOut_orMatrixOutputs_hi_hi_lo_hi_2, normSigOut_andMatrixOutputs_12_2};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_hi_hi_lo_2 = {normSigOut_andMatrixOutputs_51_2, normSigOut_andMatrixOutputs_63_2};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_hi_hi_hi_2 = {normSigOut_andMatrixOutputs_65_2, normSigOut_andMatrixOutputs_7_2};
  wire [3:0]   normSigOut_orMatrixOutputs_hi_hi_hi_2 = {normSigOut_orMatrixOutputs_hi_hi_hi_hi_2, normSigOut_orMatrixOutputs_hi_hi_hi_lo_2};
  wire [6:0]   normSigOut_orMatrixOutputs_hi_hi_2 = {normSigOut_orMatrixOutputs_hi_hi_hi_2, normSigOut_orMatrixOutputs_hi_hi_lo_2};
  wire [13:0]  normSigOut_orMatrixOutputs_hi_2 = {normSigOut_orMatrixOutputs_hi_hi_2, normSigOut_orMatrixOutputs_hi_lo_2};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_lo_lo_3 = {normSigOut_andMatrixOutputs_76_2, normSigOut_andMatrixOutputs_28_2};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_lo_hi_hi_3 = {normSigOut_andMatrixOutputs_73_2, normSigOut_andMatrixOutputs_72_2};
  wire [2:0]   normSigOut_orMatrixOutputs_lo_lo_hi_3 = {normSigOut_orMatrixOutputs_lo_lo_hi_hi_3, normSigOut_andMatrixOutputs_84_2};
  wire [4:0]   normSigOut_orMatrixOutputs_lo_lo_3 = {normSigOut_orMatrixOutputs_lo_lo_hi_3, normSigOut_orMatrixOutputs_lo_lo_lo_3};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_hi_lo_hi_3 = {normSigOut_andMatrixOutputs_44_2, normSigOut_andMatrixOutputs_49_2};
  wire [2:0]   normSigOut_orMatrixOutputs_lo_hi_lo_3 = {normSigOut_orMatrixOutputs_lo_hi_lo_hi_3, normSigOut_andMatrixOutputs_69_2};
  wire [1:0]   _GEN_0 = {normSigOut_andMatrixOutputs_66_2, normSigOut_andMatrixOutputs_57_2};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_hi_hi_hi_3;
  assign normSigOut_orMatrixOutputs_lo_hi_hi_hi_3 = _GEN_0;
  wire [1:0]   normSigOut_orMatrixOutputs_lo_hi_hi_5;
  assign normSigOut_orMatrixOutputs_lo_hi_hi_5 = _GEN_0;
  wire [2:0]   normSigOut_orMatrixOutputs_lo_hi_hi_3 = {normSigOut_orMatrixOutputs_lo_hi_hi_hi_3, normSigOut_andMatrixOutputs_18_2};
  wire [5:0]   normSigOut_orMatrixOutputs_lo_hi_3 = {normSigOut_orMatrixOutputs_lo_hi_hi_3, normSigOut_orMatrixOutputs_lo_hi_lo_3};
  wire [10:0]  normSigOut_orMatrixOutputs_lo_3 = {normSigOut_orMatrixOutputs_lo_hi_3, normSigOut_orMatrixOutputs_lo_lo_3};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_lo_lo_3 = {normSigOut_andMatrixOutputs_60_2, normSigOut_andMatrixOutputs_4_2};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_lo_hi_hi_3 = {normSigOut_andMatrixOutputs_1_2, normSigOut_andMatrixOutputs_3_2};
  wire [2:0]   normSigOut_orMatrixOutputs_hi_lo_hi_3 = {normSigOut_orMatrixOutputs_hi_lo_hi_hi_3, normSigOut_andMatrixOutputs_93_2};
  wire [4:0]   normSigOut_orMatrixOutputs_hi_lo_3 = {normSigOut_orMatrixOutputs_hi_lo_hi_3, normSigOut_orMatrixOutputs_hi_lo_lo_3};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_hi_lo_hi_3 = {normSigOut_andMatrixOutputs_86_2, normSigOut_andMatrixOutputs_27_2};
  wire [2:0]   normSigOut_orMatrixOutputs_hi_hi_lo_3 = {normSigOut_orMatrixOutputs_hi_hi_lo_hi_3, normSigOut_andMatrixOutputs_6_2};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_hi_hi_hi_3 = {normSigOut_andMatrixOutputs_41_2, normSigOut_andMatrixOutputs_83_2};
  wire [2:0]   normSigOut_orMatrixOutputs_hi_hi_hi_3 = {normSigOut_orMatrixOutputs_hi_hi_hi_hi_3, normSigOut_andMatrixOutputs_64_2};
  wire [5:0]   normSigOut_orMatrixOutputs_hi_hi_3 = {normSigOut_orMatrixOutputs_hi_hi_hi_3, normSigOut_orMatrixOutputs_hi_hi_lo_3};
  wire [10:0]  normSigOut_orMatrixOutputs_hi_3 = {normSigOut_orMatrixOutputs_hi_hi_3, normSigOut_orMatrixOutputs_hi_lo_3};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_lo_lo_4 = {normSigOut_andMatrixOutputs_21_2, normSigOut_andMatrixOutputs_36_2};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_lo_hi_4 = {normSigOut_andMatrixOutputs_69_2, normSigOut_andMatrixOutputs_5_2};
  wire [3:0]   normSigOut_orMatrixOutputs_lo_lo_4 = {normSigOut_orMatrixOutputs_lo_lo_hi_4, normSigOut_orMatrixOutputs_lo_lo_lo_4};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_hi_lo_4 = {normSigOut_andMatrixOutputs_46_2, normSigOut_andMatrixOutputs_26_2};
  wire [1:0]   _GEN_1 = {normSigOut_andMatrixOutputs_82_2, normSigOut_andMatrixOutputs_50_2};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_hi_hi_4;
  assign normSigOut_orMatrixOutputs_lo_hi_hi_4 = _GEN_1;
  wire [1:0]   normSigOut_orMatrixOutputs_lo_lo_hi_5;
  assign normSigOut_orMatrixOutputs_lo_lo_hi_5 = _GEN_1;
  wire [3:0]   normSigOut_orMatrixOutputs_lo_hi_4 = {normSigOut_orMatrixOutputs_lo_hi_hi_4, normSigOut_orMatrixOutputs_lo_hi_lo_4};
  wire [7:0]   normSigOut_orMatrixOutputs_lo_4 = {normSigOut_orMatrixOutputs_lo_hi_4, normSigOut_orMatrixOutputs_lo_lo_4};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_lo_lo_4 = {normSigOut_andMatrixOutputs_9_2, normSigOut_andMatrixOutputs_16_2};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_lo_hi_4 = {normSigOut_andMatrixOutputs_34_2, normSigOut_andMatrixOutputs_56_2};
  wire [3:0]   normSigOut_orMatrixOutputs_hi_lo_4 = {normSigOut_orMatrixOutputs_hi_lo_hi_4, normSigOut_orMatrixOutputs_hi_lo_lo_4};
  wire [1:0]   _GEN_2 = {normSigOut_andMatrixOutputs_14_2, normSigOut_andMatrixOutputs_1_2};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_hi_lo_4;
  assign normSigOut_orMatrixOutputs_hi_hi_lo_4 = _GEN_2;
  wire [1:0]   normSigOut_orMatrixOutputs_lo_hi_hi_6;
  assign normSigOut_orMatrixOutputs_lo_hi_hi_6 = _GEN_2;
  wire [1:0]   normSigOut_orMatrixOutputs_hi_hi_hi_hi_4 = {normSigOut_andMatrixOutputs_11_2, normSigOut_andMatrixOutputs_78_2};
  wire [2:0]   normSigOut_orMatrixOutputs_hi_hi_hi_4 = {normSigOut_orMatrixOutputs_hi_hi_hi_hi_4, normSigOut_andMatrixOutputs_6_2};
  wire [4:0]   normSigOut_orMatrixOutputs_hi_hi_4 = {normSigOut_orMatrixOutputs_hi_hi_hi_4, normSigOut_orMatrixOutputs_hi_hi_lo_4};
  wire [8:0]   normSigOut_orMatrixOutputs_hi_4 = {normSigOut_orMatrixOutputs_hi_hi_4, normSigOut_orMatrixOutputs_hi_lo_4};
  wire [2:0]   normSigOut_orMatrixOutputs_lo_lo_5 = {normSigOut_orMatrixOutputs_lo_lo_hi_5, normSigOut_andMatrixOutputs_31_2};
  wire [2:0]   normSigOut_orMatrixOutputs_lo_hi_5 = {normSigOut_orMatrixOutputs_lo_hi_hi_5, normSigOut_andMatrixOutputs_16_2};
  wire [5:0]   normSigOut_orMatrixOutputs_lo_5 = {normSigOut_orMatrixOutputs_lo_hi_5, normSigOut_orMatrixOutputs_lo_lo_5};
  wire [1:0]   _GEN_3 = {normSigOut_andMatrixOutputs_47_2, normSigOut_andMatrixOutputs_39_2};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_lo_hi_5;
  assign normSigOut_orMatrixOutputs_hi_lo_hi_5 = _GEN_3;
  wire [1:0]   normSigOut_orMatrixOutputs_hi_lo_hi_6;
  assign normSigOut_orMatrixOutputs_hi_lo_hi_6 = _GEN_3;
  wire [2:0]   normSigOut_orMatrixOutputs_hi_lo_5 = {normSigOut_orMatrixOutputs_hi_lo_hi_5, normSigOut_andMatrixOutputs_4_2};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_hi_hi_5 = {normSigOut_andMatrixOutputs_37_2, normSigOut_andMatrixOutputs_62_2};
  wire [2:0]   normSigOut_orMatrixOutputs_hi_hi_5 = {normSigOut_orMatrixOutputs_hi_hi_hi_5, normSigOut_andMatrixOutputs_35_2};
  wire [5:0]   normSigOut_orMatrixOutputs_hi_5 = {normSigOut_orMatrixOutputs_hi_hi_5, normSigOut_orMatrixOutputs_hi_lo_5};
  wire [2:0]   normSigOut_orMatrixOutputs_lo_lo_6 = {normSigOut_orMatrixOutputs_lo_lo_hi_6, normSigOut_andMatrixOutputs_43_2};
  wire [2:0]   normSigOut_orMatrixOutputs_lo_hi_6 = {normSigOut_orMatrixOutputs_lo_hi_hi_6, normSigOut_andMatrixOutputs_34_2};
  wire [5:0]   normSigOut_orMatrixOutputs_lo_6 = {normSigOut_orMatrixOutputs_lo_hi_6, normSigOut_orMatrixOutputs_lo_lo_6};
  wire [2:0]   normSigOut_orMatrixOutputs_hi_lo_6 = {normSigOut_orMatrixOutputs_hi_lo_hi_6, normSigOut_andMatrixOutputs_6_2};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_hi_hi_6 = {normSigOut_andMatrixOutputs_13_2, normSigOut_andMatrixOutputs_83_2};
  wire [2:0]   normSigOut_orMatrixOutputs_hi_hi_6 = {normSigOut_orMatrixOutputs_hi_hi_hi_6, normSigOut_andMatrixOutputs_35_2};
  wire [5:0]   normSigOut_orMatrixOutputs_hi_6 = {normSigOut_orMatrixOutputs_hi_hi_6, normSigOut_orMatrixOutputs_hi_lo_6};
  wire [1:0]   normSigOut_orMatrixOutputs_lo_hi_7 = {|{normSigOut_orMatrixOutputs_hi_2, normSigOut_orMatrixOutputs_lo_2}, |{normSigOut_orMatrixOutputs_hi_1, normSigOut_orMatrixOutputs_lo_1}};
  wire [2:0]   normSigOut_orMatrixOutputs_lo_7 = {normSigOut_orMatrixOutputs_lo_hi_7, |{normSigOut_orMatrixOutputs_hi, normSigOut_orMatrixOutputs_lo}};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_lo_7 = {|{normSigOut_orMatrixOutputs_hi_4, normSigOut_orMatrixOutputs_lo_4}, |{normSigOut_orMatrixOutputs_hi_3, normSigOut_orMatrixOutputs_lo_3}};
  wire [1:0]   normSigOut_orMatrixOutputs_hi_hi_7 = {|{normSigOut_orMatrixOutputs_hi_6, normSigOut_orMatrixOutputs_lo_6}, |{normSigOut_orMatrixOutputs_hi_5, normSigOut_orMatrixOutputs_lo_5}};
  wire [3:0]   normSigOut_orMatrixOutputs_hi_7 = {normSigOut_orMatrixOutputs_hi_hi_7, normSigOut_orMatrixOutputs_hi_lo_7};
  wire [6:0]   normSigOut_orMatrixOutputs = {normSigOut_orMatrixOutputs_hi_7, normSigOut_orMatrixOutputs_lo_7};
  wire [1:0]   normSigOut_invMatrixOutputs_lo_hi = normSigOut_orMatrixOutputs[2:1];
  wire [2:0]   normSigOut_invMatrixOutputs_lo = {normSigOut_invMatrixOutputs_lo_hi, normSigOut_orMatrixOutputs[0]};
  wire [1:0]   normSigOut_invMatrixOutputs_hi_lo = normSigOut_orMatrixOutputs[4:3];
  wire [1:0]   normSigOut_invMatrixOutputs_hi_hi = normSigOut_orMatrixOutputs[6:5];
  wire [3:0]   normSigOut_invMatrixOutputs_hi = {normSigOut_invMatrixOutputs_hi_hi, normSigOut_invMatrixOutputs_hi_lo};
  assign normSigOut_invMatrixOutputs = {normSigOut_invMatrixOutputs_hi, normSigOut_invMatrixOutputs_lo};
  wire [6:0]   normSigOut_plaOutput = normSigOut_invMatrixOutputs;
  wire [22:0]  normSigOut = {normSigOut_plaOutput, 16'h0};
  wire [7:0]   normExpOut = 8'hFD - normExpIn;
  wire         _outSubShift_T = normExpOut == 8'h0;
  wire         outIsSub = _outSubShift_T | (&normExpOut);
  wire [7:0]   expOut = outIsSub ? 8'h0 : normExpOut;
  wire [1:0]   outSubShift = _outSubShift_T ? 2'h1 : 2'h2;
  wire [23:0]  _sigOut_T_1 = {1'h1, normSigOut} >> outSubShift;
  wire [22:0]  sigOut = outIsSub ? _sigOut_T_1[22:0] : normSigOut;
  wire [8:0]   view__out_data_hi = {sign, expOut};
  assign out_data =
    inIsNegativeInf
      ? 32'h80000000
      : inIsPositiveInf
          ? 32'h0
          : inIsNegativeZero | roundAbnormalToNegaInf ? 32'hFF800000 : inIsPositveZero | roundAbnormalToPosInf ? 32'h7F800000 : inIsQNaN | inIsSNaN ? 32'h7FC00000 : roundAbnormalToMax ? {sign, 31'h7F7FFFFF} : {view__out_data_hi, sigOut};
  assign out_exceptionFlags = inIsSNaN ? 5'h10 : {1'h0, inIsPositveZero | inIsNegativeZero ? 4'h8 : {1'h0, roundAbnormal ? 3'h5 : 3'h0}};
endmodule

