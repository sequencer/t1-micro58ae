module VectorAdder64(
  input  [63:0] a,
                b,
  output [63:0] z,
  input  [3:0]  sew
);

  wire        as_0 = a[0];
  wire        as_1 = a[1];
  wire        as_2 = a[2];
  wire        as_3 = a[3];
  wire        as_4 = a[4];
  wire        as_5 = a[5];
  wire        as_6 = a[6];
  wire        as_7 = a[7];
  wire        as_8 = a[8];
  wire        as_9 = a[9];
  wire        as_10 = a[10];
  wire        as_11 = a[11];
  wire        as_12 = a[12];
  wire        as_13 = a[13];
  wire        as_14 = a[14];
  wire        as_15 = a[15];
  wire        as_16 = a[16];
  wire        as_17 = a[17];
  wire        as_18 = a[18];
  wire        as_19 = a[19];
  wire        as_20 = a[20];
  wire        as_21 = a[21];
  wire        as_22 = a[22];
  wire        as_23 = a[23];
  wire        as_24 = a[24];
  wire        as_25 = a[25];
  wire        as_26 = a[26];
  wire        as_27 = a[27];
  wire        as_28 = a[28];
  wire        as_29 = a[29];
  wire        as_30 = a[30];
  wire        as_31 = a[31];
  wire        as_32 = a[32];
  wire        as_33 = a[33];
  wire        as_34 = a[34];
  wire        as_35 = a[35];
  wire        as_36 = a[36];
  wire        as_37 = a[37];
  wire        as_38 = a[38];
  wire        as_39 = a[39];
  wire        as_40 = a[40];
  wire        as_41 = a[41];
  wire        as_42 = a[42];
  wire        as_43 = a[43];
  wire        as_44 = a[44];
  wire        as_45 = a[45];
  wire        as_46 = a[46];
  wire        as_47 = a[47];
  wire        as_48 = a[48];
  wire        as_49 = a[49];
  wire        as_50 = a[50];
  wire        as_51 = a[51];
  wire        as_52 = a[52];
  wire        as_53 = a[53];
  wire        as_54 = a[54];
  wire        as_55 = a[55];
  wire        as_56 = a[56];
  wire        as_57 = a[57];
  wire        as_58 = a[58];
  wire        as_59 = a[59];
  wire        as_60 = a[60];
  wire        as_61 = a[61];
  wire        as_62 = a[62];
  wire        as_63 = a[63];
  wire        bs_0 = b[0];
  wire        bs_1 = b[1];
  wire        bs_2 = b[2];
  wire        bs_3 = b[3];
  wire        bs_4 = b[4];
  wire        bs_5 = b[5];
  wire        bs_6 = b[6];
  wire        bs_7 = b[7];
  wire        bs_8 = b[8];
  wire        bs_9 = b[9];
  wire        bs_10 = b[10];
  wire        bs_11 = b[11];
  wire        bs_12 = b[12];
  wire        bs_13 = b[13];
  wire        bs_14 = b[14];
  wire        bs_15 = b[15];
  wire        bs_16 = b[16];
  wire        bs_17 = b[17];
  wire        bs_18 = b[18];
  wire        bs_19 = b[19];
  wire        bs_20 = b[20];
  wire        bs_21 = b[21];
  wire        bs_22 = b[22];
  wire        bs_23 = b[23];
  wire        bs_24 = b[24];
  wire        bs_25 = b[25];
  wire        bs_26 = b[26];
  wire        bs_27 = b[27];
  wire        bs_28 = b[28];
  wire        bs_29 = b[29];
  wire        bs_30 = b[30];
  wire        bs_31 = b[31];
  wire        bs_32 = b[32];
  wire        bs_33 = b[33];
  wire        bs_34 = b[34];
  wire        bs_35 = b[35];
  wire        bs_36 = b[36];
  wire        bs_37 = b[37];
  wire        bs_38 = b[38];
  wire        bs_39 = b[39];
  wire        bs_40 = b[40];
  wire        bs_41 = b[41];
  wire        bs_42 = b[42];
  wire        bs_43 = b[43];
  wire        bs_44 = b[44];
  wire        bs_45 = b[45];
  wire        bs_46 = b[46];
  wire        bs_47 = b[47];
  wire        bs_48 = b[48];
  wire        bs_49 = b[49];
  wire        bs_50 = b[50];
  wire        bs_51 = b[51];
  wire        bs_52 = b[52];
  wire        bs_53 = b[53];
  wire        bs_54 = b[54];
  wire        bs_55 = b[55];
  wire        bs_56 = b[56];
  wire        bs_57 = b[57];
  wire        bs_58 = b[58];
  wire        bs_59 = b[59];
  wire        bs_60 = b[60];
  wire        bs_61 = b[61];
  wire        bs_62 = b[62];
  wire        bs_63 = b[63];
  wire        pairs_0_1 = as_0 ^ bs_0;
  wire        pairs_0_2 = as_0 & bs_0;
  wire        pairs_1_1 = as_1 ^ bs_1;
  wire        pairs_1_2 = as_1 & bs_1;
  wire        pairs_2_1 = as_2 ^ bs_2;
  wire        pairs_2_2 = as_2 & bs_2;
  wire        pairs_3_1 = as_3 ^ bs_3;
  wire        pairs_3_2 = as_3 & bs_3;
  wire        pairs_4_1 = as_4 ^ bs_4;
  wire        pairs_4_2 = as_4 & bs_4;
  wire        pairs_5_1 = as_5 ^ bs_5;
  wire        pairs_5_2 = as_5 & bs_5;
  wire        pairs_6_1 = as_6 ^ bs_6;
  wire        pairs_6_2 = as_6 & bs_6;
  wire        pairs_7_1 = as_7 ^ bs_7;
  wire        pairs_7_2 = as_7 & bs_7;
  wire        pairs_8_1 = as_8 ^ bs_8;
  wire        pairs_8_2 = as_8 & bs_8;
  wire        pairs_9_1 = as_9 ^ bs_9;
  wire        pairs_9_2 = as_9 & bs_9;
  wire        pairs_10_1 = as_10 ^ bs_10;
  wire        pairs_10_2 = as_10 & bs_10;
  wire        pairs_11_1 = as_11 ^ bs_11;
  wire        pairs_11_2 = as_11 & bs_11;
  wire        pairs_12_1 = as_12 ^ bs_12;
  wire        pairs_12_2 = as_12 & bs_12;
  wire        pairs_13_1 = as_13 ^ bs_13;
  wire        pairs_13_2 = as_13 & bs_13;
  wire        pairs_14_1 = as_14 ^ bs_14;
  wire        pairs_14_2 = as_14 & bs_14;
  wire        pairs_15_1 = as_15 ^ bs_15;
  wire        pairs_15_2 = as_15 & bs_15;
  wire        pairs_16_1 = as_16 ^ bs_16;
  wire        pairs_16_2 = as_16 & bs_16;
  wire        pairs_17_1 = as_17 ^ bs_17;
  wire        pairs_17_2 = as_17 & bs_17;
  wire        pairs_18_1 = as_18 ^ bs_18;
  wire        pairs_18_2 = as_18 & bs_18;
  wire        pairs_19_1 = as_19 ^ bs_19;
  wire        pairs_19_2 = as_19 & bs_19;
  wire        pairs_20_1 = as_20 ^ bs_20;
  wire        pairs_20_2 = as_20 & bs_20;
  wire        pairs_21_1 = as_21 ^ bs_21;
  wire        pairs_21_2 = as_21 & bs_21;
  wire        pairs_22_1 = as_22 ^ bs_22;
  wire        pairs_22_2 = as_22 & bs_22;
  wire        pairs_23_1 = as_23 ^ bs_23;
  wire        pairs_23_2 = as_23 & bs_23;
  wire        pairs_24_1 = as_24 ^ bs_24;
  wire        pairs_24_2 = as_24 & bs_24;
  wire        pairs_25_1 = as_25 ^ bs_25;
  wire        pairs_25_2 = as_25 & bs_25;
  wire        pairs_26_1 = as_26 ^ bs_26;
  wire        pairs_26_2 = as_26 & bs_26;
  wire        pairs_27_1 = as_27 ^ bs_27;
  wire        pairs_27_2 = as_27 & bs_27;
  wire        pairs_28_1 = as_28 ^ bs_28;
  wire        pairs_28_2 = as_28 & bs_28;
  wire        pairs_29_1 = as_29 ^ bs_29;
  wire        pairs_29_2 = as_29 & bs_29;
  wire        pairs_30_1 = as_30 ^ bs_30;
  wire        pairs_30_2 = as_30 & bs_30;
  wire        pairs_31_1 = as_31 ^ bs_31;
  wire        pairs_31_2 = as_31 & bs_31;
  wire        pairs_32_1 = as_32 ^ bs_32;
  wire        pairs_32_2 = as_32 & bs_32;
  wire        pairs_33_1 = as_33 ^ bs_33;
  wire        pairs_33_2 = as_33 & bs_33;
  wire        pairs_34_1 = as_34 ^ bs_34;
  wire        pairs_34_2 = as_34 & bs_34;
  wire        pairs_35_1 = as_35 ^ bs_35;
  wire        pairs_35_2 = as_35 & bs_35;
  wire        pairs_36_1 = as_36 ^ bs_36;
  wire        pairs_36_2 = as_36 & bs_36;
  wire        pairs_37_1 = as_37 ^ bs_37;
  wire        pairs_37_2 = as_37 & bs_37;
  wire        pairs_38_1 = as_38 ^ bs_38;
  wire        pairs_38_2 = as_38 & bs_38;
  wire        pairs_39_1 = as_39 ^ bs_39;
  wire        pairs_39_2 = as_39 & bs_39;
  wire        pairs_40_1 = as_40 ^ bs_40;
  wire        pairs_40_2 = as_40 & bs_40;
  wire        pairs_41_1 = as_41 ^ bs_41;
  wire        pairs_41_2 = as_41 & bs_41;
  wire        pairs_42_1 = as_42 ^ bs_42;
  wire        pairs_42_2 = as_42 & bs_42;
  wire        pairs_43_1 = as_43 ^ bs_43;
  wire        pairs_43_2 = as_43 & bs_43;
  wire        pairs_44_1 = as_44 ^ bs_44;
  wire        pairs_44_2 = as_44 & bs_44;
  wire        pairs_45_1 = as_45 ^ bs_45;
  wire        pairs_45_2 = as_45 & bs_45;
  wire        pairs_46_1 = as_46 ^ bs_46;
  wire        pairs_46_2 = as_46 & bs_46;
  wire        pairs_47_1 = as_47 ^ bs_47;
  wire        pairs_47_2 = as_47 & bs_47;
  wire        pairs_48_1 = as_48 ^ bs_48;
  wire        pairs_48_2 = as_48 & bs_48;
  wire        pairs_49_1 = as_49 ^ bs_49;
  wire        pairs_49_2 = as_49 & bs_49;
  wire        pairs_50_1 = as_50 ^ bs_50;
  wire        pairs_50_2 = as_50 & bs_50;
  wire        pairs_51_1 = as_51 ^ bs_51;
  wire        pairs_51_2 = as_51 & bs_51;
  wire        pairs_52_1 = as_52 ^ bs_52;
  wire        pairs_52_2 = as_52 & bs_52;
  wire        pairs_53_1 = as_53 ^ bs_53;
  wire        pairs_53_2 = as_53 & bs_53;
  wire        pairs_54_1 = as_54 ^ bs_54;
  wire        pairs_54_2 = as_54 & bs_54;
  wire        pairs_55_1 = as_55 ^ bs_55;
  wire        pairs_55_2 = as_55 & bs_55;
  wire        pairs_56_1 = as_56 ^ bs_56;
  wire        pairs_56_2 = as_56 & bs_56;
  wire        pairs_57_1 = as_57 ^ bs_57;
  wire        pairs_57_2 = as_57 & bs_57;
  wire        pairs_58_1 = as_58 ^ bs_58;
  wire        pairs_58_2 = as_58 & bs_58;
  wire        pairs_59_1 = as_59 ^ bs_59;
  wire        pairs_59_2 = as_59 & bs_59;
  wire        pairs_60_1 = as_60 ^ bs_60;
  wire        pairs_60_2 = as_60 & bs_60;
  wire        pairs_61_1 = as_61 ^ bs_61;
  wire        pairs_61_2 = as_61 & bs_61;
  wire        pairs_62_1 = as_62 ^ bs_62;
  wire        pairs_62_2 = as_62 & bs_62;
  wire        pairs_63_1 = as_63 ^ bs_63;
  wire        pairs_63_2 = as_63 & bs_63;
  wire        tree8Leaf_layer0_0_1 = pairs_7_1 & pairs_6_1;
  wire        tree8Leaf_layer0_0_2 = pairs_7_2 | pairs_7_1 & pairs_6_2;
  wire        tree8Leaf_layer0_1_1 = pairs_5_1 & pairs_4_1;
  wire        tree8Leaf_layer0_1_2 = pairs_5_2 | pairs_5_1 & pairs_4_2;
  wire        tree8Leaf_layer0_2_1 = pairs_3_1 & pairs_2_1;
  wire        tree8Leaf_layer0_2_2 = pairs_3_2 | pairs_3_1 & pairs_2_2;
  wire        tree8Leaf_0_1_1 = pairs_1_1 & pairs_0_1;
  wire        tree8Leaf_0_1_2 = pairs_1_2 | pairs_1_1 & pairs_0_2;
  wire        tree8Leaf_layer1_0_1 = tree8Leaf_layer0_0_1 & tree8Leaf_layer0_1_1;
  wire        tree8Leaf_layer1_0_2 = tree8Leaf_layer0_0_2 | tree8Leaf_layer0_0_1 & tree8Leaf_layer0_1_2;
  wire        tree8Leaf_0_3_1 = tree8Leaf_layer0_2_1 & tree8Leaf_0_1_1;
  wire        tree8Leaf_0_3_2 = tree8Leaf_layer0_2_2 | tree8Leaf_layer0_2_1 & tree8Leaf_0_1_2;
  wire        tree8Leaf_0_2_1 = pairs_2_1 & tree8Leaf_0_1_1;
  wire        tree8Leaf_0_2_2 = pairs_2_2 | pairs_2_1 & tree8Leaf_0_1_2;
  wire        tree8Leaf_0_4_1 = pairs_4_1 & tree8Leaf_0_3_1;
  wire        tree8Leaf_0_4_2 = pairs_4_2 | pairs_4_1 & tree8Leaf_0_3_2;
  wire        tree8Leaf_0_5_1 = tree8Leaf_layer0_1_1 & tree8Leaf_0_3_1;
  wire        tree8Leaf_0_5_2 = tree8Leaf_layer0_1_2 | tree8Leaf_layer0_1_1 & tree8Leaf_0_3_2;
  wire        tree8Leaf_0_6_1 = pairs_6_1 & tree8Leaf_0_5_1;
  wire        tree8Leaf_0_6_2 = pairs_6_2 | pairs_6_1 & tree8Leaf_0_5_2;
  wire        tree8Leaf_0_7_1 = tree8Leaf_layer1_0_1 & tree8Leaf_0_3_1;
  wire        tree8Leaf_0_7_2 = tree8Leaf_layer1_0_2 | tree8Leaf_layer1_0_1 & tree8Leaf_0_3_2;
  wire        tree8Leaf_layer0_0_1_1 = pairs_15_1 & pairs_14_1;
  wire        tree8Leaf_layer0_0_2_1 = pairs_15_2 | pairs_15_1 & pairs_14_2;
  wire        tree8Leaf_layer0_1_1_1 = pairs_13_1 & pairs_12_1;
  wire        tree8Leaf_layer0_1_2_1 = pairs_13_2 | pairs_13_1 & pairs_12_2;
  wire        tree8Leaf_layer0_2_1_1 = pairs_11_1 & pairs_10_1;
  wire        tree8Leaf_layer0_2_2_1 = pairs_11_2 | pairs_11_1 & pairs_10_2;
  wire        tree8Leaf_1_1_1 = pairs_9_1 & pairs_8_1;
  wire        tree8Leaf_1_1_2 = pairs_9_2 | pairs_9_1 & pairs_8_2;
  wire        tree8Leaf_layer1_0_1_1 = tree8Leaf_layer0_0_1_1 & tree8Leaf_layer0_1_1_1;
  wire        tree8Leaf_layer1_0_2_1 = tree8Leaf_layer0_0_2_1 | tree8Leaf_layer0_0_1_1 & tree8Leaf_layer0_1_2_1;
  wire        tree8Leaf_1_3_1 = tree8Leaf_layer0_2_1_1 & tree8Leaf_1_1_1;
  wire        tree8Leaf_1_3_2 = tree8Leaf_layer0_2_2_1 | tree8Leaf_layer0_2_1_1 & tree8Leaf_1_1_2;
  wire        tree8Leaf_1_2_1 = pairs_10_1 & tree8Leaf_1_1_1;
  wire        tree8Leaf_1_2_2 = pairs_10_2 | pairs_10_1 & tree8Leaf_1_1_2;
  wire        tree8Leaf_1_4_1 = pairs_12_1 & tree8Leaf_1_3_1;
  wire        tree8Leaf_1_4_2 = pairs_12_2 | pairs_12_1 & tree8Leaf_1_3_2;
  wire        tree8Leaf_1_5_1 = tree8Leaf_layer0_1_1_1 & tree8Leaf_1_3_1;
  wire        tree8Leaf_1_5_2 = tree8Leaf_layer0_1_2_1 | tree8Leaf_layer0_1_1_1 & tree8Leaf_1_3_2;
  wire        tree8Leaf_1_6_1 = pairs_14_1 & tree8Leaf_1_5_1;
  wire        tree8Leaf_1_6_2 = pairs_14_2 | pairs_14_1 & tree8Leaf_1_5_2;
  wire        tree8Leaf_1_7_1 = tree8Leaf_layer1_0_1_1 & tree8Leaf_1_3_1;
  wire        tree8Leaf_1_7_2 = tree8Leaf_layer1_0_2_1 | tree8Leaf_layer1_0_1_1 & tree8Leaf_1_3_2;
  wire        tree8Leaf_layer0_0_1_2 = pairs_23_1 & pairs_22_1;
  wire        tree8Leaf_layer0_0_2_2 = pairs_23_2 | pairs_23_1 & pairs_22_2;
  wire        tree8Leaf_layer0_1_1_2 = pairs_21_1 & pairs_20_1;
  wire        tree8Leaf_layer0_1_2_2 = pairs_21_2 | pairs_21_1 & pairs_20_2;
  wire        tree8Leaf_layer0_2_1_2 = pairs_19_1 & pairs_18_1;
  wire        tree8Leaf_layer0_2_2_2 = pairs_19_2 | pairs_19_1 & pairs_18_2;
  wire        tree8Leaf_2_1_1 = pairs_17_1 & pairs_16_1;
  wire        tree8Leaf_2_1_2 = pairs_17_2 | pairs_17_1 & pairs_16_2;
  wire        tree8Leaf_layer1_0_1_2 = tree8Leaf_layer0_0_1_2 & tree8Leaf_layer0_1_1_2;
  wire        tree8Leaf_layer1_0_2_2 = tree8Leaf_layer0_0_2_2 | tree8Leaf_layer0_0_1_2 & tree8Leaf_layer0_1_2_2;
  wire        tree8Leaf_2_3_1 = tree8Leaf_layer0_2_1_2 & tree8Leaf_2_1_1;
  wire        tree8Leaf_2_3_2 = tree8Leaf_layer0_2_2_2 | tree8Leaf_layer0_2_1_2 & tree8Leaf_2_1_2;
  wire        tree8Leaf_2_2_1 = pairs_18_1 & tree8Leaf_2_1_1;
  wire        tree8Leaf_2_2_2 = pairs_18_2 | pairs_18_1 & tree8Leaf_2_1_2;
  wire        tree8Leaf_2_4_1 = pairs_20_1 & tree8Leaf_2_3_1;
  wire        tree8Leaf_2_4_2 = pairs_20_2 | pairs_20_1 & tree8Leaf_2_3_2;
  wire        tree8Leaf_2_5_1 = tree8Leaf_layer0_1_1_2 & tree8Leaf_2_3_1;
  wire        tree8Leaf_2_5_2 = tree8Leaf_layer0_1_2_2 | tree8Leaf_layer0_1_1_2 & tree8Leaf_2_3_2;
  wire        tree8Leaf_2_6_1 = pairs_22_1 & tree8Leaf_2_5_1;
  wire        tree8Leaf_2_6_2 = pairs_22_2 | pairs_22_1 & tree8Leaf_2_5_2;
  wire        tree8Leaf_2_7_1 = tree8Leaf_layer1_0_1_2 & tree8Leaf_2_3_1;
  wire        tree8Leaf_2_7_2 = tree8Leaf_layer1_0_2_2 | tree8Leaf_layer1_0_1_2 & tree8Leaf_2_3_2;
  wire        tree8Leaf_layer0_0_1_3 = pairs_31_1 & pairs_30_1;
  wire        tree8Leaf_layer0_0_2_3 = pairs_31_2 | pairs_31_1 & pairs_30_2;
  wire        tree8Leaf_layer0_1_1_3 = pairs_29_1 & pairs_28_1;
  wire        tree8Leaf_layer0_1_2_3 = pairs_29_2 | pairs_29_1 & pairs_28_2;
  wire        tree8Leaf_layer0_2_1_3 = pairs_27_1 & pairs_26_1;
  wire        tree8Leaf_layer0_2_2_3 = pairs_27_2 | pairs_27_1 & pairs_26_2;
  wire        tree8Leaf_3_1_1 = pairs_25_1 & pairs_24_1;
  wire        tree8Leaf_3_1_2 = pairs_25_2 | pairs_25_1 & pairs_24_2;
  wire        tree8Leaf_layer1_0_1_3 = tree8Leaf_layer0_0_1_3 & tree8Leaf_layer0_1_1_3;
  wire        tree8Leaf_layer1_0_2_3 = tree8Leaf_layer0_0_2_3 | tree8Leaf_layer0_0_1_3 & tree8Leaf_layer0_1_2_3;
  wire        tree8Leaf_3_3_1 = tree8Leaf_layer0_2_1_3 & tree8Leaf_3_1_1;
  wire        tree8Leaf_3_3_2 = tree8Leaf_layer0_2_2_3 | tree8Leaf_layer0_2_1_3 & tree8Leaf_3_1_2;
  wire        tree8Leaf_3_2_1 = pairs_26_1 & tree8Leaf_3_1_1;
  wire        tree8Leaf_3_2_2 = pairs_26_2 | pairs_26_1 & tree8Leaf_3_1_2;
  wire        tree8Leaf_3_4_1 = pairs_28_1 & tree8Leaf_3_3_1;
  wire        tree8Leaf_3_4_2 = pairs_28_2 | pairs_28_1 & tree8Leaf_3_3_2;
  wire        tree8Leaf_3_5_1 = tree8Leaf_layer0_1_1_3 & tree8Leaf_3_3_1;
  wire        tree8Leaf_3_5_2 = tree8Leaf_layer0_1_2_3 | tree8Leaf_layer0_1_1_3 & tree8Leaf_3_3_2;
  wire        tree8Leaf_3_6_1 = pairs_30_1 & tree8Leaf_3_5_1;
  wire        tree8Leaf_3_6_2 = pairs_30_2 | pairs_30_1 & tree8Leaf_3_5_2;
  wire        tree8Leaf_3_7_1 = tree8Leaf_layer1_0_1_3 & tree8Leaf_3_3_1;
  wire        tree8Leaf_3_7_2 = tree8Leaf_layer1_0_2_3 | tree8Leaf_layer1_0_1_3 & tree8Leaf_3_3_2;
  wire        tree8Leaf_layer0_0_1_4 = pairs_39_1 & pairs_38_1;
  wire        tree8Leaf_layer0_0_2_4 = pairs_39_2 | pairs_39_1 & pairs_38_2;
  wire        tree8Leaf_layer0_1_1_4 = pairs_37_1 & pairs_36_1;
  wire        tree8Leaf_layer0_1_2_4 = pairs_37_2 | pairs_37_1 & pairs_36_2;
  wire        tree8Leaf_layer0_2_1_4 = pairs_35_1 & pairs_34_1;
  wire        tree8Leaf_layer0_2_2_4 = pairs_35_2 | pairs_35_1 & pairs_34_2;
  wire        tree8Leaf_4_1_1 = pairs_33_1 & pairs_32_1;
  wire        tree8Leaf_4_1_2 = pairs_33_2 | pairs_33_1 & pairs_32_2;
  wire        tree8Leaf_layer1_0_1_4 = tree8Leaf_layer0_0_1_4 & tree8Leaf_layer0_1_1_4;
  wire        tree8Leaf_layer1_0_2_4 = tree8Leaf_layer0_0_2_4 | tree8Leaf_layer0_0_1_4 & tree8Leaf_layer0_1_2_4;
  wire        tree8Leaf_4_3_1 = tree8Leaf_layer0_2_1_4 & tree8Leaf_4_1_1;
  wire        tree8Leaf_4_3_2 = tree8Leaf_layer0_2_2_4 | tree8Leaf_layer0_2_1_4 & tree8Leaf_4_1_2;
  wire        tree8Leaf_4_2_1 = pairs_34_1 & tree8Leaf_4_1_1;
  wire        tree8Leaf_4_2_2 = pairs_34_2 | pairs_34_1 & tree8Leaf_4_1_2;
  wire        tree8Leaf_4_4_1 = pairs_36_1 & tree8Leaf_4_3_1;
  wire        tree8Leaf_4_4_2 = pairs_36_2 | pairs_36_1 & tree8Leaf_4_3_2;
  wire        tree8Leaf_4_5_1 = tree8Leaf_layer0_1_1_4 & tree8Leaf_4_3_1;
  wire        tree8Leaf_4_5_2 = tree8Leaf_layer0_1_2_4 | tree8Leaf_layer0_1_1_4 & tree8Leaf_4_3_2;
  wire        tree8Leaf_4_6_1 = pairs_38_1 & tree8Leaf_4_5_1;
  wire        tree8Leaf_4_6_2 = pairs_38_2 | pairs_38_1 & tree8Leaf_4_5_2;
  wire        tree8Leaf_4_7_1 = tree8Leaf_layer1_0_1_4 & tree8Leaf_4_3_1;
  wire        tree8Leaf_4_7_2 = tree8Leaf_layer1_0_2_4 | tree8Leaf_layer1_0_1_4 & tree8Leaf_4_3_2;
  wire        tree8Leaf_layer0_0_1_5 = pairs_47_1 & pairs_46_1;
  wire        tree8Leaf_layer0_0_2_5 = pairs_47_2 | pairs_47_1 & pairs_46_2;
  wire        tree8Leaf_layer0_1_1_5 = pairs_45_1 & pairs_44_1;
  wire        tree8Leaf_layer0_1_2_5 = pairs_45_2 | pairs_45_1 & pairs_44_2;
  wire        tree8Leaf_layer0_2_1_5 = pairs_43_1 & pairs_42_1;
  wire        tree8Leaf_layer0_2_2_5 = pairs_43_2 | pairs_43_1 & pairs_42_2;
  wire        tree8Leaf_5_1_1 = pairs_41_1 & pairs_40_1;
  wire        tree8Leaf_5_1_2 = pairs_41_2 | pairs_41_1 & pairs_40_2;
  wire        tree8Leaf_layer1_0_1_5 = tree8Leaf_layer0_0_1_5 & tree8Leaf_layer0_1_1_5;
  wire        tree8Leaf_layer1_0_2_5 = tree8Leaf_layer0_0_2_5 | tree8Leaf_layer0_0_1_5 & tree8Leaf_layer0_1_2_5;
  wire        tree8Leaf_5_3_1 = tree8Leaf_layer0_2_1_5 & tree8Leaf_5_1_1;
  wire        tree8Leaf_5_3_2 = tree8Leaf_layer0_2_2_5 | tree8Leaf_layer0_2_1_5 & tree8Leaf_5_1_2;
  wire        tree8Leaf_5_2_1 = pairs_42_1 & tree8Leaf_5_1_1;
  wire        tree8Leaf_5_2_2 = pairs_42_2 | pairs_42_1 & tree8Leaf_5_1_2;
  wire        tree8Leaf_5_4_1 = pairs_44_1 & tree8Leaf_5_3_1;
  wire        tree8Leaf_5_4_2 = pairs_44_2 | pairs_44_1 & tree8Leaf_5_3_2;
  wire        tree8Leaf_5_5_1 = tree8Leaf_layer0_1_1_5 & tree8Leaf_5_3_1;
  wire        tree8Leaf_5_5_2 = tree8Leaf_layer0_1_2_5 | tree8Leaf_layer0_1_1_5 & tree8Leaf_5_3_2;
  wire        tree8Leaf_5_6_1 = pairs_46_1 & tree8Leaf_5_5_1;
  wire        tree8Leaf_5_6_2 = pairs_46_2 | pairs_46_1 & tree8Leaf_5_5_2;
  wire        tree8Leaf_5_7_1 = tree8Leaf_layer1_0_1_5 & tree8Leaf_5_3_1;
  wire        tree8Leaf_5_7_2 = tree8Leaf_layer1_0_2_5 | tree8Leaf_layer1_0_1_5 & tree8Leaf_5_3_2;
  wire        tree8Leaf_layer0_0_1_6 = pairs_55_1 & pairs_54_1;
  wire        tree8Leaf_layer0_0_2_6 = pairs_55_2 | pairs_55_1 & pairs_54_2;
  wire        tree8Leaf_layer0_1_1_6 = pairs_53_1 & pairs_52_1;
  wire        tree8Leaf_layer0_1_2_6 = pairs_53_2 | pairs_53_1 & pairs_52_2;
  wire        tree8Leaf_layer0_2_1_6 = pairs_51_1 & pairs_50_1;
  wire        tree8Leaf_layer0_2_2_6 = pairs_51_2 | pairs_51_1 & pairs_50_2;
  wire        tree8Leaf_6_1_1 = pairs_49_1 & pairs_48_1;
  wire        tree8Leaf_6_1_2 = pairs_49_2 | pairs_49_1 & pairs_48_2;
  wire        tree8Leaf_layer1_0_1_6 = tree8Leaf_layer0_0_1_6 & tree8Leaf_layer0_1_1_6;
  wire        tree8Leaf_layer1_0_2_6 = tree8Leaf_layer0_0_2_6 | tree8Leaf_layer0_0_1_6 & tree8Leaf_layer0_1_2_6;
  wire        tree8Leaf_6_3_1 = tree8Leaf_layer0_2_1_6 & tree8Leaf_6_1_1;
  wire        tree8Leaf_6_3_2 = tree8Leaf_layer0_2_2_6 | tree8Leaf_layer0_2_1_6 & tree8Leaf_6_1_2;
  wire        tree8Leaf_6_2_1 = pairs_50_1 & tree8Leaf_6_1_1;
  wire        tree8Leaf_6_2_2 = pairs_50_2 | pairs_50_1 & tree8Leaf_6_1_2;
  wire        tree8Leaf_6_4_1 = pairs_52_1 & tree8Leaf_6_3_1;
  wire        tree8Leaf_6_4_2 = pairs_52_2 | pairs_52_1 & tree8Leaf_6_3_2;
  wire        tree8Leaf_6_5_1 = tree8Leaf_layer0_1_1_6 & tree8Leaf_6_3_1;
  wire        tree8Leaf_6_5_2 = tree8Leaf_layer0_1_2_6 | tree8Leaf_layer0_1_1_6 & tree8Leaf_6_3_2;
  wire        tree8Leaf_6_6_1 = pairs_54_1 & tree8Leaf_6_5_1;
  wire        tree8Leaf_6_6_2 = pairs_54_2 | pairs_54_1 & tree8Leaf_6_5_2;
  wire        tree8Leaf_6_7_1 = tree8Leaf_layer1_0_1_6 & tree8Leaf_6_3_1;
  wire        tree8Leaf_6_7_2 = tree8Leaf_layer1_0_2_6 | tree8Leaf_layer1_0_1_6 & tree8Leaf_6_3_2;
  wire        tree8Leaf_layer0_0_1_7 = pairs_63_1 & pairs_62_1;
  wire        tree8Leaf_layer0_0_2_7 = pairs_63_2 | pairs_63_1 & pairs_62_2;
  wire        tree8Leaf_layer0_1_1_7 = pairs_61_1 & pairs_60_1;
  wire        tree8Leaf_layer0_1_2_7 = pairs_61_2 | pairs_61_1 & pairs_60_2;
  wire        tree8Leaf_layer0_2_1_7 = pairs_59_1 & pairs_58_1;
  wire        tree8Leaf_layer0_2_2_7 = pairs_59_2 | pairs_59_1 & pairs_58_2;
  wire        tree8Leaf_7_1_1 = pairs_57_1 & pairs_56_1;
  wire        tree8Leaf_7_1_2 = pairs_57_2 | pairs_57_1 & pairs_56_2;
  wire        tree8Leaf_layer1_0_1_7 = tree8Leaf_layer0_0_1_7 & tree8Leaf_layer0_1_1_7;
  wire        tree8Leaf_layer1_0_2_7 = tree8Leaf_layer0_0_2_7 | tree8Leaf_layer0_0_1_7 & tree8Leaf_layer0_1_2_7;
  wire        tree8Leaf_7_3_1 = tree8Leaf_layer0_2_1_7 & tree8Leaf_7_1_1;
  wire        tree8Leaf_7_3_2 = tree8Leaf_layer0_2_2_7 | tree8Leaf_layer0_2_1_7 & tree8Leaf_7_1_2;
  wire        tree8Leaf_7_2_1 = pairs_58_1 & tree8Leaf_7_1_1;
  wire        tree8Leaf_7_2_2 = pairs_58_2 | pairs_58_1 & tree8Leaf_7_1_2;
  wire        tree8Leaf_7_4_1 = pairs_60_1 & tree8Leaf_7_3_1;
  wire        tree8Leaf_7_4_2 = pairs_60_2 | pairs_60_1 & tree8Leaf_7_3_2;
  wire        tree8Leaf_7_5_1 = tree8Leaf_layer0_1_1_7 & tree8Leaf_7_3_1;
  wire        tree8Leaf_7_5_2 = tree8Leaf_layer0_1_2_7 | tree8Leaf_layer0_1_1_7 & tree8Leaf_7_3_2;
  wire        tree8Leaf_7_6_1 = pairs_62_1 & tree8Leaf_7_5_1;
  wire        tree8Leaf_7_6_2 = pairs_62_2 | pairs_62_1 & tree8Leaf_7_5_2;
  wire        tree8Leaf_7_7_1 = tree8Leaf_layer1_0_1_7 & tree8Leaf_7_3_1;
  wire        tree8Leaf_7_7_2 = tree8Leaf_layer1_0_2_7 | tree8Leaf_layer1_0_1_7 & tree8Leaf_7_3_2;
  wire        tree16Leaf0_8_1 = pairs_8_1 & tree8Leaf_0_7_1;
  wire        tree16Leaf0_8_2 = pairs_8_2 | pairs_8_1 & tree8Leaf_0_7_2;
  wire        tree16Leaf0_9_1 = tree8Leaf_1_1_1 & tree8Leaf_0_7_1;
  wire        tree16Leaf0_9_2 = tree8Leaf_1_1_2 | tree8Leaf_1_1_1 & tree8Leaf_0_7_2;
  wire        tree16Leaf0_10_1 = tree8Leaf_1_2_1 & tree8Leaf_0_7_1;
  wire        tree16Leaf0_10_2 = tree8Leaf_1_2_2 | tree8Leaf_1_2_1 & tree8Leaf_0_7_2;
  wire        tree16Leaf0_11_1 = tree8Leaf_1_3_1 & tree8Leaf_0_7_1;
  wire        tree16Leaf0_11_2 = tree8Leaf_1_3_2 | tree8Leaf_1_3_1 & tree8Leaf_0_7_2;
  wire        tree16Leaf0_12_1 = tree8Leaf_1_4_1 & tree8Leaf_0_7_1;
  wire        tree16Leaf0_12_2 = tree8Leaf_1_4_2 | tree8Leaf_1_4_1 & tree8Leaf_0_7_2;
  wire        tree16Leaf0_13_1 = tree8Leaf_1_5_1 & tree8Leaf_0_7_1;
  wire        tree16Leaf0_13_2 = tree8Leaf_1_5_2 | tree8Leaf_1_5_1 & tree8Leaf_0_7_2;
  wire        tree16Leaf0_14_1 = tree8Leaf_1_6_1 & tree8Leaf_0_7_1;
  wire        tree16Leaf0_14_2 = tree8Leaf_1_6_2 | tree8Leaf_1_6_1 & tree8Leaf_0_7_2;
  wire        tree16Leaf0_15_1 = tree8Leaf_1_7_1 & tree8Leaf_0_7_1;
  wire        tree16Leaf0_15_2 = tree8Leaf_1_7_2 | tree8Leaf_1_7_1 & tree8Leaf_0_7_2;
  wire        tree16Leaf1_8_1 = pairs_24_1 & tree8Leaf_2_7_1;
  wire        tree16Leaf1_8_2 = pairs_24_2 | pairs_24_1 & tree8Leaf_2_7_2;
  wire        tree16Leaf1_9_1 = tree8Leaf_3_1_1 & tree8Leaf_2_7_1;
  wire        tree16Leaf1_9_2 = tree8Leaf_3_1_2 | tree8Leaf_3_1_1 & tree8Leaf_2_7_2;
  wire        tree16Leaf1_10_1 = tree8Leaf_3_2_1 & tree8Leaf_2_7_1;
  wire        tree16Leaf1_10_2 = tree8Leaf_3_2_2 | tree8Leaf_3_2_1 & tree8Leaf_2_7_2;
  wire        tree16Leaf1_11_1 = tree8Leaf_3_3_1 & tree8Leaf_2_7_1;
  wire        tree16Leaf1_11_2 = tree8Leaf_3_3_2 | tree8Leaf_3_3_1 & tree8Leaf_2_7_2;
  wire        tree16Leaf1_12_1 = tree8Leaf_3_4_1 & tree8Leaf_2_7_1;
  wire        tree16Leaf1_12_2 = tree8Leaf_3_4_2 | tree8Leaf_3_4_1 & tree8Leaf_2_7_2;
  wire        tree16Leaf1_13_1 = tree8Leaf_3_5_1 & tree8Leaf_2_7_1;
  wire        tree16Leaf1_13_2 = tree8Leaf_3_5_2 | tree8Leaf_3_5_1 & tree8Leaf_2_7_2;
  wire        tree16Leaf1_14_1 = tree8Leaf_3_6_1 & tree8Leaf_2_7_1;
  wire        tree16Leaf1_14_2 = tree8Leaf_3_6_2 | tree8Leaf_3_6_1 & tree8Leaf_2_7_2;
  wire        tree16Leaf1_15_1 = tree8Leaf_3_7_1 & tree8Leaf_2_7_1;
  wire        tree16Leaf1_15_2 = tree8Leaf_3_7_2 | tree8Leaf_3_7_1 & tree8Leaf_2_7_2;
  wire        tree16Leaf2_8_1 = pairs_40_1 & tree8Leaf_4_7_1;
  wire        tree16Leaf2_8_2 = pairs_40_2 | pairs_40_1 & tree8Leaf_4_7_2;
  wire        tree16Leaf2_9_1 = tree8Leaf_5_1_1 & tree8Leaf_4_7_1;
  wire        tree16Leaf2_9_2 = tree8Leaf_5_1_2 | tree8Leaf_5_1_1 & tree8Leaf_4_7_2;
  wire        tree16Leaf2_10_1 = tree8Leaf_5_2_1 & tree8Leaf_4_7_1;
  wire        tree16Leaf2_10_2 = tree8Leaf_5_2_2 | tree8Leaf_5_2_1 & tree8Leaf_4_7_2;
  wire        tree16Leaf2_11_1 = tree8Leaf_5_3_1 & tree8Leaf_4_7_1;
  wire        tree16Leaf2_11_2 = tree8Leaf_5_3_2 | tree8Leaf_5_3_1 & tree8Leaf_4_7_2;
  wire        tree16Leaf2_12_1 = tree8Leaf_5_4_1 & tree8Leaf_4_7_1;
  wire        tree16Leaf2_12_2 = tree8Leaf_5_4_2 | tree8Leaf_5_4_1 & tree8Leaf_4_7_2;
  wire        tree16Leaf2_13_1 = tree8Leaf_5_5_1 & tree8Leaf_4_7_1;
  wire        tree16Leaf2_13_2 = tree8Leaf_5_5_2 | tree8Leaf_5_5_1 & tree8Leaf_4_7_2;
  wire        tree16Leaf2_14_1 = tree8Leaf_5_6_1 & tree8Leaf_4_7_1;
  wire        tree16Leaf2_14_2 = tree8Leaf_5_6_2 | tree8Leaf_5_6_1 & tree8Leaf_4_7_2;
  wire        tree16Leaf2_15_1 = tree8Leaf_5_7_1 & tree8Leaf_4_7_1;
  wire        tree16Leaf2_15_2 = tree8Leaf_5_7_2 | tree8Leaf_5_7_1 & tree8Leaf_4_7_2;
  wire        tree16Leaf3_8_1 = pairs_56_1 & tree8Leaf_6_7_1;
  wire        tree16Leaf3_8_2 = pairs_56_2 | pairs_56_1 & tree8Leaf_6_7_2;
  wire        tree16Leaf3_9_1 = tree8Leaf_7_1_1 & tree8Leaf_6_7_1;
  wire        tree16Leaf3_9_2 = tree8Leaf_7_1_2 | tree8Leaf_7_1_1 & tree8Leaf_6_7_2;
  wire        tree16Leaf3_10_1 = tree8Leaf_7_2_1 & tree8Leaf_6_7_1;
  wire        tree16Leaf3_10_2 = tree8Leaf_7_2_2 | tree8Leaf_7_2_1 & tree8Leaf_6_7_2;
  wire        tree16Leaf3_11_1 = tree8Leaf_7_3_1 & tree8Leaf_6_7_1;
  wire        tree16Leaf3_11_2 = tree8Leaf_7_3_2 | tree8Leaf_7_3_1 & tree8Leaf_6_7_2;
  wire        tree16Leaf3_12_1 = tree8Leaf_7_4_1 & tree8Leaf_6_7_1;
  wire        tree16Leaf3_12_2 = tree8Leaf_7_4_2 | tree8Leaf_7_4_1 & tree8Leaf_6_7_2;
  wire        tree16Leaf3_13_1 = tree8Leaf_7_5_1 & tree8Leaf_6_7_1;
  wire        tree16Leaf3_13_2 = tree8Leaf_7_5_2 | tree8Leaf_7_5_1 & tree8Leaf_6_7_2;
  wire        tree16Leaf3_14_1 = tree8Leaf_7_6_1 & tree8Leaf_6_7_1;
  wire        tree16Leaf3_14_2 = tree8Leaf_7_6_2 | tree8Leaf_7_6_1 & tree8Leaf_6_7_2;
  wire        tree16Leaf3_15_1 = tree8Leaf_7_7_1 & tree8Leaf_6_7_1;
  wire        tree16Leaf3_15_2 = tree8Leaf_7_7_2 | tree8Leaf_7_7_1 & tree8Leaf_6_7_2;
  wire        tree32Leaf0_16_1 = pairs_16_1 & tree16Leaf0_15_1;
  wire        tree32Leaf0_16_2 = pairs_16_2 | pairs_16_1 & tree16Leaf0_15_2;
  wire        tree32Leaf0_17_1 = tree8Leaf_2_1_1 & tree16Leaf0_15_1;
  wire        tree32Leaf0_17_2 = tree8Leaf_2_1_2 | tree8Leaf_2_1_1 & tree16Leaf0_15_2;
  wire        tree32Leaf0_18_1 = tree8Leaf_2_2_1 & tree16Leaf0_15_1;
  wire        tree32Leaf0_18_2 = tree8Leaf_2_2_2 | tree8Leaf_2_2_1 & tree16Leaf0_15_2;
  wire        tree32Leaf0_19_1 = tree8Leaf_2_3_1 & tree16Leaf0_15_1;
  wire        tree32Leaf0_19_2 = tree8Leaf_2_3_2 | tree8Leaf_2_3_1 & tree16Leaf0_15_2;
  wire        tree32Leaf0_20_1 = tree8Leaf_2_4_1 & tree16Leaf0_15_1;
  wire        tree32Leaf0_20_2 = tree8Leaf_2_4_2 | tree8Leaf_2_4_1 & tree16Leaf0_15_2;
  wire        tree32Leaf0_21_1 = tree8Leaf_2_5_1 & tree16Leaf0_15_1;
  wire        tree32Leaf0_21_2 = tree8Leaf_2_5_2 | tree8Leaf_2_5_1 & tree16Leaf0_15_2;
  wire        tree32Leaf0_22_1 = tree8Leaf_2_6_1 & tree16Leaf0_15_1;
  wire        tree32Leaf0_22_2 = tree8Leaf_2_6_2 | tree8Leaf_2_6_1 & tree16Leaf0_15_2;
  wire        tree32Leaf0_23_1 = tree8Leaf_2_7_1 & tree16Leaf0_15_1;
  wire        tree32Leaf0_23_2 = tree8Leaf_2_7_2 | tree8Leaf_2_7_1 & tree16Leaf0_15_2;
  wire        tree32Leaf0_24_1 = tree16Leaf1_8_1 & tree16Leaf0_15_1;
  wire        tree32Leaf0_24_2 = tree16Leaf1_8_2 | tree16Leaf1_8_1 & tree16Leaf0_15_2;
  wire        tree32Leaf0_25_1 = tree16Leaf1_9_1 & tree16Leaf0_15_1;
  wire        tree32Leaf0_25_2 = tree16Leaf1_9_2 | tree16Leaf1_9_1 & tree16Leaf0_15_2;
  wire        tree32Leaf0_26_1 = tree16Leaf1_10_1 & tree16Leaf0_15_1;
  wire        tree32Leaf0_26_2 = tree16Leaf1_10_2 | tree16Leaf1_10_1 & tree16Leaf0_15_2;
  wire        tree32Leaf0_27_1 = tree16Leaf1_11_1 & tree16Leaf0_15_1;
  wire        tree32Leaf0_27_2 = tree16Leaf1_11_2 | tree16Leaf1_11_1 & tree16Leaf0_15_2;
  wire        tree32Leaf0_28_1 = tree16Leaf1_12_1 & tree16Leaf0_15_1;
  wire        tree32Leaf0_28_2 = tree16Leaf1_12_2 | tree16Leaf1_12_1 & tree16Leaf0_15_2;
  wire        tree32Leaf0_29_1 = tree16Leaf1_13_1 & tree16Leaf0_15_1;
  wire        tree32Leaf0_29_2 = tree16Leaf1_13_2 | tree16Leaf1_13_1 & tree16Leaf0_15_2;
  wire        tree32Leaf0_30_1 = tree16Leaf1_14_1 & tree16Leaf0_15_1;
  wire        tree32Leaf0_30_2 = tree16Leaf1_14_2 | tree16Leaf1_14_1 & tree16Leaf0_15_2;
  wire        tree32Leaf0_31_1 = tree16Leaf1_15_1 & tree16Leaf0_15_1;
  wire        tree32Leaf0_31_2 = tree16Leaf1_15_2 | tree16Leaf1_15_1 & tree16Leaf0_15_2;
  wire        tree32Leaf1_16_1 = pairs_48_1 & tree16Leaf2_15_1;
  wire        tree32Leaf1_16_2 = pairs_48_2 | pairs_48_1 & tree16Leaf2_15_2;
  wire        tree32Leaf1_17_1 = tree8Leaf_6_1_1 & tree16Leaf2_15_1;
  wire        tree32Leaf1_17_2 = tree8Leaf_6_1_2 | tree8Leaf_6_1_1 & tree16Leaf2_15_2;
  wire        tree32Leaf1_18_1 = tree8Leaf_6_2_1 & tree16Leaf2_15_1;
  wire        tree32Leaf1_18_2 = tree8Leaf_6_2_2 | tree8Leaf_6_2_1 & tree16Leaf2_15_2;
  wire        tree32Leaf1_19_1 = tree8Leaf_6_3_1 & tree16Leaf2_15_1;
  wire        tree32Leaf1_19_2 = tree8Leaf_6_3_2 | tree8Leaf_6_3_1 & tree16Leaf2_15_2;
  wire        tree32Leaf1_20_1 = tree8Leaf_6_4_1 & tree16Leaf2_15_1;
  wire        tree32Leaf1_20_2 = tree8Leaf_6_4_2 | tree8Leaf_6_4_1 & tree16Leaf2_15_2;
  wire        tree32Leaf1_21_1 = tree8Leaf_6_5_1 & tree16Leaf2_15_1;
  wire        tree32Leaf1_21_2 = tree8Leaf_6_5_2 | tree8Leaf_6_5_1 & tree16Leaf2_15_2;
  wire        tree32Leaf1_22_1 = tree8Leaf_6_6_1 & tree16Leaf2_15_1;
  wire        tree32Leaf1_22_2 = tree8Leaf_6_6_2 | tree8Leaf_6_6_1 & tree16Leaf2_15_2;
  wire        tree32Leaf1_23_1 = tree8Leaf_6_7_1 & tree16Leaf2_15_1;
  wire        tree32Leaf1_23_2 = tree8Leaf_6_7_2 | tree8Leaf_6_7_1 & tree16Leaf2_15_2;
  wire        tree32Leaf1_24_1 = tree16Leaf3_8_1 & tree16Leaf2_15_1;
  wire        tree32Leaf1_24_2 = tree16Leaf3_8_2 | tree16Leaf3_8_1 & tree16Leaf2_15_2;
  wire        tree32Leaf1_25_1 = tree16Leaf3_9_1 & tree16Leaf2_15_1;
  wire        tree32Leaf1_25_2 = tree16Leaf3_9_2 | tree16Leaf3_9_1 & tree16Leaf2_15_2;
  wire        tree32Leaf1_26_1 = tree16Leaf3_10_1 & tree16Leaf2_15_1;
  wire        tree32Leaf1_26_2 = tree16Leaf3_10_2 | tree16Leaf3_10_1 & tree16Leaf2_15_2;
  wire        tree32Leaf1_27_1 = tree16Leaf3_11_1 & tree16Leaf2_15_1;
  wire        tree32Leaf1_27_2 = tree16Leaf3_11_2 | tree16Leaf3_11_1 & tree16Leaf2_15_2;
  wire        tree32Leaf1_28_1 = tree16Leaf3_12_1 & tree16Leaf2_15_1;
  wire        tree32Leaf1_28_2 = tree16Leaf3_12_2 | tree16Leaf3_12_1 & tree16Leaf2_15_2;
  wire        tree32Leaf1_29_1 = tree16Leaf3_13_1 & tree16Leaf2_15_1;
  wire        tree32Leaf1_29_2 = tree16Leaf3_13_2 | tree16Leaf3_13_1 & tree16Leaf2_15_2;
  wire        tree32Leaf1_30_1 = tree16Leaf3_14_1 & tree16Leaf2_15_1;
  wire        tree32Leaf1_30_2 = tree16Leaf3_14_2 | tree16Leaf3_14_1 & tree16Leaf2_15_2;
  wire        tree32Leaf1_31_1 = tree16Leaf3_15_1 & tree16Leaf2_15_1;
  wire        tree32Leaf1_31_2 = tree16Leaf3_15_2 | tree16Leaf3_15_1 & tree16Leaf2_15_2;
  wire        tree64_32_1 = pairs_32_1 & tree32Leaf0_31_1;
  wire        tree64_32_2 = pairs_32_2 | pairs_32_1 & tree32Leaf0_31_2;
  wire        tree64_33_1 = tree8Leaf_4_1_1 & tree32Leaf0_31_1;
  wire        tree64_33_2 = tree8Leaf_4_1_2 | tree8Leaf_4_1_1 & tree32Leaf0_31_2;
  wire        tree64_34_1 = tree8Leaf_4_2_1 & tree32Leaf0_31_1;
  wire        tree64_34_2 = tree8Leaf_4_2_2 | tree8Leaf_4_2_1 & tree32Leaf0_31_2;
  wire        tree64_35_1 = tree8Leaf_4_3_1 & tree32Leaf0_31_1;
  wire        tree64_35_2 = tree8Leaf_4_3_2 | tree8Leaf_4_3_1 & tree32Leaf0_31_2;
  wire        tree64_36_1 = tree8Leaf_4_4_1 & tree32Leaf0_31_1;
  wire        tree64_36_2 = tree8Leaf_4_4_2 | tree8Leaf_4_4_1 & tree32Leaf0_31_2;
  wire        tree64_37_1 = tree8Leaf_4_5_1 & tree32Leaf0_31_1;
  wire        tree64_37_2 = tree8Leaf_4_5_2 | tree8Leaf_4_5_1 & tree32Leaf0_31_2;
  wire        tree64_38_1 = tree8Leaf_4_6_1 & tree32Leaf0_31_1;
  wire        tree64_38_2 = tree8Leaf_4_6_2 | tree8Leaf_4_6_1 & tree32Leaf0_31_2;
  wire        tree64_39_1 = tree8Leaf_4_7_1 & tree32Leaf0_31_1;
  wire        tree64_39_2 = tree8Leaf_4_7_2 | tree8Leaf_4_7_1 & tree32Leaf0_31_2;
  wire        tree64_40_1 = tree16Leaf2_8_1 & tree32Leaf0_31_1;
  wire        tree64_40_2 = tree16Leaf2_8_2 | tree16Leaf2_8_1 & tree32Leaf0_31_2;
  wire        tree64_41_1 = tree16Leaf2_9_1 & tree32Leaf0_31_1;
  wire        tree64_41_2 = tree16Leaf2_9_2 | tree16Leaf2_9_1 & tree32Leaf0_31_2;
  wire        tree64_42_1 = tree16Leaf2_10_1 & tree32Leaf0_31_1;
  wire        tree64_42_2 = tree16Leaf2_10_2 | tree16Leaf2_10_1 & tree32Leaf0_31_2;
  wire        tree64_43_1 = tree16Leaf2_11_1 & tree32Leaf0_31_1;
  wire        tree64_43_2 = tree16Leaf2_11_2 | tree16Leaf2_11_1 & tree32Leaf0_31_2;
  wire        tree64_44_1 = tree16Leaf2_12_1 & tree32Leaf0_31_1;
  wire        tree64_44_2 = tree16Leaf2_12_2 | tree16Leaf2_12_1 & tree32Leaf0_31_2;
  wire        tree64_45_1 = tree16Leaf2_13_1 & tree32Leaf0_31_1;
  wire        tree64_45_2 = tree16Leaf2_13_2 | tree16Leaf2_13_1 & tree32Leaf0_31_2;
  wire        tree64_46_1 = tree16Leaf2_14_1 & tree32Leaf0_31_1;
  wire        tree64_46_2 = tree16Leaf2_14_2 | tree16Leaf2_14_1 & tree32Leaf0_31_2;
  wire        tree64_47_1 = tree16Leaf2_15_1 & tree32Leaf0_31_1;
  wire        tree64_47_2 = tree16Leaf2_15_2 | tree16Leaf2_15_1 & tree32Leaf0_31_2;
  wire        tree64_48_1 = tree32Leaf1_16_1 & tree32Leaf0_31_1;
  wire        tree64_48_2 = tree32Leaf1_16_2 | tree32Leaf1_16_1 & tree32Leaf0_31_2;
  wire        tree64_49_1 = tree32Leaf1_17_1 & tree32Leaf0_31_1;
  wire        tree64_49_2 = tree32Leaf1_17_2 | tree32Leaf1_17_1 & tree32Leaf0_31_2;
  wire        tree64_50_1 = tree32Leaf1_18_1 & tree32Leaf0_31_1;
  wire        tree64_50_2 = tree32Leaf1_18_2 | tree32Leaf1_18_1 & tree32Leaf0_31_2;
  wire        tree64_51_1 = tree32Leaf1_19_1 & tree32Leaf0_31_1;
  wire        tree64_51_2 = tree32Leaf1_19_2 | tree32Leaf1_19_1 & tree32Leaf0_31_2;
  wire        tree64_52_1 = tree32Leaf1_20_1 & tree32Leaf0_31_1;
  wire        tree64_52_2 = tree32Leaf1_20_2 | tree32Leaf1_20_1 & tree32Leaf0_31_2;
  wire        tree64_53_1 = tree32Leaf1_21_1 & tree32Leaf0_31_1;
  wire        tree64_53_2 = tree32Leaf1_21_2 | tree32Leaf1_21_1 & tree32Leaf0_31_2;
  wire        tree64_54_1 = tree32Leaf1_22_1 & tree32Leaf0_31_1;
  wire        tree64_54_2 = tree32Leaf1_22_2 | tree32Leaf1_22_1 & tree32Leaf0_31_2;
  wire        tree64_55_1 = tree32Leaf1_23_1 & tree32Leaf0_31_1;
  wire        tree64_55_2 = tree32Leaf1_23_2 | tree32Leaf1_23_1 & tree32Leaf0_31_2;
  wire        tree64_56_1 = tree32Leaf1_24_1 & tree32Leaf0_31_1;
  wire        tree64_56_2 = tree32Leaf1_24_2 | tree32Leaf1_24_1 & tree32Leaf0_31_2;
  wire        tree64_57_1 = tree32Leaf1_25_1 & tree32Leaf0_31_1;
  wire        tree64_57_2 = tree32Leaf1_25_2 | tree32Leaf1_25_1 & tree32Leaf0_31_2;
  wire        tree64_58_1 = tree32Leaf1_26_1 & tree32Leaf0_31_1;
  wire        tree64_58_2 = tree32Leaf1_26_2 | tree32Leaf1_26_1 & tree32Leaf0_31_2;
  wire        tree64_59_1 = tree32Leaf1_27_1 & tree32Leaf0_31_1;
  wire        tree64_59_2 = tree32Leaf1_27_2 | tree32Leaf1_27_1 & tree32Leaf0_31_2;
  wire        tree64_60_1 = tree32Leaf1_28_1 & tree32Leaf0_31_1;
  wire        tree64_60_2 = tree32Leaf1_28_2 | tree32Leaf1_28_1 & tree32Leaf0_31_2;
  wire        tree64_61_1 = tree32Leaf1_29_1 & tree32Leaf0_31_1;
  wire        tree64_61_2 = tree32Leaf1_29_2 | tree32Leaf1_29_1 & tree32Leaf0_31_2;
  wire        tree64_62_1 = tree32Leaf1_30_1 & tree32Leaf0_31_1;
  wire        tree64_62_2 = tree32Leaf1_30_2 | tree32Leaf1_30_1 & tree32Leaf0_31_2;
  wire        tree64_63_1 = tree32Leaf1_31_1 & tree32Leaf0_31_1;
  wire        tree64_63_2 = tree32Leaf1_31_2 | tree32Leaf1_31_1 & tree32Leaf0_31_2;
  wire [1:0]  _GEN = {tree8Leaf_0_1_1, pairs_0_1};
  wire [1:0]  tree8P_lo_lo_lo_lo_lo;
  assign tree8P_lo_lo_lo_lo_lo = _GEN;
  wire [1:0]  tree16P_lo_lo_lo_lo_lo;
  assign tree16P_lo_lo_lo_lo_lo = _GEN;
  wire [1:0]  tree32P_lo_lo_lo_lo_lo;
  assign tree32P_lo_lo_lo_lo_lo = _GEN;
  wire [1:0]  tree64P_lo_lo_lo_lo_lo;
  assign tree64P_lo_lo_lo_lo_lo = _GEN;
  wire [1:0]  _GEN_0 = {tree8Leaf_0_3_1, tree8Leaf_0_2_1};
  wire [1:0]  tree8P_lo_lo_lo_lo_hi;
  assign tree8P_lo_lo_lo_lo_hi = _GEN_0;
  wire [1:0]  tree16P_lo_lo_lo_lo_hi;
  assign tree16P_lo_lo_lo_lo_hi = _GEN_0;
  wire [1:0]  tree32P_lo_lo_lo_lo_hi;
  assign tree32P_lo_lo_lo_lo_hi = _GEN_0;
  wire [1:0]  tree64P_lo_lo_lo_lo_hi;
  assign tree64P_lo_lo_lo_lo_hi = _GEN_0;
  wire [3:0]  tree8P_lo_lo_lo_lo = {tree8P_lo_lo_lo_lo_hi, tree8P_lo_lo_lo_lo_lo};
  wire [1:0]  _GEN_1 = {tree8Leaf_0_5_1, tree8Leaf_0_4_1};
  wire [1:0]  tree8P_lo_lo_lo_hi_lo;
  assign tree8P_lo_lo_lo_hi_lo = _GEN_1;
  wire [1:0]  tree16P_lo_lo_lo_hi_lo;
  assign tree16P_lo_lo_lo_hi_lo = _GEN_1;
  wire [1:0]  tree32P_lo_lo_lo_hi_lo;
  assign tree32P_lo_lo_lo_hi_lo = _GEN_1;
  wire [1:0]  tree64P_lo_lo_lo_hi_lo;
  assign tree64P_lo_lo_lo_hi_lo = _GEN_1;
  wire [1:0]  _GEN_2 = {tree8Leaf_0_7_1, tree8Leaf_0_6_1};
  wire [1:0]  tree8P_lo_lo_lo_hi_hi;
  assign tree8P_lo_lo_lo_hi_hi = _GEN_2;
  wire [1:0]  tree16P_lo_lo_lo_hi_hi;
  assign tree16P_lo_lo_lo_hi_hi = _GEN_2;
  wire [1:0]  tree32P_lo_lo_lo_hi_hi;
  assign tree32P_lo_lo_lo_hi_hi = _GEN_2;
  wire [1:0]  tree64P_lo_lo_lo_hi_hi;
  assign tree64P_lo_lo_lo_hi_hi = _GEN_2;
  wire [3:0]  tree8P_lo_lo_lo_hi = {tree8P_lo_lo_lo_hi_hi, tree8P_lo_lo_lo_hi_lo};
  wire [7:0]  tree8P_lo_lo_lo = {tree8P_lo_lo_lo_hi, tree8P_lo_lo_lo_lo};
  wire [1:0]  tree8P_lo_lo_hi_lo_lo = {tree8Leaf_1_1_1, pairs_8_1};
  wire [1:0]  tree8P_lo_lo_hi_lo_hi = {tree8Leaf_1_3_1, tree8Leaf_1_2_1};
  wire [3:0]  tree8P_lo_lo_hi_lo = {tree8P_lo_lo_hi_lo_hi, tree8P_lo_lo_hi_lo_lo};
  wire [1:0]  tree8P_lo_lo_hi_hi_lo = {tree8Leaf_1_5_1, tree8Leaf_1_4_1};
  wire [1:0]  tree8P_lo_lo_hi_hi_hi = {tree8Leaf_1_7_1, tree8Leaf_1_6_1};
  wire [3:0]  tree8P_lo_lo_hi_hi = {tree8P_lo_lo_hi_hi_hi, tree8P_lo_lo_hi_hi_lo};
  wire [7:0]  tree8P_lo_lo_hi = {tree8P_lo_lo_hi_hi, tree8P_lo_lo_hi_lo};
  wire [15:0] tree8P_lo_lo = {tree8P_lo_lo_hi, tree8P_lo_lo_lo};
  wire [1:0]  _GEN_3 = {tree8Leaf_2_1_1, pairs_16_1};
  wire [1:0]  tree8P_lo_hi_lo_lo_lo;
  assign tree8P_lo_hi_lo_lo_lo = _GEN_3;
  wire [1:0]  tree16P_lo_hi_lo_lo_lo;
  assign tree16P_lo_hi_lo_lo_lo = _GEN_3;
  wire [1:0]  _GEN_4 = {tree8Leaf_2_3_1, tree8Leaf_2_2_1};
  wire [1:0]  tree8P_lo_hi_lo_lo_hi;
  assign tree8P_lo_hi_lo_lo_hi = _GEN_4;
  wire [1:0]  tree16P_lo_hi_lo_lo_hi;
  assign tree16P_lo_hi_lo_lo_hi = _GEN_4;
  wire [3:0]  tree8P_lo_hi_lo_lo = {tree8P_lo_hi_lo_lo_hi, tree8P_lo_hi_lo_lo_lo};
  wire [1:0]  _GEN_5 = {tree8Leaf_2_5_1, tree8Leaf_2_4_1};
  wire [1:0]  tree8P_lo_hi_lo_hi_lo;
  assign tree8P_lo_hi_lo_hi_lo = _GEN_5;
  wire [1:0]  tree16P_lo_hi_lo_hi_lo;
  assign tree16P_lo_hi_lo_hi_lo = _GEN_5;
  wire [1:0]  _GEN_6 = {tree8Leaf_2_7_1, tree8Leaf_2_6_1};
  wire [1:0]  tree8P_lo_hi_lo_hi_hi;
  assign tree8P_lo_hi_lo_hi_hi = _GEN_6;
  wire [1:0]  tree16P_lo_hi_lo_hi_hi;
  assign tree16P_lo_hi_lo_hi_hi = _GEN_6;
  wire [3:0]  tree8P_lo_hi_lo_hi = {tree8P_lo_hi_lo_hi_hi, tree8P_lo_hi_lo_hi_lo};
  wire [7:0]  tree8P_lo_hi_lo = {tree8P_lo_hi_lo_hi, tree8P_lo_hi_lo_lo};
  wire [1:0]  tree8P_lo_hi_hi_lo_lo = {tree8Leaf_3_1_1, pairs_24_1};
  wire [1:0]  tree8P_lo_hi_hi_lo_hi = {tree8Leaf_3_3_1, tree8Leaf_3_2_1};
  wire [3:0]  tree8P_lo_hi_hi_lo = {tree8P_lo_hi_hi_lo_hi, tree8P_lo_hi_hi_lo_lo};
  wire [1:0]  tree8P_lo_hi_hi_hi_lo = {tree8Leaf_3_5_1, tree8Leaf_3_4_1};
  wire [1:0]  tree8P_lo_hi_hi_hi_hi = {tree8Leaf_3_7_1, tree8Leaf_3_6_1};
  wire [3:0]  tree8P_lo_hi_hi_hi = {tree8P_lo_hi_hi_hi_hi, tree8P_lo_hi_hi_hi_lo};
  wire [7:0]  tree8P_lo_hi_hi = {tree8P_lo_hi_hi_hi, tree8P_lo_hi_hi_lo};
  wire [15:0] tree8P_lo_hi = {tree8P_lo_hi_hi, tree8P_lo_hi_lo};
  wire [31:0] tree8P_lo = {tree8P_lo_hi, tree8P_lo_lo};
  wire [1:0]  _GEN_7 = {tree8Leaf_4_1_1, pairs_32_1};
  wire [1:0]  tree8P_hi_lo_lo_lo_lo;
  assign tree8P_hi_lo_lo_lo_lo = _GEN_7;
  wire [1:0]  tree16P_hi_lo_lo_lo_lo;
  assign tree16P_hi_lo_lo_lo_lo = _GEN_7;
  wire [1:0]  tree32P_hi_lo_lo_lo_lo;
  assign tree32P_hi_lo_lo_lo_lo = _GEN_7;
  wire [1:0]  _GEN_8 = {tree8Leaf_4_3_1, tree8Leaf_4_2_1};
  wire [1:0]  tree8P_hi_lo_lo_lo_hi;
  assign tree8P_hi_lo_lo_lo_hi = _GEN_8;
  wire [1:0]  tree16P_hi_lo_lo_lo_hi;
  assign tree16P_hi_lo_lo_lo_hi = _GEN_8;
  wire [1:0]  tree32P_hi_lo_lo_lo_hi;
  assign tree32P_hi_lo_lo_lo_hi = _GEN_8;
  wire [3:0]  tree8P_hi_lo_lo_lo = {tree8P_hi_lo_lo_lo_hi, tree8P_hi_lo_lo_lo_lo};
  wire [1:0]  _GEN_9 = {tree8Leaf_4_5_1, tree8Leaf_4_4_1};
  wire [1:0]  tree8P_hi_lo_lo_hi_lo;
  assign tree8P_hi_lo_lo_hi_lo = _GEN_9;
  wire [1:0]  tree16P_hi_lo_lo_hi_lo;
  assign tree16P_hi_lo_lo_hi_lo = _GEN_9;
  wire [1:0]  tree32P_hi_lo_lo_hi_lo;
  assign tree32P_hi_lo_lo_hi_lo = _GEN_9;
  wire [1:0]  _GEN_10 = {tree8Leaf_4_7_1, tree8Leaf_4_6_1};
  wire [1:0]  tree8P_hi_lo_lo_hi_hi;
  assign tree8P_hi_lo_lo_hi_hi = _GEN_10;
  wire [1:0]  tree16P_hi_lo_lo_hi_hi;
  assign tree16P_hi_lo_lo_hi_hi = _GEN_10;
  wire [1:0]  tree32P_hi_lo_lo_hi_hi;
  assign tree32P_hi_lo_lo_hi_hi = _GEN_10;
  wire [3:0]  tree8P_hi_lo_lo_hi = {tree8P_hi_lo_lo_hi_hi, tree8P_hi_lo_lo_hi_lo};
  wire [7:0]  tree8P_hi_lo_lo = {tree8P_hi_lo_lo_hi, tree8P_hi_lo_lo_lo};
  wire [1:0]  tree8P_hi_lo_hi_lo_lo = {tree8Leaf_5_1_1, pairs_40_1};
  wire [1:0]  tree8P_hi_lo_hi_lo_hi = {tree8Leaf_5_3_1, tree8Leaf_5_2_1};
  wire [3:0]  tree8P_hi_lo_hi_lo = {tree8P_hi_lo_hi_lo_hi, tree8P_hi_lo_hi_lo_lo};
  wire [1:0]  tree8P_hi_lo_hi_hi_lo = {tree8Leaf_5_5_1, tree8Leaf_5_4_1};
  wire [1:0]  tree8P_hi_lo_hi_hi_hi = {tree8Leaf_5_7_1, tree8Leaf_5_6_1};
  wire [3:0]  tree8P_hi_lo_hi_hi = {tree8P_hi_lo_hi_hi_hi, tree8P_hi_lo_hi_hi_lo};
  wire [7:0]  tree8P_hi_lo_hi = {tree8P_hi_lo_hi_hi, tree8P_hi_lo_hi_lo};
  wire [15:0] tree8P_hi_lo = {tree8P_hi_lo_hi, tree8P_hi_lo_lo};
  wire [1:0]  _GEN_11 = {tree8Leaf_6_1_1, pairs_48_1};
  wire [1:0]  tree8P_hi_hi_lo_lo_lo;
  assign tree8P_hi_hi_lo_lo_lo = _GEN_11;
  wire [1:0]  tree16P_hi_hi_lo_lo_lo;
  assign tree16P_hi_hi_lo_lo_lo = _GEN_11;
  wire [1:0]  _GEN_12 = {tree8Leaf_6_3_1, tree8Leaf_6_2_1};
  wire [1:0]  tree8P_hi_hi_lo_lo_hi;
  assign tree8P_hi_hi_lo_lo_hi = _GEN_12;
  wire [1:0]  tree16P_hi_hi_lo_lo_hi;
  assign tree16P_hi_hi_lo_lo_hi = _GEN_12;
  wire [3:0]  tree8P_hi_hi_lo_lo = {tree8P_hi_hi_lo_lo_hi, tree8P_hi_hi_lo_lo_lo};
  wire [1:0]  _GEN_13 = {tree8Leaf_6_5_1, tree8Leaf_6_4_1};
  wire [1:0]  tree8P_hi_hi_lo_hi_lo;
  assign tree8P_hi_hi_lo_hi_lo = _GEN_13;
  wire [1:0]  tree16P_hi_hi_lo_hi_lo;
  assign tree16P_hi_hi_lo_hi_lo = _GEN_13;
  wire [1:0]  _GEN_14 = {tree8Leaf_6_7_1, tree8Leaf_6_6_1};
  wire [1:0]  tree8P_hi_hi_lo_hi_hi;
  assign tree8P_hi_hi_lo_hi_hi = _GEN_14;
  wire [1:0]  tree16P_hi_hi_lo_hi_hi;
  assign tree16P_hi_hi_lo_hi_hi = _GEN_14;
  wire [3:0]  tree8P_hi_hi_lo_hi = {tree8P_hi_hi_lo_hi_hi, tree8P_hi_hi_lo_hi_lo};
  wire [7:0]  tree8P_hi_hi_lo = {tree8P_hi_hi_lo_hi, tree8P_hi_hi_lo_lo};
  wire [1:0]  tree8P_hi_hi_hi_lo_lo = {tree8Leaf_7_1_1, pairs_56_1};
  wire [1:0]  tree8P_hi_hi_hi_lo_hi = {tree8Leaf_7_3_1, tree8Leaf_7_2_1};
  wire [3:0]  tree8P_hi_hi_hi_lo = {tree8P_hi_hi_hi_lo_hi, tree8P_hi_hi_hi_lo_lo};
  wire [1:0]  tree8P_hi_hi_hi_hi_lo = {tree8Leaf_7_5_1, tree8Leaf_7_4_1};
  wire [1:0]  tree8P_hi_hi_hi_hi_hi = {tree8Leaf_7_7_1, tree8Leaf_7_6_1};
  wire [3:0]  tree8P_hi_hi_hi_hi = {tree8P_hi_hi_hi_hi_hi, tree8P_hi_hi_hi_hi_lo};
  wire [7:0]  tree8P_hi_hi_hi = {tree8P_hi_hi_hi_hi, tree8P_hi_hi_hi_lo};
  wire [15:0] tree8P_hi_hi = {tree8P_hi_hi_hi, tree8P_hi_hi_lo};
  wire [31:0] tree8P_hi = {tree8P_hi_hi, tree8P_hi_lo};
  wire [63:0] tree8P = {tree8P_hi, tree8P_lo};
  wire [1:0]  _GEN_15 = {tree8Leaf_0_1_2, pairs_0_2};
  wire [1:0]  tree8G_lo_lo_lo_lo_lo;
  assign tree8G_lo_lo_lo_lo_lo = _GEN_15;
  wire [1:0]  tree16G_lo_lo_lo_lo_lo;
  assign tree16G_lo_lo_lo_lo_lo = _GEN_15;
  wire [1:0]  tree32G_lo_lo_lo_lo_lo;
  assign tree32G_lo_lo_lo_lo_lo = _GEN_15;
  wire [1:0]  tree64G_lo_lo_lo_lo_lo;
  assign tree64G_lo_lo_lo_lo_lo = _GEN_15;
  wire [1:0]  _GEN_16 = {tree8Leaf_0_3_2, tree8Leaf_0_2_2};
  wire [1:0]  tree8G_lo_lo_lo_lo_hi;
  assign tree8G_lo_lo_lo_lo_hi = _GEN_16;
  wire [1:0]  tree16G_lo_lo_lo_lo_hi;
  assign tree16G_lo_lo_lo_lo_hi = _GEN_16;
  wire [1:0]  tree32G_lo_lo_lo_lo_hi;
  assign tree32G_lo_lo_lo_lo_hi = _GEN_16;
  wire [1:0]  tree64G_lo_lo_lo_lo_hi;
  assign tree64G_lo_lo_lo_lo_hi = _GEN_16;
  wire [3:0]  tree8G_lo_lo_lo_lo = {tree8G_lo_lo_lo_lo_hi, tree8G_lo_lo_lo_lo_lo};
  wire [1:0]  _GEN_17 = {tree8Leaf_0_5_2, tree8Leaf_0_4_2};
  wire [1:0]  tree8G_lo_lo_lo_hi_lo;
  assign tree8G_lo_lo_lo_hi_lo = _GEN_17;
  wire [1:0]  tree16G_lo_lo_lo_hi_lo;
  assign tree16G_lo_lo_lo_hi_lo = _GEN_17;
  wire [1:0]  tree32G_lo_lo_lo_hi_lo;
  assign tree32G_lo_lo_lo_hi_lo = _GEN_17;
  wire [1:0]  tree64G_lo_lo_lo_hi_lo;
  assign tree64G_lo_lo_lo_hi_lo = _GEN_17;
  wire [1:0]  _GEN_18 = {tree8Leaf_0_7_2, tree8Leaf_0_6_2};
  wire [1:0]  tree8G_lo_lo_lo_hi_hi;
  assign tree8G_lo_lo_lo_hi_hi = _GEN_18;
  wire [1:0]  tree16G_lo_lo_lo_hi_hi;
  assign tree16G_lo_lo_lo_hi_hi = _GEN_18;
  wire [1:0]  tree32G_lo_lo_lo_hi_hi;
  assign tree32G_lo_lo_lo_hi_hi = _GEN_18;
  wire [1:0]  tree64G_lo_lo_lo_hi_hi;
  assign tree64G_lo_lo_lo_hi_hi = _GEN_18;
  wire [3:0]  tree8G_lo_lo_lo_hi = {tree8G_lo_lo_lo_hi_hi, tree8G_lo_lo_lo_hi_lo};
  wire [7:0]  tree8G_lo_lo_lo = {tree8G_lo_lo_lo_hi, tree8G_lo_lo_lo_lo};
  wire [1:0]  tree8G_lo_lo_hi_lo_lo = {tree8Leaf_1_1_2, pairs_8_2};
  wire [1:0]  tree8G_lo_lo_hi_lo_hi = {tree8Leaf_1_3_2, tree8Leaf_1_2_2};
  wire [3:0]  tree8G_lo_lo_hi_lo = {tree8G_lo_lo_hi_lo_hi, tree8G_lo_lo_hi_lo_lo};
  wire [1:0]  tree8G_lo_lo_hi_hi_lo = {tree8Leaf_1_5_2, tree8Leaf_1_4_2};
  wire [1:0]  tree8G_lo_lo_hi_hi_hi = {tree8Leaf_1_7_2, tree8Leaf_1_6_2};
  wire [3:0]  tree8G_lo_lo_hi_hi = {tree8G_lo_lo_hi_hi_hi, tree8G_lo_lo_hi_hi_lo};
  wire [7:0]  tree8G_lo_lo_hi = {tree8G_lo_lo_hi_hi, tree8G_lo_lo_hi_lo};
  wire [15:0] tree8G_lo_lo = {tree8G_lo_lo_hi, tree8G_lo_lo_lo};
  wire [1:0]  _GEN_19 = {tree8Leaf_2_1_2, pairs_16_2};
  wire [1:0]  tree8G_lo_hi_lo_lo_lo;
  assign tree8G_lo_hi_lo_lo_lo = _GEN_19;
  wire [1:0]  tree16G_lo_hi_lo_lo_lo;
  assign tree16G_lo_hi_lo_lo_lo = _GEN_19;
  wire [1:0]  _GEN_20 = {tree8Leaf_2_3_2, tree8Leaf_2_2_2};
  wire [1:0]  tree8G_lo_hi_lo_lo_hi;
  assign tree8G_lo_hi_lo_lo_hi = _GEN_20;
  wire [1:0]  tree16G_lo_hi_lo_lo_hi;
  assign tree16G_lo_hi_lo_lo_hi = _GEN_20;
  wire [3:0]  tree8G_lo_hi_lo_lo = {tree8G_lo_hi_lo_lo_hi, tree8G_lo_hi_lo_lo_lo};
  wire [1:0]  _GEN_21 = {tree8Leaf_2_5_2, tree8Leaf_2_4_2};
  wire [1:0]  tree8G_lo_hi_lo_hi_lo;
  assign tree8G_lo_hi_lo_hi_lo = _GEN_21;
  wire [1:0]  tree16G_lo_hi_lo_hi_lo;
  assign tree16G_lo_hi_lo_hi_lo = _GEN_21;
  wire [1:0]  _GEN_22 = {tree8Leaf_2_7_2, tree8Leaf_2_6_2};
  wire [1:0]  tree8G_lo_hi_lo_hi_hi;
  assign tree8G_lo_hi_lo_hi_hi = _GEN_22;
  wire [1:0]  tree16G_lo_hi_lo_hi_hi;
  assign tree16G_lo_hi_lo_hi_hi = _GEN_22;
  wire [3:0]  tree8G_lo_hi_lo_hi = {tree8G_lo_hi_lo_hi_hi, tree8G_lo_hi_lo_hi_lo};
  wire [7:0]  tree8G_lo_hi_lo = {tree8G_lo_hi_lo_hi, tree8G_lo_hi_lo_lo};
  wire [1:0]  tree8G_lo_hi_hi_lo_lo = {tree8Leaf_3_1_2, pairs_24_2};
  wire [1:0]  tree8G_lo_hi_hi_lo_hi = {tree8Leaf_3_3_2, tree8Leaf_3_2_2};
  wire [3:0]  tree8G_lo_hi_hi_lo = {tree8G_lo_hi_hi_lo_hi, tree8G_lo_hi_hi_lo_lo};
  wire [1:0]  tree8G_lo_hi_hi_hi_lo = {tree8Leaf_3_5_2, tree8Leaf_3_4_2};
  wire [1:0]  tree8G_lo_hi_hi_hi_hi = {tree8Leaf_3_7_2, tree8Leaf_3_6_2};
  wire [3:0]  tree8G_lo_hi_hi_hi = {tree8G_lo_hi_hi_hi_hi, tree8G_lo_hi_hi_hi_lo};
  wire [7:0]  tree8G_lo_hi_hi = {tree8G_lo_hi_hi_hi, tree8G_lo_hi_hi_lo};
  wire [15:0] tree8G_lo_hi = {tree8G_lo_hi_hi, tree8G_lo_hi_lo};
  wire [31:0] tree8G_lo = {tree8G_lo_hi, tree8G_lo_lo};
  wire [1:0]  _GEN_23 = {tree8Leaf_4_1_2, pairs_32_2};
  wire [1:0]  tree8G_hi_lo_lo_lo_lo;
  assign tree8G_hi_lo_lo_lo_lo = _GEN_23;
  wire [1:0]  tree16G_hi_lo_lo_lo_lo;
  assign tree16G_hi_lo_lo_lo_lo = _GEN_23;
  wire [1:0]  tree32G_hi_lo_lo_lo_lo;
  assign tree32G_hi_lo_lo_lo_lo = _GEN_23;
  wire [1:0]  _GEN_24 = {tree8Leaf_4_3_2, tree8Leaf_4_2_2};
  wire [1:0]  tree8G_hi_lo_lo_lo_hi;
  assign tree8G_hi_lo_lo_lo_hi = _GEN_24;
  wire [1:0]  tree16G_hi_lo_lo_lo_hi;
  assign tree16G_hi_lo_lo_lo_hi = _GEN_24;
  wire [1:0]  tree32G_hi_lo_lo_lo_hi;
  assign tree32G_hi_lo_lo_lo_hi = _GEN_24;
  wire [3:0]  tree8G_hi_lo_lo_lo = {tree8G_hi_lo_lo_lo_hi, tree8G_hi_lo_lo_lo_lo};
  wire [1:0]  _GEN_25 = {tree8Leaf_4_5_2, tree8Leaf_4_4_2};
  wire [1:0]  tree8G_hi_lo_lo_hi_lo;
  assign tree8G_hi_lo_lo_hi_lo = _GEN_25;
  wire [1:0]  tree16G_hi_lo_lo_hi_lo;
  assign tree16G_hi_lo_lo_hi_lo = _GEN_25;
  wire [1:0]  tree32G_hi_lo_lo_hi_lo;
  assign tree32G_hi_lo_lo_hi_lo = _GEN_25;
  wire [1:0]  _GEN_26 = {tree8Leaf_4_7_2, tree8Leaf_4_6_2};
  wire [1:0]  tree8G_hi_lo_lo_hi_hi;
  assign tree8G_hi_lo_lo_hi_hi = _GEN_26;
  wire [1:0]  tree16G_hi_lo_lo_hi_hi;
  assign tree16G_hi_lo_lo_hi_hi = _GEN_26;
  wire [1:0]  tree32G_hi_lo_lo_hi_hi;
  assign tree32G_hi_lo_lo_hi_hi = _GEN_26;
  wire [3:0]  tree8G_hi_lo_lo_hi = {tree8G_hi_lo_lo_hi_hi, tree8G_hi_lo_lo_hi_lo};
  wire [7:0]  tree8G_hi_lo_lo = {tree8G_hi_lo_lo_hi, tree8G_hi_lo_lo_lo};
  wire [1:0]  tree8G_hi_lo_hi_lo_lo = {tree8Leaf_5_1_2, pairs_40_2};
  wire [1:0]  tree8G_hi_lo_hi_lo_hi = {tree8Leaf_5_3_2, tree8Leaf_5_2_2};
  wire [3:0]  tree8G_hi_lo_hi_lo = {tree8G_hi_lo_hi_lo_hi, tree8G_hi_lo_hi_lo_lo};
  wire [1:0]  tree8G_hi_lo_hi_hi_lo = {tree8Leaf_5_5_2, tree8Leaf_5_4_2};
  wire [1:0]  tree8G_hi_lo_hi_hi_hi = {tree8Leaf_5_7_2, tree8Leaf_5_6_2};
  wire [3:0]  tree8G_hi_lo_hi_hi = {tree8G_hi_lo_hi_hi_hi, tree8G_hi_lo_hi_hi_lo};
  wire [7:0]  tree8G_hi_lo_hi = {tree8G_hi_lo_hi_hi, tree8G_hi_lo_hi_lo};
  wire [15:0] tree8G_hi_lo = {tree8G_hi_lo_hi, tree8G_hi_lo_lo};
  wire [1:0]  _GEN_27 = {tree8Leaf_6_1_2, pairs_48_2};
  wire [1:0]  tree8G_hi_hi_lo_lo_lo;
  assign tree8G_hi_hi_lo_lo_lo = _GEN_27;
  wire [1:0]  tree16G_hi_hi_lo_lo_lo;
  assign tree16G_hi_hi_lo_lo_lo = _GEN_27;
  wire [1:0]  _GEN_28 = {tree8Leaf_6_3_2, tree8Leaf_6_2_2};
  wire [1:0]  tree8G_hi_hi_lo_lo_hi;
  assign tree8G_hi_hi_lo_lo_hi = _GEN_28;
  wire [1:0]  tree16G_hi_hi_lo_lo_hi;
  assign tree16G_hi_hi_lo_lo_hi = _GEN_28;
  wire [3:0]  tree8G_hi_hi_lo_lo = {tree8G_hi_hi_lo_lo_hi, tree8G_hi_hi_lo_lo_lo};
  wire [1:0]  _GEN_29 = {tree8Leaf_6_5_2, tree8Leaf_6_4_2};
  wire [1:0]  tree8G_hi_hi_lo_hi_lo;
  assign tree8G_hi_hi_lo_hi_lo = _GEN_29;
  wire [1:0]  tree16G_hi_hi_lo_hi_lo;
  assign tree16G_hi_hi_lo_hi_lo = _GEN_29;
  wire [1:0]  _GEN_30 = {tree8Leaf_6_7_2, tree8Leaf_6_6_2};
  wire [1:0]  tree8G_hi_hi_lo_hi_hi;
  assign tree8G_hi_hi_lo_hi_hi = _GEN_30;
  wire [1:0]  tree16G_hi_hi_lo_hi_hi;
  assign tree16G_hi_hi_lo_hi_hi = _GEN_30;
  wire [3:0]  tree8G_hi_hi_lo_hi = {tree8G_hi_hi_lo_hi_hi, tree8G_hi_hi_lo_hi_lo};
  wire [7:0]  tree8G_hi_hi_lo = {tree8G_hi_hi_lo_hi, tree8G_hi_hi_lo_lo};
  wire [1:0]  tree8G_hi_hi_hi_lo_lo = {tree8Leaf_7_1_2, pairs_56_2};
  wire [1:0]  tree8G_hi_hi_hi_lo_hi = {tree8Leaf_7_3_2, tree8Leaf_7_2_2};
  wire [3:0]  tree8G_hi_hi_hi_lo = {tree8G_hi_hi_hi_lo_hi, tree8G_hi_hi_hi_lo_lo};
  wire [1:0]  tree8G_hi_hi_hi_hi_lo = {tree8Leaf_7_5_2, tree8Leaf_7_4_2};
  wire [1:0]  tree8G_hi_hi_hi_hi_hi = {tree8Leaf_7_7_2, tree8Leaf_7_6_2};
  wire [3:0]  tree8G_hi_hi_hi_hi = {tree8G_hi_hi_hi_hi_hi, tree8G_hi_hi_hi_hi_lo};
  wire [7:0]  tree8G_hi_hi_hi = {tree8G_hi_hi_hi_hi, tree8G_hi_hi_hi_lo};
  wire [15:0] tree8G_hi_hi = {tree8G_hi_hi_hi, tree8G_hi_hi_lo};
  wire [31:0] tree8G_hi = {tree8G_hi_hi, tree8G_hi_lo};
  wire [63:0] tree8G = {tree8G_hi, tree8G_lo};
  wire [3:0]  tree16P_lo_lo_lo_lo = {tree16P_lo_lo_lo_lo_hi, tree16P_lo_lo_lo_lo_lo};
  wire [3:0]  tree16P_lo_lo_lo_hi = {tree16P_lo_lo_lo_hi_hi, tree16P_lo_lo_lo_hi_lo};
  wire [7:0]  tree16P_lo_lo_lo = {tree16P_lo_lo_lo_hi, tree16P_lo_lo_lo_lo};
  wire [1:0]  _GEN_31 = {tree16Leaf0_9_1, tree16Leaf0_8_1};
  wire [1:0]  tree16P_lo_lo_hi_lo_lo;
  assign tree16P_lo_lo_hi_lo_lo = _GEN_31;
  wire [1:0]  tree32P_lo_lo_hi_lo_lo;
  assign tree32P_lo_lo_hi_lo_lo = _GEN_31;
  wire [1:0]  tree64P_lo_lo_hi_lo_lo;
  assign tree64P_lo_lo_hi_lo_lo = _GEN_31;
  wire [1:0]  _GEN_32 = {tree16Leaf0_11_1, tree16Leaf0_10_1};
  wire [1:0]  tree16P_lo_lo_hi_lo_hi;
  assign tree16P_lo_lo_hi_lo_hi = _GEN_32;
  wire [1:0]  tree32P_lo_lo_hi_lo_hi;
  assign tree32P_lo_lo_hi_lo_hi = _GEN_32;
  wire [1:0]  tree64P_lo_lo_hi_lo_hi;
  assign tree64P_lo_lo_hi_lo_hi = _GEN_32;
  wire [3:0]  tree16P_lo_lo_hi_lo = {tree16P_lo_lo_hi_lo_hi, tree16P_lo_lo_hi_lo_lo};
  wire [1:0]  _GEN_33 = {tree16Leaf0_13_1, tree16Leaf0_12_1};
  wire [1:0]  tree16P_lo_lo_hi_hi_lo;
  assign tree16P_lo_lo_hi_hi_lo = _GEN_33;
  wire [1:0]  tree32P_lo_lo_hi_hi_lo;
  assign tree32P_lo_lo_hi_hi_lo = _GEN_33;
  wire [1:0]  tree64P_lo_lo_hi_hi_lo;
  assign tree64P_lo_lo_hi_hi_lo = _GEN_33;
  wire [1:0]  _GEN_34 = {tree16Leaf0_15_1, tree16Leaf0_14_1};
  wire [1:0]  tree16P_lo_lo_hi_hi_hi;
  assign tree16P_lo_lo_hi_hi_hi = _GEN_34;
  wire [1:0]  tree32P_lo_lo_hi_hi_hi;
  assign tree32P_lo_lo_hi_hi_hi = _GEN_34;
  wire [1:0]  tree64P_lo_lo_hi_hi_hi;
  assign tree64P_lo_lo_hi_hi_hi = _GEN_34;
  wire [3:0]  tree16P_lo_lo_hi_hi = {tree16P_lo_lo_hi_hi_hi, tree16P_lo_lo_hi_hi_lo};
  wire [7:0]  tree16P_lo_lo_hi = {tree16P_lo_lo_hi_hi, tree16P_lo_lo_hi_lo};
  wire [15:0] tree16P_lo_lo = {tree16P_lo_lo_hi, tree16P_lo_lo_lo};
  wire [3:0]  tree16P_lo_hi_lo_lo = {tree16P_lo_hi_lo_lo_hi, tree16P_lo_hi_lo_lo_lo};
  wire [3:0]  tree16P_lo_hi_lo_hi = {tree16P_lo_hi_lo_hi_hi, tree16P_lo_hi_lo_hi_lo};
  wire [7:0]  tree16P_lo_hi_lo = {tree16P_lo_hi_lo_hi, tree16P_lo_hi_lo_lo};
  wire [1:0]  tree16P_lo_hi_hi_lo_lo = {tree16Leaf1_9_1, tree16Leaf1_8_1};
  wire [1:0]  tree16P_lo_hi_hi_lo_hi = {tree16Leaf1_11_1, tree16Leaf1_10_1};
  wire [3:0]  tree16P_lo_hi_hi_lo = {tree16P_lo_hi_hi_lo_hi, tree16P_lo_hi_hi_lo_lo};
  wire [1:0]  tree16P_lo_hi_hi_hi_lo = {tree16Leaf1_13_1, tree16Leaf1_12_1};
  wire [1:0]  tree16P_lo_hi_hi_hi_hi = {tree16Leaf1_15_1, tree16Leaf1_14_1};
  wire [3:0]  tree16P_lo_hi_hi_hi = {tree16P_lo_hi_hi_hi_hi, tree16P_lo_hi_hi_hi_lo};
  wire [7:0]  tree16P_lo_hi_hi = {tree16P_lo_hi_hi_hi, tree16P_lo_hi_hi_lo};
  wire [15:0] tree16P_lo_hi = {tree16P_lo_hi_hi, tree16P_lo_hi_lo};
  wire [31:0] tree16P_lo = {tree16P_lo_hi, tree16P_lo_lo};
  wire [3:0]  tree16P_hi_lo_lo_lo = {tree16P_hi_lo_lo_lo_hi, tree16P_hi_lo_lo_lo_lo};
  wire [3:0]  tree16P_hi_lo_lo_hi = {tree16P_hi_lo_lo_hi_hi, tree16P_hi_lo_lo_hi_lo};
  wire [7:0]  tree16P_hi_lo_lo = {tree16P_hi_lo_lo_hi, tree16P_hi_lo_lo_lo};
  wire [1:0]  _GEN_35 = {tree16Leaf2_9_1, tree16Leaf2_8_1};
  wire [1:0]  tree16P_hi_lo_hi_lo_lo;
  assign tree16P_hi_lo_hi_lo_lo = _GEN_35;
  wire [1:0]  tree32P_hi_lo_hi_lo_lo;
  assign tree32P_hi_lo_hi_lo_lo = _GEN_35;
  wire [1:0]  _GEN_36 = {tree16Leaf2_11_1, tree16Leaf2_10_1};
  wire [1:0]  tree16P_hi_lo_hi_lo_hi;
  assign tree16P_hi_lo_hi_lo_hi = _GEN_36;
  wire [1:0]  tree32P_hi_lo_hi_lo_hi;
  assign tree32P_hi_lo_hi_lo_hi = _GEN_36;
  wire [3:0]  tree16P_hi_lo_hi_lo = {tree16P_hi_lo_hi_lo_hi, tree16P_hi_lo_hi_lo_lo};
  wire [1:0]  _GEN_37 = {tree16Leaf2_13_1, tree16Leaf2_12_1};
  wire [1:0]  tree16P_hi_lo_hi_hi_lo;
  assign tree16P_hi_lo_hi_hi_lo = _GEN_37;
  wire [1:0]  tree32P_hi_lo_hi_hi_lo;
  assign tree32P_hi_lo_hi_hi_lo = _GEN_37;
  wire [1:0]  _GEN_38 = {tree16Leaf2_15_1, tree16Leaf2_14_1};
  wire [1:0]  tree16P_hi_lo_hi_hi_hi;
  assign tree16P_hi_lo_hi_hi_hi = _GEN_38;
  wire [1:0]  tree32P_hi_lo_hi_hi_hi;
  assign tree32P_hi_lo_hi_hi_hi = _GEN_38;
  wire [3:0]  tree16P_hi_lo_hi_hi = {tree16P_hi_lo_hi_hi_hi, tree16P_hi_lo_hi_hi_lo};
  wire [7:0]  tree16P_hi_lo_hi = {tree16P_hi_lo_hi_hi, tree16P_hi_lo_hi_lo};
  wire [15:0] tree16P_hi_lo = {tree16P_hi_lo_hi, tree16P_hi_lo_lo};
  wire [3:0]  tree16P_hi_hi_lo_lo = {tree16P_hi_hi_lo_lo_hi, tree16P_hi_hi_lo_lo_lo};
  wire [3:0]  tree16P_hi_hi_lo_hi = {tree16P_hi_hi_lo_hi_hi, tree16P_hi_hi_lo_hi_lo};
  wire [7:0]  tree16P_hi_hi_lo = {tree16P_hi_hi_lo_hi, tree16P_hi_hi_lo_lo};
  wire [1:0]  tree16P_hi_hi_hi_lo_lo = {tree16Leaf3_9_1, tree16Leaf3_8_1};
  wire [1:0]  tree16P_hi_hi_hi_lo_hi = {tree16Leaf3_11_1, tree16Leaf3_10_1};
  wire [3:0]  tree16P_hi_hi_hi_lo = {tree16P_hi_hi_hi_lo_hi, tree16P_hi_hi_hi_lo_lo};
  wire [1:0]  tree16P_hi_hi_hi_hi_lo = {tree16Leaf3_13_1, tree16Leaf3_12_1};
  wire [1:0]  tree16P_hi_hi_hi_hi_hi = {tree16Leaf3_15_1, tree16Leaf3_14_1};
  wire [3:0]  tree16P_hi_hi_hi_hi = {tree16P_hi_hi_hi_hi_hi, tree16P_hi_hi_hi_hi_lo};
  wire [7:0]  tree16P_hi_hi_hi = {tree16P_hi_hi_hi_hi, tree16P_hi_hi_hi_lo};
  wire [15:0] tree16P_hi_hi = {tree16P_hi_hi_hi, tree16P_hi_hi_lo};
  wire [31:0] tree16P_hi = {tree16P_hi_hi, tree16P_hi_lo};
  wire [63:0] tree16P = {tree16P_hi, tree16P_lo};
  wire [3:0]  tree16G_lo_lo_lo_lo = {tree16G_lo_lo_lo_lo_hi, tree16G_lo_lo_lo_lo_lo};
  wire [3:0]  tree16G_lo_lo_lo_hi = {tree16G_lo_lo_lo_hi_hi, tree16G_lo_lo_lo_hi_lo};
  wire [7:0]  tree16G_lo_lo_lo = {tree16G_lo_lo_lo_hi, tree16G_lo_lo_lo_lo};
  wire [1:0]  _GEN_39 = {tree16Leaf0_9_2, tree16Leaf0_8_2};
  wire [1:0]  tree16G_lo_lo_hi_lo_lo;
  assign tree16G_lo_lo_hi_lo_lo = _GEN_39;
  wire [1:0]  tree32G_lo_lo_hi_lo_lo;
  assign tree32G_lo_lo_hi_lo_lo = _GEN_39;
  wire [1:0]  tree64G_lo_lo_hi_lo_lo;
  assign tree64G_lo_lo_hi_lo_lo = _GEN_39;
  wire [1:0]  _GEN_40 = {tree16Leaf0_11_2, tree16Leaf0_10_2};
  wire [1:0]  tree16G_lo_lo_hi_lo_hi;
  assign tree16G_lo_lo_hi_lo_hi = _GEN_40;
  wire [1:0]  tree32G_lo_lo_hi_lo_hi;
  assign tree32G_lo_lo_hi_lo_hi = _GEN_40;
  wire [1:0]  tree64G_lo_lo_hi_lo_hi;
  assign tree64G_lo_lo_hi_lo_hi = _GEN_40;
  wire [3:0]  tree16G_lo_lo_hi_lo = {tree16G_lo_lo_hi_lo_hi, tree16G_lo_lo_hi_lo_lo};
  wire [1:0]  _GEN_41 = {tree16Leaf0_13_2, tree16Leaf0_12_2};
  wire [1:0]  tree16G_lo_lo_hi_hi_lo;
  assign tree16G_lo_lo_hi_hi_lo = _GEN_41;
  wire [1:0]  tree32G_lo_lo_hi_hi_lo;
  assign tree32G_lo_lo_hi_hi_lo = _GEN_41;
  wire [1:0]  tree64G_lo_lo_hi_hi_lo;
  assign tree64G_lo_lo_hi_hi_lo = _GEN_41;
  wire [1:0]  _GEN_42 = {tree16Leaf0_15_2, tree16Leaf0_14_2};
  wire [1:0]  tree16G_lo_lo_hi_hi_hi;
  assign tree16G_lo_lo_hi_hi_hi = _GEN_42;
  wire [1:0]  tree32G_lo_lo_hi_hi_hi;
  assign tree32G_lo_lo_hi_hi_hi = _GEN_42;
  wire [1:0]  tree64G_lo_lo_hi_hi_hi;
  assign tree64G_lo_lo_hi_hi_hi = _GEN_42;
  wire [3:0]  tree16G_lo_lo_hi_hi = {tree16G_lo_lo_hi_hi_hi, tree16G_lo_lo_hi_hi_lo};
  wire [7:0]  tree16G_lo_lo_hi = {tree16G_lo_lo_hi_hi, tree16G_lo_lo_hi_lo};
  wire [15:0] tree16G_lo_lo = {tree16G_lo_lo_hi, tree16G_lo_lo_lo};
  wire [3:0]  tree16G_lo_hi_lo_lo = {tree16G_lo_hi_lo_lo_hi, tree16G_lo_hi_lo_lo_lo};
  wire [3:0]  tree16G_lo_hi_lo_hi = {tree16G_lo_hi_lo_hi_hi, tree16G_lo_hi_lo_hi_lo};
  wire [7:0]  tree16G_lo_hi_lo = {tree16G_lo_hi_lo_hi, tree16G_lo_hi_lo_lo};
  wire [1:0]  tree16G_lo_hi_hi_lo_lo = {tree16Leaf1_9_2, tree16Leaf1_8_2};
  wire [1:0]  tree16G_lo_hi_hi_lo_hi = {tree16Leaf1_11_2, tree16Leaf1_10_2};
  wire [3:0]  tree16G_lo_hi_hi_lo = {tree16G_lo_hi_hi_lo_hi, tree16G_lo_hi_hi_lo_lo};
  wire [1:0]  tree16G_lo_hi_hi_hi_lo = {tree16Leaf1_13_2, tree16Leaf1_12_2};
  wire [1:0]  tree16G_lo_hi_hi_hi_hi = {tree16Leaf1_15_2, tree16Leaf1_14_2};
  wire [3:0]  tree16G_lo_hi_hi_hi = {tree16G_lo_hi_hi_hi_hi, tree16G_lo_hi_hi_hi_lo};
  wire [7:0]  tree16G_lo_hi_hi = {tree16G_lo_hi_hi_hi, tree16G_lo_hi_hi_lo};
  wire [15:0] tree16G_lo_hi = {tree16G_lo_hi_hi, tree16G_lo_hi_lo};
  wire [31:0] tree16G_lo = {tree16G_lo_hi, tree16G_lo_lo};
  wire [3:0]  tree16G_hi_lo_lo_lo = {tree16G_hi_lo_lo_lo_hi, tree16G_hi_lo_lo_lo_lo};
  wire [3:0]  tree16G_hi_lo_lo_hi = {tree16G_hi_lo_lo_hi_hi, tree16G_hi_lo_lo_hi_lo};
  wire [7:0]  tree16G_hi_lo_lo = {tree16G_hi_lo_lo_hi, tree16G_hi_lo_lo_lo};
  wire [1:0]  _GEN_43 = {tree16Leaf2_9_2, tree16Leaf2_8_2};
  wire [1:0]  tree16G_hi_lo_hi_lo_lo;
  assign tree16G_hi_lo_hi_lo_lo = _GEN_43;
  wire [1:0]  tree32G_hi_lo_hi_lo_lo;
  assign tree32G_hi_lo_hi_lo_lo = _GEN_43;
  wire [1:0]  _GEN_44 = {tree16Leaf2_11_2, tree16Leaf2_10_2};
  wire [1:0]  tree16G_hi_lo_hi_lo_hi;
  assign tree16G_hi_lo_hi_lo_hi = _GEN_44;
  wire [1:0]  tree32G_hi_lo_hi_lo_hi;
  assign tree32G_hi_lo_hi_lo_hi = _GEN_44;
  wire [3:0]  tree16G_hi_lo_hi_lo = {tree16G_hi_lo_hi_lo_hi, tree16G_hi_lo_hi_lo_lo};
  wire [1:0]  _GEN_45 = {tree16Leaf2_13_2, tree16Leaf2_12_2};
  wire [1:0]  tree16G_hi_lo_hi_hi_lo;
  assign tree16G_hi_lo_hi_hi_lo = _GEN_45;
  wire [1:0]  tree32G_hi_lo_hi_hi_lo;
  assign tree32G_hi_lo_hi_hi_lo = _GEN_45;
  wire [1:0]  _GEN_46 = {tree16Leaf2_15_2, tree16Leaf2_14_2};
  wire [1:0]  tree16G_hi_lo_hi_hi_hi;
  assign tree16G_hi_lo_hi_hi_hi = _GEN_46;
  wire [1:0]  tree32G_hi_lo_hi_hi_hi;
  assign tree32G_hi_lo_hi_hi_hi = _GEN_46;
  wire [3:0]  tree16G_hi_lo_hi_hi = {tree16G_hi_lo_hi_hi_hi, tree16G_hi_lo_hi_hi_lo};
  wire [7:0]  tree16G_hi_lo_hi = {tree16G_hi_lo_hi_hi, tree16G_hi_lo_hi_lo};
  wire [15:0] tree16G_hi_lo = {tree16G_hi_lo_hi, tree16G_hi_lo_lo};
  wire [3:0]  tree16G_hi_hi_lo_lo = {tree16G_hi_hi_lo_lo_hi, tree16G_hi_hi_lo_lo_lo};
  wire [3:0]  tree16G_hi_hi_lo_hi = {tree16G_hi_hi_lo_hi_hi, tree16G_hi_hi_lo_hi_lo};
  wire [7:0]  tree16G_hi_hi_lo = {tree16G_hi_hi_lo_hi, tree16G_hi_hi_lo_lo};
  wire [1:0]  tree16G_hi_hi_hi_lo_lo = {tree16Leaf3_9_2, tree16Leaf3_8_2};
  wire [1:0]  tree16G_hi_hi_hi_lo_hi = {tree16Leaf3_11_2, tree16Leaf3_10_2};
  wire [3:0]  tree16G_hi_hi_hi_lo = {tree16G_hi_hi_hi_lo_hi, tree16G_hi_hi_hi_lo_lo};
  wire [1:0]  tree16G_hi_hi_hi_hi_lo = {tree16Leaf3_13_2, tree16Leaf3_12_2};
  wire [1:0]  tree16G_hi_hi_hi_hi_hi = {tree16Leaf3_15_2, tree16Leaf3_14_2};
  wire [3:0]  tree16G_hi_hi_hi_hi = {tree16G_hi_hi_hi_hi_hi, tree16G_hi_hi_hi_hi_lo};
  wire [7:0]  tree16G_hi_hi_hi = {tree16G_hi_hi_hi_hi, tree16G_hi_hi_hi_lo};
  wire [15:0] tree16G_hi_hi = {tree16G_hi_hi_hi, tree16G_hi_hi_lo};
  wire [31:0] tree16G_hi = {tree16G_hi_hi, tree16G_hi_lo};
  wire [63:0] tree16G = {tree16G_hi, tree16G_lo};
  wire [3:0]  tree32P_lo_lo_lo_lo = {tree32P_lo_lo_lo_lo_hi, tree32P_lo_lo_lo_lo_lo};
  wire [3:0]  tree32P_lo_lo_lo_hi = {tree32P_lo_lo_lo_hi_hi, tree32P_lo_lo_lo_hi_lo};
  wire [7:0]  tree32P_lo_lo_lo = {tree32P_lo_lo_lo_hi, tree32P_lo_lo_lo_lo};
  wire [3:0]  tree32P_lo_lo_hi_lo = {tree32P_lo_lo_hi_lo_hi, tree32P_lo_lo_hi_lo_lo};
  wire [3:0]  tree32P_lo_lo_hi_hi = {tree32P_lo_lo_hi_hi_hi, tree32P_lo_lo_hi_hi_lo};
  wire [7:0]  tree32P_lo_lo_hi = {tree32P_lo_lo_hi_hi, tree32P_lo_lo_hi_lo};
  wire [15:0] tree32P_lo_lo = {tree32P_lo_lo_hi, tree32P_lo_lo_lo};
  wire [1:0]  _GEN_47 = {tree32Leaf0_17_1, tree32Leaf0_16_1};
  wire [1:0]  tree32P_lo_hi_lo_lo_lo;
  assign tree32P_lo_hi_lo_lo_lo = _GEN_47;
  wire [1:0]  tree64P_lo_hi_lo_lo_lo;
  assign tree64P_lo_hi_lo_lo_lo = _GEN_47;
  wire [1:0]  _GEN_48 = {tree32Leaf0_19_1, tree32Leaf0_18_1};
  wire [1:0]  tree32P_lo_hi_lo_lo_hi;
  assign tree32P_lo_hi_lo_lo_hi = _GEN_48;
  wire [1:0]  tree64P_lo_hi_lo_lo_hi;
  assign tree64P_lo_hi_lo_lo_hi = _GEN_48;
  wire [3:0]  tree32P_lo_hi_lo_lo = {tree32P_lo_hi_lo_lo_hi, tree32P_lo_hi_lo_lo_lo};
  wire [1:0]  _GEN_49 = {tree32Leaf0_21_1, tree32Leaf0_20_1};
  wire [1:0]  tree32P_lo_hi_lo_hi_lo;
  assign tree32P_lo_hi_lo_hi_lo = _GEN_49;
  wire [1:0]  tree64P_lo_hi_lo_hi_lo;
  assign tree64P_lo_hi_lo_hi_lo = _GEN_49;
  wire [1:0]  _GEN_50 = {tree32Leaf0_23_1, tree32Leaf0_22_1};
  wire [1:0]  tree32P_lo_hi_lo_hi_hi;
  assign tree32P_lo_hi_lo_hi_hi = _GEN_50;
  wire [1:0]  tree64P_lo_hi_lo_hi_hi;
  assign tree64P_lo_hi_lo_hi_hi = _GEN_50;
  wire [3:0]  tree32P_lo_hi_lo_hi = {tree32P_lo_hi_lo_hi_hi, tree32P_lo_hi_lo_hi_lo};
  wire [7:0]  tree32P_lo_hi_lo = {tree32P_lo_hi_lo_hi, tree32P_lo_hi_lo_lo};
  wire [1:0]  _GEN_51 = {tree32Leaf0_25_1, tree32Leaf0_24_1};
  wire [1:0]  tree32P_lo_hi_hi_lo_lo;
  assign tree32P_lo_hi_hi_lo_lo = _GEN_51;
  wire [1:0]  tree64P_lo_hi_hi_lo_lo;
  assign tree64P_lo_hi_hi_lo_lo = _GEN_51;
  wire [1:0]  _GEN_52 = {tree32Leaf0_27_1, tree32Leaf0_26_1};
  wire [1:0]  tree32P_lo_hi_hi_lo_hi;
  assign tree32P_lo_hi_hi_lo_hi = _GEN_52;
  wire [1:0]  tree64P_lo_hi_hi_lo_hi;
  assign tree64P_lo_hi_hi_lo_hi = _GEN_52;
  wire [3:0]  tree32P_lo_hi_hi_lo = {tree32P_lo_hi_hi_lo_hi, tree32P_lo_hi_hi_lo_lo};
  wire [1:0]  _GEN_53 = {tree32Leaf0_29_1, tree32Leaf0_28_1};
  wire [1:0]  tree32P_lo_hi_hi_hi_lo;
  assign tree32P_lo_hi_hi_hi_lo = _GEN_53;
  wire [1:0]  tree64P_lo_hi_hi_hi_lo;
  assign tree64P_lo_hi_hi_hi_lo = _GEN_53;
  wire [1:0]  _GEN_54 = {tree32Leaf0_31_1, tree32Leaf0_30_1};
  wire [1:0]  tree32P_lo_hi_hi_hi_hi;
  assign tree32P_lo_hi_hi_hi_hi = _GEN_54;
  wire [1:0]  tree64P_lo_hi_hi_hi_hi;
  assign tree64P_lo_hi_hi_hi_hi = _GEN_54;
  wire [3:0]  tree32P_lo_hi_hi_hi = {tree32P_lo_hi_hi_hi_hi, tree32P_lo_hi_hi_hi_lo};
  wire [7:0]  tree32P_lo_hi_hi = {tree32P_lo_hi_hi_hi, tree32P_lo_hi_hi_lo};
  wire [15:0] tree32P_lo_hi = {tree32P_lo_hi_hi, tree32P_lo_hi_lo};
  wire [31:0] tree32P_lo = {tree32P_lo_hi, tree32P_lo_lo};
  wire [3:0]  tree32P_hi_lo_lo_lo = {tree32P_hi_lo_lo_lo_hi, tree32P_hi_lo_lo_lo_lo};
  wire [3:0]  tree32P_hi_lo_lo_hi = {tree32P_hi_lo_lo_hi_hi, tree32P_hi_lo_lo_hi_lo};
  wire [7:0]  tree32P_hi_lo_lo = {tree32P_hi_lo_lo_hi, tree32P_hi_lo_lo_lo};
  wire [3:0]  tree32P_hi_lo_hi_lo = {tree32P_hi_lo_hi_lo_hi, tree32P_hi_lo_hi_lo_lo};
  wire [3:0]  tree32P_hi_lo_hi_hi = {tree32P_hi_lo_hi_hi_hi, tree32P_hi_lo_hi_hi_lo};
  wire [7:0]  tree32P_hi_lo_hi = {tree32P_hi_lo_hi_hi, tree32P_hi_lo_hi_lo};
  wire [15:0] tree32P_hi_lo = {tree32P_hi_lo_hi, tree32P_hi_lo_lo};
  wire [1:0]  tree32P_hi_hi_lo_lo_lo = {tree32Leaf1_17_1, tree32Leaf1_16_1};
  wire [1:0]  tree32P_hi_hi_lo_lo_hi = {tree32Leaf1_19_1, tree32Leaf1_18_1};
  wire [3:0]  tree32P_hi_hi_lo_lo = {tree32P_hi_hi_lo_lo_hi, tree32P_hi_hi_lo_lo_lo};
  wire [1:0]  tree32P_hi_hi_lo_hi_lo = {tree32Leaf1_21_1, tree32Leaf1_20_1};
  wire [1:0]  tree32P_hi_hi_lo_hi_hi = {tree32Leaf1_23_1, tree32Leaf1_22_1};
  wire [3:0]  tree32P_hi_hi_lo_hi = {tree32P_hi_hi_lo_hi_hi, tree32P_hi_hi_lo_hi_lo};
  wire [7:0]  tree32P_hi_hi_lo = {tree32P_hi_hi_lo_hi, tree32P_hi_hi_lo_lo};
  wire [1:0]  tree32P_hi_hi_hi_lo_lo = {tree32Leaf1_25_1, tree32Leaf1_24_1};
  wire [1:0]  tree32P_hi_hi_hi_lo_hi = {tree32Leaf1_27_1, tree32Leaf1_26_1};
  wire [3:0]  tree32P_hi_hi_hi_lo = {tree32P_hi_hi_hi_lo_hi, tree32P_hi_hi_hi_lo_lo};
  wire [1:0]  tree32P_hi_hi_hi_hi_lo = {tree32Leaf1_29_1, tree32Leaf1_28_1};
  wire [1:0]  tree32P_hi_hi_hi_hi_hi = {tree32Leaf1_31_1, tree32Leaf1_30_1};
  wire [3:0]  tree32P_hi_hi_hi_hi = {tree32P_hi_hi_hi_hi_hi, tree32P_hi_hi_hi_hi_lo};
  wire [7:0]  tree32P_hi_hi_hi = {tree32P_hi_hi_hi_hi, tree32P_hi_hi_hi_lo};
  wire [15:0] tree32P_hi_hi = {tree32P_hi_hi_hi, tree32P_hi_hi_lo};
  wire [31:0] tree32P_hi = {tree32P_hi_hi, tree32P_hi_lo};
  wire [63:0] tree32P = {tree32P_hi, tree32P_lo};
  wire [3:0]  tree32G_lo_lo_lo_lo = {tree32G_lo_lo_lo_lo_hi, tree32G_lo_lo_lo_lo_lo};
  wire [3:0]  tree32G_lo_lo_lo_hi = {tree32G_lo_lo_lo_hi_hi, tree32G_lo_lo_lo_hi_lo};
  wire [7:0]  tree32G_lo_lo_lo = {tree32G_lo_lo_lo_hi, tree32G_lo_lo_lo_lo};
  wire [3:0]  tree32G_lo_lo_hi_lo = {tree32G_lo_lo_hi_lo_hi, tree32G_lo_lo_hi_lo_lo};
  wire [3:0]  tree32G_lo_lo_hi_hi = {tree32G_lo_lo_hi_hi_hi, tree32G_lo_lo_hi_hi_lo};
  wire [7:0]  tree32G_lo_lo_hi = {tree32G_lo_lo_hi_hi, tree32G_lo_lo_hi_lo};
  wire [15:0] tree32G_lo_lo = {tree32G_lo_lo_hi, tree32G_lo_lo_lo};
  wire [1:0]  _GEN_55 = {tree32Leaf0_17_2, tree32Leaf0_16_2};
  wire [1:0]  tree32G_lo_hi_lo_lo_lo;
  assign tree32G_lo_hi_lo_lo_lo = _GEN_55;
  wire [1:0]  tree64G_lo_hi_lo_lo_lo;
  assign tree64G_lo_hi_lo_lo_lo = _GEN_55;
  wire [1:0]  _GEN_56 = {tree32Leaf0_19_2, tree32Leaf0_18_2};
  wire [1:0]  tree32G_lo_hi_lo_lo_hi;
  assign tree32G_lo_hi_lo_lo_hi = _GEN_56;
  wire [1:0]  tree64G_lo_hi_lo_lo_hi;
  assign tree64G_lo_hi_lo_lo_hi = _GEN_56;
  wire [3:0]  tree32G_lo_hi_lo_lo = {tree32G_lo_hi_lo_lo_hi, tree32G_lo_hi_lo_lo_lo};
  wire [1:0]  _GEN_57 = {tree32Leaf0_21_2, tree32Leaf0_20_2};
  wire [1:0]  tree32G_lo_hi_lo_hi_lo;
  assign tree32G_lo_hi_lo_hi_lo = _GEN_57;
  wire [1:0]  tree64G_lo_hi_lo_hi_lo;
  assign tree64G_lo_hi_lo_hi_lo = _GEN_57;
  wire [1:0]  _GEN_58 = {tree32Leaf0_23_2, tree32Leaf0_22_2};
  wire [1:0]  tree32G_lo_hi_lo_hi_hi;
  assign tree32G_lo_hi_lo_hi_hi = _GEN_58;
  wire [1:0]  tree64G_lo_hi_lo_hi_hi;
  assign tree64G_lo_hi_lo_hi_hi = _GEN_58;
  wire [3:0]  tree32G_lo_hi_lo_hi = {tree32G_lo_hi_lo_hi_hi, tree32G_lo_hi_lo_hi_lo};
  wire [7:0]  tree32G_lo_hi_lo = {tree32G_lo_hi_lo_hi, tree32G_lo_hi_lo_lo};
  wire [1:0]  _GEN_59 = {tree32Leaf0_25_2, tree32Leaf0_24_2};
  wire [1:0]  tree32G_lo_hi_hi_lo_lo;
  assign tree32G_lo_hi_hi_lo_lo = _GEN_59;
  wire [1:0]  tree64G_lo_hi_hi_lo_lo;
  assign tree64G_lo_hi_hi_lo_lo = _GEN_59;
  wire [1:0]  _GEN_60 = {tree32Leaf0_27_2, tree32Leaf0_26_2};
  wire [1:0]  tree32G_lo_hi_hi_lo_hi;
  assign tree32G_lo_hi_hi_lo_hi = _GEN_60;
  wire [1:0]  tree64G_lo_hi_hi_lo_hi;
  assign tree64G_lo_hi_hi_lo_hi = _GEN_60;
  wire [3:0]  tree32G_lo_hi_hi_lo = {tree32G_lo_hi_hi_lo_hi, tree32G_lo_hi_hi_lo_lo};
  wire [1:0]  _GEN_61 = {tree32Leaf0_29_2, tree32Leaf0_28_2};
  wire [1:0]  tree32G_lo_hi_hi_hi_lo;
  assign tree32G_lo_hi_hi_hi_lo = _GEN_61;
  wire [1:0]  tree64G_lo_hi_hi_hi_lo;
  assign tree64G_lo_hi_hi_hi_lo = _GEN_61;
  wire [1:0]  _GEN_62 = {tree32Leaf0_31_2, tree32Leaf0_30_2};
  wire [1:0]  tree32G_lo_hi_hi_hi_hi;
  assign tree32G_lo_hi_hi_hi_hi = _GEN_62;
  wire [1:0]  tree64G_lo_hi_hi_hi_hi;
  assign tree64G_lo_hi_hi_hi_hi = _GEN_62;
  wire [3:0]  tree32G_lo_hi_hi_hi = {tree32G_lo_hi_hi_hi_hi, tree32G_lo_hi_hi_hi_lo};
  wire [7:0]  tree32G_lo_hi_hi = {tree32G_lo_hi_hi_hi, tree32G_lo_hi_hi_lo};
  wire [15:0] tree32G_lo_hi = {tree32G_lo_hi_hi, tree32G_lo_hi_lo};
  wire [31:0] tree32G_lo = {tree32G_lo_hi, tree32G_lo_lo};
  wire [3:0]  tree32G_hi_lo_lo_lo = {tree32G_hi_lo_lo_lo_hi, tree32G_hi_lo_lo_lo_lo};
  wire [3:0]  tree32G_hi_lo_lo_hi = {tree32G_hi_lo_lo_hi_hi, tree32G_hi_lo_lo_hi_lo};
  wire [7:0]  tree32G_hi_lo_lo = {tree32G_hi_lo_lo_hi, tree32G_hi_lo_lo_lo};
  wire [3:0]  tree32G_hi_lo_hi_lo = {tree32G_hi_lo_hi_lo_hi, tree32G_hi_lo_hi_lo_lo};
  wire [3:0]  tree32G_hi_lo_hi_hi = {tree32G_hi_lo_hi_hi_hi, tree32G_hi_lo_hi_hi_lo};
  wire [7:0]  tree32G_hi_lo_hi = {tree32G_hi_lo_hi_hi, tree32G_hi_lo_hi_lo};
  wire [15:0] tree32G_hi_lo = {tree32G_hi_lo_hi, tree32G_hi_lo_lo};
  wire [1:0]  tree32G_hi_hi_lo_lo_lo = {tree32Leaf1_17_2, tree32Leaf1_16_2};
  wire [1:0]  tree32G_hi_hi_lo_lo_hi = {tree32Leaf1_19_2, tree32Leaf1_18_2};
  wire [3:0]  tree32G_hi_hi_lo_lo = {tree32G_hi_hi_lo_lo_hi, tree32G_hi_hi_lo_lo_lo};
  wire [1:0]  tree32G_hi_hi_lo_hi_lo = {tree32Leaf1_21_2, tree32Leaf1_20_2};
  wire [1:0]  tree32G_hi_hi_lo_hi_hi = {tree32Leaf1_23_2, tree32Leaf1_22_2};
  wire [3:0]  tree32G_hi_hi_lo_hi = {tree32G_hi_hi_lo_hi_hi, tree32G_hi_hi_lo_hi_lo};
  wire [7:0]  tree32G_hi_hi_lo = {tree32G_hi_hi_lo_hi, tree32G_hi_hi_lo_lo};
  wire [1:0]  tree32G_hi_hi_hi_lo_lo = {tree32Leaf1_25_2, tree32Leaf1_24_2};
  wire [1:0]  tree32G_hi_hi_hi_lo_hi = {tree32Leaf1_27_2, tree32Leaf1_26_2};
  wire [3:0]  tree32G_hi_hi_hi_lo = {tree32G_hi_hi_hi_lo_hi, tree32G_hi_hi_hi_lo_lo};
  wire [1:0]  tree32G_hi_hi_hi_hi_lo = {tree32Leaf1_29_2, tree32Leaf1_28_2};
  wire [1:0]  tree32G_hi_hi_hi_hi_hi = {tree32Leaf1_31_2, tree32Leaf1_30_2};
  wire [3:0]  tree32G_hi_hi_hi_hi = {tree32G_hi_hi_hi_hi_hi, tree32G_hi_hi_hi_hi_lo};
  wire [7:0]  tree32G_hi_hi_hi = {tree32G_hi_hi_hi_hi, tree32G_hi_hi_hi_lo};
  wire [15:0] tree32G_hi_hi = {tree32G_hi_hi_hi, tree32G_hi_hi_lo};
  wire [31:0] tree32G_hi = {tree32G_hi_hi, tree32G_hi_lo};
  wire [63:0] tree32G = {tree32G_hi, tree32G_lo};
  wire [3:0]  tree64P_lo_lo_lo_lo = {tree64P_lo_lo_lo_lo_hi, tree64P_lo_lo_lo_lo_lo};
  wire [3:0]  tree64P_lo_lo_lo_hi = {tree64P_lo_lo_lo_hi_hi, tree64P_lo_lo_lo_hi_lo};
  wire [7:0]  tree64P_lo_lo_lo = {tree64P_lo_lo_lo_hi, tree64P_lo_lo_lo_lo};
  wire [3:0]  tree64P_lo_lo_hi_lo = {tree64P_lo_lo_hi_lo_hi, tree64P_lo_lo_hi_lo_lo};
  wire [3:0]  tree64P_lo_lo_hi_hi = {tree64P_lo_lo_hi_hi_hi, tree64P_lo_lo_hi_hi_lo};
  wire [7:0]  tree64P_lo_lo_hi = {tree64P_lo_lo_hi_hi, tree64P_lo_lo_hi_lo};
  wire [15:0] tree64P_lo_lo = {tree64P_lo_lo_hi, tree64P_lo_lo_lo};
  wire [3:0]  tree64P_lo_hi_lo_lo = {tree64P_lo_hi_lo_lo_hi, tree64P_lo_hi_lo_lo_lo};
  wire [3:0]  tree64P_lo_hi_lo_hi = {tree64P_lo_hi_lo_hi_hi, tree64P_lo_hi_lo_hi_lo};
  wire [7:0]  tree64P_lo_hi_lo = {tree64P_lo_hi_lo_hi, tree64P_lo_hi_lo_lo};
  wire [3:0]  tree64P_lo_hi_hi_lo = {tree64P_lo_hi_hi_lo_hi, tree64P_lo_hi_hi_lo_lo};
  wire [3:0]  tree64P_lo_hi_hi_hi = {tree64P_lo_hi_hi_hi_hi, tree64P_lo_hi_hi_hi_lo};
  wire [7:0]  tree64P_lo_hi_hi = {tree64P_lo_hi_hi_hi, tree64P_lo_hi_hi_lo};
  wire [15:0] tree64P_lo_hi = {tree64P_lo_hi_hi, tree64P_lo_hi_lo};
  wire [31:0] tree64P_lo = {tree64P_lo_hi, tree64P_lo_lo};
  wire [1:0]  tree64P_hi_lo_lo_lo_lo = {tree64_33_1, tree64_32_1};
  wire [1:0]  tree64P_hi_lo_lo_lo_hi = {tree64_35_1, tree64_34_1};
  wire [3:0]  tree64P_hi_lo_lo_lo = {tree64P_hi_lo_lo_lo_hi, tree64P_hi_lo_lo_lo_lo};
  wire [1:0]  tree64P_hi_lo_lo_hi_lo = {tree64_37_1, tree64_36_1};
  wire [1:0]  tree64P_hi_lo_lo_hi_hi = {tree64_39_1, tree64_38_1};
  wire [3:0]  tree64P_hi_lo_lo_hi = {tree64P_hi_lo_lo_hi_hi, tree64P_hi_lo_lo_hi_lo};
  wire [7:0]  tree64P_hi_lo_lo = {tree64P_hi_lo_lo_hi, tree64P_hi_lo_lo_lo};
  wire [1:0]  tree64P_hi_lo_hi_lo_lo = {tree64_41_1, tree64_40_1};
  wire [1:0]  tree64P_hi_lo_hi_lo_hi = {tree64_43_1, tree64_42_1};
  wire [3:0]  tree64P_hi_lo_hi_lo = {tree64P_hi_lo_hi_lo_hi, tree64P_hi_lo_hi_lo_lo};
  wire [1:0]  tree64P_hi_lo_hi_hi_lo = {tree64_45_1, tree64_44_1};
  wire [1:0]  tree64P_hi_lo_hi_hi_hi = {tree64_47_1, tree64_46_1};
  wire [3:0]  tree64P_hi_lo_hi_hi = {tree64P_hi_lo_hi_hi_hi, tree64P_hi_lo_hi_hi_lo};
  wire [7:0]  tree64P_hi_lo_hi = {tree64P_hi_lo_hi_hi, tree64P_hi_lo_hi_lo};
  wire [15:0] tree64P_hi_lo = {tree64P_hi_lo_hi, tree64P_hi_lo_lo};
  wire [1:0]  tree64P_hi_hi_lo_lo_lo = {tree64_49_1, tree64_48_1};
  wire [1:0]  tree64P_hi_hi_lo_lo_hi = {tree64_51_1, tree64_50_1};
  wire [3:0]  tree64P_hi_hi_lo_lo = {tree64P_hi_hi_lo_lo_hi, tree64P_hi_hi_lo_lo_lo};
  wire [1:0]  tree64P_hi_hi_lo_hi_lo = {tree64_53_1, tree64_52_1};
  wire [1:0]  tree64P_hi_hi_lo_hi_hi = {tree64_55_1, tree64_54_1};
  wire [3:0]  tree64P_hi_hi_lo_hi = {tree64P_hi_hi_lo_hi_hi, tree64P_hi_hi_lo_hi_lo};
  wire [7:0]  tree64P_hi_hi_lo = {tree64P_hi_hi_lo_hi, tree64P_hi_hi_lo_lo};
  wire [1:0]  tree64P_hi_hi_hi_lo_lo = {tree64_57_1, tree64_56_1};
  wire [1:0]  tree64P_hi_hi_hi_lo_hi = {tree64_59_1, tree64_58_1};
  wire [3:0]  tree64P_hi_hi_hi_lo = {tree64P_hi_hi_hi_lo_hi, tree64P_hi_hi_hi_lo_lo};
  wire [1:0]  tree64P_hi_hi_hi_hi_lo = {tree64_61_1, tree64_60_1};
  wire [1:0]  tree64P_hi_hi_hi_hi_hi = {tree64_63_1, tree64_62_1};
  wire [3:0]  tree64P_hi_hi_hi_hi = {tree64P_hi_hi_hi_hi_hi, tree64P_hi_hi_hi_hi_lo};
  wire [7:0]  tree64P_hi_hi_hi = {tree64P_hi_hi_hi_hi, tree64P_hi_hi_hi_lo};
  wire [15:0] tree64P_hi_hi = {tree64P_hi_hi_hi, tree64P_hi_hi_lo};
  wire [31:0] tree64P_hi = {tree64P_hi_hi, tree64P_hi_lo};
  wire [63:0] tree64P = {tree64P_hi, tree64P_lo};
  wire [3:0]  tree64G_lo_lo_lo_lo = {tree64G_lo_lo_lo_lo_hi, tree64G_lo_lo_lo_lo_lo};
  wire [3:0]  tree64G_lo_lo_lo_hi = {tree64G_lo_lo_lo_hi_hi, tree64G_lo_lo_lo_hi_lo};
  wire [7:0]  tree64G_lo_lo_lo = {tree64G_lo_lo_lo_hi, tree64G_lo_lo_lo_lo};
  wire [3:0]  tree64G_lo_lo_hi_lo = {tree64G_lo_lo_hi_lo_hi, tree64G_lo_lo_hi_lo_lo};
  wire [3:0]  tree64G_lo_lo_hi_hi = {tree64G_lo_lo_hi_hi_hi, tree64G_lo_lo_hi_hi_lo};
  wire [7:0]  tree64G_lo_lo_hi = {tree64G_lo_lo_hi_hi, tree64G_lo_lo_hi_lo};
  wire [15:0] tree64G_lo_lo = {tree64G_lo_lo_hi, tree64G_lo_lo_lo};
  wire [3:0]  tree64G_lo_hi_lo_lo = {tree64G_lo_hi_lo_lo_hi, tree64G_lo_hi_lo_lo_lo};
  wire [3:0]  tree64G_lo_hi_lo_hi = {tree64G_lo_hi_lo_hi_hi, tree64G_lo_hi_lo_hi_lo};
  wire [7:0]  tree64G_lo_hi_lo = {tree64G_lo_hi_lo_hi, tree64G_lo_hi_lo_lo};
  wire [3:0]  tree64G_lo_hi_hi_lo = {tree64G_lo_hi_hi_lo_hi, tree64G_lo_hi_hi_lo_lo};
  wire [3:0]  tree64G_lo_hi_hi_hi = {tree64G_lo_hi_hi_hi_hi, tree64G_lo_hi_hi_hi_lo};
  wire [7:0]  tree64G_lo_hi_hi = {tree64G_lo_hi_hi_hi, tree64G_lo_hi_hi_lo};
  wire [15:0] tree64G_lo_hi = {tree64G_lo_hi_hi, tree64G_lo_hi_lo};
  wire [31:0] tree64G_lo = {tree64G_lo_hi, tree64G_lo_lo};
  wire [1:0]  tree64G_hi_lo_lo_lo_lo = {tree64_33_2, tree64_32_2};
  wire [1:0]  tree64G_hi_lo_lo_lo_hi = {tree64_35_2, tree64_34_2};
  wire [3:0]  tree64G_hi_lo_lo_lo = {tree64G_hi_lo_lo_lo_hi, tree64G_hi_lo_lo_lo_lo};
  wire [1:0]  tree64G_hi_lo_lo_hi_lo = {tree64_37_2, tree64_36_2};
  wire [1:0]  tree64G_hi_lo_lo_hi_hi = {tree64_39_2, tree64_38_2};
  wire [3:0]  tree64G_hi_lo_lo_hi = {tree64G_hi_lo_lo_hi_hi, tree64G_hi_lo_lo_hi_lo};
  wire [7:0]  tree64G_hi_lo_lo = {tree64G_hi_lo_lo_hi, tree64G_hi_lo_lo_lo};
  wire [1:0]  tree64G_hi_lo_hi_lo_lo = {tree64_41_2, tree64_40_2};
  wire [1:0]  tree64G_hi_lo_hi_lo_hi = {tree64_43_2, tree64_42_2};
  wire [3:0]  tree64G_hi_lo_hi_lo = {tree64G_hi_lo_hi_lo_hi, tree64G_hi_lo_hi_lo_lo};
  wire [1:0]  tree64G_hi_lo_hi_hi_lo = {tree64_45_2, tree64_44_2};
  wire [1:0]  tree64G_hi_lo_hi_hi_hi = {tree64_47_2, tree64_46_2};
  wire [3:0]  tree64G_hi_lo_hi_hi = {tree64G_hi_lo_hi_hi_hi, tree64G_hi_lo_hi_hi_lo};
  wire [7:0]  tree64G_hi_lo_hi = {tree64G_hi_lo_hi_hi, tree64G_hi_lo_hi_lo};
  wire [15:0] tree64G_hi_lo = {tree64G_hi_lo_hi, tree64G_hi_lo_lo};
  wire [1:0]  tree64G_hi_hi_lo_lo_lo = {tree64_49_2, tree64_48_2};
  wire [1:0]  tree64G_hi_hi_lo_lo_hi = {tree64_51_2, tree64_50_2};
  wire [3:0]  tree64G_hi_hi_lo_lo = {tree64G_hi_hi_lo_lo_hi, tree64G_hi_hi_lo_lo_lo};
  wire [1:0]  tree64G_hi_hi_lo_hi_lo = {tree64_53_2, tree64_52_2};
  wire [1:0]  tree64G_hi_hi_lo_hi_hi = {tree64_55_2, tree64_54_2};
  wire [3:0]  tree64G_hi_hi_lo_hi = {tree64G_hi_hi_lo_hi_hi, tree64G_hi_hi_lo_hi_lo};
  wire [7:0]  tree64G_hi_hi_lo = {tree64G_hi_hi_lo_hi, tree64G_hi_hi_lo_lo};
  wire [1:0]  tree64G_hi_hi_hi_lo_lo = {tree64_57_2, tree64_56_2};
  wire [1:0]  tree64G_hi_hi_hi_lo_hi = {tree64_59_2, tree64_58_2};
  wire [3:0]  tree64G_hi_hi_hi_lo = {tree64G_hi_hi_hi_lo_hi, tree64G_hi_hi_hi_lo_lo};
  wire [1:0]  tree64G_hi_hi_hi_hi_lo = {tree64_61_2, tree64_60_2};
  wire [1:0]  tree64G_hi_hi_hi_hi_hi = {tree64_63_2, tree64_62_2};
  wire [3:0]  tree64G_hi_hi_hi_hi = {tree64G_hi_hi_hi_hi_hi, tree64G_hi_hi_hi_hi_lo};
  wire [7:0]  tree64G_hi_hi_hi = {tree64G_hi_hi_hi_hi, tree64G_hi_hi_hi_lo};
  wire [15:0] tree64G_hi_hi = {tree64G_hi_hi_hi, tree64G_hi_hi_lo};
  wire [31:0] tree64G_hi = {tree64G_hi_hi, tree64G_hi_lo};
  wire [63:0] tree64G = {tree64G_hi, tree64G_lo};
  wire [63:0] treeP = (sew[0] ? tree8P : 64'h0) | (sew[1] ? tree16P : 64'h0) | (sew[2] ? tree32P : 64'h0) | (sew[3] ? tree64P : 64'h0);
  wire [63:0] treeG = (sew[0] ? tree8G : 64'h0) | (sew[1] ? tree16G : 64'h0) | (sew[2] ? tree32G : 64'h0) | (sew[3] ? tree64G : 64'h0);
  wire        tree_0_1 = treeP[0];
  wire        tree_1_1 = treeP[1];
  wire        tree_2_1 = treeP[2];
  wire        tree_3_1 = treeP[3];
  wire        tree_4_1 = treeP[4];
  wire        tree_5_1 = treeP[5];
  wire        tree_6_1 = treeP[6];
  wire        tree_7_1 = treeP[7];
  wire        tree_8_1 = treeP[8];
  wire        tree_9_1 = treeP[9];
  wire        tree_10_1 = treeP[10];
  wire        tree_11_1 = treeP[11];
  wire        tree_12_1 = treeP[12];
  wire        tree_13_1 = treeP[13];
  wire        tree_14_1 = treeP[14];
  wire        tree_15_1 = treeP[15];
  wire        tree_16_1 = treeP[16];
  wire        tree_17_1 = treeP[17];
  wire        tree_18_1 = treeP[18];
  wire        tree_19_1 = treeP[19];
  wire        tree_20_1 = treeP[20];
  wire        tree_21_1 = treeP[21];
  wire        tree_22_1 = treeP[22];
  wire        tree_23_1 = treeP[23];
  wire        tree_24_1 = treeP[24];
  wire        tree_25_1 = treeP[25];
  wire        tree_26_1 = treeP[26];
  wire        tree_27_1 = treeP[27];
  wire        tree_28_1 = treeP[28];
  wire        tree_29_1 = treeP[29];
  wire        tree_30_1 = treeP[30];
  wire        tree_31_1 = treeP[31];
  wire        tree_32_1 = treeP[32];
  wire        tree_33_1 = treeP[33];
  wire        tree_34_1 = treeP[34];
  wire        tree_35_1 = treeP[35];
  wire        tree_36_1 = treeP[36];
  wire        tree_37_1 = treeP[37];
  wire        tree_38_1 = treeP[38];
  wire        tree_39_1 = treeP[39];
  wire        tree_40_1 = treeP[40];
  wire        tree_41_1 = treeP[41];
  wire        tree_42_1 = treeP[42];
  wire        tree_43_1 = treeP[43];
  wire        tree_44_1 = treeP[44];
  wire        tree_45_1 = treeP[45];
  wire        tree_46_1 = treeP[46];
  wire        tree_47_1 = treeP[47];
  wire        tree_48_1 = treeP[48];
  wire        tree_49_1 = treeP[49];
  wire        tree_50_1 = treeP[50];
  wire        tree_51_1 = treeP[51];
  wire        tree_52_1 = treeP[52];
  wire        tree_53_1 = treeP[53];
  wire        tree_54_1 = treeP[54];
  wire        tree_55_1 = treeP[55];
  wire        tree_56_1 = treeP[56];
  wire        tree_57_1 = treeP[57];
  wire        tree_58_1 = treeP[58];
  wire        tree_59_1 = treeP[59];
  wire        tree_60_1 = treeP[60];
  wire        tree_61_1 = treeP[61];
  wire        tree_62_1 = treeP[62];
  wire        tree_63_1 = treeP[63];
  wire        tree_0_2 = treeG[0];
  wire        tree_1_2 = treeG[1];
  wire        tree_2_2 = treeG[2];
  wire        tree_3_2 = treeG[3];
  wire        tree_4_2 = treeG[4];
  wire        tree_5_2 = treeG[5];
  wire        tree_6_2 = treeG[6];
  wire        tree_7_2 = treeG[7];
  wire        tree_8_2 = treeG[8];
  wire        tree_9_2 = treeG[9];
  wire        tree_10_2 = treeG[10];
  wire        tree_11_2 = treeG[11];
  wire        tree_12_2 = treeG[12];
  wire        tree_13_2 = treeG[13];
  wire        tree_14_2 = treeG[14];
  wire        tree_15_2 = treeG[15];
  wire        tree_16_2 = treeG[16];
  wire        tree_17_2 = treeG[17];
  wire        tree_18_2 = treeG[18];
  wire        tree_19_2 = treeG[19];
  wire        tree_20_2 = treeG[20];
  wire        tree_21_2 = treeG[21];
  wire        tree_22_2 = treeG[22];
  wire        tree_23_2 = treeG[23];
  wire        tree_24_2 = treeG[24];
  wire        tree_25_2 = treeG[25];
  wire        tree_26_2 = treeG[26];
  wire        tree_27_2 = treeG[27];
  wire        tree_28_2 = treeG[28];
  wire        tree_29_2 = treeG[29];
  wire        tree_30_2 = treeG[30];
  wire        tree_31_2 = treeG[31];
  wire        tree_32_2 = treeG[32];
  wire        tree_33_2 = treeG[33];
  wire        tree_34_2 = treeG[34];
  wire        tree_35_2 = treeG[35];
  wire        tree_36_2 = treeG[36];
  wire        tree_37_2 = treeG[37];
  wire        tree_38_2 = treeG[38];
  wire        tree_39_2 = treeG[39];
  wire        tree_40_2 = treeG[40];
  wire        tree_41_2 = treeG[41];
  wire        tree_42_2 = treeG[42];
  wire        tree_43_2 = treeG[43];
  wire        tree_44_2 = treeG[44];
  wire        tree_45_2 = treeG[45];
  wire        tree_46_2 = treeG[46];
  wire        tree_47_2 = treeG[47];
  wire        tree_48_2 = treeG[48];
  wire        tree_49_2 = treeG[49];
  wire        tree_50_2 = treeG[50];
  wire        tree_51_2 = treeG[51];
  wire        tree_52_2 = treeG[52];
  wire        tree_53_2 = treeG[53];
  wire        tree_54_2 = treeG[54];
  wire        tree_55_2 = treeG[55];
  wire        tree_56_2 = treeG[56];
  wire        tree_57_2 = treeG[57];
  wire        tree_58_2 = treeG[58];
  wire        tree_59_2 = treeG[59];
  wire        tree_60_2 = treeG[60];
  wire        tree_61_2 = treeG[61];
  wire        tree_62_2 = treeG[62];
  wire        tree_63_2 = treeG[63];
  wire [1:0]  carryResult_cbank_lo_lo = {tree_1_2, tree_0_2};
  wire [1:0]  carryResult_cbank_lo_hi = {tree_3_2, tree_2_2};
  wire [3:0]  carryResult_cbank_lo = {carryResult_cbank_lo_hi, carryResult_cbank_lo_lo};
  wire [1:0]  carryResult_cbank_hi_lo = {tree_5_2, tree_4_2};
  wire [1:0]  carryResult_cbank_hi_hi = {tree_7_2, tree_6_2};
  wire [3:0]  carryResult_cbank_hi = {carryResult_cbank_hi_hi, carryResult_cbank_hi_lo};
  wire [7:0]  carryResult_cbank_0 = {carryResult_cbank_hi, carryResult_cbank_lo};
  wire [1:0]  carryResult_cbank_lo_lo_1 = {tree_9_2, tree_8_2};
  wire [1:0]  carryResult_cbank_lo_hi_1 = {tree_11_2, tree_10_2};
  wire [3:0]  carryResult_cbank_lo_1 = {carryResult_cbank_lo_hi_1, carryResult_cbank_lo_lo_1};
  wire [1:0]  carryResult_cbank_hi_lo_1 = {tree_13_2, tree_12_2};
  wire [1:0]  carryResult_cbank_hi_hi_1 = {tree_15_2, tree_14_2};
  wire [3:0]  carryResult_cbank_hi_1 = {carryResult_cbank_hi_hi_1, carryResult_cbank_hi_lo_1};
  wire [7:0]  carryResult_cbank_1 = {carryResult_cbank_hi_1, carryResult_cbank_lo_1};
  wire [1:0]  carryResult_cbank_lo_lo_2 = {tree_17_2, tree_16_2};
  wire [1:0]  carryResult_cbank_lo_hi_2 = {tree_19_2, tree_18_2};
  wire [3:0]  carryResult_cbank_lo_2 = {carryResult_cbank_lo_hi_2, carryResult_cbank_lo_lo_2};
  wire [1:0]  carryResult_cbank_hi_lo_2 = {tree_21_2, tree_20_2};
  wire [1:0]  carryResult_cbank_hi_hi_2 = {tree_23_2, tree_22_2};
  wire [3:0]  carryResult_cbank_hi_2 = {carryResult_cbank_hi_hi_2, carryResult_cbank_hi_lo_2};
  wire [7:0]  carryResult_cbank_2 = {carryResult_cbank_hi_2, carryResult_cbank_lo_2};
  wire [1:0]  carryResult_cbank_lo_lo_3 = {tree_25_2, tree_24_2};
  wire [1:0]  carryResult_cbank_lo_hi_3 = {tree_27_2, tree_26_2};
  wire [3:0]  carryResult_cbank_lo_3 = {carryResult_cbank_lo_hi_3, carryResult_cbank_lo_lo_3};
  wire [1:0]  carryResult_cbank_hi_lo_3 = {tree_29_2, tree_28_2};
  wire [1:0]  carryResult_cbank_hi_hi_3 = {tree_31_2, tree_30_2};
  wire [3:0]  carryResult_cbank_hi_3 = {carryResult_cbank_hi_hi_3, carryResult_cbank_hi_lo_3};
  wire [7:0]  carryResult_cbank_3 = {carryResult_cbank_hi_3, carryResult_cbank_lo_3};
  wire [1:0]  carryResult_cbank_lo_lo_4 = {tree_33_2, tree_32_2};
  wire [1:0]  carryResult_cbank_lo_hi_4 = {tree_35_2, tree_34_2};
  wire [3:0]  carryResult_cbank_lo_4 = {carryResult_cbank_lo_hi_4, carryResult_cbank_lo_lo_4};
  wire [1:0]  carryResult_cbank_hi_lo_4 = {tree_37_2, tree_36_2};
  wire [1:0]  carryResult_cbank_hi_hi_4 = {tree_39_2, tree_38_2};
  wire [3:0]  carryResult_cbank_hi_4 = {carryResult_cbank_hi_hi_4, carryResult_cbank_hi_lo_4};
  wire [7:0]  carryResult_cbank_4 = {carryResult_cbank_hi_4, carryResult_cbank_lo_4};
  wire [1:0]  carryResult_cbank_lo_lo_5 = {tree_41_2, tree_40_2};
  wire [1:0]  carryResult_cbank_lo_hi_5 = {tree_43_2, tree_42_2};
  wire [3:0]  carryResult_cbank_lo_5 = {carryResult_cbank_lo_hi_5, carryResult_cbank_lo_lo_5};
  wire [1:0]  carryResult_cbank_hi_lo_5 = {tree_45_2, tree_44_2};
  wire [1:0]  carryResult_cbank_hi_hi_5 = {tree_47_2, tree_46_2};
  wire [3:0]  carryResult_cbank_hi_5 = {carryResult_cbank_hi_hi_5, carryResult_cbank_hi_lo_5};
  wire [7:0]  carryResult_cbank_5 = {carryResult_cbank_hi_5, carryResult_cbank_lo_5};
  wire [1:0]  carryResult_cbank_lo_lo_6 = {tree_49_2, tree_48_2};
  wire [1:0]  carryResult_cbank_lo_hi_6 = {tree_51_2, tree_50_2};
  wire [3:0]  carryResult_cbank_lo_6 = {carryResult_cbank_lo_hi_6, carryResult_cbank_lo_lo_6};
  wire [1:0]  carryResult_cbank_hi_lo_6 = {tree_53_2, tree_52_2};
  wire [1:0]  carryResult_cbank_hi_hi_6 = {tree_55_2, tree_54_2};
  wire [3:0]  carryResult_cbank_hi_6 = {carryResult_cbank_hi_hi_6, carryResult_cbank_hi_lo_6};
  wire [7:0]  carryResult_cbank_6 = {carryResult_cbank_hi_6, carryResult_cbank_lo_6};
  wire [1:0]  carryResult_cbank_lo_lo_7 = {tree_57_2, tree_56_2};
  wire [1:0]  carryResult_cbank_lo_hi_7 = {tree_59_2, tree_58_2};
  wire [3:0]  carryResult_cbank_lo_7 = {carryResult_cbank_lo_hi_7, carryResult_cbank_lo_lo_7};
  wire [1:0]  carryResult_cbank_hi_lo_7 = {tree_61_2, tree_60_2};
  wire [1:0]  carryResult_cbank_hi_hi_7 = {tree_63_2, tree_62_2};
  wire [3:0]  carryResult_cbank_hi_7 = {carryResult_cbank_hi_hi_7, carryResult_cbank_hi_lo_7};
  wire [7:0]  carryResult_cbank_7 = {carryResult_cbank_hi_7, carryResult_cbank_lo_7};
  wire [15:0] carryResult_lo_lo = {carryResult_cbank_1, carryResult_cbank_0};
  wire [15:0] carryResult_lo_hi = {carryResult_cbank_3, carryResult_cbank_2};
  wire [31:0] carryResult_lo = {carryResult_lo_hi, carryResult_lo_lo};
  wire [15:0] carryResult_hi_lo = {carryResult_cbank_5, carryResult_cbank_4};
  wire [15:0] carryResult_hi_hi = {carryResult_cbank_7, carryResult_cbank_6};
  wire [31:0] carryResult_hi = {carryResult_hi_hi, carryResult_hi_lo};
  wire [63:0] carryResult = {carryResult_hi, carryResult_lo};
  wire        cout64 = carryResult[63];
  wire [7:0]  cout8 = {cout64, carryResult[55], carryResult[47], carryResult[39], carryResult[31], carryResult[23], carryResult[15], carryResult[7]};
  wire [3:0]  cout16 = {cout64, carryResult[47], carryResult[31], carryResult[15]};
  wire [1:0]  cout32 = {cout64, carryResult[31]};
  wire [7:0]  carryInSele =
    (sew[1] ? {carryResult[55], 1'h0, carryResult[39], 1'h0, carryResult[23], 1'h0, carryResult[7], 1'h0} : 8'h0)
    | (sew[2] ? {carryResult[55], carryResult[47], carryResult[39], 1'h0, carryResult[23], carryResult[15], carryResult[7], 1'h0} : 8'h0)
    | (sew[3] ? {carryResult[55], carryResult[47], carryResult[39], carryResult[31], carryResult[23], carryResult[15], carryResult[7], 1'h0} : 8'h0);
  wire [7:0]  cs_lo_lo_lo = {carryResult[6:0], carryInSele[0]};
  wire [7:0]  cs_lo_lo_hi = {carryResult[14:8], carryInSele[1]};
  wire [15:0] cs_lo_lo = {cs_lo_lo_hi, cs_lo_lo_lo};
  wire [7:0]  cs_lo_hi_lo = {carryResult[22:16], carryInSele[2]};
  wire [7:0]  cs_lo_hi_hi = {carryResult[30:24], carryInSele[3]};
  wire [15:0] cs_lo_hi = {cs_lo_hi_hi, cs_lo_hi_lo};
  wire [31:0] cs_lo = {cs_lo_hi, cs_lo_lo};
  wire [7:0]  cs_hi_lo_lo = {carryResult[38:32], carryInSele[4]};
  wire [7:0]  cs_hi_lo_hi = {carryResult[46:40], carryInSele[5]};
  wire [15:0] cs_hi_lo = {cs_hi_lo_hi, cs_hi_lo_lo};
  wire [7:0]  cs_hi_hi_lo = {carryResult[54:48], carryInSele[6]};
  wire [7:0]  cs_hi_hi_hi = {carryResult[62:56], carryInSele[7]};
  wire [15:0] cs_hi_hi = {cs_hi_hi_hi, cs_hi_hi_lo};
  wire [31:0] cs_hi = {cs_hi_hi, cs_hi_lo};
  wire [63:0] cs = {cs_hi, cs_lo};
  wire [1:0]  ps_lo_lo_lo_lo_lo = {pairs_1_1, pairs_0_1};
  wire [1:0]  ps_lo_lo_lo_lo_hi = {pairs_3_1, pairs_2_1};
  wire [3:0]  ps_lo_lo_lo_lo = {ps_lo_lo_lo_lo_hi, ps_lo_lo_lo_lo_lo};
  wire [1:0]  ps_lo_lo_lo_hi_lo = {pairs_5_1, pairs_4_1};
  wire [1:0]  ps_lo_lo_lo_hi_hi = {pairs_7_1, pairs_6_1};
  wire [3:0]  ps_lo_lo_lo_hi = {ps_lo_lo_lo_hi_hi, ps_lo_lo_lo_hi_lo};
  wire [7:0]  ps_lo_lo_lo = {ps_lo_lo_lo_hi, ps_lo_lo_lo_lo};
  wire [1:0]  ps_lo_lo_hi_lo_lo = {pairs_9_1, pairs_8_1};
  wire [1:0]  ps_lo_lo_hi_lo_hi = {pairs_11_1, pairs_10_1};
  wire [3:0]  ps_lo_lo_hi_lo = {ps_lo_lo_hi_lo_hi, ps_lo_lo_hi_lo_lo};
  wire [1:0]  ps_lo_lo_hi_hi_lo = {pairs_13_1, pairs_12_1};
  wire [1:0]  ps_lo_lo_hi_hi_hi = {pairs_15_1, pairs_14_1};
  wire [3:0]  ps_lo_lo_hi_hi = {ps_lo_lo_hi_hi_hi, ps_lo_lo_hi_hi_lo};
  wire [7:0]  ps_lo_lo_hi = {ps_lo_lo_hi_hi, ps_lo_lo_hi_lo};
  wire [15:0] ps_lo_lo = {ps_lo_lo_hi, ps_lo_lo_lo};
  wire [1:0]  ps_lo_hi_lo_lo_lo = {pairs_17_1, pairs_16_1};
  wire [1:0]  ps_lo_hi_lo_lo_hi = {pairs_19_1, pairs_18_1};
  wire [3:0]  ps_lo_hi_lo_lo = {ps_lo_hi_lo_lo_hi, ps_lo_hi_lo_lo_lo};
  wire [1:0]  ps_lo_hi_lo_hi_lo = {pairs_21_1, pairs_20_1};
  wire [1:0]  ps_lo_hi_lo_hi_hi = {pairs_23_1, pairs_22_1};
  wire [3:0]  ps_lo_hi_lo_hi = {ps_lo_hi_lo_hi_hi, ps_lo_hi_lo_hi_lo};
  wire [7:0]  ps_lo_hi_lo = {ps_lo_hi_lo_hi, ps_lo_hi_lo_lo};
  wire [1:0]  ps_lo_hi_hi_lo_lo = {pairs_25_1, pairs_24_1};
  wire [1:0]  ps_lo_hi_hi_lo_hi = {pairs_27_1, pairs_26_1};
  wire [3:0]  ps_lo_hi_hi_lo = {ps_lo_hi_hi_lo_hi, ps_lo_hi_hi_lo_lo};
  wire [1:0]  ps_lo_hi_hi_hi_lo = {pairs_29_1, pairs_28_1};
  wire [1:0]  ps_lo_hi_hi_hi_hi = {pairs_31_1, pairs_30_1};
  wire [3:0]  ps_lo_hi_hi_hi = {ps_lo_hi_hi_hi_hi, ps_lo_hi_hi_hi_lo};
  wire [7:0]  ps_lo_hi_hi = {ps_lo_hi_hi_hi, ps_lo_hi_hi_lo};
  wire [15:0] ps_lo_hi = {ps_lo_hi_hi, ps_lo_hi_lo};
  wire [31:0] ps_lo = {ps_lo_hi, ps_lo_lo};
  wire [1:0]  ps_hi_lo_lo_lo_lo = {pairs_33_1, pairs_32_1};
  wire [1:0]  ps_hi_lo_lo_lo_hi = {pairs_35_1, pairs_34_1};
  wire [3:0]  ps_hi_lo_lo_lo = {ps_hi_lo_lo_lo_hi, ps_hi_lo_lo_lo_lo};
  wire [1:0]  ps_hi_lo_lo_hi_lo = {pairs_37_1, pairs_36_1};
  wire [1:0]  ps_hi_lo_lo_hi_hi = {pairs_39_1, pairs_38_1};
  wire [3:0]  ps_hi_lo_lo_hi = {ps_hi_lo_lo_hi_hi, ps_hi_lo_lo_hi_lo};
  wire [7:0]  ps_hi_lo_lo = {ps_hi_lo_lo_hi, ps_hi_lo_lo_lo};
  wire [1:0]  ps_hi_lo_hi_lo_lo = {pairs_41_1, pairs_40_1};
  wire [1:0]  ps_hi_lo_hi_lo_hi = {pairs_43_1, pairs_42_1};
  wire [3:0]  ps_hi_lo_hi_lo = {ps_hi_lo_hi_lo_hi, ps_hi_lo_hi_lo_lo};
  wire [1:0]  ps_hi_lo_hi_hi_lo = {pairs_45_1, pairs_44_1};
  wire [1:0]  ps_hi_lo_hi_hi_hi = {pairs_47_1, pairs_46_1};
  wire [3:0]  ps_hi_lo_hi_hi = {ps_hi_lo_hi_hi_hi, ps_hi_lo_hi_hi_lo};
  wire [7:0]  ps_hi_lo_hi = {ps_hi_lo_hi_hi, ps_hi_lo_hi_lo};
  wire [15:0] ps_hi_lo = {ps_hi_lo_hi, ps_hi_lo_lo};
  wire [1:0]  ps_hi_hi_lo_lo_lo = {pairs_49_1, pairs_48_1};
  wire [1:0]  ps_hi_hi_lo_lo_hi = {pairs_51_1, pairs_50_1};
  wire [3:0]  ps_hi_hi_lo_lo = {ps_hi_hi_lo_lo_hi, ps_hi_hi_lo_lo_lo};
  wire [1:0]  ps_hi_hi_lo_hi_lo = {pairs_53_1, pairs_52_1};
  wire [1:0]  ps_hi_hi_lo_hi_hi = {pairs_55_1, pairs_54_1};
  wire [3:0]  ps_hi_hi_lo_hi = {ps_hi_hi_lo_hi_hi, ps_hi_hi_lo_hi_lo};
  wire [7:0]  ps_hi_hi_lo = {ps_hi_hi_lo_hi, ps_hi_hi_lo_lo};
  wire [1:0]  ps_hi_hi_hi_lo_lo = {pairs_57_1, pairs_56_1};
  wire [1:0]  ps_hi_hi_hi_lo_hi = {pairs_59_1, pairs_58_1};
  wire [3:0]  ps_hi_hi_hi_lo = {ps_hi_hi_hi_lo_hi, ps_hi_hi_hi_lo_lo};
  wire [1:0]  ps_hi_hi_hi_hi_lo = {pairs_61_1, pairs_60_1};
  wire [1:0]  ps_hi_hi_hi_hi_hi = {pairs_63_1, pairs_62_1};
  wire [3:0]  ps_hi_hi_hi_hi = {ps_hi_hi_hi_hi_hi, ps_hi_hi_hi_hi_lo};
  wire [7:0]  ps_hi_hi_hi = {ps_hi_hi_hi_hi, ps_hi_hi_hi_lo};
  wire [15:0] ps_hi_hi = {ps_hi_hi_hi, ps_hi_hi_lo};
  wire [31:0] ps_hi = {ps_hi_hi, ps_hi_lo};
  wire [63:0] ps = {ps_hi, ps_lo};
  assign z = ps ^ cs;
endmodule

