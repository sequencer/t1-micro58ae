module MaskUnitReadCrossBar(
  output       input_0_ready,
  input        input_0_valid,
  input  [4:0] input_0_bits_vs,
  input  [1:0] input_0_bits_offset,
  input  [3:0] input_0_bits_readLane,
  input  [1:0] input_0_bits_dataOffset,
  output       input_1_ready,
  input        input_1_valid,
  input  [4:0] input_1_bits_vs,
  input  [1:0] input_1_bits_offset,
  input  [3:0] input_1_bits_readLane,
  input  [1:0] input_1_bits_dataOffset,
  output       input_2_ready,
  input        input_2_valid,
  input  [4:0] input_2_bits_vs,
  input  [1:0] input_2_bits_offset,
  input  [3:0] input_2_bits_readLane,
  input  [1:0] input_2_bits_dataOffset,
  output       input_3_ready,
  input        input_3_valid,
  input  [4:0] input_3_bits_vs,
  input  [1:0] input_3_bits_offset,
  input  [3:0] input_3_bits_readLane,
  input  [1:0] input_3_bits_dataOffset,
  output       input_4_ready,
  input        input_4_valid,
  input  [4:0] input_4_bits_vs,
  input  [1:0] input_4_bits_offset,
  input  [3:0] input_4_bits_readLane,
  input  [1:0] input_4_bits_dataOffset,
  output       input_5_ready,
  input        input_5_valid,
  input  [4:0] input_5_bits_vs,
  input  [1:0] input_5_bits_offset,
  input  [3:0] input_5_bits_readLane,
  input  [1:0] input_5_bits_dataOffset,
  output       input_6_ready,
  input        input_6_valid,
  input  [4:0] input_6_bits_vs,
  input  [1:0] input_6_bits_offset,
  input  [3:0] input_6_bits_readLane,
  input  [1:0] input_6_bits_dataOffset,
  output       input_7_ready,
  input        input_7_valid,
  input  [4:0] input_7_bits_vs,
  input  [1:0] input_7_bits_offset,
  input  [3:0] input_7_bits_readLane,
  input  [1:0] input_7_bits_dataOffset,
  output       input_8_ready,
  input        input_8_valid,
  input  [4:0] input_8_bits_vs,
  input  [1:0] input_8_bits_offset,
  input  [3:0] input_8_bits_readLane,
  input  [1:0] input_8_bits_dataOffset,
  output       input_9_ready,
  input        input_9_valid,
  input  [4:0] input_9_bits_vs,
  input  [1:0] input_9_bits_offset,
  input  [3:0] input_9_bits_readLane,
  input  [1:0] input_9_bits_dataOffset,
  output       input_10_ready,
  input        input_10_valid,
  input  [4:0] input_10_bits_vs,
  input  [1:0] input_10_bits_offset,
  input  [3:0] input_10_bits_readLane,
  input  [1:0] input_10_bits_dataOffset,
  output       input_11_ready,
  input        input_11_valid,
  input  [4:0] input_11_bits_vs,
  input  [1:0] input_11_bits_offset,
  input  [3:0] input_11_bits_readLane,
  input  [1:0] input_11_bits_dataOffset,
  output       input_12_ready,
  input        input_12_valid,
  input  [4:0] input_12_bits_vs,
  input  [1:0] input_12_bits_offset,
  input  [3:0] input_12_bits_readLane,
  input  [1:0] input_12_bits_dataOffset,
  output       input_13_ready,
  input        input_13_valid,
  input  [4:0] input_13_bits_vs,
  input  [1:0] input_13_bits_offset,
  input  [3:0] input_13_bits_readLane,
  input  [1:0] input_13_bits_dataOffset,
  output       input_14_ready,
  input        input_14_valid,
  input  [4:0] input_14_bits_vs,
  input  [1:0] input_14_bits_offset,
  input  [3:0] input_14_bits_readLane,
  input  [1:0] input_14_bits_dataOffset,
  output       input_15_ready,
  input        input_15_valid,
  input  [4:0] input_15_bits_vs,
  input  [1:0] input_15_bits_offset,
  input  [3:0] input_15_bits_readLane,
  input  [1:0] input_15_bits_dataOffset,
  input        output_0_ready,
  output       output_0_valid,
  output [4:0] output_0_bits_vs,
  output [1:0] output_0_bits_offset,
  output [3:0] output_0_bits_writeIndex,
  output [1:0] output_0_bits_dataOffset,
  input        output_1_ready,
  output       output_1_valid,
  output [4:0] output_1_bits_vs,
  output [1:0] output_1_bits_offset,
  output [3:0] output_1_bits_writeIndex,
  output [1:0] output_1_bits_dataOffset,
  input        output_2_ready,
  output       output_2_valid,
  output [4:0] output_2_bits_vs,
  output [1:0] output_2_bits_offset,
  output [3:0] output_2_bits_writeIndex,
  output [1:0] output_2_bits_dataOffset,
  input        output_3_ready,
  output       output_3_valid,
  output [4:0] output_3_bits_vs,
  output [1:0] output_3_bits_offset,
  output [3:0] output_3_bits_writeIndex,
  output [1:0] output_3_bits_dataOffset,
  input        output_4_ready,
  output       output_4_valid,
  output [4:0] output_4_bits_vs,
  output [1:0] output_4_bits_offset,
  output [3:0] output_4_bits_writeIndex,
  output [1:0] output_4_bits_dataOffset,
  input        output_5_ready,
  output       output_5_valid,
  output [4:0] output_5_bits_vs,
  output [1:0] output_5_bits_offset,
  output [3:0] output_5_bits_writeIndex,
  output [1:0] output_5_bits_dataOffset,
  input        output_6_ready,
  output       output_6_valid,
  output [4:0] output_6_bits_vs,
  output [1:0] output_6_bits_offset,
  output [3:0] output_6_bits_writeIndex,
  output [1:0] output_6_bits_dataOffset,
  input        output_7_ready,
  output       output_7_valid,
  output [4:0] output_7_bits_vs,
  output [1:0] output_7_bits_offset,
  output [3:0] output_7_bits_writeIndex,
  output [1:0] output_7_bits_dataOffset,
  input        output_8_ready,
  output       output_8_valid,
  output [4:0] output_8_bits_vs,
  output [1:0] output_8_bits_offset,
  output [3:0] output_8_bits_writeIndex,
  output [1:0] output_8_bits_dataOffset,
  input        output_9_ready,
  output       output_9_valid,
  output [4:0] output_9_bits_vs,
  output [1:0] output_9_bits_offset,
  output [3:0] output_9_bits_writeIndex,
  output [1:0] output_9_bits_dataOffset,
  input        output_10_ready,
  output       output_10_valid,
  output [4:0] output_10_bits_vs,
  output [1:0] output_10_bits_offset,
  output [3:0] output_10_bits_writeIndex,
  output [1:0] output_10_bits_dataOffset,
  input        output_11_ready,
  output       output_11_valid,
  output [4:0] output_11_bits_vs,
  output [1:0] output_11_bits_offset,
  output [3:0] output_11_bits_writeIndex,
  output [1:0] output_11_bits_dataOffset,
  input        output_12_ready,
  output       output_12_valid,
  output [4:0] output_12_bits_vs,
  output [1:0] output_12_bits_offset,
  output [3:0] output_12_bits_writeIndex,
  output [1:0] output_12_bits_dataOffset,
  input        output_13_ready,
  output       output_13_valid,
  output [4:0] output_13_bits_vs,
  output [1:0] output_13_bits_offset,
  output [3:0] output_13_bits_writeIndex,
  output [1:0] output_13_bits_dataOffset,
  input        output_14_ready,
  output       output_14_valid,
  output [4:0] output_14_bits_vs,
  output [1:0] output_14_bits_offset,
  output [3:0] output_14_bits_writeIndex,
  output [1:0] output_14_bits_dataOffset,
  input        output_15_ready,
  output       output_15_valid,
  output [4:0] output_15_bits_vs,
  output [1:0] output_15_bits_offset,
  output [3:0] output_15_bits_writeIndex,
  output [1:0] output_15_bits_dataOffset
);

  wire        input_0_valid_0 = input_0_valid;
  wire [4:0]  input_0_bits_vs_0 = input_0_bits_vs;
  wire [1:0]  input_0_bits_offset_0 = input_0_bits_offset;
  wire [3:0]  input_0_bits_readLane_0 = input_0_bits_readLane;
  wire [1:0]  input_0_bits_dataOffset_0 = input_0_bits_dataOffset;
  wire        input_1_valid_0 = input_1_valid;
  wire [4:0]  input_1_bits_vs_0 = input_1_bits_vs;
  wire [1:0]  input_1_bits_offset_0 = input_1_bits_offset;
  wire [3:0]  input_1_bits_readLane_0 = input_1_bits_readLane;
  wire [1:0]  input_1_bits_dataOffset_0 = input_1_bits_dataOffset;
  wire        input_2_valid_0 = input_2_valid;
  wire [4:0]  input_2_bits_vs_0 = input_2_bits_vs;
  wire [1:0]  input_2_bits_offset_0 = input_2_bits_offset;
  wire [3:0]  input_2_bits_readLane_0 = input_2_bits_readLane;
  wire [1:0]  input_2_bits_dataOffset_0 = input_2_bits_dataOffset;
  wire        input_3_valid_0 = input_3_valid;
  wire [4:0]  input_3_bits_vs_0 = input_3_bits_vs;
  wire [1:0]  input_3_bits_offset_0 = input_3_bits_offset;
  wire [3:0]  input_3_bits_readLane_0 = input_3_bits_readLane;
  wire [1:0]  input_3_bits_dataOffset_0 = input_3_bits_dataOffset;
  wire        input_4_valid_0 = input_4_valid;
  wire [4:0]  input_4_bits_vs_0 = input_4_bits_vs;
  wire [1:0]  input_4_bits_offset_0 = input_4_bits_offset;
  wire [3:0]  input_4_bits_readLane_0 = input_4_bits_readLane;
  wire [1:0]  input_4_bits_dataOffset_0 = input_4_bits_dataOffset;
  wire        input_5_valid_0 = input_5_valid;
  wire [4:0]  input_5_bits_vs_0 = input_5_bits_vs;
  wire [1:0]  input_5_bits_offset_0 = input_5_bits_offset;
  wire [3:0]  input_5_bits_readLane_0 = input_5_bits_readLane;
  wire [1:0]  input_5_bits_dataOffset_0 = input_5_bits_dataOffset;
  wire        input_6_valid_0 = input_6_valid;
  wire [4:0]  input_6_bits_vs_0 = input_6_bits_vs;
  wire [1:0]  input_6_bits_offset_0 = input_6_bits_offset;
  wire [3:0]  input_6_bits_readLane_0 = input_6_bits_readLane;
  wire [1:0]  input_6_bits_dataOffset_0 = input_6_bits_dataOffset;
  wire        input_7_valid_0 = input_7_valid;
  wire [4:0]  input_7_bits_vs_0 = input_7_bits_vs;
  wire [1:0]  input_7_bits_offset_0 = input_7_bits_offset;
  wire [3:0]  input_7_bits_readLane_0 = input_7_bits_readLane;
  wire [1:0]  input_7_bits_dataOffset_0 = input_7_bits_dataOffset;
  wire        input_8_valid_0 = input_8_valid;
  wire [4:0]  input_8_bits_vs_0 = input_8_bits_vs;
  wire [1:0]  input_8_bits_offset_0 = input_8_bits_offset;
  wire [3:0]  input_8_bits_readLane_0 = input_8_bits_readLane;
  wire [1:0]  input_8_bits_dataOffset_0 = input_8_bits_dataOffset;
  wire        input_9_valid_0 = input_9_valid;
  wire [4:0]  input_9_bits_vs_0 = input_9_bits_vs;
  wire [1:0]  input_9_bits_offset_0 = input_9_bits_offset;
  wire [3:0]  input_9_bits_readLane_0 = input_9_bits_readLane;
  wire [1:0]  input_9_bits_dataOffset_0 = input_9_bits_dataOffset;
  wire        input_10_valid_0 = input_10_valid;
  wire [4:0]  input_10_bits_vs_0 = input_10_bits_vs;
  wire [1:0]  input_10_bits_offset_0 = input_10_bits_offset;
  wire [3:0]  input_10_bits_readLane_0 = input_10_bits_readLane;
  wire [1:0]  input_10_bits_dataOffset_0 = input_10_bits_dataOffset;
  wire        input_11_valid_0 = input_11_valid;
  wire [4:0]  input_11_bits_vs_0 = input_11_bits_vs;
  wire [1:0]  input_11_bits_offset_0 = input_11_bits_offset;
  wire [3:0]  input_11_bits_readLane_0 = input_11_bits_readLane;
  wire [1:0]  input_11_bits_dataOffset_0 = input_11_bits_dataOffset;
  wire        input_12_valid_0 = input_12_valid;
  wire [4:0]  input_12_bits_vs_0 = input_12_bits_vs;
  wire [1:0]  input_12_bits_offset_0 = input_12_bits_offset;
  wire [3:0]  input_12_bits_readLane_0 = input_12_bits_readLane;
  wire [1:0]  input_12_bits_dataOffset_0 = input_12_bits_dataOffset;
  wire        input_13_valid_0 = input_13_valid;
  wire [4:0]  input_13_bits_vs_0 = input_13_bits_vs;
  wire [1:0]  input_13_bits_offset_0 = input_13_bits_offset;
  wire [3:0]  input_13_bits_readLane_0 = input_13_bits_readLane;
  wire [1:0]  input_13_bits_dataOffset_0 = input_13_bits_dataOffset;
  wire        input_14_valid_0 = input_14_valid;
  wire [4:0]  input_14_bits_vs_0 = input_14_bits_vs;
  wire [1:0]  input_14_bits_offset_0 = input_14_bits_offset;
  wire [3:0]  input_14_bits_readLane_0 = input_14_bits_readLane;
  wire [1:0]  input_14_bits_dataOffset_0 = input_14_bits_dataOffset;
  wire        input_15_valid_0 = input_15_valid;
  wire [4:0]  input_15_bits_vs_0 = input_15_bits_vs;
  wire [1:0]  input_15_bits_offset_0 = input_15_bits_offset;
  wire [3:0]  input_15_bits_readLane_0 = input_15_bits_readLane;
  wire [1:0]  input_15_bits_dataOffset_0 = input_15_bits_dataOffset;
  wire        output_0_ready_0 = output_0_ready;
  wire        output_1_ready_0 = output_1_ready;
  wire        output_2_ready_0 = output_2_ready;
  wire        output_3_ready_0 = output_3_ready;
  wire        output_4_ready_0 = output_4_ready;
  wire        output_5_ready_0 = output_5_ready;
  wire        output_6_ready_0 = output_6_ready;
  wire        output_7_ready_0 = output_7_ready;
  wire        output_8_ready_0 = output_8_ready;
  wire        output_9_ready_0 = output_9_ready;
  wire        output_10_ready_0 = output_10_ready;
  wire        output_11_ready_0 = output_11_ready;
  wire        output_12_ready_0 = output_12_ready;
  wire        output_13_ready_0 = output_13_ready;
  wire        output_14_ready_0 = output_14_ready;
  wire        output_15_ready_0 = output_15_ready;
  wire [3:0]  input_15_bits_requestIndex = 4'hF;
  wire [3:0]  input_14_bits_requestIndex = 4'hE;
  wire [3:0]  input_13_bits_requestIndex = 4'hD;
  wire [3:0]  input_12_bits_requestIndex = 4'hC;
  wire [3:0]  input_11_bits_requestIndex = 4'hB;
  wire [3:0]  input_10_bits_requestIndex = 4'hA;
  wire [3:0]  input_9_bits_requestIndex = 4'h9;
  wire [3:0]  input_8_bits_requestIndex = 4'h8;
  wire [3:0]  input_7_bits_requestIndex = 4'h7;
  wire [3:0]  input_6_bits_requestIndex = 4'h6;
  wire [3:0]  input_5_bits_requestIndex = 4'h5;
  wire [3:0]  input_4_bits_requestIndex = 4'h4;
  wire [3:0]  input_3_bits_requestIndex = 4'h3;
  wire [3:0]  input_2_bits_requestIndex = 4'h2;
  wire [3:0]  input_1_bits_requestIndex = 4'h1;
  wire [3:0]  input_0_bits_requestIndex = 4'h0;
  wire [4:0]  selectReq_bits_vs;
  wire [1:0]  selectReq_bits_offset;
  wire [3:0]  selectReq_bits_requestIndex;
  wire [1:0]  selectReq_bits_dataOffset;
  wire [4:0]  selectReq_1_bits_vs;
  wire [1:0]  selectReq_1_bits_offset;
  wire [3:0]  selectReq_1_bits_requestIndex;
  wire [1:0]  selectReq_1_bits_dataOffset;
  wire [4:0]  selectReq_2_bits_vs;
  wire [1:0]  selectReq_2_bits_offset;
  wire [3:0]  selectReq_2_bits_requestIndex;
  wire [1:0]  selectReq_2_bits_dataOffset;
  wire [4:0]  selectReq_3_bits_vs;
  wire [1:0]  selectReq_3_bits_offset;
  wire [3:0]  selectReq_3_bits_requestIndex;
  wire [1:0]  selectReq_3_bits_dataOffset;
  wire [4:0]  selectReq_4_bits_vs;
  wire [1:0]  selectReq_4_bits_offset;
  wire [3:0]  selectReq_4_bits_requestIndex;
  wire [1:0]  selectReq_4_bits_dataOffset;
  wire [4:0]  selectReq_5_bits_vs;
  wire [1:0]  selectReq_5_bits_offset;
  wire [3:0]  selectReq_5_bits_requestIndex;
  wire [1:0]  selectReq_5_bits_dataOffset;
  wire [4:0]  selectReq_6_bits_vs;
  wire [1:0]  selectReq_6_bits_offset;
  wire [3:0]  selectReq_6_bits_requestIndex;
  wire [1:0]  selectReq_6_bits_dataOffset;
  wire [4:0]  selectReq_7_bits_vs;
  wire [1:0]  selectReq_7_bits_offset;
  wire [3:0]  selectReq_7_bits_requestIndex;
  wire [1:0]  selectReq_7_bits_dataOffset;
  wire [4:0]  selectReq_8_bits_vs;
  wire [1:0]  selectReq_8_bits_offset;
  wire [3:0]  selectReq_8_bits_requestIndex;
  wire [1:0]  selectReq_8_bits_dataOffset;
  wire [4:0]  selectReq_9_bits_vs;
  wire [1:0]  selectReq_9_bits_offset;
  wire [3:0]  selectReq_9_bits_requestIndex;
  wire [1:0]  selectReq_9_bits_dataOffset;
  wire [4:0]  selectReq_10_bits_vs;
  wire [1:0]  selectReq_10_bits_offset;
  wire [3:0]  selectReq_10_bits_requestIndex;
  wire [1:0]  selectReq_10_bits_dataOffset;
  wire [4:0]  selectReq_11_bits_vs;
  wire [1:0]  selectReq_11_bits_offset;
  wire [3:0]  selectReq_11_bits_requestIndex;
  wire [1:0]  selectReq_11_bits_dataOffset;
  wire [4:0]  selectReq_12_bits_vs;
  wire [1:0]  selectReq_12_bits_offset;
  wire [3:0]  selectReq_12_bits_requestIndex;
  wire [1:0]  selectReq_12_bits_dataOffset;
  wire [4:0]  selectReq_13_bits_vs;
  wire [1:0]  selectReq_13_bits_offset;
  wire [3:0]  selectReq_13_bits_requestIndex;
  wire [1:0]  selectReq_13_bits_dataOffset;
  wire [4:0]  selectReq_14_bits_vs;
  wire [1:0]  selectReq_14_bits_offset;
  wire [3:0]  selectReq_14_bits_requestIndex;
  wire [1:0]  selectReq_14_bits_dataOffset;
  wire [4:0]  selectReq_15_bits_vs;
  wire [1:0]  selectReq_15_bits_offset;
  wire [3:0]  selectReq_15_bits_requestIndex;
  wire [1:0]  selectReq_15_bits_dataOffset;
  wire [15:0] requestReadLane = 16'h1 << input_0_bits_readLane_0;
  wire        free = |requestReadLane;
  wire        outReady =
    requestReadLane[0] & output_0_ready_0 | requestReadLane[1] & output_1_ready_0 | requestReadLane[2] & output_2_ready_0 | requestReadLane[3] & output_3_ready_0 | requestReadLane[4] & output_4_ready_0 | requestReadLane[5]
    & output_5_ready_0 | requestReadLane[6] & output_6_ready_0 | requestReadLane[7] & output_7_ready_0 | requestReadLane[8] & output_8_ready_0 | requestReadLane[9] & output_9_ready_0 | requestReadLane[10] & output_10_ready_0
    | requestReadLane[11] & output_11_ready_0 | requestReadLane[12] & output_12_ready_0 | requestReadLane[13] & output_13_ready_0 | requestReadLane[14] & output_14_ready_0 | requestReadLane[15] & output_15_ready_0;
  wire        input_0_ready_0 = free & outReady;
  wire [15:0] inputSelect1H_0 = input_0_valid_0 & free ? requestReadLane : 16'h0;
  wire [15:0] requestReadLane_1 = 16'h1 << input_1_bits_readLane_0;
  wire        free_1 = |(requestReadLane_1 & ~inputSelect1H_0);
  wire        outReady_1 =
    requestReadLane_1[0] & output_0_ready_0 | requestReadLane_1[1] & output_1_ready_0 | requestReadLane_1[2] & output_2_ready_0 | requestReadLane_1[3] & output_3_ready_0 | requestReadLane_1[4] & output_4_ready_0 | requestReadLane_1[5]
    & output_5_ready_0 | requestReadLane_1[6] & output_6_ready_0 | requestReadLane_1[7] & output_7_ready_0 | requestReadLane_1[8] & output_8_ready_0 | requestReadLane_1[9] & output_9_ready_0 | requestReadLane_1[10] & output_10_ready_0
    | requestReadLane_1[11] & output_11_ready_0 | requestReadLane_1[12] & output_12_ready_0 | requestReadLane_1[13] & output_13_ready_0 | requestReadLane_1[14] & output_14_ready_0 | requestReadLane_1[15] & output_15_ready_0;
  wire        input_1_ready_0 = free_1 & outReady_1;
  wire [15:0] inputSelect1H_1 = input_1_valid_0 & free_1 ? requestReadLane_1 : 16'h0;
  wire [15:0] _GEN = inputSelect1H_0 | inputSelect1H_1;
  wire [15:0] requestReadLane_2 = 16'h1 << input_2_bits_readLane_0;
  wire        free_2 = |(requestReadLane_2 & ~_GEN);
  wire        outReady_2 =
    requestReadLane_2[0] & output_0_ready_0 | requestReadLane_2[1] & output_1_ready_0 | requestReadLane_2[2] & output_2_ready_0 | requestReadLane_2[3] & output_3_ready_0 | requestReadLane_2[4] & output_4_ready_0 | requestReadLane_2[5]
    & output_5_ready_0 | requestReadLane_2[6] & output_6_ready_0 | requestReadLane_2[7] & output_7_ready_0 | requestReadLane_2[8] & output_8_ready_0 | requestReadLane_2[9] & output_9_ready_0 | requestReadLane_2[10] & output_10_ready_0
    | requestReadLane_2[11] & output_11_ready_0 | requestReadLane_2[12] & output_12_ready_0 | requestReadLane_2[13] & output_13_ready_0 | requestReadLane_2[14] & output_14_ready_0 | requestReadLane_2[15] & output_15_ready_0;
  wire        input_2_ready_0 = free_2 & outReady_2;
  wire [15:0] inputSelect1H_2 = input_2_valid_0 & free_2 ? requestReadLane_2 : 16'h0;
  wire [15:0] _GEN_0 = _GEN | inputSelect1H_2;
  wire [15:0] requestReadLane_3 = 16'h1 << input_3_bits_readLane_0;
  wire        free_3 = |(requestReadLane_3 & ~_GEN_0);
  wire        outReady_3 =
    requestReadLane_3[0] & output_0_ready_0 | requestReadLane_3[1] & output_1_ready_0 | requestReadLane_3[2] & output_2_ready_0 | requestReadLane_3[3] & output_3_ready_0 | requestReadLane_3[4] & output_4_ready_0 | requestReadLane_3[5]
    & output_5_ready_0 | requestReadLane_3[6] & output_6_ready_0 | requestReadLane_3[7] & output_7_ready_0 | requestReadLane_3[8] & output_8_ready_0 | requestReadLane_3[9] & output_9_ready_0 | requestReadLane_3[10] & output_10_ready_0
    | requestReadLane_3[11] & output_11_ready_0 | requestReadLane_3[12] & output_12_ready_0 | requestReadLane_3[13] & output_13_ready_0 | requestReadLane_3[14] & output_14_ready_0 | requestReadLane_3[15] & output_15_ready_0;
  wire        input_3_ready_0 = free_3 & outReady_3;
  wire [15:0] inputSelect1H_3 = input_3_valid_0 & free_3 ? requestReadLane_3 : 16'h0;
  wire [15:0] _GEN_1 = _GEN_0 | inputSelect1H_3;
  wire [15:0] requestReadLane_4 = 16'h1 << input_4_bits_readLane_0;
  wire        free_4 = |(requestReadLane_4 & ~_GEN_1);
  wire        outReady_4 =
    requestReadLane_4[0] & output_0_ready_0 | requestReadLane_4[1] & output_1_ready_0 | requestReadLane_4[2] & output_2_ready_0 | requestReadLane_4[3] & output_3_ready_0 | requestReadLane_4[4] & output_4_ready_0 | requestReadLane_4[5]
    & output_5_ready_0 | requestReadLane_4[6] & output_6_ready_0 | requestReadLane_4[7] & output_7_ready_0 | requestReadLane_4[8] & output_8_ready_0 | requestReadLane_4[9] & output_9_ready_0 | requestReadLane_4[10] & output_10_ready_0
    | requestReadLane_4[11] & output_11_ready_0 | requestReadLane_4[12] & output_12_ready_0 | requestReadLane_4[13] & output_13_ready_0 | requestReadLane_4[14] & output_14_ready_0 | requestReadLane_4[15] & output_15_ready_0;
  wire        input_4_ready_0 = free_4 & outReady_4;
  wire [15:0] inputSelect1H_4 = input_4_valid_0 & free_4 ? requestReadLane_4 : 16'h0;
  wire [15:0] _GEN_2 = _GEN_1 | inputSelect1H_4;
  wire [15:0] requestReadLane_5 = 16'h1 << input_5_bits_readLane_0;
  wire        free_5 = |(requestReadLane_5 & ~_GEN_2);
  wire        outReady_5 =
    requestReadLane_5[0] & output_0_ready_0 | requestReadLane_5[1] & output_1_ready_0 | requestReadLane_5[2] & output_2_ready_0 | requestReadLane_5[3] & output_3_ready_0 | requestReadLane_5[4] & output_4_ready_0 | requestReadLane_5[5]
    & output_5_ready_0 | requestReadLane_5[6] & output_6_ready_0 | requestReadLane_5[7] & output_7_ready_0 | requestReadLane_5[8] & output_8_ready_0 | requestReadLane_5[9] & output_9_ready_0 | requestReadLane_5[10] & output_10_ready_0
    | requestReadLane_5[11] & output_11_ready_0 | requestReadLane_5[12] & output_12_ready_0 | requestReadLane_5[13] & output_13_ready_0 | requestReadLane_5[14] & output_14_ready_0 | requestReadLane_5[15] & output_15_ready_0;
  wire        input_5_ready_0 = free_5 & outReady_5;
  wire [15:0] inputSelect1H_5 = input_5_valid_0 & free_5 ? requestReadLane_5 : 16'h0;
  wire [15:0] _GEN_3 = _GEN_2 | inputSelect1H_5;
  wire [15:0] requestReadLane_6 = 16'h1 << input_6_bits_readLane_0;
  wire        free_6 = |(requestReadLane_6 & ~_GEN_3);
  wire        outReady_6 =
    requestReadLane_6[0] & output_0_ready_0 | requestReadLane_6[1] & output_1_ready_0 | requestReadLane_6[2] & output_2_ready_0 | requestReadLane_6[3] & output_3_ready_0 | requestReadLane_6[4] & output_4_ready_0 | requestReadLane_6[5]
    & output_5_ready_0 | requestReadLane_6[6] & output_6_ready_0 | requestReadLane_6[7] & output_7_ready_0 | requestReadLane_6[8] & output_8_ready_0 | requestReadLane_6[9] & output_9_ready_0 | requestReadLane_6[10] & output_10_ready_0
    | requestReadLane_6[11] & output_11_ready_0 | requestReadLane_6[12] & output_12_ready_0 | requestReadLane_6[13] & output_13_ready_0 | requestReadLane_6[14] & output_14_ready_0 | requestReadLane_6[15] & output_15_ready_0;
  wire        input_6_ready_0 = free_6 & outReady_6;
  wire [15:0] inputSelect1H_6 = input_6_valid_0 & free_6 ? requestReadLane_6 : 16'h0;
  wire [15:0] _GEN_4 = _GEN_3 | inputSelect1H_6;
  wire [15:0] requestReadLane_7 = 16'h1 << input_7_bits_readLane_0;
  wire        free_7 = |(requestReadLane_7 & ~_GEN_4);
  wire        outReady_7 =
    requestReadLane_7[0] & output_0_ready_0 | requestReadLane_7[1] & output_1_ready_0 | requestReadLane_7[2] & output_2_ready_0 | requestReadLane_7[3] & output_3_ready_0 | requestReadLane_7[4] & output_4_ready_0 | requestReadLane_7[5]
    & output_5_ready_0 | requestReadLane_7[6] & output_6_ready_0 | requestReadLane_7[7] & output_7_ready_0 | requestReadLane_7[8] & output_8_ready_0 | requestReadLane_7[9] & output_9_ready_0 | requestReadLane_7[10] & output_10_ready_0
    | requestReadLane_7[11] & output_11_ready_0 | requestReadLane_7[12] & output_12_ready_0 | requestReadLane_7[13] & output_13_ready_0 | requestReadLane_7[14] & output_14_ready_0 | requestReadLane_7[15] & output_15_ready_0;
  wire        input_7_ready_0 = free_7 & outReady_7;
  wire [15:0] inputSelect1H_7 = input_7_valid_0 & free_7 ? requestReadLane_7 : 16'h0;
  wire [15:0] _GEN_5 = _GEN_4 | inputSelect1H_7;
  wire [15:0] requestReadLane_8 = 16'h1 << input_8_bits_readLane_0;
  wire        free_8 = |(requestReadLane_8 & ~_GEN_5);
  wire        outReady_8 =
    requestReadLane_8[0] & output_0_ready_0 | requestReadLane_8[1] & output_1_ready_0 | requestReadLane_8[2] & output_2_ready_0 | requestReadLane_8[3] & output_3_ready_0 | requestReadLane_8[4] & output_4_ready_0 | requestReadLane_8[5]
    & output_5_ready_0 | requestReadLane_8[6] & output_6_ready_0 | requestReadLane_8[7] & output_7_ready_0 | requestReadLane_8[8] & output_8_ready_0 | requestReadLane_8[9] & output_9_ready_0 | requestReadLane_8[10] & output_10_ready_0
    | requestReadLane_8[11] & output_11_ready_0 | requestReadLane_8[12] & output_12_ready_0 | requestReadLane_8[13] & output_13_ready_0 | requestReadLane_8[14] & output_14_ready_0 | requestReadLane_8[15] & output_15_ready_0;
  wire        input_8_ready_0 = free_8 & outReady_8;
  wire [15:0] inputSelect1H_8 = input_8_valid_0 & free_8 ? requestReadLane_8 : 16'h0;
  wire [15:0] _GEN_6 = _GEN_5 | inputSelect1H_8;
  wire [15:0] requestReadLane_9 = 16'h1 << input_9_bits_readLane_0;
  wire        free_9 = |(requestReadLane_9 & ~_GEN_6);
  wire        outReady_9 =
    requestReadLane_9[0] & output_0_ready_0 | requestReadLane_9[1] & output_1_ready_0 | requestReadLane_9[2] & output_2_ready_0 | requestReadLane_9[3] & output_3_ready_0 | requestReadLane_9[4] & output_4_ready_0 | requestReadLane_9[5]
    & output_5_ready_0 | requestReadLane_9[6] & output_6_ready_0 | requestReadLane_9[7] & output_7_ready_0 | requestReadLane_9[8] & output_8_ready_0 | requestReadLane_9[9] & output_9_ready_0 | requestReadLane_9[10] & output_10_ready_0
    | requestReadLane_9[11] & output_11_ready_0 | requestReadLane_9[12] & output_12_ready_0 | requestReadLane_9[13] & output_13_ready_0 | requestReadLane_9[14] & output_14_ready_0 | requestReadLane_9[15] & output_15_ready_0;
  wire        input_9_ready_0 = free_9 & outReady_9;
  wire [15:0] inputSelect1H_9 = input_9_valid_0 & free_9 ? requestReadLane_9 : 16'h0;
  wire [15:0] _GEN_7 = _GEN_6 | inputSelect1H_9;
  wire [15:0] requestReadLane_10 = 16'h1 << input_10_bits_readLane_0;
  wire        free_10 = |(requestReadLane_10 & ~_GEN_7);
  wire        outReady_10 =
    requestReadLane_10[0] & output_0_ready_0 | requestReadLane_10[1] & output_1_ready_0 | requestReadLane_10[2] & output_2_ready_0 | requestReadLane_10[3] & output_3_ready_0 | requestReadLane_10[4] & output_4_ready_0 | requestReadLane_10[5]
    & output_5_ready_0 | requestReadLane_10[6] & output_6_ready_0 | requestReadLane_10[7] & output_7_ready_0 | requestReadLane_10[8] & output_8_ready_0 | requestReadLane_10[9] & output_9_ready_0 | requestReadLane_10[10] & output_10_ready_0
    | requestReadLane_10[11] & output_11_ready_0 | requestReadLane_10[12] & output_12_ready_0 | requestReadLane_10[13] & output_13_ready_0 | requestReadLane_10[14] & output_14_ready_0 | requestReadLane_10[15] & output_15_ready_0;
  wire        input_10_ready_0 = free_10 & outReady_10;
  wire [15:0] inputSelect1H_10 = input_10_valid_0 & free_10 ? requestReadLane_10 : 16'h0;
  wire [15:0] _GEN_8 = _GEN_7 | inputSelect1H_10;
  wire [15:0] requestReadLane_11 = 16'h1 << input_11_bits_readLane_0;
  wire        free_11 = |(requestReadLane_11 & ~_GEN_8);
  wire        outReady_11 =
    requestReadLane_11[0] & output_0_ready_0 | requestReadLane_11[1] & output_1_ready_0 | requestReadLane_11[2] & output_2_ready_0 | requestReadLane_11[3] & output_3_ready_0 | requestReadLane_11[4] & output_4_ready_0 | requestReadLane_11[5]
    & output_5_ready_0 | requestReadLane_11[6] & output_6_ready_0 | requestReadLane_11[7] & output_7_ready_0 | requestReadLane_11[8] & output_8_ready_0 | requestReadLane_11[9] & output_9_ready_0 | requestReadLane_11[10] & output_10_ready_0
    | requestReadLane_11[11] & output_11_ready_0 | requestReadLane_11[12] & output_12_ready_0 | requestReadLane_11[13] & output_13_ready_0 | requestReadLane_11[14] & output_14_ready_0 | requestReadLane_11[15] & output_15_ready_0;
  wire        input_11_ready_0 = free_11 & outReady_11;
  wire [15:0] inputSelect1H_11 = input_11_valid_0 & free_11 ? requestReadLane_11 : 16'h0;
  wire [15:0] _GEN_9 = _GEN_8 | inputSelect1H_11;
  wire [15:0] requestReadLane_12 = 16'h1 << input_12_bits_readLane_0;
  wire        free_12 = |(requestReadLane_12 & ~_GEN_9);
  wire        outReady_12 =
    requestReadLane_12[0] & output_0_ready_0 | requestReadLane_12[1] & output_1_ready_0 | requestReadLane_12[2] & output_2_ready_0 | requestReadLane_12[3] & output_3_ready_0 | requestReadLane_12[4] & output_4_ready_0 | requestReadLane_12[5]
    & output_5_ready_0 | requestReadLane_12[6] & output_6_ready_0 | requestReadLane_12[7] & output_7_ready_0 | requestReadLane_12[8] & output_8_ready_0 | requestReadLane_12[9] & output_9_ready_0 | requestReadLane_12[10] & output_10_ready_0
    | requestReadLane_12[11] & output_11_ready_0 | requestReadLane_12[12] & output_12_ready_0 | requestReadLane_12[13] & output_13_ready_0 | requestReadLane_12[14] & output_14_ready_0 | requestReadLane_12[15] & output_15_ready_0;
  wire        input_12_ready_0 = free_12 & outReady_12;
  wire [15:0] inputSelect1H_12 = input_12_valid_0 & free_12 ? requestReadLane_12 : 16'h0;
  wire [15:0] _GEN_10 = _GEN_9 | inputSelect1H_12;
  wire [15:0] requestReadLane_13 = 16'h1 << input_13_bits_readLane_0;
  wire        free_13 = |(requestReadLane_13 & ~_GEN_10);
  wire        outReady_13 =
    requestReadLane_13[0] & output_0_ready_0 | requestReadLane_13[1] & output_1_ready_0 | requestReadLane_13[2] & output_2_ready_0 | requestReadLane_13[3] & output_3_ready_0 | requestReadLane_13[4] & output_4_ready_0 | requestReadLane_13[5]
    & output_5_ready_0 | requestReadLane_13[6] & output_6_ready_0 | requestReadLane_13[7] & output_7_ready_0 | requestReadLane_13[8] & output_8_ready_0 | requestReadLane_13[9] & output_9_ready_0 | requestReadLane_13[10] & output_10_ready_0
    | requestReadLane_13[11] & output_11_ready_0 | requestReadLane_13[12] & output_12_ready_0 | requestReadLane_13[13] & output_13_ready_0 | requestReadLane_13[14] & output_14_ready_0 | requestReadLane_13[15] & output_15_ready_0;
  wire        input_13_ready_0 = free_13 & outReady_13;
  wire [15:0] inputSelect1H_13 = input_13_valid_0 & free_13 ? requestReadLane_13 : 16'h0;
  wire [15:0] _GEN_11 = _GEN_10 | inputSelect1H_13;
  wire [15:0] requestReadLane_14 = 16'h1 << input_14_bits_readLane_0;
  wire        free_14 = |(requestReadLane_14 & ~_GEN_11);
  wire        outReady_14 =
    requestReadLane_14[0] & output_0_ready_0 | requestReadLane_14[1] & output_1_ready_0 | requestReadLane_14[2] & output_2_ready_0 | requestReadLane_14[3] & output_3_ready_0 | requestReadLane_14[4] & output_4_ready_0 | requestReadLane_14[5]
    & output_5_ready_0 | requestReadLane_14[6] & output_6_ready_0 | requestReadLane_14[7] & output_7_ready_0 | requestReadLane_14[8] & output_8_ready_0 | requestReadLane_14[9] & output_9_ready_0 | requestReadLane_14[10] & output_10_ready_0
    | requestReadLane_14[11] & output_11_ready_0 | requestReadLane_14[12] & output_12_ready_0 | requestReadLane_14[13] & output_13_ready_0 | requestReadLane_14[14] & output_14_ready_0 | requestReadLane_14[15] & output_15_ready_0;
  wire        input_14_ready_0 = free_14 & outReady_14;
  wire [15:0] inputSelect1H_14 = input_14_valid_0 & free_14 ? requestReadLane_14 : 16'h0;
  wire [15:0] requestReadLane_15 = 16'h1 << input_15_bits_readLane_0;
  wire        free_15 = |(requestReadLane_15 & ~(_GEN_11 | inputSelect1H_14));
  wire        outReady_15 =
    requestReadLane_15[0] & output_0_ready_0 | requestReadLane_15[1] & output_1_ready_0 | requestReadLane_15[2] & output_2_ready_0 | requestReadLane_15[3] & output_3_ready_0 | requestReadLane_15[4] & output_4_ready_0 | requestReadLane_15[5]
    & output_5_ready_0 | requestReadLane_15[6] & output_6_ready_0 | requestReadLane_15[7] & output_7_ready_0 | requestReadLane_15[8] & output_8_ready_0 | requestReadLane_15[9] & output_9_ready_0 | requestReadLane_15[10] & output_10_ready_0
    | requestReadLane_15[11] & output_11_ready_0 | requestReadLane_15[12] & output_12_ready_0 | requestReadLane_15[13] & output_13_ready_0 | requestReadLane_15[14] & output_14_ready_0 | requestReadLane_15[15] & output_15_ready_0;
  wire        input_15_ready_0 = free_15 & outReady_15;
  wire [15:0] inputSelect1H_15 = input_15_valid_0 & free_15 ? requestReadLane_15 : 16'h0;
  wire [1:0]  tryToRead_lo_lo_lo = {inputSelect1H_1[0], inputSelect1H_0[0]};
  wire [1:0]  tryToRead_lo_lo_hi = {inputSelect1H_3[0], inputSelect1H_2[0]};
  wire [3:0]  tryToRead_lo_lo = {tryToRead_lo_lo_hi, tryToRead_lo_lo_lo};
  wire [1:0]  tryToRead_lo_hi_lo = {inputSelect1H_5[0], inputSelect1H_4[0]};
  wire [1:0]  tryToRead_lo_hi_hi = {inputSelect1H_7[0], inputSelect1H_6[0]};
  wire [3:0]  tryToRead_lo_hi = {tryToRead_lo_hi_hi, tryToRead_lo_hi_lo};
  wire [7:0]  tryToRead_lo = {tryToRead_lo_hi, tryToRead_lo_lo};
  wire [1:0]  tryToRead_hi_lo_lo = {inputSelect1H_9[0], inputSelect1H_8[0]};
  wire [1:0]  tryToRead_hi_lo_hi = {inputSelect1H_11[0], inputSelect1H_10[0]};
  wire [3:0]  tryToRead_hi_lo = {tryToRead_hi_lo_hi, tryToRead_hi_lo_lo};
  wire [1:0]  tryToRead_hi_hi_lo = {inputSelect1H_13[0], inputSelect1H_12[0]};
  wire [1:0]  tryToRead_hi_hi_hi = {inputSelect1H_15[0], inputSelect1H_14[0]};
  wire [3:0]  tryToRead_hi_hi = {tryToRead_hi_hi_hi, tryToRead_hi_hi_lo};
  wire [7:0]  tryToRead_hi = {tryToRead_hi_hi, tryToRead_hi_lo};
  wire [15:0] tryToRead = {tryToRead_hi, tryToRead_lo};
  wire        output_0_valid_0 = |tryToRead;
  wire [4:0]  output_0_bits_vs_0 = selectReq_bits_vs;
  wire [1:0]  output_0_bits_offset_0 = selectReq_bits_offset;
  wire [3:0]  output_0_bits_writeIndex_0 = selectReq_bits_requestIndex;
  wire [1:0]  output_0_bits_dataOffset_0 = selectReq_bits_dataOffset;
  assign selectReq_bits_dataOffset =
    (tryToRead[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead[15] ? input_15_bits_dataOffset_0 : 2'h0);
  assign selectReq_bits_requestIndex =
    {3'h0, tryToRead[1]} | {2'h0, tryToRead[2], 1'h0} | (tryToRead[3] ? 4'h3 : 4'h0) | {1'h0, tryToRead[4], 2'h0} | (tryToRead[5] ? 4'h5 : 4'h0) | (tryToRead[6] ? 4'h6 : 4'h0) | (tryToRead[7] ? 4'h7 : 4'h0) | {tryToRead[8], 3'h0}
    | (tryToRead[9] ? 4'h9 : 4'h0) | (tryToRead[10] ? 4'hA : 4'h0) | (tryToRead[11] ? 4'hB : 4'h0) | (tryToRead[12] ? 4'hC : 4'h0) | (tryToRead[13] ? 4'hD : 4'h0) | (tryToRead[14] ? 4'hE : 4'h0) | {4{tryToRead[15]}};
  wire [3:0]  selectReq_bits_readLane =
    (tryToRead[0] ? input_0_bits_readLane_0 : 4'h0) | (tryToRead[1] ? input_1_bits_readLane_0 : 4'h0) | (tryToRead[2] ? input_2_bits_readLane_0 : 4'h0) | (tryToRead[3] ? input_3_bits_readLane_0 : 4'h0)
    | (tryToRead[4] ? input_4_bits_readLane_0 : 4'h0) | (tryToRead[5] ? input_5_bits_readLane_0 : 4'h0) | (tryToRead[6] ? input_6_bits_readLane_0 : 4'h0) | (tryToRead[7] ? input_7_bits_readLane_0 : 4'h0)
    | (tryToRead[8] ? input_8_bits_readLane_0 : 4'h0) | (tryToRead[9] ? input_9_bits_readLane_0 : 4'h0) | (tryToRead[10] ? input_10_bits_readLane_0 : 4'h0) | (tryToRead[11] ? input_11_bits_readLane_0 : 4'h0)
    | (tryToRead[12] ? input_12_bits_readLane_0 : 4'h0) | (tryToRead[13] ? input_13_bits_readLane_0 : 4'h0) | (tryToRead[14] ? input_14_bits_readLane_0 : 4'h0) | (tryToRead[15] ? input_15_bits_readLane_0 : 4'h0);
  assign selectReq_bits_offset =
    (tryToRead[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead[7] ? input_7_bits_offset_0 : 2'h0)
    | (tryToRead[8] ? input_8_bits_offset_0 : 2'h0) | (tryToRead[9] ? input_9_bits_offset_0 : 2'h0) | (tryToRead[10] ? input_10_bits_offset_0 : 2'h0) | (tryToRead[11] ? input_11_bits_offset_0 : 2'h0)
    | (tryToRead[12] ? input_12_bits_offset_0 : 2'h0) | (tryToRead[13] ? input_13_bits_offset_0 : 2'h0) | (tryToRead[14] ? input_14_bits_offset_0 : 2'h0) | (tryToRead[15] ? input_15_bits_offset_0 : 2'h0);
  assign selectReq_bits_vs =
    (tryToRead[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead[13] ? input_13_bits_vs_0 : 5'h0) | (tryToRead[14] ? input_14_bits_vs_0 : 5'h0)
    | (tryToRead[15] ? input_15_bits_vs_0 : 5'h0);
  wire        selectReq_valid =
    tryToRead[0] & input_0_valid_0 | tryToRead[1] & input_1_valid_0 | tryToRead[2] & input_2_valid_0 | tryToRead[3] & input_3_valid_0 | tryToRead[4] & input_4_valid_0 | tryToRead[5] & input_5_valid_0 | tryToRead[6] & input_6_valid_0
    | tryToRead[7] & input_7_valid_0 | tryToRead[8] & input_8_valid_0 | tryToRead[9] & input_9_valid_0 | tryToRead[10] & input_10_valid_0 | tryToRead[11] & input_11_valid_0 | tryToRead[12] & input_12_valid_0 | tryToRead[13]
    & input_13_valid_0 | tryToRead[14] & input_14_valid_0 | tryToRead[15] & input_15_valid_0;
  wire        selectReq_ready =
    tryToRead[0] & input_0_ready_0 | tryToRead[1] & input_1_ready_0 | tryToRead[2] & input_2_ready_0 | tryToRead[3] & input_3_ready_0 | tryToRead[4] & input_4_ready_0 | tryToRead[5] & input_5_ready_0 | tryToRead[6] & input_6_ready_0
    | tryToRead[7] & input_7_ready_0 | tryToRead[8] & input_8_ready_0 | tryToRead[9] & input_9_ready_0 | tryToRead[10] & input_10_ready_0 | tryToRead[11] & input_11_ready_0 | tryToRead[12] & input_12_ready_0 | tryToRead[13]
    & input_13_ready_0 | tryToRead[14] & input_14_ready_0 | tryToRead[15] & input_15_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_1 = {inputSelect1H_1[1], inputSelect1H_0[1]};
  wire [1:0]  tryToRead_lo_lo_hi_1 = {inputSelect1H_3[1], inputSelect1H_2[1]};
  wire [3:0]  tryToRead_lo_lo_1 = {tryToRead_lo_lo_hi_1, tryToRead_lo_lo_lo_1};
  wire [1:0]  tryToRead_lo_hi_lo_1 = {inputSelect1H_5[1], inputSelect1H_4[1]};
  wire [1:0]  tryToRead_lo_hi_hi_1 = {inputSelect1H_7[1], inputSelect1H_6[1]};
  wire [3:0]  tryToRead_lo_hi_1 = {tryToRead_lo_hi_hi_1, tryToRead_lo_hi_lo_1};
  wire [7:0]  tryToRead_lo_1 = {tryToRead_lo_hi_1, tryToRead_lo_lo_1};
  wire [1:0]  tryToRead_hi_lo_lo_1 = {inputSelect1H_9[1], inputSelect1H_8[1]};
  wire [1:0]  tryToRead_hi_lo_hi_1 = {inputSelect1H_11[1], inputSelect1H_10[1]};
  wire [3:0]  tryToRead_hi_lo_1 = {tryToRead_hi_lo_hi_1, tryToRead_hi_lo_lo_1};
  wire [1:0]  tryToRead_hi_hi_lo_1 = {inputSelect1H_13[1], inputSelect1H_12[1]};
  wire [1:0]  tryToRead_hi_hi_hi_1 = {inputSelect1H_15[1], inputSelect1H_14[1]};
  wire [3:0]  tryToRead_hi_hi_1 = {tryToRead_hi_hi_hi_1, tryToRead_hi_hi_lo_1};
  wire [7:0]  tryToRead_hi_1 = {tryToRead_hi_hi_1, tryToRead_hi_lo_1};
  wire [15:0] tryToRead_1 = {tryToRead_hi_1, tryToRead_lo_1};
  wire        output_1_valid_0 = |tryToRead_1;
  wire [4:0]  output_1_bits_vs_0 = selectReq_1_bits_vs;
  wire [1:0]  output_1_bits_offset_0 = selectReq_1_bits_offset;
  wire [3:0]  output_1_bits_writeIndex_0 = selectReq_1_bits_requestIndex;
  wire [1:0]  output_1_bits_dataOffset_0 = selectReq_1_bits_dataOffset;
  assign selectReq_1_bits_dataOffset =
    (tryToRead_1[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_1[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_1[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_1[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_1[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_1[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_1[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_1[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_1[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_1[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_1[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_1[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_1[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_1[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_1[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_1[15] ? input_15_bits_dataOffset_0 : 2'h0);
  assign selectReq_1_bits_requestIndex =
    {3'h0, tryToRead_1[1]} | {2'h0, tryToRead_1[2], 1'h0} | (tryToRead_1[3] ? 4'h3 : 4'h0) | {1'h0, tryToRead_1[4], 2'h0} | (tryToRead_1[5] ? 4'h5 : 4'h0) | (tryToRead_1[6] ? 4'h6 : 4'h0) | (tryToRead_1[7] ? 4'h7 : 4'h0)
    | {tryToRead_1[8], 3'h0} | (tryToRead_1[9] ? 4'h9 : 4'h0) | (tryToRead_1[10] ? 4'hA : 4'h0) | (tryToRead_1[11] ? 4'hB : 4'h0) | (tryToRead_1[12] ? 4'hC : 4'h0) | (tryToRead_1[13] ? 4'hD : 4'h0) | (tryToRead_1[14] ? 4'hE : 4'h0)
    | {4{tryToRead_1[15]}};
  wire [3:0]  selectReq_1_bits_readLane =
    (tryToRead_1[0] ? input_0_bits_readLane_0 : 4'h0) | (tryToRead_1[1] ? input_1_bits_readLane_0 : 4'h0) | (tryToRead_1[2] ? input_2_bits_readLane_0 : 4'h0) | (tryToRead_1[3] ? input_3_bits_readLane_0 : 4'h0)
    | (tryToRead_1[4] ? input_4_bits_readLane_0 : 4'h0) | (tryToRead_1[5] ? input_5_bits_readLane_0 : 4'h0) | (tryToRead_1[6] ? input_6_bits_readLane_0 : 4'h0) | (tryToRead_1[7] ? input_7_bits_readLane_0 : 4'h0)
    | (tryToRead_1[8] ? input_8_bits_readLane_0 : 4'h0) | (tryToRead_1[9] ? input_9_bits_readLane_0 : 4'h0) | (tryToRead_1[10] ? input_10_bits_readLane_0 : 4'h0) | (tryToRead_1[11] ? input_11_bits_readLane_0 : 4'h0)
    | (tryToRead_1[12] ? input_12_bits_readLane_0 : 4'h0) | (tryToRead_1[13] ? input_13_bits_readLane_0 : 4'h0) | (tryToRead_1[14] ? input_14_bits_readLane_0 : 4'h0) | (tryToRead_1[15] ? input_15_bits_readLane_0 : 4'h0);
  assign selectReq_1_bits_offset =
    (tryToRead_1[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead_1[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead_1[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead_1[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead_1[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead_1[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead_1[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead_1[7] ? input_7_bits_offset_0 : 2'h0)
    | (tryToRead_1[8] ? input_8_bits_offset_0 : 2'h0) | (tryToRead_1[9] ? input_9_bits_offset_0 : 2'h0) | (tryToRead_1[10] ? input_10_bits_offset_0 : 2'h0) | (tryToRead_1[11] ? input_11_bits_offset_0 : 2'h0)
    | (tryToRead_1[12] ? input_12_bits_offset_0 : 2'h0) | (tryToRead_1[13] ? input_13_bits_offset_0 : 2'h0) | (tryToRead_1[14] ? input_14_bits_offset_0 : 2'h0) | (tryToRead_1[15] ? input_15_bits_offset_0 : 2'h0);
  assign selectReq_1_bits_vs =
    (tryToRead_1[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_1[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_1[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_1[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_1[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_1[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_1[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_1[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_1[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_1[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_1[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_1[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_1[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_1[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_1[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_1[15] ? input_15_bits_vs_0 : 5'h0);
  wire        selectReq_1_valid =
    tryToRead_1[0] & input_0_valid_0 | tryToRead_1[1] & input_1_valid_0 | tryToRead_1[2] & input_2_valid_0 | tryToRead_1[3] & input_3_valid_0 | tryToRead_1[4] & input_4_valid_0 | tryToRead_1[5] & input_5_valid_0 | tryToRead_1[6]
    & input_6_valid_0 | tryToRead_1[7] & input_7_valid_0 | tryToRead_1[8] & input_8_valid_0 | tryToRead_1[9] & input_9_valid_0 | tryToRead_1[10] & input_10_valid_0 | tryToRead_1[11] & input_11_valid_0 | tryToRead_1[12] & input_12_valid_0
    | tryToRead_1[13] & input_13_valid_0 | tryToRead_1[14] & input_14_valid_0 | tryToRead_1[15] & input_15_valid_0;
  wire        selectReq_1_ready =
    tryToRead_1[0] & input_0_ready_0 | tryToRead_1[1] & input_1_ready_0 | tryToRead_1[2] & input_2_ready_0 | tryToRead_1[3] & input_3_ready_0 | tryToRead_1[4] & input_4_ready_0 | tryToRead_1[5] & input_5_ready_0 | tryToRead_1[6]
    & input_6_ready_0 | tryToRead_1[7] & input_7_ready_0 | tryToRead_1[8] & input_8_ready_0 | tryToRead_1[9] & input_9_ready_0 | tryToRead_1[10] & input_10_ready_0 | tryToRead_1[11] & input_11_ready_0 | tryToRead_1[12] & input_12_ready_0
    | tryToRead_1[13] & input_13_ready_0 | tryToRead_1[14] & input_14_ready_0 | tryToRead_1[15] & input_15_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_2 = {inputSelect1H_1[2], inputSelect1H_0[2]};
  wire [1:0]  tryToRead_lo_lo_hi_2 = {inputSelect1H_3[2], inputSelect1H_2[2]};
  wire [3:0]  tryToRead_lo_lo_2 = {tryToRead_lo_lo_hi_2, tryToRead_lo_lo_lo_2};
  wire [1:0]  tryToRead_lo_hi_lo_2 = {inputSelect1H_5[2], inputSelect1H_4[2]};
  wire [1:0]  tryToRead_lo_hi_hi_2 = {inputSelect1H_7[2], inputSelect1H_6[2]};
  wire [3:0]  tryToRead_lo_hi_2 = {tryToRead_lo_hi_hi_2, tryToRead_lo_hi_lo_2};
  wire [7:0]  tryToRead_lo_2 = {tryToRead_lo_hi_2, tryToRead_lo_lo_2};
  wire [1:0]  tryToRead_hi_lo_lo_2 = {inputSelect1H_9[2], inputSelect1H_8[2]};
  wire [1:0]  tryToRead_hi_lo_hi_2 = {inputSelect1H_11[2], inputSelect1H_10[2]};
  wire [3:0]  tryToRead_hi_lo_2 = {tryToRead_hi_lo_hi_2, tryToRead_hi_lo_lo_2};
  wire [1:0]  tryToRead_hi_hi_lo_2 = {inputSelect1H_13[2], inputSelect1H_12[2]};
  wire [1:0]  tryToRead_hi_hi_hi_2 = {inputSelect1H_15[2], inputSelect1H_14[2]};
  wire [3:0]  tryToRead_hi_hi_2 = {tryToRead_hi_hi_hi_2, tryToRead_hi_hi_lo_2};
  wire [7:0]  tryToRead_hi_2 = {tryToRead_hi_hi_2, tryToRead_hi_lo_2};
  wire [15:0] tryToRead_2 = {tryToRead_hi_2, tryToRead_lo_2};
  wire        output_2_valid_0 = |tryToRead_2;
  wire [4:0]  output_2_bits_vs_0 = selectReq_2_bits_vs;
  wire [1:0]  output_2_bits_offset_0 = selectReq_2_bits_offset;
  wire [3:0]  output_2_bits_writeIndex_0 = selectReq_2_bits_requestIndex;
  wire [1:0]  output_2_bits_dataOffset_0 = selectReq_2_bits_dataOffset;
  assign selectReq_2_bits_dataOffset =
    (tryToRead_2[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_2[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_2[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_2[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_2[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_2[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_2[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_2[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_2[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_2[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_2[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_2[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_2[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_2[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_2[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_2[15] ? input_15_bits_dataOffset_0 : 2'h0);
  assign selectReq_2_bits_requestIndex =
    {3'h0, tryToRead_2[1]} | {2'h0, tryToRead_2[2], 1'h0} | (tryToRead_2[3] ? 4'h3 : 4'h0) | {1'h0, tryToRead_2[4], 2'h0} | (tryToRead_2[5] ? 4'h5 : 4'h0) | (tryToRead_2[6] ? 4'h6 : 4'h0) | (tryToRead_2[7] ? 4'h7 : 4'h0)
    | {tryToRead_2[8], 3'h0} | (tryToRead_2[9] ? 4'h9 : 4'h0) | (tryToRead_2[10] ? 4'hA : 4'h0) | (tryToRead_2[11] ? 4'hB : 4'h0) | (tryToRead_2[12] ? 4'hC : 4'h0) | (tryToRead_2[13] ? 4'hD : 4'h0) | (tryToRead_2[14] ? 4'hE : 4'h0)
    | {4{tryToRead_2[15]}};
  wire [3:0]  selectReq_2_bits_readLane =
    (tryToRead_2[0] ? input_0_bits_readLane_0 : 4'h0) | (tryToRead_2[1] ? input_1_bits_readLane_0 : 4'h0) | (tryToRead_2[2] ? input_2_bits_readLane_0 : 4'h0) | (tryToRead_2[3] ? input_3_bits_readLane_0 : 4'h0)
    | (tryToRead_2[4] ? input_4_bits_readLane_0 : 4'h0) | (tryToRead_2[5] ? input_5_bits_readLane_0 : 4'h0) | (tryToRead_2[6] ? input_6_bits_readLane_0 : 4'h0) | (tryToRead_2[7] ? input_7_bits_readLane_0 : 4'h0)
    | (tryToRead_2[8] ? input_8_bits_readLane_0 : 4'h0) | (tryToRead_2[9] ? input_9_bits_readLane_0 : 4'h0) | (tryToRead_2[10] ? input_10_bits_readLane_0 : 4'h0) | (tryToRead_2[11] ? input_11_bits_readLane_0 : 4'h0)
    | (tryToRead_2[12] ? input_12_bits_readLane_0 : 4'h0) | (tryToRead_2[13] ? input_13_bits_readLane_0 : 4'h0) | (tryToRead_2[14] ? input_14_bits_readLane_0 : 4'h0) | (tryToRead_2[15] ? input_15_bits_readLane_0 : 4'h0);
  assign selectReq_2_bits_offset =
    (tryToRead_2[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead_2[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead_2[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead_2[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead_2[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead_2[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead_2[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead_2[7] ? input_7_bits_offset_0 : 2'h0)
    | (tryToRead_2[8] ? input_8_bits_offset_0 : 2'h0) | (tryToRead_2[9] ? input_9_bits_offset_0 : 2'h0) | (tryToRead_2[10] ? input_10_bits_offset_0 : 2'h0) | (tryToRead_2[11] ? input_11_bits_offset_0 : 2'h0)
    | (tryToRead_2[12] ? input_12_bits_offset_0 : 2'h0) | (tryToRead_2[13] ? input_13_bits_offset_0 : 2'h0) | (tryToRead_2[14] ? input_14_bits_offset_0 : 2'h0) | (tryToRead_2[15] ? input_15_bits_offset_0 : 2'h0);
  assign selectReq_2_bits_vs =
    (tryToRead_2[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_2[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_2[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_2[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_2[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_2[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_2[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_2[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_2[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_2[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_2[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_2[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_2[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_2[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_2[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_2[15] ? input_15_bits_vs_0 : 5'h0);
  wire        selectReq_2_valid =
    tryToRead_2[0] & input_0_valid_0 | tryToRead_2[1] & input_1_valid_0 | tryToRead_2[2] & input_2_valid_0 | tryToRead_2[3] & input_3_valid_0 | tryToRead_2[4] & input_4_valid_0 | tryToRead_2[5] & input_5_valid_0 | tryToRead_2[6]
    & input_6_valid_0 | tryToRead_2[7] & input_7_valid_0 | tryToRead_2[8] & input_8_valid_0 | tryToRead_2[9] & input_9_valid_0 | tryToRead_2[10] & input_10_valid_0 | tryToRead_2[11] & input_11_valid_0 | tryToRead_2[12] & input_12_valid_0
    | tryToRead_2[13] & input_13_valid_0 | tryToRead_2[14] & input_14_valid_0 | tryToRead_2[15] & input_15_valid_0;
  wire        selectReq_2_ready =
    tryToRead_2[0] & input_0_ready_0 | tryToRead_2[1] & input_1_ready_0 | tryToRead_2[2] & input_2_ready_0 | tryToRead_2[3] & input_3_ready_0 | tryToRead_2[4] & input_4_ready_0 | tryToRead_2[5] & input_5_ready_0 | tryToRead_2[6]
    & input_6_ready_0 | tryToRead_2[7] & input_7_ready_0 | tryToRead_2[8] & input_8_ready_0 | tryToRead_2[9] & input_9_ready_0 | tryToRead_2[10] & input_10_ready_0 | tryToRead_2[11] & input_11_ready_0 | tryToRead_2[12] & input_12_ready_0
    | tryToRead_2[13] & input_13_ready_0 | tryToRead_2[14] & input_14_ready_0 | tryToRead_2[15] & input_15_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_3 = {inputSelect1H_1[3], inputSelect1H_0[3]};
  wire [1:0]  tryToRead_lo_lo_hi_3 = {inputSelect1H_3[3], inputSelect1H_2[3]};
  wire [3:0]  tryToRead_lo_lo_3 = {tryToRead_lo_lo_hi_3, tryToRead_lo_lo_lo_3};
  wire [1:0]  tryToRead_lo_hi_lo_3 = {inputSelect1H_5[3], inputSelect1H_4[3]};
  wire [1:0]  tryToRead_lo_hi_hi_3 = {inputSelect1H_7[3], inputSelect1H_6[3]};
  wire [3:0]  tryToRead_lo_hi_3 = {tryToRead_lo_hi_hi_3, tryToRead_lo_hi_lo_3};
  wire [7:0]  tryToRead_lo_3 = {tryToRead_lo_hi_3, tryToRead_lo_lo_3};
  wire [1:0]  tryToRead_hi_lo_lo_3 = {inputSelect1H_9[3], inputSelect1H_8[3]};
  wire [1:0]  tryToRead_hi_lo_hi_3 = {inputSelect1H_11[3], inputSelect1H_10[3]};
  wire [3:0]  tryToRead_hi_lo_3 = {tryToRead_hi_lo_hi_3, tryToRead_hi_lo_lo_3};
  wire [1:0]  tryToRead_hi_hi_lo_3 = {inputSelect1H_13[3], inputSelect1H_12[3]};
  wire [1:0]  tryToRead_hi_hi_hi_3 = {inputSelect1H_15[3], inputSelect1H_14[3]};
  wire [3:0]  tryToRead_hi_hi_3 = {tryToRead_hi_hi_hi_3, tryToRead_hi_hi_lo_3};
  wire [7:0]  tryToRead_hi_3 = {tryToRead_hi_hi_3, tryToRead_hi_lo_3};
  wire [15:0] tryToRead_3 = {tryToRead_hi_3, tryToRead_lo_3};
  wire        output_3_valid_0 = |tryToRead_3;
  wire [4:0]  output_3_bits_vs_0 = selectReq_3_bits_vs;
  wire [1:0]  output_3_bits_offset_0 = selectReq_3_bits_offset;
  wire [3:0]  output_3_bits_writeIndex_0 = selectReq_3_bits_requestIndex;
  wire [1:0]  output_3_bits_dataOffset_0 = selectReq_3_bits_dataOffset;
  assign selectReq_3_bits_dataOffset =
    (tryToRead_3[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_3[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_3[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_3[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_3[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_3[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_3[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_3[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_3[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_3[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_3[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_3[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_3[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_3[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_3[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_3[15] ? input_15_bits_dataOffset_0 : 2'h0);
  assign selectReq_3_bits_requestIndex =
    {3'h0, tryToRead_3[1]} | {2'h0, tryToRead_3[2], 1'h0} | (tryToRead_3[3] ? 4'h3 : 4'h0) | {1'h0, tryToRead_3[4], 2'h0} | (tryToRead_3[5] ? 4'h5 : 4'h0) | (tryToRead_3[6] ? 4'h6 : 4'h0) | (tryToRead_3[7] ? 4'h7 : 4'h0)
    | {tryToRead_3[8], 3'h0} | (tryToRead_3[9] ? 4'h9 : 4'h0) | (tryToRead_3[10] ? 4'hA : 4'h0) | (tryToRead_3[11] ? 4'hB : 4'h0) | (tryToRead_3[12] ? 4'hC : 4'h0) | (tryToRead_3[13] ? 4'hD : 4'h0) | (tryToRead_3[14] ? 4'hE : 4'h0)
    | {4{tryToRead_3[15]}};
  wire [3:0]  selectReq_3_bits_readLane =
    (tryToRead_3[0] ? input_0_bits_readLane_0 : 4'h0) | (tryToRead_3[1] ? input_1_bits_readLane_0 : 4'h0) | (tryToRead_3[2] ? input_2_bits_readLane_0 : 4'h0) | (tryToRead_3[3] ? input_3_bits_readLane_0 : 4'h0)
    | (tryToRead_3[4] ? input_4_bits_readLane_0 : 4'h0) | (tryToRead_3[5] ? input_5_bits_readLane_0 : 4'h0) | (tryToRead_3[6] ? input_6_bits_readLane_0 : 4'h0) | (tryToRead_3[7] ? input_7_bits_readLane_0 : 4'h0)
    | (tryToRead_3[8] ? input_8_bits_readLane_0 : 4'h0) | (tryToRead_3[9] ? input_9_bits_readLane_0 : 4'h0) | (tryToRead_3[10] ? input_10_bits_readLane_0 : 4'h0) | (tryToRead_3[11] ? input_11_bits_readLane_0 : 4'h0)
    | (tryToRead_3[12] ? input_12_bits_readLane_0 : 4'h0) | (tryToRead_3[13] ? input_13_bits_readLane_0 : 4'h0) | (tryToRead_3[14] ? input_14_bits_readLane_0 : 4'h0) | (tryToRead_3[15] ? input_15_bits_readLane_0 : 4'h0);
  assign selectReq_3_bits_offset =
    (tryToRead_3[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead_3[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead_3[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead_3[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead_3[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead_3[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead_3[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead_3[7] ? input_7_bits_offset_0 : 2'h0)
    | (tryToRead_3[8] ? input_8_bits_offset_0 : 2'h0) | (tryToRead_3[9] ? input_9_bits_offset_0 : 2'h0) | (tryToRead_3[10] ? input_10_bits_offset_0 : 2'h0) | (tryToRead_3[11] ? input_11_bits_offset_0 : 2'h0)
    | (tryToRead_3[12] ? input_12_bits_offset_0 : 2'h0) | (tryToRead_3[13] ? input_13_bits_offset_0 : 2'h0) | (tryToRead_3[14] ? input_14_bits_offset_0 : 2'h0) | (tryToRead_3[15] ? input_15_bits_offset_0 : 2'h0);
  assign selectReq_3_bits_vs =
    (tryToRead_3[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_3[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_3[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_3[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_3[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_3[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_3[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_3[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_3[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_3[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_3[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_3[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_3[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_3[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_3[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_3[15] ? input_15_bits_vs_0 : 5'h0);
  wire        selectReq_3_valid =
    tryToRead_3[0] & input_0_valid_0 | tryToRead_3[1] & input_1_valid_0 | tryToRead_3[2] & input_2_valid_0 | tryToRead_3[3] & input_3_valid_0 | tryToRead_3[4] & input_4_valid_0 | tryToRead_3[5] & input_5_valid_0 | tryToRead_3[6]
    & input_6_valid_0 | tryToRead_3[7] & input_7_valid_0 | tryToRead_3[8] & input_8_valid_0 | tryToRead_3[9] & input_9_valid_0 | tryToRead_3[10] & input_10_valid_0 | tryToRead_3[11] & input_11_valid_0 | tryToRead_3[12] & input_12_valid_0
    | tryToRead_3[13] & input_13_valid_0 | tryToRead_3[14] & input_14_valid_0 | tryToRead_3[15] & input_15_valid_0;
  wire        selectReq_3_ready =
    tryToRead_3[0] & input_0_ready_0 | tryToRead_3[1] & input_1_ready_0 | tryToRead_3[2] & input_2_ready_0 | tryToRead_3[3] & input_3_ready_0 | tryToRead_3[4] & input_4_ready_0 | tryToRead_3[5] & input_5_ready_0 | tryToRead_3[6]
    & input_6_ready_0 | tryToRead_3[7] & input_7_ready_0 | tryToRead_3[8] & input_8_ready_0 | tryToRead_3[9] & input_9_ready_0 | tryToRead_3[10] & input_10_ready_0 | tryToRead_3[11] & input_11_ready_0 | tryToRead_3[12] & input_12_ready_0
    | tryToRead_3[13] & input_13_ready_0 | tryToRead_3[14] & input_14_ready_0 | tryToRead_3[15] & input_15_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_4 = {inputSelect1H_1[4], inputSelect1H_0[4]};
  wire [1:0]  tryToRead_lo_lo_hi_4 = {inputSelect1H_3[4], inputSelect1H_2[4]};
  wire [3:0]  tryToRead_lo_lo_4 = {tryToRead_lo_lo_hi_4, tryToRead_lo_lo_lo_4};
  wire [1:0]  tryToRead_lo_hi_lo_4 = {inputSelect1H_5[4], inputSelect1H_4[4]};
  wire [1:0]  tryToRead_lo_hi_hi_4 = {inputSelect1H_7[4], inputSelect1H_6[4]};
  wire [3:0]  tryToRead_lo_hi_4 = {tryToRead_lo_hi_hi_4, tryToRead_lo_hi_lo_4};
  wire [7:0]  tryToRead_lo_4 = {tryToRead_lo_hi_4, tryToRead_lo_lo_4};
  wire [1:0]  tryToRead_hi_lo_lo_4 = {inputSelect1H_9[4], inputSelect1H_8[4]};
  wire [1:0]  tryToRead_hi_lo_hi_4 = {inputSelect1H_11[4], inputSelect1H_10[4]};
  wire [3:0]  tryToRead_hi_lo_4 = {tryToRead_hi_lo_hi_4, tryToRead_hi_lo_lo_4};
  wire [1:0]  tryToRead_hi_hi_lo_4 = {inputSelect1H_13[4], inputSelect1H_12[4]};
  wire [1:0]  tryToRead_hi_hi_hi_4 = {inputSelect1H_15[4], inputSelect1H_14[4]};
  wire [3:0]  tryToRead_hi_hi_4 = {tryToRead_hi_hi_hi_4, tryToRead_hi_hi_lo_4};
  wire [7:0]  tryToRead_hi_4 = {tryToRead_hi_hi_4, tryToRead_hi_lo_4};
  wire [15:0] tryToRead_4 = {tryToRead_hi_4, tryToRead_lo_4};
  wire        output_4_valid_0 = |tryToRead_4;
  wire [4:0]  output_4_bits_vs_0 = selectReq_4_bits_vs;
  wire [1:0]  output_4_bits_offset_0 = selectReq_4_bits_offset;
  wire [3:0]  output_4_bits_writeIndex_0 = selectReq_4_bits_requestIndex;
  wire [1:0]  output_4_bits_dataOffset_0 = selectReq_4_bits_dataOffset;
  assign selectReq_4_bits_dataOffset =
    (tryToRead_4[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_4[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_4[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_4[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_4[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_4[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_4[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_4[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_4[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_4[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_4[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_4[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_4[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_4[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_4[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_4[15] ? input_15_bits_dataOffset_0 : 2'h0);
  assign selectReq_4_bits_requestIndex =
    {3'h0, tryToRead_4[1]} | {2'h0, tryToRead_4[2], 1'h0} | (tryToRead_4[3] ? 4'h3 : 4'h0) | {1'h0, tryToRead_4[4], 2'h0} | (tryToRead_4[5] ? 4'h5 : 4'h0) | (tryToRead_4[6] ? 4'h6 : 4'h0) | (tryToRead_4[7] ? 4'h7 : 4'h0)
    | {tryToRead_4[8], 3'h0} | (tryToRead_4[9] ? 4'h9 : 4'h0) | (tryToRead_4[10] ? 4'hA : 4'h0) | (tryToRead_4[11] ? 4'hB : 4'h0) | (tryToRead_4[12] ? 4'hC : 4'h0) | (tryToRead_4[13] ? 4'hD : 4'h0) | (tryToRead_4[14] ? 4'hE : 4'h0)
    | {4{tryToRead_4[15]}};
  wire [3:0]  selectReq_4_bits_readLane =
    (tryToRead_4[0] ? input_0_bits_readLane_0 : 4'h0) | (tryToRead_4[1] ? input_1_bits_readLane_0 : 4'h0) | (tryToRead_4[2] ? input_2_bits_readLane_0 : 4'h0) | (tryToRead_4[3] ? input_3_bits_readLane_0 : 4'h0)
    | (tryToRead_4[4] ? input_4_bits_readLane_0 : 4'h0) | (tryToRead_4[5] ? input_5_bits_readLane_0 : 4'h0) | (tryToRead_4[6] ? input_6_bits_readLane_0 : 4'h0) | (tryToRead_4[7] ? input_7_bits_readLane_0 : 4'h0)
    | (tryToRead_4[8] ? input_8_bits_readLane_0 : 4'h0) | (tryToRead_4[9] ? input_9_bits_readLane_0 : 4'h0) | (tryToRead_4[10] ? input_10_bits_readLane_0 : 4'h0) | (tryToRead_4[11] ? input_11_bits_readLane_0 : 4'h0)
    | (tryToRead_4[12] ? input_12_bits_readLane_0 : 4'h0) | (tryToRead_4[13] ? input_13_bits_readLane_0 : 4'h0) | (tryToRead_4[14] ? input_14_bits_readLane_0 : 4'h0) | (tryToRead_4[15] ? input_15_bits_readLane_0 : 4'h0);
  assign selectReq_4_bits_offset =
    (tryToRead_4[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead_4[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead_4[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead_4[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead_4[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead_4[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead_4[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead_4[7] ? input_7_bits_offset_0 : 2'h0)
    | (tryToRead_4[8] ? input_8_bits_offset_0 : 2'h0) | (tryToRead_4[9] ? input_9_bits_offset_0 : 2'h0) | (tryToRead_4[10] ? input_10_bits_offset_0 : 2'h0) | (tryToRead_4[11] ? input_11_bits_offset_0 : 2'h0)
    | (tryToRead_4[12] ? input_12_bits_offset_0 : 2'h0) | (tryToRead_4[13] ? input_13_bits_offset_0 : 2'h0) | (tryToRead_4[14] ? input_14_bits_offset_0 : 2'h0) | (tryToRead_4[15] ? input_15_bits_offset_0 : 2'h0);
  assign selectReq_4_bits_vs =
    (tryToRead_4[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_4[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_4[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_4[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_4[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_4[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_4[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_4[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_4[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_4[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_4[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_4[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_4[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_4[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_4[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_4[15] ? input_15_bits_vs_0 : 5'h0);
  wire        selectReq_4_valid =
    tryToRead_4[0] & input_0_valid_0 | tryToRead_4[1] & input_1_valid_0 | tryToRead_4[2] & input_2_valid_0 | tryToRead_4[3] & input_3_valid_0 | tryToRead_4[4] & input_4_valid_0 | tryToRead_4[5] & input_5_valid_0 | tryToRead_4[6]
    & input_6_valid_0 | tryToRead_4[7] & input_7_valid_0 | tryToRead_4[8] & input_8_valid_0 | tryToRead_4[9] & input_9_valid_0 | tryToRead_4[10] & input_10_valid_0 | tryToRead_4[11] & input_11_valid_0 | tryToRead_4[12] & input_12_valid_0
    | tryToRead_4[13] & input_13_valid_0 | tryToRead_4[14] & input_14_valid_0 | tryToRead_4[15] & input_15_valid_0;
  wire        selectReq_4_ready =
    tryToRead_4[0] & input_0_ready_0 | tryToRead_4[1] & input_1_ready_0 | tryToRead_4[2] & input_2_ready_0 | tryToRead_4[3] & input_3_ready_0 | tryToRead_4[4] & input_4_ready_0 | tryToRead_4[5] & input_5_ready_0 | tryToRead_4[6]
    & input_6_ready_0 | tryToRead_4[7] & input_7_ready_0 | tryToRead_4[8] & input_8_ready_0 | tryToRead_4[9] & input_9_ready_0 | tryToRead_4[10] & input_10_ready_0 | tryToRead_4[11] & input_11_ready_0 | tryToRead_4[12] & input_12_ready_0
    | tryToRead_4[13] & input_13_ready_0 | tryToRead_4[14] & input_14_ready_0 | tryToRead_4[15] & input_15_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_5 = {inputSelect1H_1[5], inputSelect1H_0[5]};
  wire [1:0]  tryToRead_lo_lo_hi_5 = {inputSelect1H_3[5], inputSelect1H_2[5]};
  wire [3:0]  tryToRead_lo_lo_5 = {tryToRead_lo_lo_hi_5, tryToRead_lo_lo_lo_5};
  wire [1:0]  tryToRead_lo_hi_lo_5 = {inputSelect1H_5[5], inputSelect1H_4[5]};
  wire [1:0]  tryToRead_lo_hi_hi_5 = {inputSelect1H_7[5], inputSelect1H_6[5]};
  wire [3:0]  tryToRead_lo_hi_5 = {tryToRead_lo_hi_hi_5, tryToRead_lo_hi_lo_5};
  wire [7:0]  tryToRead_lo_5 = {tryToRead_lo_hi_5, tryToRead_lo_lo_5};
  wire [1:0]  tryToRead_hi_lo_lo_5 = {inputSelect1H_9[5], inputSelect1H_8[5]};
  wire [1:0]  tryToRead_hi_lo_hi_5 = {inputSelect1H_11[5], inputSelect1H_10[5]};
  wire [3:0]  tryToRead_hi_lo_5 = {tryToRead_hi_lo_hi_5, tryToRead_hi_lo_lo_5};
  wire [1:0]  tryToRead_hi_hi_lo_5 = {inputSelect1H_13[5], inputSelect1H_12[5]};
  wire [1:0]  tryToRead_hi_hi_hi_5 = {inputSelect1H_15[5], inputSelect1H_14[5]};
  wire [3:0]  tryToRead_hi_hi_5 = {tryToRead_hi_hi_hi_5, tryToRead_hi_hi_lo_5};
  wire [7:0]  tryToRead_hi_5 = {tryToRead_hi_hi_5, tryToRead_hi_lo_5};
  wire [15:0] tryToRead_5 = {tryToRead_hi_5, tryToRead_lo_5};
  wire        output_5_valid_0 = |tryToRead_5;
  wire [4:0]  output_5_bits_vs_0 = selectReq_5_bits_vs;
  wire [1:0]  output_5_bits_offset_0 = selectReq_5_bits_offset;
  wire [3:0]  output_5_bits_writeIndex_0 = selectReq_5_bits_requestIndex;
  wire [1:0]  output_5_bits_dataOffset_0 = selectReq_5_bits_dataOffset;
  assign selectReq_5_bits_dataOffset =
    (tryToRead_5[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_5[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_5[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_5[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_5[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_5[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_5[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_5[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_5[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_5[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_5[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_5[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_5[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_5[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_5[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_5[15] ? input_15_bits_dataOffset_0 : 2'h0);
  assign selectReq_5_bits_requestIndex =
    {3'h0, tryToRead_5[1]} | {2'h0, tryToRead_5[2], 1'h0} | (tryToRead_5[3] ? 4'h3 : 4'h0) | {1'h0, tryToRead_5[4], 2'h0} | (tryToRead_5[5] ? 4'h5 : 4'h0) | (tryToRead_5[6] ? 4'h6 : 4'h0) | (tryToRead_5[7] ? 4'h7 : 4'h0)
    | {tryToRead_5[8], 3'h0} | (tryToRead_5[9] ? 4'h9 : 4'h0) | (tryToRead_5[10] ? 4'hA : 4'h0) | (tryToRead_5[11] ? 4'hB : 4'h0) | (tryToRead_5[12] ? 4'hC : 4'h0) | (tryToRead_5[13] ? 4'hD : 4'h0) | (tryToRead_5[14] ? 4'hE : 4'h0)
    | {4{tryToRead_5[15]}};
  wire [3:0]  selectReq_5_bits_readLane =
    (tryToRead_5[0] ? input_0_bits_readLane_0 : 4'h0) | (tryToRead_5[1] ? input_1_bits_readLane_0 : 4'h0) | (tryToRead_5[2] ? input_2_bits_readLane_0 : 4'h0) | (tryToRead_5[3] ? input_3_bits_readLane_0 : 4'h0)
    | (tryToRead_5[4] ? input_4_bits_readLane_0 : 4'h0) | (tryToRead_5[5] ? input_5_bits_readLane_0 : 4'h0) | (tryToRead_5[6] ? input_6_bits_readLane_0 : 4'h0) | (tryToRead_5[7] ? input_7_bits_readLane_0 : 4'h0)
    | (tryToRead_5[8] ? input_8_bits_readLane_0 : 4'h0) | (tryToRead_5[9] ? input_9_bits_readLane_0 : 4'h0) | (tryToRead_5[10] ? input_10_bits_readLane_0 : 4'h0) | (tryToRead_5[11] ? input_11_bits_readLane_0 : 4'h0)
    | (tryToRead_5[12] ? input_12_bits_readLane_0 : 4'h0) | (tryToRead_5[13] ? input_13_bits_readLane_0 : 4'h0) | (tryToRead_5[14] ? input_14_bits_readLane_0 : 4'h0) | (tryToRead_5[15] ? input_15_bits_readLane_0 : 4'h0);
  assign selectReq_5_bits_offset =
    (tryToRead_5[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead_5[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead_5[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead_5[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead_5[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead_5[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead_5[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead_5[7] ? input_7_bits_offset_0 : 2'h0)
    | (tryToRead_5[8] ? input_8_bits_offset_0 : 2'h0) | (tryToRead_5[9] ? input_9_bits_offset_0 : 2'h0) | (tryToRead_5[10] ? input_10_bits_offset_0 : 2'h0) | (tryToRead_5[11] ? input_11_bits_offset_0 : 2'h0)
    | (tryToRead_5[12] ? input_12_bits_offset_0 : 2'h0) | (tryToRead_5[13] ? input_13_bits_offset_0 : 2'h0) | (tryToRead_5[14] ? input_14_bits_offset_0 : 2'h0) | (tryToRead_5[15] ? input_15_bits_offset_0 : 2'h0);
  assign selectReq_5_bits_vs =
    (tryToRead_5[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_5[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_5[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_5[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_5[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_5[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_5[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_5[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_5[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_5[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_5[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_5[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_5[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_5[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_5[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_5[15] ? input_15_bits_vs_0 : 5'h0);
  wire        selectReq_5_valid =
    tryToRead_5[0] & input_0_valid_0 | tryToRead_5[1] & input_1_valid_0 | tryToRead_5[2] & input_2_valid_0 | tryToRead_5[3] & input_3_valid_0 | tryToRead_5[4] & input_4_valid_0 | tryToRead_5[5] & input_5_valid_0 | tryToRead_5[6]
    & input_6_valid_0 | tryToRead_5[7] & input_7_valid_0 | tryToRead_5[8] & input_8_valid_0 | tryToRead_5[9] & input_9_valid_0 | tryToRead_5[10] & input_10_valid_0 | tryToRead_5[11] & input_11_valid_0 | tryToRead_5[12] & input_12_valid_0
    | tryToRead_5[13] & input_13_valid_0 | tryToRead_5[14] & input_14_valid_0 | tryToRead_5[15] & input_15_valid_0;
  wire        selectReq_5_ready =
    tryToRead_5[0] & input_0_ready_0 | tryToRead_5[1] & input_1_ready_0 | tryToRead_5[2] & input_2_ready_0 | tryToRead_5[3] & input_3_ready_0 | tryToRead_5[4] & input_4_ready_0 | tryToRead_5[5] & input_5_ready_0 | tryToRead_5[6]
    & input_6_ready_0 | tryToRead_5[7] & input_7_ready_0 | tryToRead_5[8] & input_8_ready_0 | tryToRead_5[9] & input_9_ready_0 | tryToRead_5[10] & input_10_ready_0 | tryToRead_5[11] & input_11_ready_0 | tryToRead_5[12] & input_12_ready_0
    | tryToRead_5[13] & input_13_ready_0 | tryToRead_5[14] & input_14_ready_0 | tryToRead_5[15] & input_15_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_6 = {inputSelect1H_1[6], inputSelect1H_0[6]};
  wire [1:0]  tryToRead_lo_lo_hi_6 = {inputSelect1H_3[6], inputSelect1H_2[6]};
  wire [3:0]  tryToRead_lo_lo_6 = {tryToRead_lo_lo_hi_6, tryToRead_lo_lo_lo_6};
  wire [1:0]  tryToRead_lo_hi_lo_6 = {inputSelect1H_5[6], inputSelect1H_4[6]};
  wire [1:0]  tryToRead_lo_hi_hi_6 = {inputSelect1H_7[6], inputSelect1H_6[6]};
  wire [3:0]  tryToRead_lo_hi_6 = {tryToRead_lo_hi_hi_6, tryToRead_lo_hi_lo_6};
  wire [7:0]  tryToRead_lo_6 = {tryToRead_lo_hi_6, tryToRead_lo_lo_6};
  wire [1:0]  tryToRead_hi_lo_lo_6 = {inputSelect1H_9[6], inputSelect1H_8[6]};
  wire [1:0]  tryToRead_hi_lo_hi_6 = {inputSelect1H_11[6], inputSelect1H_10[6]};
  wire [3:0]  tryToRead_hi_lo_6 = {tryToRead_hi_lo_hi_6, tryToRead_hi_lo_lo_6};
  wire [1:0]  tryToRead_hi_hi_lo_6 = {inputSelect1H_13[6], inputSelect1H_12[6]};
  wire [1:0]  tryToRead_hi_hi_hi_6 = {inputSelect1H_15[6], inputSelect1H_14[6]};
  wire [3:0]  tryToRead_hi_hi_6 = {tryToRead_hi_hi_hi_6, tryToRead_hi_hi_lo_6};
  wire [7:0]  tryToRead_hi_6 = {tryToRead_hi_hi_6, tryToRead_hi_lo_6};
  wire [15:0] tryToRead_6 = {tryToRead_hi_6, tryToRead_lo_6};
  wire        output_6_valid_0 = |tryToRead_6;
  wire [4:0]  output_6_bits_vs_0 = selectReq_6_bits_vs;
  wire [1:0]  output_6_bits_offset_0 = selectReq_6_bits_offset;
  wire [3:0]  output_6_bits_writeIndex_0 = selectReq_6_bits_requestIndex;
  wire [1:0]  output_6_bits_dataOffset_0 = selectReq_6_bits_dataOffset;
  assign selectReq_6_bits_dataOffset =
    (tryToRead_6[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_6[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_6[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_6[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_6[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_6[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_6[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_6[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_6[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_6[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_6[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_6[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_6[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_6[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_6[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_6[15] ? input_15_bits_dataOffset_0 : 2'h0);
  assign selectReq_6_bits_requestIndex =
    {3'h0, tryToRead_6[1]} | {2'h0, tryToRead_6[2], 1'h0} | (tryToRead_6[3] ? 4'h3 : 4'h0) | {1'h0, tryToRead_6[4], 2'h0} | (tryToRead_6[5] ? 4'h5 : 4'h0) | (tryToRead_6[6] ? 4'h6 : 4'h0) | (tryToRead_6[7] ? 4'h7 : 4'h0)
    | {tryToRead_6[8], 3'h0} | (tryToRead_6[9] ? 4'h9 : 4'h0) | (tryToRead_6[10] ? 4'hA : 4'h0) | (tryToRead_6[11] ? 4'hB : 4'h0) | (tryToRead_6[12] ? 4'hC : 4'h0) | (tryToRead_6[13] ? 4'hD : 4'h0) | (tryToRead_6[14] ? 4'hE : 4'h0)
    | {4{tryToRead_6[15]}};
  wire [3:0]  selectReq_6_bits_readLane =
    (tryToRead_6[0] ? input_0_bits_readLane_0 : 4'h0) | (tryToRead_6[1] ? input_1_bits_readLane_0 : 4'h0) | (tryToRead_6[2] ? input_2_bits_readLane_0 : 4'h0) | (tryToRead_6[3] ? input_3_bits_readLane_0 : 4'h0)
    | (tryToRead_6[4] ? input_4_bits_readLane_0 : 4'h0) | (tryToRead_6[5] ? input_5_bits_readLane_0 : 4'h0) | (tryToRead_6[6] ? input_6_bits_readLane_0 : 4'h0) | (tryToRead_6[7] ? input_7_bits_readLane_0 : 4'h0)
    | (tryToRead_6[8] ? input_8_bits_readLane_0 : 4'h0) | (tryToRead_6[9] ? input_9_bits_readLane_0 : 4'h0) | (tryToRead_6[10] ? input_10_bits_readLane_0 : 4'h0) | (tryToRead_6[11] ? input_11_bits_readLane_0 : 4'h0)
    | (tryToRead_6[12] ? input_12_bits_readLane_0 : 4'h0) | (tryToRead_6[13] ? input_13_bits_readLane_0 : 4'h0) | (tryToRead_6[14] ? input_14_bits_readLane_0 : 4'h0) | (tryToRead_6[15] ? input_15_bits_readLane_0 : 4'h0);
  assign selectReq_6_bits_offset =
    (tryToRead_6[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead_6[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead_6[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead_6[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead_6[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead_6[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead_6[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead_6[7] ? input_7_bits_offset_0 : 2'h0)
    | (tryToRead_6[8] ? input_8_bits_offset_0 : 2'h0) | (tryToRead_6[9] ? input_9_bits_offset_0 : 2'h0) | (tryToRead_6[10] ? input_10_bits_offset_0 : 2'h0) | (tryToRead_6[11] ? input_11_bits_offset_0 : 2'h0)
    | (tryToRead_6[12] ? input_12_bits_offset_0 : 2'h0) | (tryToRead_6[13] ? input_13_bits_offset_0 : 2'h0) | (tryToRead_6[14] ? input_14_bits_offset_0 : 2'h0) | (tryToRead_6[15] ? input_15_bits_offset_0 : 2'h0);
  assign selectReq_6_bits_vs =
    (tryToRead_6[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_6[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_6[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_6[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_6[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_6[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_6[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_6[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_6[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_6[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_6[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_6[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_6[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_6[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_6[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_6[15] ? input_15_bits_vs_0 : 5'h0);
  wire        selectReq_6_valid =
    tryToRead_6[0] & input_0_valid_0 | tryToRead_6[1] & input_1_valid_0 | tryToRead_6[2] & input_2_valid_0 | tryToRead_6[3] & input_3_valid_0 | tryToRead_6[4] & input_4_valid_0 | tryToRead_6[5] & input_5_valid_0 | tryToRead_6[6]
    & input_6_valid_0 | tryToRead_6[7] & input_7_valid_0 | tryToRead_6[8] & input_8_valid_0 | tryToRead_6[9] & input_9_valid_0 | tryToRead_6[10] & input_10_valid_0 | tryToRead_6[11] & input_11_valid_0 | tryToRead_6[12] & input_12_valid_0
    | tryToRead_6[13] & input_13_valid_0 | tryToRead_6[14] & input_14_valid_0 | tryToRead_6[15] & input_15_valid_0;
  wire        selectReq_6_ready =
    tryToRead_6[0] & input_0_ready_0 | tryToRead_6[1] & input_1_ready_0 | tryToRead_6[2] & input_2_ready_0 | tryToRead_6[3] & input_3_ready_0 | tryToRead_6[4] & input_4_ready_0 | tryToRead_6[5] & input_5_ready_0 | tryToRead_6[6]
    & input_6_ready_0 | tryToRead_6[7] & input_7_ready_0 | tryToRead_6[8] & input_8_ready_0 | tryToRead_6[9] & input_9_ready_0 | tryToRead_6[10] & input_10_ready_0 | tryToRead_6[11] & input_11_ready_0 | tryToRead_6[12] & input_12_ready_0
    | tryToRead_6[13] & input_13_ready_0 | tryToRead_6[14] & input_14_ready_0 | tryToRead_6[15] & input_15_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_7 = {inputSelect1H_1[7], inputSelect1H_0[7]};
  wire [1:0]  tryToRead_lo_lo_hi_7 = {inputSelect1H_3[7], inputSelect1H_2[7]};
  wire [3:0]  tryToRead_lo_lo_7 = {tryToRead_lo_lo_hi_7, tryToRead_lo_lo_lo_7};
  wire [1:0]  tryToRead_lo_hi_lo_7 = {inputSelect1H_5[7], inputSelect1H_4[7]};
  wire [1:0]  tryToRead_lo_hi_hi_7 = {inputSelect1H_7[7], inputSelect1H_6[7]};
  wire [3:0]  tryToRead_lo_hi_7 = {tryToRead_lo_hi_hi_7, tryToRead_lo_hi_lo_7};
  wire [7:0]  tryToRead_lo_7 = {tryToRead_lo_hi_7, tryToRead_lo_lo_7};
  wire [1:0]  tryToRead_hi_lo_lo_7 = {inputSelect1H_9[7], inputSelect1H_8[7]};
  wire [1:0]  tryToRead_hi_lo_hi_7 = {inputSelect1H_11[7], inputSelect1H_10[7]};
  wire [3:0]  tryToRead_hi_lo_7 = {tryToRead_hi_lo_hi_7, tryToRead_hi_lo_lo_7};
  wire [1:0]  tryToRead_hi_hi_lo_7 = {inputSelect1H_13[7], inputSelect1H_12[7]};
  wire [1:0]  tryToRead_hi_hi_hi_7 = {inputSelect1H_15[7], inputSelect1H_14[7]};
  wire [3:0]  tryToRead_hi_hi_7 = {tryToRead_hi_hi_hi_7, tryToRead_hi_hi_lo_7};
  wire [7:0]  tryToRead_hi_7 = {tryToRead_hi_hi_7, tryToRead_hi_lo_7};
  wire [15:0] tryToRead_7 = {tryToRead_hi_7, tryToRead_lo_7};
  wire        output_7_valid_0 = |tryToRead_7;
  wire [4:0]  output_7_bits_vs_0 = selectReq_7_bits_vs;
  wire [1:0]  output_7_bits_offset_0 = selectReq_7_bits_offset;
  wire [3:0]  output_7_bits_writeIndex_0 = selectReq_7_bits_requestIndex;
  wire [1:0]  output_7_bits_dataOffset_0 = selectReq_7_bits_dataOffset;
  assign selectReq_7_bits_dataOffset =
    (tryToRead_7[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_7[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_7[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_7[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_7[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_7[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_7[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_7[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_7[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_7[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_7[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_7[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_7[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_7[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_7[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_7[15] ? input_15_bits_dataOffset_0 : 2'h0);
  assign selectReq_7_bits_requestIndex =
    {3'h0, tryToRead_7[1]} | {2'h0, tryToRead_7[2], 1'h0} | (tryToRead_7[3] ? 4'h3 : 4'h0) | {1'h0, tryToRead_7[4], 2'h0} | (tryToRead_7[5] ? 4'h5 : 4'h0) | (tryToRead_7[6] ? 4'h6 : 4'h0) | (tryToRead_7[7] ? 4'h7 : 4'h0)
    | {tryToRead_7[8], 3'h0} | (tryToRead_7[9] ? 4'h9 : 4'h0) | (tryToRead_7[10] ? 4'hA : 4'h0) | (tryToRead_7[11] ? 4'hB : 4'h0) | (tryToRead_7[12] ? 4'hC : 4'h0) | (tryToRead_7[13] ? 4'hD : 4'h0) | (tryToRead_7[14] ? 4'hE : 4'h0)
    | {4{tryToRead_7[15]}};
  wire [3:0]  selectReq_7_bits_readLane =
    (tryToRead_7[0] ? input_0_bits_readLane_0 : 4'h0) | (tryToRead_7[1] ? input_1_bits_readLane_0 : 4'h0) | (tryToRead_7[2] ? input_2_bits_readLane_0 : 4'h0) | (tryToRead_7[3] ? input_3_bits_readLane_0 : 4'h0)
    | (tryToRead_7[4] ? input_4_bits_readLane_0 : 4'h0) | (tryToRead_7[5] ? input_5_bits_readLane_0 : 4'h0) | (tryToRead_7[6] ? input_6_bits_readLane_0 : 4'h0) | (tryToRead_7[7] ? input_7_bits_readLane_0 : 4'h0)
    | (tryToRead_7[8] ? input_8_bits_readLane_0 : 4'h0) | (tryToRead_7[9] ? input_9_bits_readLane_0 : 4'h0) | (tryToRead_7[10] ? input_10_bits_readLane_0 : 4'h0) | (tryToRead_7[11] ? input_11_bits_readLane_0 : 4'h0)
    | (tryToRead_7[12] ? input_12_bits_readLane_0 : 4'h0) | (tryToRead_7[13] ? input_13_bits_readLane_0 : 4'h0) | (tryToRead_7[14] ? input_14_bits_readLane_0 : 4'h0) | (tryToRead_7[15] ? input_15_bits_readLane_0 : 4'h0);
  assign selectReq_7_bits_offset =
    (tryToRead_7[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead_7[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead_7[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead_7[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead_7[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead_7[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead_7[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead_7[7] ? input_7_bits_offset_0 : 2'h0)
    | (tryToRead_7[8] ? input_8_bits_offset_0 : 2'h0) | (tryToRead_7[9] ? input_9_bits_offset_0 : 2'h0) | (tryToRead_7[10] ? input_10_bits_offset_0 : 2'h0) | (tryToRead_7[11] ? input_11_bits_offset_0 : 2'h0)
    | (tryToRead_7[12] ? input_12_bits_offset_0 : 2'h0) | (tryToRead_7[13] ? input_13_bits_offset_0 : 2'h0) | (tryToRead_7[14] ? input_14_bits_offset_0 : 2'h0) | (tryToRead_7[15] ? input_15_bits_offset_0 : 2'h0);
  assign selectReq_7_bits_vs =
    (tryToRead_7[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_7[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_7[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_7[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_7[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_7[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_7[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_7[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_7[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_7[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_7[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_7[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_7[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_7[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_7[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_7[15] ? input_15_bits_vs_0 : 5'h0);
  wire        selectReq_7_valid =
    tryToRead_7[0] & input_0_valid_0 | tryToRead_7[1] & input_1_valid_0 | tryToRead_7[2] & input_2_valid_0 | tryToRead_7[3] & input_3_valid_0 | tryToRead_7[4] & input_4_valid_0 | tryToRead_7[5] & input_5_valid_0 | tryToRead_7[6]
    & input_6_valid_0 | tryToRead_7[7] & input_7_valid_0 | tryToRead_7[8] & input_8_valid_0 | tryToRead_7[9] & input_9_valid_0 | tryToRead_7[10] & input_10_valid_0 | tryToRead_7[11] & input_11_valid_0 | tryToRead_7[12] & input_12_valid_0
    | tryToRead_7[13] & input_13_valid_0 | tryToRead_7[14] & input_14_valid_0 | tryToRead_7[15] & input_15_valid_0;
  wire        selectReq_7_ready =
    tryToRead_7[0] & input_0_ready_0 | tryToRead_7[1] & input_1_ready_0 | tryToRead_7[2] & input_2_ready_0 | tryToRead_7[3] & input_3_ready_0 | tryToRead_7[4] & input_4_ready_0 | tryToRead_7[5] & input_5_ready_0 | tryToRead_7[6]
    & input_6_ready_0 | tryToRead_7[7] & input_7_ready_0 | tryToRead_7[8] & input_8_ready_0 | tryToRead_7[9] & input_9_ready_0 | tryToRead_7[10] & input_10_ready_0 | tryToRead_7[11] & input_11_ready_0 | tryToRead_7[12] & input_12_ready_0
    | tryToRead_7[13] & input_13_ready_0 | tryToRead_7[14] & input_14_ready_0 | tryToRead_7[15] & input_15_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_8 = {inputSelect1H_1[8], inputSelect1H_0[8]};
  wire [1:0]  tryToRead_lo_lo_hi_8 = {inputSelect1H_3[8], inputSelect1H_2[8]};
  wire [3:0]  tryToRead_lo_lo_8 = {tryToRead_lo_lo_hi_8, tryToRead_lo_lo_lo_8};
  wire [1:0]  tryToRead_lo_hi_lo_8 = {inputSelect1H_5[8], inputSelect1H_4[8]};
  wire [1:0]  tryToRead_lo_hi_hi_8 = {inputSelect1H_7[8], inputSelect1H_6[8]};
  wire [3:0]  tryToRead_lo_hi_8 = {tryToRead_lo_hi_hi_8, tryToRead_lo_hi_lo_8};
  wire [7:0]  tryToRead_lo_8 = {tryToRead_lo_hi_8, tryToRead_lo_lo_8};
  wire [1:0]  tryToRead_hi_lo_lo_8 = {inputSelect1H_9[8], inputSelect1H_8[8]};
  wire [1:0]  tryToRead_hi_lo_hi_8 = {inputSelect1H_11[8], inputSelect1H_10[8]};
  wire [3:0]  tryToRead_hi_lo_8 = {tryToRead_hi_lo_hi_8, tryToRead_hi_lo_lo_8};
  wire [1:0]  tryToRead_hi_hi_lo_8 = {inputSelect1H_13[8], inputSelect1H_12[8]};
  wire [1:0]  tryToRead_hi_hi_hi_8 = {inputSelect1H_15[8], inputSelect1H_14[8]};
  wire [3:0]  tryToRead_hi_hi_8 = {tryToRead_hi_hi_hi_8, tryToRead_hi_hi_lo_8};
  wire [7:0]  tryToRead_hi_8 = {tryToRead_hi_hi_8, tryToRead_hi_lo_8};
  wire [15:0] tryToRead_8 = {tryToRead_hi_8, tryToRead_lo_8};
  wire        output_8_valid_0 = |tryToRead_8;
  wire [4:0]  output_8_bits_vs_0 = selectReq_8_bits_vs;
  wire [1:0]  output_8_bits_offset_0 = selectReq_8_bits_offset;
  wire [3:0]  output_8_bits_writeIndex_0 = selectReq_8_bits_requestIndex;
  wire [1:0]  output_8_bits_dataOffset_0 = selectReq_8_bits_dataOffset;
  assign selectReq_8_bits_dataOffset =
    (tryToRead_8[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_8[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_8[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_8[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_8[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_8[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_8[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_8[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_8[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_8[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_8[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_8[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_8[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_8[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_8[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_8[15] ? input_15_bits_dataOffset_0 : 2'h0);
  assign selectReq_8_bits_requestIndex =
    {3'h0, tryToRead_8[1]} | {2'h0, tryToRead_8[2], 1'h0} | (tryToRead_8[3] ? 4'h3 : 4'h0) | {1'h0, tryToRead_8[4], 2'h0} | (tryToRead_8[5] ? 4'h5 : 4'h0) | (tryToRead_8[6] ? 4'h6 : 4'h0) | (tryToRead_8[7] ? 4'h7 : 4'h0)
    | {tryToRead_8[8], 3'h0} | (tryToRead_8[9] ? 4'h9 : 4'h0) | (tryToRead_8[10] ? 4'hA : 4'h0) | (tryToRead_8[11] ? 4'hB : 4'h0) | (tryToRead_8[12] ? 4'hC : 4'h0) | (tryToRead_8[13] ? 4'hD : 4'h0) | (tryToRead_8[14] ? 4'hE : 4'h0)
    | {4{tryToRead_8[15]}};
  wire [3:0]  selectReq_8_bits_readLane =
    (tryToRead_8[0] ? input_0_bits_readLane_0 : 4'h0) | (tryToRead_8[1] ? input_1_bits_readLane_0 : 4'h0) | (tryToRead_8[2] ? input_2_bits_readLane_0 : 4'h0) | (tryToRead_8[3] ? input_3_bits_readLane_0 : 4'h0)
    | (tryToRead_8[4] ? input_4_bits_readLane_0 : 4'h0) | (tryToRead_8[5] ? input_5_bits_readLane_0 : 4'h0) | (tryToRead_8[6] ? input_6_bits_readLane_0 : 4'h0) | (tryToRead_8[7] ? input_7_bits_readLane_0 : 4'h0)
    | (tryToRead_8[8] ? input_8_bits_readLane_0 : 4'h0) | (tryToRead_8[9] ? input_9_bits_readLane_0 : 4'h0) | (tryToRead_8[10] ? input_10_bits_readLane_0 : 4'h0) | (tryToRead_8[11] ? input_11_bits_readLane_0 : 4'h0)
    | (tryToRead_8[12] ? input_12_bits_readLane_0 : 4'h0) | (tryToRead_8[13] ? input_13_bits_readLane_0 : 4'h0) | (tryToRead_8[14] ? input_14_bits_readLane_0 : 4'h0) | (tryToRead_8[15] ? input_15_bits_readLane_0 : 4'h0);
  assign selectReq_8_bits_offset =
    (tryToRead_8[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead_8[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead_8[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead_8[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead_8[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead_8[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead_8[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead_8[7] ? input_7_bits_offset_0 : 2'h0)
    | (tryToRead_8[8] ? input_8_bits_offset_0 : 2'h0) | (tryToRead_8[9] ? input_9_bits_offset_0 : 2'h0) | (tryToRead_8[10] ? input_10_bits_offset_0 : 2'h0) | (tryToRead_8[11] ? input_11_bits_offset_0 : 2'h0)
    | (tryToRead_8[12] ? input_12_bits_offset_0 : 2'h0) | (tryToRead_8[13] ? input_13_bits_offset_0 : 2'h0) | (tryToRead_8[14] ? input_14_bits_offset_0 : 2'h0) | (tryToRead_8[15] ? input_15_bits_offset_0 : 2'h0);
  assign selectReq_8_bits_vs =
    (tryToRead_8[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_8[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_8[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_8[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_8[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_8[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_8[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_8[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_8[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_8[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_8[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_8[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_8[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_8[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_8[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_8[15] ? input_15_bits_vs_0 : 5'h0);
  wire        selectReq_8_valid =
    tryToRead_8[0] & input_0_valid_0 | tryToRead_8[1] & input_1_valid_0 | tryToRead_8[2] & input_2_valid_0 | tryToRead_8[3] & input_3_valid_0 | tryToRead_8[4] & input_4_valid_0 | tryToRead_8[5] & input_5_valid_0 | tryToRead_8[6]
    & input_6_valid_0 | tryToRead_8[7] & input_7_valid_0 | tryToRead_8[8] & input_8_valid_0 | tryToRead_8[9] & input_9_valid_0 | tryToRead_8[10] & input_10_valid_0 | tryToRead_8[11] & input_11_valid_0 | tryToRead_8[12] & input_12_valid_0
    | tryToRead_8[13] & input_13_valid_0 | tryToRead_8[14] & input_14_valid_0 | tryToRead_8[15] & input_15_valid_0;
  wire        selectReq_8_ready =
    tryToRead_8[0] & input_0_ready_0 | tryToRead_8[1] & input_1_ready_0 | tryToRead_8[2] & input_2_ready_0 | tryToRead_8[3] & input_3_ready_0 | tryToRead_8[4] & input_4_ready_0 | tryToRead_8[5] & input_5_ready_0 | tryToRead_8[6]
    & input_6_ready_0 | tryToRead_8[7] & input_7_ready_0 | tryToRead_8[8] & input_8_ready_0 | tryToRead_8[9] & input_9_ready_0 | tryToRead_8[10] & input_10_ready_0 | tryToRead_8[11] & input_11_ready_0 | tryToRead_8[12] & input_12_ready_0
    | tryToRead_8[13] & input_13_ready_0 | tryToRead_8[14] & input_14_ready_0 | tryToRead_8[15] & input_15_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_9 = {inputSelect1H_1[9], inputSelect1H_0[9]};
  wire [1:0]  tryToRead_lo_lo_hi_9 = {inputSelect1H_3[9], inputSelect1H_2[9]};
  wire [3:0]  tryToRead_lo_lo_9 = {tryToRead_lo_lo_hi_9, tryToRead_lo_lo_lo_9};
  wire [1:0]  tryToRead_lo_hi_lo_9 = {inputSelect1H_5[9], inputSelect1H_4[9]};
  wire [1:0]  tryToRead_lo_hi_hi_9 = {inputSelect1H_7[9], inputSelect1H_6[9]};
  wire [3:0]  tryToRead_lo_hi_9 = {tryToRead_lo_hi_hi_9, tryToRead_lo_hi_lo_9};
  wire [7:0]  tryToRead_lo_9 = {tryToRead_lo_hi_9, tryToRead_lo_lo_9};
  wire [1:0]  tryToRead_hi_lo_lo_9 = {inputSelect1H_9[9], inputSelect1H_8[9]};
  wire [1:0]  tryToRead_hi_lo_hi_9 = {inputSelect1H_11[9], inputSelect1H_10[9]};
  wire [3:0]  tryToRead_hi_lo_9 = {tryToRead_hi_lo_hi_9, tryToRead_hi_lo_lo_9};
  wire [1:0]  tryToRead_hi_hi_lo_9 = {inputSelect1H_13[9], inputSelect1H_12[9]};
  wire [1:0]  tryToRead_hi_hi_hi_9 = {inputSelect1H_15[9], inputSelect1H_14[9]};
  wire [3:0]  tryToRead_hi_hi_9 = {tryToRead_hi_hi_hi_9, tryToRead_hi_hi_lo_9};
  wire [7:0]  tryToRead_hi_9 = {tryToRead_hi_hi_9, tryToRead_hi_lo_9};
  wire [15:0] tryToRead_9 = {tryToRead_hi_9, tryToRead_lo_9};
  wire        output_9_valid_0 = |tryToRead_9;
  wire [4:0]  output_9_bits_vs_0 = selectReq_9_bits_vs;
  wire [1:0]  output_9_bits_offset_0 = selectReq_9_bits_offset;
  wire [3:0]  output_9_bits_writeIndex_0 = selectReq_9_bits_requestIndex;
  wire [1:0]  output_9_bits_dataOffset_0 = selectReq_9_bits_dataOffset;
  assign selectReq_9_bits_dataOffset =
    (tryToRead_9[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_9[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_9[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_9[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_9[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_9[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_9[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_9[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_9[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_9[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_9[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_9[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_9[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_9[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_9[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_9[15] ? input_15_bits_dataOffset_0 : 2'h0);
  assign selectReq_9_bits_requestIndex =
    {3'h0, tryToRead_9[1]} | {2'h0, tryToRead_9[2], 1'h0} | (tryToRead_9[3] ? 4'h3 : 4'h0) | {1'h0, tryToRead_9[4], 2'h0} | (tryToRead_9[5] ? 4'h5 : 4'h0) | (tryToRead_9[6] ? 4'h6 : 4'h0) | (tryToRead_9[7] ? 4'h7 : 4'h0)
    | {tryToRead_9[8], 3'h0} | (tryToRead_9[9] ? 4'h9 : 4'h0) | (tryToRead_9[10] ? 4'hA : 4'h0) | (tryToRead_9[11] ? 4'hB : 4'h0) | (tryToRead_9[12] ? 4'hC : 4'h0) | (tryToRead_9[13] ? 4'hD : 4'h0) | (tryToRead_9[14] ? 4'hE : 4'h0)
    | {4{tryToRead_9[15]}};
  wire [3:0]  selectReq_9_bits_readLane =
    (tryToRead_9[0] ? input_0_bits_readLane_0 : 4'h0) | (tryToRead_9[1] ? input_1_bits_readLane_0 : 4'h0) | (tryToRead_9[2] ? input_2_bits_readLane_0 : 4'h0) | (tryToRead_9[3] ? input_3_bits_readLane_0 : 4'h0)
    | (tryToRead_9[4] ? input_4_bits_readLane_0 : 4'h0) | (tryToRead_9[5] ? input_5_bits_readLane_0 : 4'h0) | (tryToRead_9[6] ? input_6_bits_readLane_0 : 4'h0) | (tryToRead_9[7] ? input_7_bits_readLane_0 : 4'h0)
    | (tryToRead_9[8] ? input_8_bits_readLane_0 : 4'h0) | (tryToRead_9[9] ? input_9_bits_readLane_0 : 4'h0) | (tryToRead_9[10] ? input_10_bits_readLane_0 : 4'h0) | (tryToRead_9[11] ? input_11_bits_readLane_0 : 4'h0)
    | (tryToRead_9[12] ? input_12_bits_readLane_0 : 4'h0) | (tryToRead_9[13] ? input_13_bits_readLane_0 : 4'h0) | (tryToRead_9[14] ? input_14_bits_readLane_0 : 4'h0) | (tryToRead_9[15] ? input_15_bits_readLane_0 : 4'h0);
  assign selectReq_9_bits_offset =
    (tryToRead_9[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead_9[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead_9[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead_9[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead_9[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead_9[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead_9[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead_9[7] ? input_7_bits_offset_0 : 2'h0)
    | (tryToRead_9[8] ? input_8_bits_offset_0 : 2'h0) | (tryToRead_9[9] ? input_9_bits_offset_0 : 2'h0) | (tryToRead_9[10] ? input_10_bits_offset_0 : 2'h0) | (tryToRead_9[11] ? input_11_bits_offset_0 : 2'h0)
    | (tryToRead_9[12] ? input_12_bits_offset_0 : 2'h0) | (tryToRead_9[13] ? input_13_bits_offset_0 : 2'h0) | (tryToRead_9[14] ? input_14_bits_offset_0 : 2'h0) | (tryToRead_9[15] ? input_15_bits_offset_0 : 2'h0);
  assign selectReq_9_bits_vs =
    (tryToRead_9[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_9[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_9[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_9[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_9[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_9[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_9[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_9[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_9[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_9[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_9[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_9[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_9[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_9[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_9[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_9[15] ? input_15_bits_vs_0 : 5'h0);
  wire        selectReq_9_valid =
    tryToRead_9[0] & input_0_valid_0 | tryToRead_9[1] & input_1_valid_0 | tryToRead_9[2] & input_2_valid_0 | tryToRead_9[3] & input_3_valid_0 | tryToRead_9[4] & input_4_valid_0 | tryToRead_9[5] & input_5_valid_0 | tryToRead_9[6]
    & input_6_valid_0 | tryToRead_9[7] & input_7_valid_0 | tryToRead_9[8] & input_8_valid_0 | tryToRead_9[9] & input_9_valid_0 | tryToRead_9[10] & input_10_valid_0 | tryToRead_9[11] & input_11_valid_0 | tryToRead_9[12] & input_12_valid_0
    | tryToRead_9[13] & input_13_valid_0 | tryToRead_9[14] & input_14_valid_0 | tryToRead_9[15] & input_15_valid_0;
  wire        selectReq_9_ready =
    tryToRead_9[0] & input_0_ready_0 | tryToRead_9[1] & input_1_ready_0 | tryToRead_9[2] & input_2_ready_0 | tryToRead_9[3] & input_3_ready_0 | tryToRead_9[4] & input_4_ready_0 | tryToRead_9[5] & input_5_ready_0 | tryToRead_9[6]
    & input_6_ready_0 | tryToRead_9[7] & input_7_ready_0 | tryToRead_9[8] & input_8_ready_0 | tryToRead_9[9] & input_9_ready_0 | tryToRead_9[10] & input_10_ready_0 | tryToRead_9[11] & input_11_ready_0 | tryToRead_9[12] & input_12_ready_0
    | tryToRead_9[13] & input_13_ready_0 | tryToRead_9[14] & input_14_ready_0 | tryToRead_9[15] & input_15_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_10 = {inputSelect1H_1[10], inputSelect1H_0[10]};
  wire [1:0]  tryToRead_lo_lo_hi_10 = {inputSelect1H_3[10], inputSelect1H_2[10]};
  wire [3:0]  tryToRead_lo_lo_10 = {tryToRead_lo_lo_hi_10, tryToRead_lo_lo_lo_10};
  wire [1:0]  tryToRead_lo_hi_lo_10 = {inputSelect1H_5[10], inputSelect1H_4[10]};
  wire [1:0]  tryToRead_lo_hi_hi_10 = {inputSelect1H_7[10], inputSelect1H_6[10]};
  wire [3:0]  tryToRead_lo_hi_10 = {tryToRead_lo_hi_hi_10, tryToRead_lo_hi_lo_10};
  wire [7:0]  tryToRead_lo_10 = {tryToRead_lo_hi_10, tryToRead_lo_lo_10};
  wire [1:0]  tryToRead_hi_lo_lo_10 = {inputSelect1H_9[10], inputSelect1H_8[10]};
  wire [1:0]  tryToRead_hi_lo_hi_10 = {inputSelect1H_11[10], inputSelect1H_10[10]};
  wire [3:0]  tryToRead_hi_lo_10 = {tryToRead_hi_lo_hi_10, tryToRead_hi_lo_lo_10};
  wire [1:0]  tryToRead_hi_hi_lo_10 = {inputSelect1H_13[10], inputSelect1H_12[10]};
  wire [1:0]  tryToRead_hi_hi_hi_10 = {inputSelect1H_15[10], inputSelect1H_14[10]};
  wire [3:0]  tryToRead_hi_hi_10 = {tryToRead_hi_hi_hi_10, tryToRead_hi_hi_lo_10};
  wire [7:0]  tryToRead_hi_10 = {tryToRead_hi_hi_10, tryToRead_hi_lo_10};
  wire [15:0] tryToRead_10 = {tryToRead_hi_10, tryToRead_lo_10};
  wire        output_10_valid_0 = |tryToRead_10;
  wire [4:0]  output_10_bits_vs_0 = selectReq_10_bits_vs;
  wire [1:0]  output_10_bits_offset_0 = selectReq_10_bits_offset;
  wire [3:0]  output_10_bits_writeIndex_0 = selectReq_10_bits_requestIndex;
  wire [1:0]  output_10_bits_dataOffset_0 = selectReq_10_bits_dataOffset;
  assign selectReq_10_bits_dataOffset =
    (tryToRead_10[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_10[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_10[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_10[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_10[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_10[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_10[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_10[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_10[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_10[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_10[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_10[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_10[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_10[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_10[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_10[15] ? input_15_bits_dataOffset_0 : 2'h0);
  assign selectReq_10_bits_requestIndex =
    {3'h0, tryToRead_10[1]} | {2'h0, tryToRead_10[2], 1'h0} | (tryToRead_10[3] ? 4'h3 : 4'h0) | {1'h0, tryToRead_10[4], 2'h0} | (tryToRead_10[5] ? 4'h5 : 4'h0) | (tryToRead_10[6] ? 4'h6 : 4'h0) | (tryToRead_10[7] ? 4'h7 : 4'h0)
    | {tryToRead_10[8], 3'h0} | (tryToRead_10[9] ? 4'h9 : 4'h0) | (tryToRead_10[10] ? 4'hA : 4'h0) | (tryToRead_10[11] ? 4'hB : 4'h0) | (tryToRead_10[12] ? 4'hC : 4'h0) | (tryToRead_10[13] ? 4'hD : 4'h0) | (tryToRead_10[14] ? 4'hE : 4'h0)
    | {4{tryToRead_10[15]}};
  wire [3:0]  selectReq_10_bits_readLane =
    (tryToRead_10[0] ? input_0_bits_readLane_0 : 4'h0) | (tryToRead_10[1] ? input_1_bits_readLane_0 : 4'h0) | (tryToRead_10[2] ? input_2_bits_readLane_0 : 4'h0) | (tryToRead_10[3] ? input_3_bits_readLane_0 : 4'h0)
    | (tryToRead_10[4] ? input_4_bits_readLane_0 : 4'h0) | (tryToRead_10[5] ? input_5_bits_readLane_0 : 4'h0) | (tryToRead_10[6] ? input_6_bits_readLane_0 : 4'h0) | (tryToRead_10[7] ? input_7_bits_readLane_0 : 4'h0)
    | (tryToRead_10[8] ? input_8_bits_readLane_0 : 4'h0) | (tryToRead_10[9] ? input_9_bits_readLane_0 : 4'h0) | (tryToRead_10[10] ? input_10_bits_readLane_0 : 4'h0) | (tryToRead_10[11] ? input_11_bits_readLane_0 : 4'h0)
    | (tryToRead_10[12] ? input_12_bits_readLane_0 : 4'h0) | (tryToRead_10[13] ? input_13_bits_readLane_0 : 4'h0) | (tryToRead_10[14] ? input_14_bits_readLane_0 : 4'h0) | (tryToRead_10[15] ? input_15_bits_readLane_0 : 4'h0);
  assign selectReq_10_bits_offset =
    (tryToRead_10[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead_10[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead_10[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead_10[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead_10[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead_10[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead_10[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead_10[7] ? input_7_bits_offset_0 : 2'h0)
    | (tryToRead_10[8] ? input_8_bits_offset_0 : 2'h0) | (tryToRead_10[9] ? input_9_bits_offset_0 : 2'h0) | (tryToRead_10[10] ? input_10_bits_offset_0 : 2'h0) | (tryToRead_10[11] ? input_11_bits_offset_0 : 2'h0)
    | (tryToRead_10[12] ? input_12_bits_offset_0 : 2'h0) | (tryToRead_10[13] ? input_13_bits_offset_0 : 2'h0) | (tryToRead_10[14] ? input_14_bits_offset_0 : 2'h0) | (tryToRead_10[15] ? input_15_bits_offset_0 : 2'h0);
  assign selectReq_10_bits_vs =
    (tryToRead_10[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_10[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_10[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_10[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_10[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_10[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_10[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_10[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_10[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_10[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_10[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_10[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_10[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_10[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_10[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_10[15] ? input_15_bits_vs_0 : 5'h0);
  wire        selectReq_10_valid =
    tryToRead_10[0] & input_0_valid_0 | tryToRead_10[1] & input_1_valid_0 | tryToRead_10[2] & input_2_valid_0 | tryToRead_10[3] & input_3_valid_0 | tryToRead_10[4] & input_4_valid_0 | tryToRead_10[5] & input_5_valid_0 | tryToRead_10[6]
    & input_6_valid_0 | tryToRead_10[7] & input_7_valid_0 | tryToRead_10[8] & input_8_valid_0 | tryToRead_10[9] & input_9_valid_0 | tryToRead_10[10] & input_10_valid_0 | tryToRead_10[11] & input_11_valid_0 | tryToRead_10[12]
    & input_12_valid_0 | tryToRead_10[13] & input_13_valid_0 | tryToRead_10[14] & input_14_valid_0 | tryToRead_10[15] & input_15_valid_0;
  wire        selectReq_10_ready =
    tryToRead_10[0] & input_0_ready_0 | tryToRead_10[1] & input_1_ready_0 | tryToRead_10[2] & input_2_ready_0 | tryToRead_10[3] & input_3_ready_0 | tryToRead_10[4] & input_4_ready_0 | tryToRead_10[5] & input_5_ready_0 | tryToRead_10[6]
    & input_6_ready_0 | tryToRead_10[7] & input_7_ready_0 | tryToRead_10[8] & input_8_ready_0 | tryToRead_10[9] & input_9_ready_0 | tryToRead_10[10] & input_10_ready_0 | tryToRead_10[11] & input_11_ready_0 | tryToRead_10[12]
    & input_12_ready_0 | tryToRead_10[13] & input_13_ready_0 | tryToRead_10[14] & input_14_ready_0 | tryToRead_10[15] & input_15_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_11 = {inputSelect1H_1[11], inputSelect1H_0[11]};
  wire [1:0]  tryToRead_lo_lo_hi_11 = {inputSelect1H_3[11], inputSelect1H_2[11]};
  wire [3:0]  tryToRead_lo_lo_11 = {tryToRead_lo_lo_hi_11, tryToRead_lo_lo_lo_11};
  wire [1:0]  tryToRead_lo_hi_lo_11 = {inputSelect1H_5[11], inputSelect1H_4[11]};
  wire [1:0]  tryToRead_lo_hi_hi_11 = {inputSelect1H_7[11], inputSelect1H_6[11]};
  wire [3:0]  tryToRead_lo_hi_11 = {tryToRead_lo_hi_hi_11, tryToRead_lo_hi_lo_11};
  wire [7:0]  tryToRead_lo_11 = {tryToRead_lo_hi_11, tryToRead_lo_lo_11};
  wire [1:0]  tryToRead_hi_lo_lo_11 = {inputSelect1H_9[11], inputSelect1H_8[11]};
  wire [1:0]  tryToRead_hi_lo_hi_11 = {inputSelect1H_11[11], inputSelect1H_10[11]};
  wire [3:0]  tryToRead_hi_lo_11 = {tryToRead_hi_lo_hi_11, tryToRead_hi_lo_lo_11};
  wire [1:0]  tryToRead_hi_hi_lo_11 = {inputSelect1H_13[11], inputSelect1H_12[11]};
  wire [1:0]  tryToRead_hi_hi_hi_11 = {inputSelect1H_15[11], inputSelect1H_14[11]};
  wire [3:0]  tryToRead_hi_hi_11 = {tryToRead_hi_hi_hi_11, tryToRead_hi_hi_lo_11};
  wire [7:0]  tryToRead_hi_11 = {tryToRead_hi_hi_11, tryToRead_hi_lo_11};
  wire [15:0] tryToRead_11 = {tryToRead_hi_11, tryToRead_lo_11};
  wire        output_11_valid_0 = |tryToRead_11;
  wire [4:0]  output_11_bits_vs_0 = selectReq_11_bits_vs;
  wire [1:0]  output_11_bits_offset_0 = selectReq_11_bits_offset;
  wire [3:0]  output_11_bits_writeIndex_0 = selectReq_11_bits_requestIndex;
  wire [1:0]  output_11_bits_dataOffset_0 = selectReq_11_bits_dataOffset;
  assign selectReq_11_bits_dataOffset =
    (tryToRead_11[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_11[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_11[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_11[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_11[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_11[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_11[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_11[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_11[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_11[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_11[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_11[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_11[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_11[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_11[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_11[15] ? input_15_bits_dataOffset_0 : 2'h0);
  assign selectReq_11_bits_requestIndex =
    {3'h0, tryToRead_11[1]} | {2'h0, tryToRead_11[2], 1'h0} | (tryToRead_11[3] ? 4'h3 : 4'h0) | {1'h0, tryToRead_11[4], 2'h0} | (tryToRead_11[5] ? 4'h5 : 4'h0) | (tryToRead_11[6] ? 4'h6 : 4'h0) | (tryToRead_11[7] ? 4'h7 : 4'h0)
    | {tryToRead_11[8], 3'h0} | (tryToRead_11[9] ? 4'h9 : 4'h0) | (tryToRead_11[10] ? 4'hA : 4'h0) | (tryToRead_11[11] ? 4'hB : 4'h0) | (tryToRead_11[12] ? 4'hC : 4'h0) | (tryToRead_11[13] ? 4'hD : 4'h0) | (tryToRead_11[14] ? 4'hE : 4'h0)
    | {4{tryToRead_11[15]}};
  wire [3:0]  selectReq_11_bits_readLane =
    (tryToRead_11[0] ? input_0_bits_readLane_0 : 4'h0) | (tryToRead_11[1] ? input_1_bits_readLane_0 : 4'h0) | (tryToRead_11[2] ? input_2_bits_readLane_0 : 4'h0) | (tryToRead_11[3] ? input_3_bits_readLane_0 : 4'h0)
    | (tryToRead_11[4] ? input_4_bits_readLane_0 : 4'h0) | (tryToRead_11[5] ? input_5_bits_readLane_0 : 4'h0) | (tryToRead_11[6] ? input_6_bits_readLane_0 : 4'h0) | (tryToRead_11[7] ? input_7_bits_readLane_0 : 4'h0)
    | (tryToRead_11[8] ? input_8_bits_readLane_0 : 4'h0) | (tryToRead_11[9] ? input_9_bits_readLane_0 : 4'h0) | (tryToRead_11[10] ? input_10_bits_readLane_0 : 4'h0) | (tryToRead_11[11] ? input_11_bits_readLane_0 : 4'h0)
    | (tryToRead_11[12] ? input_12_bits_readLane_0 : 4'h0) | (tryToRead_11[13] ? input_13_bits_readLane_0 : 4'h0) | (tryToRead_11[14] ? input_14_bits_readLane_0 : 4'h0) | (tryToRead_11[15] ? input_15_bits_readLane_0 : 4'h0);
  assign selectReq_11_bits_offset =
    (tryToRead_11[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead_11[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead_11[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead_11[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead_11[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead_11[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead_11[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead_11[7] ? input_7_bits_offset_0 : 2'h0)
    | (tryToRead_11[8] ? input_8_bits_offset_0 : 2'h0) | (tryToRead_11[9] ? input_9_bits_offset_0 : 2'h0) | (tryToRead_11[10] ? input_10_bits_offset_0 : 2'h0) | (tryToRead_11[11] ? input_11_bits_offset_0 : 2'h0)
    | (tryToRead_11[12] ? input_12_bits_offset_0 : 2'h0) | (tryToRead_11[13] ? input_13_bits_offset_0 : 2'h0) | (tryToRead_11[14] ? input_14_bits_offset_0 : 2'h0) | (tryToRead_11[15] ? input_15_bits_offset_0 : 2'h0);
  assign selectReq_11_bits_vs =
    (tryToRead_11[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_11[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_11[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_11[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_11[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_11[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_11[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_11[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_11[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_11[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_11[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_11[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_11[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_11[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_11[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_11[15] ? input_15_bits_vs_0 : 5'h0);
  wire        selectReq_11_valid =
    tryToRead_11[0] & input_0_valid_0 | tryToRead_11[1] & input_1_valid_0 | tryToRead_11[2] & input_2_valid_0 | tryToRead_11[3] & input_3_valid_0 | tryToRead_11[4] & input_4_valid_0 | tryToRead_11[5] & input_5_valid_0 | tryToRead_11[6]
    & input_6_valid_0 | tryToRead_11[7] & input_7_valid_0 | tryToRead_11[8] & input_8_valid_0 | tryToRead_11[9] & input_9_valid_0 | tryToRead_11[10] & input_10_valid_0 | tryToRead_11[11] & input_11_valid_0 | tryToRead_11[12]
    & input_12_valid_0 | tryToRead_11[13] & input_13_valid_0 | tryToRead_11[14] & input_14_valid_0 | tryToRead_11[15] & input_15_valid_0;
  wire        selectReq_11_ready =
    tryToRead_11[0] & input_0_ready_0 | tryToRead_11[1] & input_1_ready_0 | tryToRead_11[2] & input_2_ready_0 | tryToRead_11[3] & input_3_ready_0 | tryToRead_11[4] & input_4_ready_0 | tryToRead_11[5] & input_5_ready_0 | tryToRead_11[6]
    & input_6_ready_0 | tryToRead_11[7] & input_7_ready_0 | tryToRead_11[8] & input_8_ready_0 | tryToRead_11[9] & input_9_ready_0 | tryToRead_11[10] & input_10_ready_0 | tryToRead_11[11] & input_11_ready_0 | tryToRead_11[12]
    & input_12_ready_0 | tryToRead_11[13] & input_13_ready_0 | tryToRead_11[14] & input_14_ready_0 | tryToRead_11[15] & input_15_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_12 = {inputSelect1H_1[12], inputSelect1H_0[12]};
  wire [1:0]  tryToRead_lo_lo_hi_12 = {inputSelect1H_3[12], inputSelect1H_2[12]};
  wire [3:0]  tryToRead_lo_lo_12 = {tryToRead_lo_lo_hi_12, tryToRead_lo_lo_lo_12};
  wire [1:0]  tryToRead_lo_hi_lo_12 = {inputSelect1H_5[12], inputSelect1H_4[12]};
  wire [1:0]  tryToRead_lo_hi_hi_12 = {inputSelect1H_7[12], inputSelect1H_6[12]};
  wire [3:0]  tryToRead_lo_hi_12 = {tryToRead_lo_hi_hi_12, tryToRead_lo_hi_lo_12};
  wire [7:0]  tryToRead_lo_12 = {tryToRead_lo_hi_12, tryToRead_lo_lo_12};
  wire [1:0]  tryToRead_hi_lo_lo_12 = {inputSelect1H_9[12], inputSelect1H_8[12]};
  wire [1:0]  tryToRead_hi_lo_hi_12 = {inputSelect1H_11[12], inputSelect1H_10[12]};
  wire [3:0]  tryToRead_hi_lo_12 = {tryToRead_hi_lo_hi_12, tryToRead_hi_lo_lo_12};
  wire [1:0]  tryToRead_hi_hi_lo_12 = {inputSelect1H_13[12], inputSelect1H_12[12]};
  wire [1:0]  tryToRead_hi_hi_hi_12 = {inputSelect1H_15[12], inputSelect1H_14[12]};
  wire [3:0]  tryToRead_hi_hi_12 = {tryToRead_hi_hi_hi_12, tryToRead_hi_hi_lo_12};
  wire [7:0]  tryToRead_hi_12 = {tryToRead_hi_hi_12, tryToRead_hi_lo_12};
  wire [15:0] tryToRead_12 = {tryToRead_hi_12, tryToRead_lo_12};
  wire        output_12_valid_0 = |tryToRead_12;
  wire [4:0]  output_12_bits_vs_0 = selectReq_12_bits_vs;
  wire [1:0]  output_12_bits_offset_0 = selectReq_12_bits_offset;
  wire [3:0]  output_12_bits_writeIndex_0 = selectReq_12_bits_requestIndex;
  wire [1:0]  output_12_bits_dataOffset_0 = selectReq_12_bits_dataOffset;
  assign selectReq_12_bits_dataOffset =
    (tryToRead_12[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_12[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_12[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_12[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_12[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_12[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_12[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_12[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_12[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_12[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_12[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_12[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_12[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_12[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_12[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_12[15] ? input_15_bits_dataOffset_0 : 2'h0);
  assign selectReq_12_bits_requestIndex =
    {3'h0, tryToRead_12[1]} | {2'h0, tryToRead_12[2], 1'h0} | (tryToRead_12[3] ? 4'h3 : 4'h0) | {1'h0, tryToRead_12[4], 2'h0} | (tryToRead_12[5] ? 4'h5 : 4'h0) | (tryToRead_12[6] ? 4'h6 : 4'h0) | (tryToRead_12[7] ? 4'h7 : 4'h0)
    | {tryToRead_12[8], 3'h0} | (tryToRead_12[9] ? 4'h9 : 4'h0) | (tryToRead_12[10] ? 4'hA : 4'h0) | (tryToRead_12[11] ? 4'hB : 4'h0) | (tryToRead_12[12] ? 4'hC : 4'h0) | (tryToRead_12[13] ? 4'hD : 4'h0) | (tryToRead_12[14] ? 4'hE : 4'h0)
    | {4{tryToRead_12[15]}};
  wire [3:0]  selectReq_12_bits_readLane =
    (tryToRead_12[0] ? input_0_bits_readLane_0 : 4'h0) | (tryToRead_12[1] ? input_1_bits_readLane_0 : 4'h0) | (tryToRead_12[2] ? input_2_bits_readLane_0 : 4'h0) | (tryToRead_12[3] ? input_3_bits_readLane_0 : 4'h0)
    | (tryToRead_12[4] ? input_4_bits_readLane_0 : 4'h0) | (tryToRead_12[5] ? input_5_bits_readLane_0 : 4'h0) | (tryToRead_12[6] ? input_6_bits_readLane_0 : 4'h0) | (tryToRead_12[7] ? input_7_bits_readLane_0 : 4'h0)
    | (tryToRead_12[8] ? input_8_bits_readLane_0 : 4'h0) | (tryToRead_12[9] ? input_9_bits_readLane_0 : 4'h0) | (tryToRead_12[10] ? input_10_bits_readLane_0 : 4'h0) | (tryToRead_12[11] ? input_11_bits_readLane_0 : 4'h0)
    | (tryToRead_12[12] ? input_12_bits_readLane_0 : 4'h0) | (tryToRead_12[13] ? input_13_bits_readLane_0 : 4'h0) | (tryToRead_12[14] ? input_14_bits_readLane_0 : 4'h0) | (tryToRead_12[15] ? input_15_bits_readLane_0 : 4'h0);
  assign selectReq_12_bits_offset =
    (tryToRead_12[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead_12[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead_12[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead_12[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead_12[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead_12[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead_12[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead_12[7] ? input_7_bits_offset_0 : 2'h0)
    | (tryToRead_12[8] ? input_8_bits_offset_0 : 2'h0) | (tryToRead_12[9] ? input_9_bits_offset_0 : 2'h0) | (tryToRead_12[10] ? input_10_bits_offset_0 : 2'h0) | (tryToRead_12[11] ? input_11_bits_offset_0 : 2'h0)
    | (tryToRead_12[12] ? input_12_bits_offset_0 : 2'h0) | (tryToRead_12[13] ? input_13_bits_offset_0 : 2'h0) | (tryToRead_12[14] ? input_14_bits_offset_0 : 2'h0) | (tryToRead_12[15] ? input_15_bits_offset_0 : 2'h0);
  assign selectReq_12_bits_vs =
    (tryToRead_12[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_12[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_12[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_12[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_12[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_12[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_12[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_12[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_12[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_12[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_12[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_12[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_12[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_12[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_12[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_12[15] ? input_15_bits_vs_0 : 5'h0);
  wire        selectReq_12_valid =
    tryToRead_12[0] & input_0_valid_0 | tryToRead_12[1] & input_1_valid_0 | tryToRead_12[2] & input_2_valid_0 | tryToRead_12[3] & input_3_valid_0 | tryToRead_12[4] & input_4_valid_0 | tryToRead_12[5] & input_5_valid_0 | tryToRead_12[6]
    & input_6_valid_0 | tryToRead_12[7] & input_7_valid_0 | tryToRead_12[8] & input_8_valid_0 | tryToRead_12[9] & input_9_valid_0 | tryToRead_12[10] & input_10_valid_0 | tryToRead_12[11] & input_11_valid_0 | tryToRead_12[12]
    & input_12_valid_0 | tryToRead_12[13] & input_13_valid_0 | tryToRead_12[14] & input_14_valid_0 | tryToRead_12[15] & input_15_valid_0;
  wire        selectReq_12_ready =
    tryToRead_12[0] & input_0_ready_0 | tryToRead_12[1] & input_1_ready_0 | tryToRead_12[2] & input_2_ready_0 | tryToRead_12[3] & input_3_ready_0 | tryToRead_12[4] & input_4_ready_0 | tryToRead_12[5] & input_5_ready_0 | tryToRead_12[6]
    & input_6_ready_0 | tryToRead_12[7] & input_7_ready_0 | tryToRead_12[8] & input_8_ready_0 | tryToRead_12[9] & input_9_ready_0 | tryToRead_12[10] & input_10_ready_0 | tryToRead_12[11] & input_11_ready_0 | tryToRead_12[12]
    & input_12_ready_0 | tryToRead_12[13] & input_13_ready_0 | tryToRead_12[14] & input_14_ready_0 | tryToRead_12[15] & input_15_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_13 = {inputSelect1H_1[13], inputSelect1H_0[13]};
  wire [1:0]  tryToRead_lo_lo_hi_13 = {inputSelect1H_3[13], inputSelect1H_2[13]};
  wire [3:0]  tryToRead_lo_lo_13 = {tryToRead_lo_lo_hi_13, tryToRead_lo_lo_lo_13};
  wire [1:0]  tryToRead_lo_hi_lo_13 = {inputSelect1H_5[13], inputSelect1H_4[13]};
  wire [1:0]  tryToRead_lo_hi_hi_13 = {inputSelect1H_7[13], inputSelect1H_6[13]};
  wire [3:0]  tryToRead_lo_hi_13 = {tryToRead_lo_hi_hi_13, tryToRead_lo_hi_lo_13};
  wire [7:0]  tryToRead_lo_13 = {tryToRead_lo_hi_13, tryToRead_lo_lo_13};
  wire [1:0]  tryToRead_hi_lo_lo_13 = {inputSelect1H_9[13], inputSelect1H_8[13]};
  wire [1:0]  tryToRead_hi_lo_hi_13 = {inputSelect1H_11[13], inputSelect1H_10[13]};
  wire [3:0]  tryToRead_hi_lo_13 = {tryToRead_hi_lo_hi_13, tryToRead_hi_lo_lo_13};
  wire [1:0]  tryToRead_hi_hi_lo_13 = {inputSelect1H_13[13], inputSelect1H_12[13]};
  wire [1:0]  tryToRead_hi_hi_hi_13 = {inputSelect1H_15[13], inputSelect1H_14[13]};
  wire [3:0]  tryToRead_hi_hi_13 = {tryToRead_hi_hi_hi_13, tryToRead_hi_hi_lo_13};
  wire [7:0]  tryToRead_hi_13 = {tryToRead_hi_hi_13, tryToRead_hi_lo_13};
  wire [15:0] tryToRead_13 = {tryToRead_hi_13, tryToRead_lo_13};
  wire        output_13_valid_0 = |tryToRead_13;
  wire [4:0]  output_13_bits_vs_0 = selectReq_13_bits_vs;
  wire [1:0]  output_13_bits_offset_0 = selectReq_13_bits_offset;
  wire [3:0]  output_13_bits_writeIndex_0 = selectReq_13_bits_requestIndex;
  wire [1:0]  output_13_bits_dataOffset_0 = selectReq_13_bits_dataOffset;
  assign selectReq_13_bits_dataOffset =
    (tryToRead_13[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_13[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_13[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_13[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_13[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_13[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_13[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_13[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_13[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_13[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_13[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_13[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_13[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_13[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_13[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_13[15] ? input_15_bits_dataOffset_0 : 2'h0);
  assign selectReq_13_bits_requestIndex =
    {3'h0, tryToRead_13[1]} | {2'h0, tryToRead_13[2], 1'h0} | (tryToRead_13[3] ? 4'h3 : 4'h0) | {1'h0, tryToRead_13[4], 2'h0} | (tryToRead_13[5] ? 4'h5 : 4'h0) | (tryToRead_13[6] ? 4'h6 : 4'h0) | (tryToRead_13[7] ? 4'h7 : 4'h0)
    | {tryToRead_13[8], 3'h0} | (tryToRead_13[9] ? 4'h9 : 4'h0) | (tryToRead_13[10] ? 4'hA : 4'h0) | (tryToRead_13[11] ? 4'hB : 4'h0) | (tryToRead_13[12] ? 4'hC : 4'h0) | (tryToRead_13[13] ? 4'hD : 4'h0) | (tryToRead_13[14] ? 4'hE : 4'h0)
    | {4{tryToRead_13[15]}};
  wire [3:0]  selectReq_13_bits_readLane =
    (tryToRead_13[0] ? input_0_bits_readLane_0 : 4'h0) | (tryToRead_13[1] ? input_1_bits_readLane_0 : 4'h0) | (tryToRead_13[2] ? input_2_bits_readLane_0 : 4'h0) | (tryToRead_13[3] ? input_3_bits_readLane_0 : 4'h0)
    | (tryToRead_13[4] ? input_4_bits_readLane_0 : 4'h0) | (tryToRead_13[5] ? input_5_bits_readLane_0 : 4'h0) | (tryToRead_13[6] ? input_6_bits_readLane_0 : 4'h0) | (tryToRead_13[7] ? input_7_bits_readLane_0 : 4'h0)
    | (tryToRead_13[8] ? input_8_bits_readLane_0 : 4'h0) | (tryToRead_13[9] ? input_9_bits_readLane_0 : 4'h0) | (tryToRead_13[10] ? input_10_bits_readLane_0 : 4'h0) | (tryToRead_13[11] ? input_11_bits_readLane_0 : 4'h0)
    | (tryToRead_13[12] ? input_12_bits_readLane_0 : 4'h0) | (tryToRead_13[13] ? input_13_bits_readLane_0 : 4'h0) | (tryToRead_13[14] ? input_14_bits_readLane_0 : 4'h0) | (tryToRead_13[15] ? input_15_bits_readLane_0 : 4'h0);
  assign selectReq_13_bits_offset =
    (tryToRead_13[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead_13[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead_13[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead_13[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead_13[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead_13[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead_13[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead_13[7] ? input_7_bits_offset_0 : 2'h0)
    | (tryToRead_13[8] ? input_8_bits_offset_0 : 2'h0) | (tryToRead_13[9] ? input_9_bits_offset_0 : 2'h0) | (tryToRead_13[10] ? input_10_bits_offset_0 : 2'h0) | (tryToRead_13[11] ? input_11_bits_offset_0 : 2'h0)
    | (tryToRead_13[12] ? input_12_bits_offset_0 : 2'h0) | (tryToRead_13[13] ? input_13_bits_offset_0 : 2'h0) | (tryToRead_13[14] ? input_14_bits_offset_0 : 2'h0) | (tryToRead_13[15] ? input_15_bits_offset_0 : 2'h0);
  assign selectReq_13_bits_vs =
    (tryToRead_13[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_13[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_13[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_13[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_13[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_13[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_13[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_13[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_13[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_13[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_13[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_13[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_13[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_13[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_13[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_13[15] ? input_15_bits_vs_0 : 5'h0);
  wire        selectReq_13_valid =
    tryToRead_13[0] & input_0_valid_0 | tryToRead_13[1] & input_1_valid_0 | tryToRead_13[2] & input_2_valid_0 | tryToRead_13[3] & input_3_valid_0 | tryToRead_13[4] & input_4_valid_0 | tryToRead_13[5] & input_5_valid_0 | tryToRead_13[6]
    & input_6_valid_0 | tryToRead_13[7] & input_7_valid_0 | tryToRead_13[8] & input_8_valid_0 | tryToRead_13[9] & input_9_valid_0 | tryToRead_13[10] & input_10_valid_0 | tryToRead_13[11] & input_11_valid_0 | tryToRead_13[12]
    & input_12_valid_0 | tryToRead_13[13] & input_13_valid_0 | tryToRead_13[14] & input_14_valid_0 | tryToRead_13[15] & input_15_valid_0;
  wire        selectReq_13_ready =
    tryToRead_13[0] & input_0_ready_0 | tryToRead_13[1] & input_1_ready_0 | tryToRead_13[2] & input_2_ready_0 | tryToRead_13[3] & input_3_ready_0 | tryToRead_13[4] & input_4_ready_0 | tryToRead_13[5] & input_5_ready_0 | tryToRead_13[6]
    & input_6_ready_0 | tryToRead_13[7] & input_7_ready_0 | tryToRead_13[8] & input_8_ready_0 | tryToRead_13[9] & input_9_ready_0 | tryToRead_13[10] & input_10_ready_0 | tryToRead_13[11] & input_11_ready_0 | tryToRead_13[12]
    & input_12_ready_0 | tryToRead_13[13] & input_13_ready_0 | tryToRead_13[14] & input_14_ready_0 | tryToRead_13[15] & input_15_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_14 = {inputSelect1H_1[14], inputSelect1H_0[14]};
  wire [1:0]  tryToRead_lo_lo_hi_14 = {inputSelect1H_3[14], inputSelect1H_2[14]};
  wire [3:0]  tryToRead_lo_lo_14 = {tryToRead_lo_lo_hi_14, tryToRead_lo_lo_lo_14};
  wire [1:0]  tryToRead_lo_hi_lo_14 = {inputSelect1H_5[14], inputSelect1H_4[14]};
  wire [1:0]  tryToRead_lo_hi_hi_14 = {inputSelect1H_7[14], inputSelect1H_6[14]};
  wire [3:0]  tryToRead_lo_hi_14 = {tryToRead_lo_hi_hi_14, tryToRead_lo_hi_lo_14};
  wire [7:0]  tryToRead_lo_14 = {tryToRead_lo_hi_14, tryToRead_lo_lo_14};
  wire [1:0]  tryToRead_hi_lo_lo_14 = {inputSelect1H_9[14], inputSelect1H_8[14]};
  wire [1:0]  tryToRead_hi_lo_hi_14 = {inputSelect1H_11[14], inputSelect1H_10[14]};
  wire [3:0]  tryToRead_hi_lo_14 = {tryToRead_hi_lo_hi_14, tryToRead_hi_lo_lo_14};
  wire [1:0]  tryToRead_hi_hi_lo_14 = {inputSelect1H_13[14], inputSelect1H_12[14]};
  wire [1:0]  tryToRead_hi_hi_hi_14 = {inputSelect1H_15[14], inputSelect1H_14[14]};
  wire [3:0]  tryToRead_hi_hi_14 = {tryToRead_hi_hi_hi_14, tryToRead_hi_hi_lo_14};
  wire [7:0]  tryToRead_hi_14 = {tryToRead_hi_hi_14, tryToRead_hi_lo_14};
  wire [15:0] tryToRead_14 = {tryToRead_hi_14, tryToRead_lo_14};
  wire        output_14_valid_0 = |tryToRead_14;
  wire [4:0]  output_14_bits_vs_0 = selectReq_14_bits_vs;
  wire [1:0]  output_14_bits_offset_0 = selectReq_14_bits_offset;
  wire [3:0]  output_14_bits_writeIndex_0 = selectReq_14_bits_requestIndex;
  wire [1:0]  output_14_bits_dataOffset_0 = selectReq_14_bits_dataOffset;
  assign selectReq_14_bits_dataOffset =
    (tryToRead_14[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_14[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_14[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_14[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_14[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_14[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_14[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_14[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_14[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_14[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_14[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_14[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_14[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_14[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_14[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_14[15] ? input_15_bits_dataOffset_0 : 2'h0);
  assign selectReq_14_bits_requestIndex =
    {3'h0, tryToRead_14[1]} | {2'h0, tryToRead_14[2], 1'h0} | (tryToRead_14[3] ? 4'h3 : 4'h0) | {1'h0, tryToRead_14[4], 2'h0} | (tryToRead_14[5] ? 4'h5 : 4'h0) | (tryToRead_14[6] ? 4'h6 : 4'h0) | (tryToRead_14[7] ? 4'h7 : 4'h0)
    | {tryToRead_14[8], 3'h0} | (tryToRead_14[9] ? 4'h9 : 4'h0) | (tryToRead_14[10] ? 4'hA : 4'h0) | (tryToRead_14[11] ? 4'hB : 4'h0) | (tryToRead_14[12] ? 4'hC : 4'h0) | (tryToRead_14[13] ? 4'hD : 4'h0) | (tryToRead_14[14] ? 4'hE : 4'h0)
    | {4{tryToRead_14[15]}};
  wire [3:0]  selectReq_14_bits_readLane =
    (tryToRead_14[0] ? input_0_bits_readLane_0 : 4'h0) | (tryToRead_14[1] ? input_1_bits_readLane_0 : 4'h0) | (tryToRead_14[2] ? input_2_bits_readLane_0 : 4'h0) | (tryToRead_14[3] ? input_3_bits_readLane_0 : 4'h0)
    | (tryToRead_14[4] ? input_4_bits_readLane_0 : 4'h0) | (tryToRead_14[5] ? input_5_bits_readLane_0 : 4'h0) | (tryToRead_14[6] ? input_6_bits_readLane_0 : 4'h0) | (tryToRead_14[7] ? input_7_bits_readLane_0 : 4'h0)
    | (tryToRead_14[8] ? input_8_bits_readLane_0 : 4'h0) | (tryToRead_14[9] ? input_9_bits_readLane_0 : 4'h0) | (tryToRead_14[10] ? input_10_bits_readLane_0 : 4'h0) | (tryToRead_14[11] ? input_11_bits_readLane_0 : 4'h0)
    | (tryToRead_14[12] ? input_12_bits_readLane_0 : 4'h0) | (tryToRead_14[13] ? input_13_bits_readLane_0 : 4'h0) | (tryToRead_14[14] ? input_14_bits_readLane_0 : 4'h0) | (tryToRead_14[15] ? input_15_bits_readLane_0 : 4'h0);
  assign selectReq_14_bits_offset =
    (tryToRead_14[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead_14[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead_14[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead_14[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead_14[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead_14[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead_14[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead_14[7] ? input_7_bits_offset_0 : 2'h0)
    | (tryToRead_14[8] ? input_8_bits_offset_0 : 2'h0) | (tryToRead_14[9] ? input_9_bits_offset_0 : 2'h0) | (tryToRead_14[10] ? input_10_bits_offset_0 : 2'h0) | (tryToRead_14[11] ? input_11_bits_offset_0 : 2'h0)
    | (tryToRead_14[12] ? input_12_bits_offset_0 : 2'h0) | (tryToRead_14[13] ? input_13_bits_offset_0 : 2'h0) | (tryToRead_14[14] ? input_14_bits_offset_0 : 2'h0) | (tryToRead_14[15] ? input_15_bits_offset_0 : 2'h0);
  assign selectReq_14_bits_vs =
    (tryToRead_14[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_14[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_14[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_14[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_14[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_14[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_14[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_14[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_14[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_14[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_14[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_14[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_14[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_14[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_14[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_14[15] ? input_15_bits_vs_0 : 5'h0);
  wire        selectReq_14_valid =
    tryToRead_14[0] & input_0_valid_0 | tryToRead_14[1] & input_1_valid_0 | tryToRead_14[2] & input_2_valid_0 | tryToRead_14[3] & input_3_valid_0 | tryToRead_14[4] & input_4_valid_0 | tryToRead_14[5] & input_5_valid_0 | tryToRead_14[6]
    & input_6_valid_0 | tryToRead_14[7] & input_7_valid_0 | tryToRead_14[8] & input_8_valid_0 | tryToRead_14[9] & input_9_valid_0 | tryToRead_14[10] & input_10_valid_0 | tryToRead_14[11] & input_11_valid_0 | tryToRead_14[12]
    & input_12_valid_0 | tryToRead_14[13] & input_13_valid_0 | tryToRead_14[14] & input_14_valid_0 | tryToRead_14[15] & input_15_valid_0;
  wire        selectReq_14_ready =
    tryToRead_14[0] & input_0_ready_0 | tryToRead_14[1] & input_1_ready_0 | tryToRead_14[2] & input_2_ready_0 | tryToRead_14[3] & input_3_ready_0 | tryToRead_14[4] & input_4_ready_0 | tryToRead_14[5] & input_5_ready_0 | tryToRead_14[6]
    & input_6_ready_0 | tryToRead_14[7] & input_7_ready_0 | tryToRead_14[8] & input_8_ready_0 | tryToRead_14[9] & input_9_ready_0 | tryToRead_14[10] & input_10_ready_0 | tryToRead_14[11] & input_11_ready_0 | tryToRead_14[12]
    & input_12_ready_0 | tryToRead_14[13] & input_13_ready_0 | tryToRead_14[14] & input_14_ready_0 | tryToRead_14[15] & input_15_ready_0;
  wire [1:0]  tryToRead_lo_lo_lo_15 = {inputSelect1H_1[15], inputSelect1H_0[15]};
  wire [1:0]  tryToRead_lo_lo_hi_15 = {inputSelect1H_3[15], inputSelect1H_2[15]};
  wire [3:0]  tryToRead_lo_lo_15 = {tryToRead_lo_lo_hi_15, tryToRead_lo_lo_lo_15};
  wire [1:0]  tryToRead_lo_hi_lo_15 = {inputSelect1H_5[15], inputSelect1H_4[15]};
  wire [1:0]  tryToRead_lo_hi_hi_15 = {inputSelect1H_7[15], inputSelect1H_6[15]};
  wire [3:0]  tryToRead_lo_hi_15 = {tryToRead_lo_hi_hi_15, tryToRead_lo_hi_lo_15};
  wire [7:0]  tryToRead_lo_15 = {tryToRead_lo_hi_15, tryToRead_lo_lo_15};
  wire [1:0]  tryToRead_hi_lo_lo_15 = {inputSelect1H_9[15], inputSelect1H_8[15]};
  wire [1:0]  tryToRead_hi_lo_hi_15 = {inputSelect1H_11[15], inputSelect1H_10[15]};
  wire [3:0]  tryToRead_hi_lo_15 = {tryToRead_hi_lo_hi_15, tryToRead_hi_lo_lo_15};
  wire [1:0]  tryToRead_hi_hi_lo_15 = {inputSelect1H_13[15], inputSelect1H_12[15]};
  wire [1:0]  tryToRead_hi_hi_hi_15 = {inputSelect1H_15[15], inputSelect1H_14[15]};
  wire [3:0]  tryToRead_hi_hi_15 = {tryToRead_hi_hi_hi_15, tryToRead_hi_hi_lo_15};
  wire [7:0]  tryToRead_hi_15 = {tryToRead_hi_hi_15, tryToRead_hi_lo_15};
  wire [15:0] tryToRead_15 = {tryToRead_hi_15, tryToRead_lo_15};
  wire        output_15_valid_0 = |tryToRead_15;
  wire [4:0]  output_15_bits_vs_0 = selectReq_15_bits_vs;
  wire [1:0]  output_15_bits_offset_0 = selectReq_15_bits_offset;
  wire [3:0]  output_15_bits_writeIndex_0 = selectReq_15_bits_requestIndex;
  wire [1:0]  output_15_bits_dataOffset_0 = selectReq_15_bits_dataOffset;
  assign selectReq_15_bits_dataOffset =
    (tryToRead_15[0] ? input_0_bits_dataOffset_0 : 2'h0) | (tryToRead_15[1] ? input_1_bits_dataOffset_0 : 2'h0) | (tryToRead_15[2] ? input_2_bits_dataOffset_0 : 2'h0) | (tryToRead_15[3] ? input_3_bits_dataOffset_0 : 2'h0)
    | (tryToRead_15[4] ? input_4_bits_dataOffset_0 : 2'h0) | (tryToRead_15[5] ? input_5_bits_dataOffset_0 : 2'h0) | (tryToRead_15[6] ? input_6_bits_dataOffset_0 : 2'h0) | (tryToRead_15[7] ? input_7_bits_dataOffset_0 : 2'h0)
    | (tryToRead_15[8] ? input_8_bits_dataOffset_0 : 2'h0) | (tryToRead_15[9] ? input_9_bits_dataOffset_0 : 2'h0) | (tryToRead_15[10] ? input_10_bits_dataOffset_0 : 2'h0) | (tryToRead_15[11] ? input_11_bits_dataOffset_0 : 2'h0)
    | (tryToRead_15[12] ? input_12_bits_dataOffset_0 : 2'h0) | (tryToRead_15[13] ? input_13_bits_dataOffset_0 : 2'h0) | (tryToRead_15[14] ? input_14_bits_dataOffset_0 : 2'h0) | (tryToRead_15[15] ? input_15_bits_dataOffset_0 : 2'h0);
  assign selectReq_15_bits_requestIndex =
    {3'h0, tryToRead_15[1]} | {2'h0, tryToRead_15[2], 1'h0} | (tryToRead_15[3] ? 4'h3 : 4'h0) | {1'h0, tryToRead_15[4], 2'h0} | (tryToRead_15[5] ? 4'h5 : 4'h0) | (tryToRead_15[6] ? 4'h6 : 4'h0) | (tryToRead_15[7] ? 4'h7 : 4'h0)
    | {tryToRead_15[8], 3'h0} | (tryToRead_15[9] ? 4'h9 : 4'h0) | (tryToRead_15[10] ? 4'hA : 4'h0) | (tryToRead_15[11] ? 4'hB : 4'h0) | (tryToRead_15[12] ? 4'hC : 4'h0) | (tryToRead_15[13] ? 4'hD : 4'h0) | (tryToRead_15[14] ? 4'hE : 4'h0)
    | {4{tryToRead_15[15]}};
  wire [3:0]  selectReq_15_bits_readLane =
    (tryToRead_15[0] ? input_0_bits_readLane_0 : 4'h0) | (tryToRead_15[1] ? input_1_bits_readLane_0 : 4'h0) | (tryToRead_15[2] ? input_2_bits_readLane_0 : 4'h0) | (tryToRead_15[3] ? input_3_bits_readLane_0 : 4'h0)
    | (tryToRead_15[4] ? input_4_bits_readLane_0 : 4'h0) | (tryToRead_15[5] ? input_5_bits_readLane_0 : 4'h0) | (tryToRead_15[6] ? input_6_bits_readLane_0 : 4'h0) | (tryToRead_15[7] ? input_7_bits_readLane_0 : 4'h0)
    | (tryToRead_15[8] ? input_8_bits_readLane_0 : 4'h0) | (tryToRead_15[9] ? input_9_bits_readLane_0 : 4'h0) | (tryToRead_15[10] ? input_10_bits_readLane_0 : 4'h0) | (tryToRead_15[11] ? input_11_bits_readLane_0 : 4'h0)
    | (tryToRead_15[12] ? input_12_bits_readLane_0 : 4'h0) | (tryToRead_15[13] ? input_13_bits_readLane_0 : 4'h0) | (tryToRead_15[14] ? input_14_bits_readLane_0 : 4'h0) | (tryToRead_15[15] ? input_15_bits_readLane_0 : 4'h0);
  assign selectReq_15_bits_offset =
    (tryToRead_15[0] ? input_0_bits_offset_0 : 2'h0) | (tryToRead_15[1] ? input_1_bits_offset_0 : 2'h0) | (tryToRead_15[2] ? input_2_bits_offset_0 : 2'h0) | (tryToRead_15[3] ? input_3_bits_offset_0 : 2'h0)
    | (tryToRead_15[4] ? input_4_bits_offset_0 : 2'h0) | (tryToRead_15[5] ? input_5_bits_offset_0 : 2'h0) | (tryToRead_15[6] ? input_6_bits_offset_0 : 2'h0) | (tryToRead_15[7] ? input_7_bits_offset_0 : 2'h0)
    | (tryToRead_15[8] ? input_8_bits_offset_0 : 2'h0) | (tryToRead_15[9] ? input_9_bits_offset_0 : 2'h0) | (tryToRead_15[10] ? input_10_bits_offset_0 : 2'h0) | (tryToRead_15[11] ? input_11_bits_offset_0 : 2'h0)
    | (tryToRead_15[12] ? input_12_bits_offset_0 : 2'h0) | (tryToRead_15[13] ? input_13_bits_offset_0 : 2'h0) | (tryToRead_15[14] ? input_14_bits_offset_0 : 2'h0) | (tryToRead_15[15] ? input_15_bits_offset_0 : 2'h0);
  assign selectReq_15_bits_vs =
    (tryToRead_15[0] ? input_0_bits_vs_0 : 5'h0) | (tryToRead_15[1] ? input_1_bits_vs_0 : 5'h0) | (tryToRead_15[2] ? input_2_bits_vs_0 : 5'h0) | (tryToRead_15[3] ? input_3_bits_vs_0 : 5'h0) | (tryToRead_15[4] ? input_4_bits_vs_0 : 5'h0)
    | (tryToRead_15[5] ? input_5_bits_vs_0 : 5'h0) | (tryToRead_15[6] ? input_6_bits_vs_0 : 5'h0) | (tryToRead_15[7] ? input_7_bits_vs_0 : 5'h0) | (tryToRead_15[8] ? input_8_bits_vs_0 : 5'h0) | (tryToRead_15[9] ? input_9_bits_vs_0 : 5'h0)
    | (tryToRead_15[10] ? input_10_bits_vs_0 : 5'h0) | (tryToRead_15[11] ? input_11_bits_vs_0 : 5'h0) | (tryToRead_15[12] ? input_12_bits_vs_0 : 5'h0) | (tryToRead_15[13] ? input_13_bits_vs_0 : 5'h0)
    | (tryToRead_15[14] ? input_14_bits_vs_0 : 5'h0) | (tryToRead_15[15] ? input_15_bits_vs_0 : 5'h0);
  wire        selectReq_15_valid =
    tryToRead_15[0] & input_0_valid_0 | tryToRead_15[1] & input_1_valid_0 | tryToRead_15[2] & input_2_valid_0 | tryToRead_15[3] & input_3_valid_0 | tryToRead_15[4] & input_4_valid_0 | tryToRead_15[5] & input_5_valid_0 | tryToRead_15[6]
    & input_6_valid_0 | tryToRead_15[7] & input_7_valid_0 | tryToRead_15[8] & input_8_valid_0 | tryToRead_15[9] & input_9_valid_0 | tryToRead_15[10] & input_10_valid_0 | tryToRead_15[11] & input_11_valid_0 | tryToRead_15[12]
    & input_12_valid_0 | tryToRead_15[13] & input_13_valid_0 | tryToRead_15[14] & input_14_valid_0 | tryToRead_15[15] & input_15_valid_0;
  wire        selectReq_15_ready =
    tryToRead_15[0] & input_0_ready_0 | tryToRead_15[1] & input_1_ready_0 | tryToRead_15[2] & input_2_ready_0 | tryToRead_15[3] & input_3_ready_0 | tryToRead_15[4] & input_4_ready_0 | tryToRead_15[5] & input_5_ready_0 | tryToRead_15[6]
    & input_6_ready_0 | tryToRead_15[7] & input_7_ready_0 | tryToRead_15[8] & input_8_ready_0 | tryToRead_15[9] & input_9_ready_0 | tryToRead_15[10] & input_10_ready_0 | tryToRead_15[11] & input_11_ready_0 | tryToRead_15[12]
    & input_12_ready_0 | tryToRead_15[13] & input_13_ready_0 | tryToRead_15[14] & input_14_ready_0 | tryToRead_15[15] & input_15_ready_0;
  assign input_0_ready = input_0_ready_0;
  assign input_1_ready = input_1_ready_0;
  assign input_2_ready = input_2_ready_0;
  assign input_3_ready = input_3_ready_0;
  assign input_4_ready = input_4_ready_0;
  assign input_5_ready = input_5_ready_0;
  assign input_6_ready = input_6_ready_0;
  assign input_7_ready = input_7_ready_0;
  assign input_8_ready = input_8_ready_0;
  assign input_9_ready = input_9_ready_0;
  assign input_10_ready = input_10_ready_0;
  assign input_11_ready = input_11_ready_0;
  assign input_12_ready = input_12_ready_0;
  assign input_13_ready = input_13_ready_0;
  assign input_14_ready = input_14_ready_0;
  assign input_15_ready = input_15_ready_0;
  assign output_0_valid = output_0_valid_0;
  assign output_0_bits_vs = output_0_bits_vs_0;
  assign output_0_bits_offset = output_0_bits_offset_0;
  assign output_0_bits_writeIndex = output_0_bits_writeIndex_0;
  assign output_0_bits_dataOffset = output_0_bits_dataOffset_0;
  assign output_1_valid = output_1_valid_0;
  assign output_1_bits_vs = output_1_bits_vs_0;
  assign output_1_bits_offset = output_1_bits_offset_0;
  assign output_1_bits_writeIndex = output_1_bits_writeIndex_0;
  assign output_1_bits_dataOffset = output_1_bits_dataOffset_0;
  assign output_2_valid = output_2_valid_0;
  assign output_2_bits_vs = output_2_bits_vs_0;
  assign output_2_bits_offset = output_2_bits_offset_0;
  assign output_2_bits_writeIndex = output_2_bits_writeIndex_0;
  assign output_2_bits_dataOffset = output_2_bits_dataOffset_0;
  assign output_3_valid = output_3_valid_0;
  assign output_3_bits_vs = output_3_bits_vs_0;
  assign output_3_bits_offset = output_3_bits_offset_0;
  assign output_3_bits_writeIndex = output_3_bits_writeIndex_0;
  assign output_3_bits_dataOffset = output_3_bits_dataOffset_0;
  assign output_4_valid = output_4_valid_0;
  assign output_4_bits_vs = output_4_bits_vs_0;
  assign output_4_bits_offset = output_4_bits_offset_0;
  assign output_4_bits_writeIndex = output_4_bits_writeIndex_0;
  assign output_4_bits_dataOffset = output_4_bits_dataOffset_0;
  assign output_5_valid = output_5_valid_0;
  assign output_5_bits_vs = output_5_bits_vs_0;
  assign output_5_bits_offset = output_5_bits_offset_0;
  assign output_5_bits_writeIndex = output_5_bits_writeIndex_0;
  assign output_5_bits_dataOffset = output_5_bits_dataOffset_0;
  assign output_6_valid = output_6_valid_0;
  assign output_6_bits_vs = output_6_bits_vs_0;
  assign output_6_bits_offset = output_6_bits_offset_0;
  assign output_6_bits_writeIndex = output_6_bits_writeIndex_0;
  assign output_6_bits_dataOffset = output_6_bits_dataOffset_0;
  assign output_7_valid = output_7_valid_0;
  assign output_7_bits_vs = output_7_bits_vs_0;
  assign output_7_bits_offset = output_7_bits_offset_0;
  assign output_7_bits_writeIndex = output_7_bits_writeIndex_0;
  assign output_7_bits_dataOffset = output_7_bits_dataOffset_0;
  assign output_8_valid = output_8_valid_0;
  assign output_8_bits_vs = output_8_bits_vs_0;
  assign output_8_bits_offset = output_8_bits_offset_0;
  assign output_8_bits_writeIndex = output_8_bits_writeIndex_0;
  assign output_8_bits_dataOffset = output_8_bits_dataOffset_0;
  assign output_9_valid = output_9_valid_0;
  assign output_9_bits_vs = output_9_bits_vs_0;
  assign output_9_bits_offset = output_9_bits_offset_0;
  assign output_9_bits_writeIndex = output_9_bits_writeIndex_0;
  assign output_9_bits_dataOffset = output_9_bits_dataOffset_0;
  assign output_10_valid = output_10_valid_0;
  assign output_10_bits_vs = output_10_bits_vs_0;
  assign output_10_bits_offset = output_10_bits_offset_0;
  assign output_10_bits_writeIndex = output_10_bits_writeIndex_0;
  assign output_10_bits_dataOffset = output_10_bits_dataOffset_0;
  assign output_11_valid = output_11_valid_0;
  assign output_11_bits_vs = output_11_bits_vs_0;
  assign output_11_bits_offset = output_11_bits_offset_0;
  assign output_11_bits_writeIndex = output_11_bits_writeIndex_0;
  assign output_11_bits_dataOffset = output_11_bits_dataOffset_0;
  assign output_12_valid = output_12_valid_0;
  assign output_12_bits_vs = output_12_bits_vs_0;
  assign output_12_bits_offset = output_12_bits_offset_0;
  assign output_12_bits_writeIndex = output_12_bits_writeIndex_0;
  assign output_12_bits_dataOffset = output_12_bits_dataOffset_0;
  assign output_13_valid = output_13_valid_0;
  assign output_13_bits_vs = output_13_bits_vs_0;
  assign output_13_bits_offset = output_13_bits_offset_0;
  assign output_13_bits_writeIndex = output_13_bits_writeIndex_0;
  assign output_13_bits_dataOffset = output_13_bits_dataOffset_0;
  assign output_14_valid = output_14_valid_0;
  assign output_14_bits_vs = output_14_bits_vs_0;
  assign output_14_bits_offset = output_14_bits_offset_0;
  assign output_14_bits_writeIndex = output_14_bits_writeIndex_0;
  assign output_14_bits_dataOffset = output_14_bits_dataOffset_0;
  assign output_15_valid = output_15_valid_0;
  assign output_15_bits_vs = output_15_bits_vs_0;
  assign output_15_bits_offset = output_15_bits_offset_0;
  assign output_15_bits_writeIndex = output_15_bits_writeIndex_0;
  assign output_15_bits_dataOffset = output_15_bits_dataOffset_0;
endmodule

