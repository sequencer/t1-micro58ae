
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module MaskUnit(
  input         clock,
                reset,
                instReq_valid,
  input  [2:0]  instReq_bits_instructionIndex,
  input         instReq_bits_decodeResult_specialSlot,
  input  [4:0]  instReq_bits_decodeResult_topUop,
  input         instReq_bits_decodeResult_popCount,
                instReq_bits_decodeResult_ffo,
                instReq_bits_decodeResult_average,
                instReq_bits_decodeResult_reverse,
                instReq_bits_decodeResult_dontNeedExecuteInLane,
                instReq_bits_decodeResult_scheduler,
                instReq_bits_decodeResult_sReadVD,
                instReq_bits_decodeResult_vtype,
                instReq_bits_decodeResult_sWrite,
                instReq_bits_decodeResult_crossRead,
                instReq_bits_decodeResult_crossWrite,
                instReq_bits_decodeResult_maskUnit,
                instReq_bits_decodeResult_special,
                instReq_bits_decodeResult_saturate,
                instReq_bits_decodeResult_vwmacc,
                instReq_bits_decodeResult_readOnly,
                instReq_bits_decodeResult_maskSource,
                instReq_bits_decodeResult_maskDestination,
                instReq_bits_decodeResult_maskLogic,
  input  [3:0]  instReq_bits_decodeResult_uop,
  input         instReq_bits_decodeResult_iota,
                instReq_bits_decodeResult_mv,
                instReq_bits_decodeResult_extend,
                instReq_bits_decodeResult_unOrderWrite,
                instReq_bits_decodeResult_compress,
                instReq_bits_decodeResult_gather16,
                instReq_bits_decodeResult_gather,
                instReq_bits_decodeResult_slid,
                instReq_bits_decodeResult_targetRd,
                instReq_bits_decodeResult_widenReduce,
                instReq_bits_decodeResult_red,
                instReq_bits_decodeResult_nr,
                instReq_bits_decodeResult_itype,
                instReq_bits_decodeResult_unsigned1,
                instReq_bits_decodeResult_unsigned0,
                instReq_bits_decodeResult_other,
                instReq_bits_decodeResult_multiCycle,
                instReq_bits_decodeResult_divider,
                instReq_bits_decodeResult_multiplier,
                instReq_bits_decodeResult_shift,
                instReq_bits_decodeResult_adder,
                instReq_bits_decodeResult_logic,
  input  [31:0] instReq_bits_readFromScala,
  input  [1:0]  instReq_bits_sew,
  input  [2:0]  instReq_bits_vlmul,
  input         instReq_bits_maskType,
  input  [2:0]  instReq_bits_vxrm,
  input  [4:0]  instReq_bits_vs2,
                instReq_bits_vs1,
                instReq_bits_vd,
  input  [11:0] instReq_bits_vl,
  input         exeReq_0_valid,
  input  [31:0] exeReq_0_bits_source1,
                exeReq_0_bits_source2,
  input  [2:0]  exeReq_0_bits_index,
  input         exeReq_0_bits_ffo,
                exeReq_1_valid,
  input  [31:0] exeReq_1_bits_source1,
                exeReq_1_bits_source2,
  input  [2:0]  exeReq_1_bits_index,
  input         exeReq_1_bits_ffo,
                exeReq_2_valid,
  input  [31:0] exeReq_2_bits_source1,
                exeReq_2_bits_source2,
  input  [2:0]  exeReq_2_bits_index,
  input         exeReq_2_bits_ffo,
                exeReq_3_valid,
  input  [31:0] exeReq_3_bits_source1,
                exeReq_3_bits_source2,
  input  [2:0]  exeReq_3_bits_index,
  input         exeReq_3_bits_ffo,
                exeReq_4_valid,
  input  [31:0] exeReq_4_bits_source1,
                exeReq_4_bits_source2,
  input  [2:0]  exeReq_4_bits_index,
  input         exeReq_4_bits_ffo,
                exeReq_5_valid,
  input  [31:0] exeReq_5_bits_source1,
                exeReq_5_bits_source2,
  input  [2:0]  exeReq_5_bits_index,
  input         exeReq_5_bits_ffo,
                exeReq_6_valid,
  input  [31:0] exeReq_6_bits_source1,
                exeReq_6_bits_source2,
  input  [2:0]  exeReq_6_bits_index,
  input         exeReq_6_bits_ffo,
                exeReq_7_valid,
  input  [31:0] exeReq_7_bits_source1,
                exeReq_7_bits_source2,
  input  [2:0]  exeReq_7_bits_index,
  input         exeReq_7_bits_ffo,
                exeReq_8_valid,
  input  [31:0] exeReq_8_bits_source1,
                exeReq_8_bits_source2,
  input  [2:0]  exeReq_8_bits_index,
  input         exeReq_8_bits_ffo,
                exeReq_9_valid,
  input  [31:0] exeReq_9_bits_source1,
                exeReq_9_bits_source2,
  input  [2:0]  exeReq_9_bits_index,
  input         exeReq_9_bits_ffo,
                exeReq_10_valid,
  input  [31:0] exeReq_10_bits_source1,
                exeReq_10_bits_source2,
  input  [2:0]  exeReq_10_bits_index,
  input         exeReq_10_bits_ffo,
                exeReq_11_valid,
  input  [31:0] exeReq_11_bits_source1,
                exeReq_11_bits_source2,
  input  [2:0]  exeReq_11_bits_index,
  input         exeReq_11_bits_ffo,
                exeReq_12_valid,
  input  [31:0] exeReq_12_bits_source1,
                exeReq_12_bits_source2,
  input  [2:0]  exeReq_12_bits_index,
  input         exeReq_12_bits_ffo,
                exeReq_13_valid,
  input  [31:0] exeReq_13_bits_source1,
                exeReq_13_bits_source2,
  input  [2:0]  exeReq_13_bits_index,
  input         exeReq_13_bits_ffo,
                exeReq_14_valid,
  input  [31:0] exeReq_14_bits_source1,
                exeReq_14_bits_source2,
  input  [2:0]  exeReq_14_bits_index,
  input         exeReq_14_bits_ffo,
                exeReq_15_valid,
  input  [31:0] exeReq_15_bits_source1,
                exeReq_15_bits_source2,
  input  [2:0]  exeReq_15_bits_index,
  input         exeReq_15_bits_ffo,
                exeReq_16_valid,
  input  [31:0] exeReq_16_bits_source1,
                exeReq_16_bits_source2,
  input  [2:0]  exeReq_16_bits_index,
  input         exeReq_16_bits_ffo,
                exeReq_17_valid,
  input  [31:0] exeReq_17_bits_source1,
                exeReq_17_bits_source2,
  input  [2:0]  exeReq_17_bits_index,
  input         exeReq_17_bits_ffo,
                exeReq_18_valid,
  input  [31:0] exeReq_18_bits_source1,
                exeReq_18_bits_source2,
  input  [2:0]  exeReq_18_bits_index,
  input         exeReq_18_bits_ffo,
                exeReq_19_valid,
  input  [31:0] exeReq_19_bits_source1,
                exeReq_19_bits_source2,
  input  [2:0]  exeReq_19_bits_index,
  input         exeReq_19_bits_ffo,
                exeReq_20_valid,
  input  [31:0] exeReq_20_bits_source1,
                exeReq_20_bits_source2,
  input  [2:0]  exeReq_20_bits_index,
  input         exeReq_20_bits_ffo,
                exeReq_21_valid,
  input  [31:0] exeReq_21_bits_source1,
                exeReq_21_bits_source2,
  input  [2:0]  exeReq_21_bits_index,
  input         exeReq_21_bits_ffo,
                exeReq_22_valid,
  input  [31:0] exeReq_22_bits_source1,
                exeReq_22_bits_source2,
  input  [2:0]  exeReq_22_bits_index,
  input         exeReq_22_bits_ffo,
                exeReq_23_valid,
  input  [31:0] exeReq_23_bits_source1,
                exeReq_23_bits_source2,
  input  [2:0]  exeReq_23_bits_index,
  input         exeReq_23_bits_ffo,
                exeReq_24_valid,
  input  [31:0] exeReq_24_bits_source1,
                exeReq_24_bits_source2,
  input  [2:0]  exeReq_24_bits_index,
  input         exeReq_24_bits_ffo,
                exeReq_25_valid,
  input  [31:0] exeReq_25_bits_source1,
                exeReq_25_bits_source2,
  input  [2:0]  exeReq_25_bits_index,
  input         exeReq_25_bits_ffo,
                exeReq_26_valid,
  input  [31:0] exeReq_26_bits_source1,
                exeReq_26_bits_source2,
  input  [2:0]  exeReq_26_bits_index,
  input         exeReq_26_bits_ffo,
                exeReq_27_valid,
  input  [31:0] exeReq_27_bits_source1,
                exeReq_27_bits_source2,
  input  [2:0]  exeReq_27_bits_index,
  input         exeReq_27_bits_ffo,
                exeReq_28_valid,
  input  [31:0] exeReq_28_bits_source1,
                exeReq_28_bits_source2,
  input  [2:0]  exeReq_28_bits_index,
  input         exeReq_28_bits_ffo,
                exeReq_29_valid,
  input  [31:0] exeReq_29_bits_source1,
                exeReq_29_bits_source2,
  input  [2:0]  exeReq_29_bits_index,
  input         exeReq_29_bits_ffo,
                exeReq_30_valid,
  input  [31:0] exeReq_30_bits_source1,
                exeReq_30_bits_source2,
  input  [2:0]  exeReq_30_bits_index,
  input         exeReq_30_bits_ffo,
                exeReq_31_valid,
  input  [31:0] exeReq_31_bits_source1,
                exeReq_31_bits_source2,
  input  [2:0]  exeReq_31_bits_index,
  input         exeReq_31_bits_ffo,
                exeResp_0_ready,
  output        exeResp_0_valid,
  output [4:0]  exeResp_0_bits_vd,
  output        exeResp_0_bits_offset,
  output [3:0]  exeResp_0_bits_mask,
  output [31:0] exeResp_0_bits_data,
  output [2:0]  exeResp_0_bits_instructionIndex,
  input         exeResp_1_ready,
  output        exeResp_1_valid,
  output [4:0]  exeResp_1_bits_vd,
  output        exeResp_1_bits_offset,
  output [3:0]  exeResp_1_bits_mask,
  output [31:0] exeResp_1_bits_data,
  output [2:0]  exeResp_1_bits_instructionIndex,
  input         exeResp_2_ready,
  output        exeResp_2_valid,
  output [4:0]  exeResp_2_bits_vd,
  output        exeResp_2_bits_offset,
  output [3:0]  exeResp_2_bits_mask,
  output [31:0] exeResp_2_bits_data,
  output [2:0]  exeResp_2_bits_instructionIndex,
  input         exeResp_3_ready,
  output        exeResp_3_valid,
  output [4:0]  exeResp_3_bits_vd,
  output        exeResp_3_bits_offset,
  output [3:0]  exeResp_3_bits_mask,
  output [31:0] exeResp_3_bits_data,
  output [2:0]  exeResp_3_bits_instructionIndex,
  input         exeResp_4_ready,
  output        exeResp_4_valid,
  output [4:0]  exeResp_4_bits_vd,
  output        exeResp_4_bits_offset,
  output [3:0]  exeResp_4_bits_mask,
  output [31:0] exeResp_4_bits_data,
  output [2:0]  exeResp_4_bits_instructionIndex,
  input         exeResp_5_ready,
  output        exeResp_5_valid,
  output [4:0]  exeResp_5_bits_vd,
  output        exeResp_5_bits_offset,
  output [3:0]  exeResp_5_bits_mask,
  output [31:0] exeResp_5_bits_data,
  output [2:0]  exeResp_5_bits_instructionIndex,
  input         exeResp_6_ready,
  output        exeResp_6_valid,
  output [4:0]  exeResp_6_bits_vd,
  output        exeResp_6_bits_offset,
  output [3:0]  exeResp_6_bits_mask,
  output [31:0] exeResp_6_bits_data,
  output [2:0]  exeResp_6_bits_instructionIndex,
  input         exeResp_7_ready,
  output        exeResp_7_valid,
  output [4:0]  exeResp_7_bits_vd,
  output        exeResp_7_bits_offset,
  output [3:0]  exeResp_7_bits_mask,
  output [31:0] exeResp_7_bits_data,
  output [2:0]  exeResp_7_bits_instructionIndex,
  input         exeResp_8_ready,
  output        exeResp_8_valid,
  output [4:0]  exeResp_8_bits_vd,
  output        exeResp_8_bits_offset,
  output [3:0]  exeResp_8_bits_mask,
  output [31:0] exeResp_8_bits_data,
  output [2:0]  exeResp_8_bits_instructionIndex,
  input         exeResp_9_ready,
  output        exeResp_9_valid,
  output [4:0]  exeResp_9_bits_vd,
  output        exeResp_9_bits_offset,
  output [3:0]  exeResp_9_bits_mask,
  output [31:0] exeResp_9_bits_data,
  output [2:0]  exeResp_9_bits_instructionIndex,
  input         exeResp_10_ready,
  output        exeResp_10_valid,
  output [4:0]  exeResp_10_bits_vd,
  output        exeResp_10_bits_offset,
  output [3:0]  exeResp_10_bits_mask,
  output [31:0] exeResp_10_bits_data,
  output [2:0]  exeResp_10_bits_instructionIndex,
  input         exeResp_11_ready,
  output        exeResp_11_valid,
  output [4:0]  exeResp_11_bits_vd,
  output        exeResp_11_bits_offset,
  output [3:0]  exeResp_11_bits_mask,
  output [31:0] exeResp_11_bits_data,
  output [2:0]  exeResp_11_bits_instructionIndex,
  input         exeResp_12_ready,
  output        exeResp_12_valid,
  output [4:0]  exeResp_12_bits_vd,
  output        exeResp_12_bits_offset,
  output [3:0]  exeResp_12_bits_mask,
  output [31:0] exeResp_12_bits_data,
  output [2:0]  exeResp_12_bits_instructionIndex,
  input         exeResp_13_ready,
  output        exeResp_13_valid,
  output [4:0]  exeResp_13_bits_vd,
  output        exeResp_13_bits_offset,
  output [3:0]  exeResp_13_bits_mask,
  output [31:0] exeResp_13_bits_data,
  output [2:0]  exeResp_13_bits_instructionIndex,
  input         exeResp_14_ready,
  output        exeResp_14_valid,
  output [4:0]  exeResp_14_bits_vd,
  output        exeResp_14_bits_offset,
  output [3:0]  exeResp_14_bits_mask,
  output [31:0] exeResp_14_bits_data,
  output [2:0]  exeResp_14_bits_instructionIndex,
  input         exeResp_15_ready,
  output        exeResp_15_valid,
  output [4:0]  exeResp_15_bits_vd,
  output        exeResp_15_bits_offset,
  output [3:0]  exeResp_15_bits_mask,
  output [31:0] exeResp_15_bits_data,
  output [2:0]  exeResp_15_bits_instructionIndex,
  input         exeResp_16_ready,
  output        exeResp_16_valid,
  output [4:0]  exeResp_16_bits_vd,
  output        exeResp_16_bits_offset,
  output [3:0]  exeResp_16_bits_mask,
  output [31:0] exeResp_16_bits_data,
  output [2:0]  exeResp_16_bits_instructionIndex,
  input         exeResp_17_ready,
  output        exeResp_17_valid,
  output [4:0]  exeResp_17_bits_vd,
  output        exeResp_17_bits_offset,
  output [3:0]  exeResp_17_bits_mask,
  output [31:0] exeResp_17_bits_data,
  output [2:0]  exeResp_17_bits_instructionIndex,
  input         exeResp_18_ready,
  output        exeResp_18_valid,
  output [4:0]  exeResp_18_bits_vd,
  output        exeResp_18_bits_offset,
  output [3:0]  exeResp_18_bits_mask,
  output [31:0] exeResp_18_bits_data,
  output [2:0]  exeResp_18_bits_instructionIndex,
  input         exeResp_19_ready,
  output        exeResp_19_valid,
  output [4:0]  exeResp_19_bits_vd,
  output        exeResp_19_bits_offset,
  output [3:0]  exeResp_19_bits_mask,
  output [31:0] exeResp_19_bits_data,
  output [2:0]  exeResp_19_bits_instructionIndex,
  input         exeResp_20_ready,
  output        exeResp_20_valid,
  output [4:0]  exeResp_20_bits_vd,
  output        exeResp_20_bits_offset,
  output [3:0]  exeResp_20_bits_mask,
  output [31:0] exeResp_20_bits_data,
  output [2:0]  exeResp_20_bits_instructionIndex,
  input         exeResp_21_ready,
  output        exeResp_21_valid,
  output [4:0]  exeResp_21_bits_vd,
  output        exeResp_21_bits_offset,
  output [3:0]  exeResp_21_bits_mask,
  output [31:0] exeResp_21_bits_data,
  output [2:0]  exeResp_21_bits_instructionIndex,
  input         exeResp_22_ready,
  output        exeResp_22_valid,
  output [4:0]  exeResp_22_bits_vd,
  output        exeResp_22_bits_offset,
  output [3:0]  exeResp_22_bits_mask,
  output [31:0] exeResp_22_bits_data,
  output [2:0]  exeResp_22_bits_instructionIndex,
  input         exeResp_23_ready,
  output        exeResp_23_valid,
  output [4:0]  exeResp_23_bits_vd,
  output        exeResp_23_bits_offset,
  output [3:0]  exeResp_23_bits_mask,
  output [31:0] exeResp_23_bits_data,
  output [2:0]  exeResp_23_bits_instructionIndex,
  input         exeResp_24_ready,
  output        exeResp_24_valid,
  output [4:0]  exeResp_24_bits_vd,
  output        exeResp_24_bits_offset,
  output [3:0]  exeResp_24_bits_mask,
  output [31:0] exeResp_24_bits_data,
  output [2:0]  exeResp_24_bits_instructionIndex,
  input         exeResp_25_ready,
  output        exeResp_25_valid,
  output [4:0]  exeResp_25_bits_vd,
  output        exeResp_25_bits_offset,
  output [3:0]  exeResp_25_bits_mask,
  output [31:0] exeResp_25_bits_data,
  output [2:0]  exeResp_25_bits_instructionIndex,
  input         exeResp_26_ready,
  output        exeResp_26_valid,
  output [4:0]  exeResp_26_bits_vd,
  output        exeResp_26_bits_offset,
  output [3:0]  exeResp_26_bits_mask,
  output [31:0] exeResp_26_bits_data,
  output [2:0]  exeResp_26_bits_instructionIndex,
  input         exeResp_27_ready,
  output        exeResp_27_valid,
  output [4:0]  exeResp_27_bits_vd,
  output        exeResp_27_bits_offset,
  output [3:0]  exeResp_27_bits_mask,
  output [31:0] exeResp_27_bits_data,
  output [2:0]  exeResp_27_bits_instructionIndex,
  input         exeResp_28_ready,
  output        exeResp_28_valid,
  output [4:0]  exeResp_28_bits_vd,
  output        exeResp_28_bits_offset,
  output [3:0]  exeResp_28_bits_mask,
  output [31:0] exeResp_28_bits_data,
  output [2:0]  exeResp_28_bits_instructionIndex,
  input         exeResp_29_ready,
  output        exeResp_29_valid,
  output [4:0]  exeResp_29_bits_vd,
  output        exeResp_29_bits_offset,
  output [3:0]  exeResp_29_bits_mask,
  output [31:0] exeResp_29_bits_data,
  output [2:0]  exeResp_29_bits_instructionIndex,
  input         exeResp_30_ready,
  output        exeResp_30_valid,
  output [4:0]  exeResp_30_bits_vd,
  output        exeResp_30_bits_offset,
  output [3:0]  exeResp_30_bits_mask,
  output [31:0] exeResp_30_bits_data,
  output [2:0]  exeResp_30_bits_instructionIndex,
  input         exeResp_31_ready,
  output        exeResp_31_valid,
  output [4:0]  exeResp_31_bits_vd,
  output        exeResp_31_bits_offset,
  output [3:0]  exeResp_31_bits_mask,
  output [31:0] exeResp_31_bits_data,
  output [2:0]  exeResp_31_bits_instructionIndex,
  input         writeRelease_0,
                writeRelease_1,
                writeRelease_2,
                writeRelease_3,
                writeRelease_4,
                writeRelease_5,
                writeRelease_6,
                writeRelease_7,
                writeRelease_8,
                writeRelease_9,
                writeRelease_10,
                writeRelease_11,
                writeRelease_12,
                writeRelease_13,
                writeRelease_14,
                writeRelease_15,
                writeRelease_16,
                writeRelease_17,
                writeRelease_18,
                writeRelease_19,
                writeRelease_20,
                writeRelease_21,
                writeRelease_22,
                writeRelease_23,
                writeRelease_24,
                writeRelease_25,
                writeRelease_26,
                writeRelease_27,
                writeRelease_28,
                writeRelease_29,
                writeRelease_30,
                writeRelease_31,
  output        tokenIO_0_maskRequestRelease,
                tokenIO_1_maskRequestRelease,
                tokenIO_2_maskRequestRelease,
                tokenIO_3_maskRequestRelease,
                tokenIO_4_maskRequestRelease,
                tokenIO_5_maskRequestRelease,
                tokenIO_6_maskRequestRelease,
                tokenIO_7_maskRequestRelease,
                tokenIO_8_maskRequestRelease,
                tokenIO_9_maskRequestRelease,
                tokenIO_10_maskRequestRelease,
                tokenIO_11_maskRequestRelease,
                tokenIO_12_maskRequestRelease,
                tokenIO_13_maskRequestRelease,
                tokenIO_14_maskRequestRelease,
                tokenIO_15_maskRequestRelease,
                tokenIO_16_maskRequestRelease,
                tokenIO_17_maskRequestRelease,
                tokenIO_18_maskRequestRelease,
                tokenIO_19_maskRequestRelease,
                tokenIO_20_maskRequestRelease,
                tokenIO_21_maskRequestRelease,
                tokenIO_22_maskRequestRelease,
                tokenIO_23_maskRequestRelease,
                tokenIO_24_maskRequestRelease,
                tokenIO_25_maskRequestRelease,
                tokenIO_26_maskRequestRelease,
                tokenIO_27_maskRequestRelease,
                tokenIO_28_maskRequestRelease,
                tokenIO_29_maskRequestRelease,
                tokenIO_30_maskRequestRelease,
                tokenIO_31_maskRequestRelease,
  input         readChannel_0_ready,
  output        readChannel_0_valid,
  output [4:0]  readChannel_0_bits_vs,
  output        readChannel_0_bits_offset,
  output [2:0]  readChannel_0_bits_instructionIndex,
  input         readChannel_1_ready,
  output        readChannel_1_valid,
  output [4:0]  readChannel_1_bits_vs,
  output        readChannel_1_bits_offset,
  output [2:0]  readChannel_1_bits_instructionIndex,
  input         readChannel_2_ready,
  output        readChannel_2_valid,
  output [4:0]  readChannel_2_bits_vs,
  output        readChannel_2_bits_offset,
  output [2:0]  readChannel_2_bits_instructionIndex,
  input         readChannel_3_ready,
  output        readChannel_3_valid,
  output [4:0]  readChannel_3_bits_vs,
  output        readChannel_3_bits_offset,
  output [2:0]  readChannel_3_bits_instructionIndex,
  input         readChannel_4_ready,
  output        readChannel_4_valid,
  output [4:0]  readChannel_4_bits_vs,
  output        readChannel_4_bits_offset,
  output [2:0]  readChannel_4_bits_instructionIndex,
  input         readChannel_5_ready,
  output        readChannel_5_valid,
  output [4:0]  readChannel_5_bits_vs,
  output        readChannel_5_bits_offset,
  output [2:0]  readChannel_5_bits_instructionIndex,
  input         readChannel_6_ready,
  output        readChannel_6_valid,
  output [4:0]  readChannel_6_bits_vs,
  output        readChannel_6_bits_offset,
  output [2:0]  readChannel_6_bits_instructionIndex,
  input         readChannel_7_ready,
  output        readChannel_7_valid,
  output [4:0]  readChannel_7_bits_vs,
  output        readChannel_7_bits_offset,
  output [2:0]  readChannel_7_bits_instructionIndex,
  input         readChannel_8_ready,
  output        readChannel_8_valid,
  output [4:0]  readChannel_8_bits_vs,
  output        readChannel_8_bits_offset,
  output [2:0]  readChannel_8_bits_instructionIndex,
  input         readChannel_9_ready,
  output        readChannel_9_valid,
  output [4:0]  readChannel_9_bits_vs,
  output        readChannel_9_bits_offset,
  output [2:0]  readChannel_9_bits_instructionIndex,
  input         readChannel_10_ready,
  output        readChannel_10_valid,
  output [4:0]  readChannel_10_bits_vs,
  output        readChannel_10_bits_offset,
  output [2:0]  readChannel_10_bits_instructionIndex,
  input         readChannel_11_ready,
  output        readChannel_11_valid,
  output [4:0]  readChannel_11_bits_vs,
  output        readChannel_11_bits_offset,
  output [2:0]  readChannel_11_bits_instructionIndex,
  input         readChannel_12_ready,
  output        readChannel_12_valid,
  output [4:0]  readChannel_12_bits_vs,
  output        readChannel_12_bits_offset,
  output [2:0]  readChannel_12_bits_instructionIndex,
  input         readChannel_13_ready,
  output        readChannel_13_valid,
  output [4:0]  readChannel_13_bits_vs,
  output        readChannel_13_bits_offset,
  output [2:0]  readChannel_13_bits_instructionIndex,
  input         readChannel_14_ready,
  output        readChannel_14_valid,
  output [4:0]  readChannel_14_bits_vs,
  output        readChannel_14_bits_offset,
  output [2:0]  readChannel_14_bits_instructionIndex,
  input         readChannel_15_ready,
  output        readChannel_15_valid,
  output [4:0]  readChannel_15_bits_vs,
  output        readChannel_15_bits_offset,
  output [2:0]  readChannel_15_bits_instructionIndex,
  input         readChannel_16_ready,
  output        readChannel_16_valid,
  output [4:0]  readChannel_16_bits_vs,
  output        readChannel_16_bits_offset,
  output [2:0]  readChannel_16_bits_instructionIndex,
  input         readChannel_17_ready,
  output        readChannel_17_valid,
  output [4:0]  readChannel_17_bits_vs,
  output        readChannel_17_bits_offset,
  output [2:0]  readChannel_17_bits_instructionIndex,
  input         readChannel_18_ready,
  output        readChannel_18_valid,
  output [4:0]  readChannel_18_bits_vs,
  output        readChannel_18_bits_offset,
  output [2:0]  readChannel_18_bits_instructionIndex,
  input         readChannel_19_ready,
  output        readChannel_19_valid,
  output [4:0]  readChannel_19_bits_vs,
  output        readChannel_19_bits_offset,
  output [2:0]  readChannel_19_bits_instructionIndex,
  input         readChannel_20_ready,
  output        readChannel_20_valid,
  output [4:0]  readChannel_20_bits_vs,
  output        readChannel_20_bits_offset,
  output [2:0]  readChannel_20_bits_instructionIndex,
  input         readChannel_21_ready,
  output        readChannel_21_valid,
  output [4:0]  readChannel_21_bits_vs,
  output        readChannel_21_bits_offset,
  output [2:0]  readChannel_21_bits_instructionIndex,
  input         readChannel_22_ready,
  output        readChannel_22_valid,
  output [4:0]  readChannel_22_bits_vs,
  output        readChannel_22_bits_offset,
  output [2:0]  readChannel_22_bits_instructionIndex,
  input         readChannel_23_ready,
  output        readChannel_23_valid,
  output [4:0]  readChannel_23_bits_vs,
  output        readChannel_23_bits_offset,
  output [2:0]  readChannel_23_bits_instructionIndex,
  input         readChannel_24_ready,
  output        readChannel_24_valid,
  output [4:0]  readChannel_24_bits_vs,
  output        readChannel_24_bits_offset,
  output [2:0]  readChannel_24_bits_instructionIndex,
  input         readChannel_25_ready,
  output        readChannel_25_valid,
  output [4:0]  readChannel_25_bits_vs,
  output        readChannel_25_bits_offset,
  output [2:0]  readChannel_25_bits_instructionIndex,
  input         readChannel_26_ready,
  output        readChannel_26_valid,
  output [4:0]  readChannel_26_bits_vs,
  output        readChannel_26_bits_offset,
  output [2:0]  readChannel_26_bits_instructionIndex,
  input         readChannel_27_ready,
  output        readChannel_27_valid,
  output [4:0]  readChannel_27_bits_vs,
  output        readChannel_27_bits_offset,
  output [2:0]  readChannel_27_bits_instructionIndex,
  input         readChannel_28_ready,
  output        readChannel_28_valid,
  output [4:0]  readChannel_28_bits_vs,
  output        readChannel_28_bits_offset,
  output [2:0]  readChannel_28_bits_instructionIndex,
  input         readChannel_29_ready,
  output        readChannel_29_valid,
  output [4:0]  readChannel_29_bits_vs,
  output        readChannel_29_bits_offset,
  output [2:0]  readChannel_29_bits_instructionIndex,
  input         readChannel_30_ready,
  output        readChannel_30_valid,
  output [4:0]  readChannel_30_bits_vs,
  output        readChannel_30_bits_offset,
  output [2:0]  readChannel_30_bits_instructionIndex,
  input         readChannel_31_ready,
  output        readChannel_31_valid,
  output [4:0]  readChannel_31_bits_vs,
  output        readChannel_31_bits_offset,
  output [2:0]  readChannel_31_bits_instructionIndex,
  input         readResult_0_valid,
  input  [31:0] readResult_0_bits,
  input         readResult_1_valid,
  input  [31:0] readResult_1_bits,
  input         readResult_2_valid,
  input  [31:0] readResult_2_bits,
  input         readResult_3_valid,
  input  [31:0] readResult_3_bits,
  input         readResult_4_valid,
  input  [31:0] readResult_4_bits,
  input         readResult_5_valid,
  input  [31:0] readResult_5_bits,
  input         readResult_6_valid,
  input  [31:0] readResult_6_bits,
  input         readResult_7_valid,
  input  [31:0] readResult_7_bits,
  input         readResult_8_valid,
  input  [31:0] readResult_8_bits,
  input         readResult_9_valid,
  input  [31:0] readResult_9_bits,
  input         readResult_10_valid,
  input  [31:0] readResult_10_bits,
  input         readResult_11_valid,
  input  [31:0] readResult_11_bits,
  input         readResult_12_valid,
  input  [31:0] readResult_12_bits,
  input         readResult_13_valid,
  input  [31:0] readResult_13_bits,
  input         readResult_14_valid,
  input  [31:0] readResult_14_bits,
  input         readResult_15_valid,
  input  [31:0] readResult_15_bits,
  input         readResult_16_valid,
  input  [31:0] readResult_16_bits,
  input         readResult_17_valid,
  input  [31:0] readResult_17_bits,
  input         readResult_18_valid,
  input  [31:0] readResult_18_bits,
  input         readResult_19_valid,
  input  [31:0] readResult_19_bits,
  input         readResult_20_valid,
  input  [31:0] readResult_20_bits,
  input         readResult_21_valid,
  input  [31:0] readResult_21_bits,
  input         readResult_22_valid,
  input  [31:0] readResult_22_bits,
  input         readResult_23_valid,
  input  [31:0] readResult_23_bits,
  input         readResult_24_valid,
  input  [31:0] readResult_24_bits,
  input         readResult_25_valid,
  input  [31:0] readResult_25_bits,
  input         readResult_26_valid,
  input  [31:0] readResult_26_bits,
  input         readResult_27_valid,
  input  [31:0] readResult_27_bits,
  input         readResult_28_valid,
  input  [31:0] readResult_28_bits,
  input         readResult_29_valid,
  input  [31:0] readResult_29_bits,
  input         readResult_30_valid,
  input  [31:0] readResult_30_bits,
  input         readResult_31_valid,
  input  [31:0] readResult_31_bits,
  output [7:0]  lastReport,
  output [31:0] laneMaskInput_0,
                laneMaskInput_1,
                laneMaskInput_2,
                laneMaskInput_3,
                laneMaskInput_4,
                laneMaskInput_5,
                laneMaskInput_6,
                laneMaskInput_7,
                laneMaskInput_8,
                laneMaskInput_9,
                laneMaskInput_10,
                laneMaskInput_11,
                laneMaskInput_12,
                laneMaskInput_13,
                laneMaskInput_14,
                laneMaskInput_15,
                laneMaskInput_16,
                laneMaskInput_17,
                laneMaskInput_18,
                laneMaskInput_19,
                laneMaskInput_20,
                laneMaskInput_21,
                laneMaskInput_22,
                laneMaskInput_23,
                laneMaskInput_24,
                laneMaskInput_25,
                laneMaskInput_26,
                laneMaskInput_27,
                laneMaskInput_28,
                laneMaskInput_29,
                laneMaskInput_30,
                laneMaskInput_31,
  input  [5:0]  laneMaskSelect_0,
                laneMaskSelect_1,
                laneMaskSelect_2,
                laneMaskSelect_3,
                laneMaskSelect_4,
                laneMaskSelect_5,
                laneMaskSelect_6,
                laneMaskSelect_7,
                laneMaskSelect_8,
                laneMaskSelect_9,
                laneMaskSelect_10,
                laneMaskSelect_11,
                laneMaskSelect_12,
                laneMaskSelect_13,
                laneMaskSelect_14,
                laneMaskSelect_15,
                laneMaskSelect_16,
                laneMaskSelect_17,
                laneMaskSelect_18,
                laneMaskSelect_19,
                laneMaskSelect_20,
                laneMaskSelect_21,
                laneMaskSelect_22,
                laneMaskSelect_23,
                laneMaskSelect_24,
                laneMaskSelect_25,
                laneMaskSelect_26,
                laneMaskSelect_27,
                laneMaskSelect_28,
                laneMaskSelect_29,
                laneMaskSelect_30,
                laneMaskSelect_31,
  input  [1:0]  laneMaskSewSelect_0,
                laneMaskSewSelect_1,
                laneMaskSewSelect_2,
                laneMaskSewSelect_3,
                laneMaskSewSelect_4,
                laneMaskSewSelect_5,
                laneMaskSewSelect_6,
                laneMaskSewSelect_7,
                laneMaskSewSelect_8,
                laneMaskSewSelect_9,
                laneMaskSewSelect_10,
                laneMaskSewSelect_11,
                laneMaskSewSelect_12,
                laneMaskSewSelect_13,
                laneMaskSewSelect_14,
                laneMaskSewSelect_15,
                laneMaskSewSelect_16,
                laneMaskSewSelect_17,
                laneMaskSewSelect_18,
                laneMaskSewSelect_19,
                laneMaskSewSelect_20,
                laneMaskSewSelect_21,
                laneMaskSewSelect_22,
                laneMaskSewSelect_23,
                laneMaskSewSelect_24,
                laneMaskSewSelect_25,
                laneMaskSewSelect_26,
                laneMaskSewSelect_27,
                laneMaskSewSelect_28,
                laneMaskSewSelect_29,
                laneMaskSewSelect_30,
                laneMaskSewSelect_31,
  input         v0UpdateVec_0_valid,
  input  [31:0] v0UpdateVec_0_bits_data,
  input         v0UpdateVec_0_bits_offset,
  input  [3:0]  v0UpdateVec_0_bits_mask,
  input         v0UpdateVec_1_valid,
  input  [31:0] v0UpdateVec_1_bits_data,
  input         v0UpdateVec_1_bits_offset,
  input  [3:0]  v0UpdateVec_1_bits_mask,
  input         v0UpdateVec_2_valid,
  input  [31:0] v0UpdateVec_2_bits_data,
  input         v0UpdateVec_2_bits_offset,
  input  [3:0]  v0UpdateVec_2_bits_mask,
  input         v0UpdateVec_3_valid,
  input  [31:0] v0UpdateVec_3_bits_data,
  input         v0UpdateVec_3_bits_offset,
  input  [3:0]  v0UpdateVec_3_bits_mask,
  input         v0UpdateVec_4_valid,
  input  [31:0] v0UpdateVec_4_bits_data,
  input         v0UpdateVec_4_bits_offset,
  input  [3:0]  v0UpdateVec_4_bits_mask,
  input         v0UpdateVec_5_valid,
  input  [31:0] v0UpdateVec_5_bits_data,
  input         v0UpdateVec_5_bits_offset,
  input  [3:0]  v0UpdateVec_5_bits_mask,
  input         v0UpdateVec_6_valid,
  input  [31:0] v0UpdateVec_6_bits_data,
  input         v0UpdateVec_6_bits_offset,
  input  [3:0]  v0UpdateVec_6_bits_mask,
  input         v0UpdateVec_7_valid,
  input  [31:0] v0UpdateVec_7_bits_data,
  input         v0UpdateVec_7_bits_offset,
  input  [3:0]  v0UpdateVec_7_bits_mask,
  input         v0UpdateVec_8_valid,
  input  [31:0] v0UpdateVec_8_bits_data,
  input         v0UpdateVec_8_bits_offset,
  input  [3:0]  v0UpdateVec_8_bits_mask,
  input         v0UpdateVec_9_valid,
  input  [31:0] v0UpdateVec_9_bits_data,
  input         v0UpdateVec_9_bits_offset,
  input  [3:0]  v0UpdateVec_9_bits_mask,
  input         v0UpdateVec_10_valid,
  input  [31:0] v0UpdateVec_10_bits_data,
  input         v0UpdateVec_10_bits_offset,
  input  [3:0]  v0UpdateVec_10_bits_mask,
  input         v0UpdateVec_11_valid,
  input  [31:0] v0UpdateVec_11_bits_data,
  input         v0UpdateVec_11_bits_offset,
  input  [3:0]  v0UpdateVec_11_bits_mask,
  input         v0UpdateVec_12_valid,
  input  [31:0] v0UpdateVec_12_bits_data,
  input         v0UpdateVec_12_bits_offset,
  input  [3:0]  v0UpdateVec_12_bits_mask,
  input         v0UpdateVec_13_valid,
  input  [31:0] v0UpdateVec_13_bits_data,
  input         v0UpdateVec_13_bits_offset,
  input  [3:0]  v0UpdateVec_13_bits_mask,
  input         v0UpdateVec_14_valid,
  input  [31:0] v0UpdateVec_14_bits_data,
  input         v0UpdateVec_14_bits_offset,
  input  [3:0]  v0UpdateVec_14_bits_mask,
  input         v0UpdateVec_15_valid,
  input  [31:0] v0UpdateVec_15_bits_data,
  input         v0UpdateVec_15_bits_offset,
  input  [3:0]  v0UpdateVec_15_bits_mask,
  input         v0UpdateVec_16_valid,
  input  [31:0] v0UpdateVec_16_bits_data,
  input         v0UpdateVec_16_bits_offset,
  input  [3:0]  v0UpdateVec_16_bits_mask,
  input         v0UpdateVec_17_valid,
  input  [31:0] v0UpdateVec_17_bits_data,
  input         v0UpdateVec_17_bits_offset,
  input  [3:0]  v0UpdateVec_17_bits_mask,
  input         v0UpdateVec_18_valid,
  input  [31:0] v0UpdateVec_18_bits_data,
  input         v0UpdateVec_18_bits_offset,
  input  [3:0]  v0UpdateVec_18_bits_mask,
  input         v0UpdateVec_19_valid,
  input  [31:0] v0UpdateVec_19_bits_data,
  input         v0UpdateVec_19_bits_offset,
  input  [3:0]  v0UpdateVec_19_bits_mask,
  input         v0UpdateVec_20_valid,
  input  [31:0] v0UpdateVec_20_bits_data,
  input         v0UpdateVec_20_bits_offset,
  input  [3:0]  v0UpdateVec_20_bits_mask,
  input         v0UpdateVec_21_valid,
  input  [31:0] v0UpdateVec_21_bits_data,
  input         v0UpdateVec_21_bits_offset,
  input  [3:0]  v0UpdateVec_21_bits_mask,
  input         v0UpdateVec_22_valid,
  input  [31:0] v0UpdateVec_22_bits_data,
  input         v0UpdateVec_22_bits_offset,
  input  [3:0]  v0UpdateVec_22_bits_mask,
  input         v0UpdateVec_23_valid,
  input  [31:0] v0UpdateVec_23_bits_data,
  input         v0UpdateVec_23_bits_offset,
  input  [3:0]  v0UpdateVec_23_bits_mask,
  input         v0UpdateVec_24_valid,
  input  [31:0] v0UpdateVec_24_bits_data,
  input         v0UpdateVec_24_bits_offset,
  input  [3:0]  v0UpdateVec_24_bits_mask,
  input         v0UpdateVec_25_valid,
  input  [31:0] v0UpdateVec_25_bits_data,
  input         v0UpdateVec_25_bits_offset,
  input  [3:0]  v0UpdateVec_25_bits_mask,
  input         v0UpdateVec_26_valid,
  input  [31:0] v0UpdateVec_26_bits_data,
  input         v0UpdateVec_26_bits_offset,
  input  [3:0]  v0UpdateVec_26_bits_mask,
  input         v0UpdateVec_27_valid,
  input  [31:0] v0UpdateVec_27_bits_data,
  input         v0UpdateVec_27_bits_offset,
  input  [3:0]  v0UpdateVec_27_bits_mask,
  input         v0UpdateVec_28_valid,
  input  [31:0] v0UpdateVec_28_bits_data,
  input         v0UpdateVec_28_bits_offset,
  input  [3:0]  v0UpdateVec_28_bits_mask,
  input         v0UpdateVec_29_valid,
  input  [31:0] v0UpdateVec_29_bits_data,
  input         v0UpdateVec_29_bits_offset,
  input  [3:0]  v0UpdateVec_29_bits_mask,
  input         v0UpdateVec_30_valid,
  input  [31:0] v0UpdateVec_30_bits_data,
  input         v0UpdateVec_30_bits_offset,
  input  [3:0]  v0UpdateVec_30_bits_mask,
  input         v0UpdateVec_31_valid,
  input  [31:0] v0UpdateVec_31_bits_data,
  input         v0UpdateVec_31_bits_offset,
  input  [3:0]  v0UpdateVec_31_bits_mask,
  output [31:0] writeRDData,
  input         gatherData_ready,
  output        gatherData_valid,
  output [31:0] gatherData_bits,
  input         gatherRead
);

  wire               readCrossBar_input_31_valid;
  wire               readCrossBar_input_30_valid;
  wire               readCrossBar_input_29_valid;
  wire               readCrossBar_input_28_valid;
  wire               readCrossBar_input_27_valid;
  wire               readCrossBar_input_26_valid;
  wire               readCrossBar_input_25_valid;
  wire               readCrossBar_input_24_valid;
  wire               readCrossBar_input_23_valid;
  wire               readCrossBar_input_22_valid;
  wire               readCrossBar_input_21_valid;
  wire               readCrossBar_input_20_valid;
  wire               readCrossBar_input_19_valid;
  wire               readCrossBar_input_18_valid;
  wire               readCrossBar_input_17_valid;
  wire               readCrossBar_input_16_valid;
  wire               readCrossBar_input_15_valid;
  wire               readCrossBar_input_14_valid;
  wire               readCrossBar_input_13_valid;
  wire               readCrossBar_input_12_valid;
  wire               readCrossBar_input_11_valid;
  wire               readCrossBar_input_10_valid;
  wire               readCrossBar_input_9_valid;
  wire               readCrossBar_input_8_valid;
  wire               readCrossBar_input_7_valid;
  wire               readCrossBar_input_6_valid;
  wire               readCrossBar_input_5_valid;
  wire               readCrossBar_input_4_valid;
  wire               readCrossBar_input_3_valid;
  wire               readCrossBar_input_2_valid;
  wire               readCrossBar_input_1_valid;
  wire               readCrossBar_input_0_valid;
  wire               _writeQueue_fifo_31_empty;
  wire               _writeQueue_fifo_31_full;
  wire               _writeQueue_fifo_31_error;
  wire [49:0]        _writeQueue_fifo_31_data_out;
  wire               _writeQueue_fifo_30_empty;
  wire               _writeQueue_fifo_30_full;
  wire               _writeQueue_fifo_30_error;
  wire [49:0]        _writeQueue_fifo_30_data_out;
  wire               _writeQueue_fifo_29_empty;
  wire               _writeQueue_fifo_29_full;
  wire               _writeQueue_fifo_29_error;
  wire [49:0]        _writeQueue_fifo_29_data_out;
  wire               _writeQueue_fifo_28_empty;
  wire               _writeQueue_fifo_28_full;
  wire               _writeQueue_fifo_28_error;
  wire [49:0]        _writeQueue_fifo_28_data_out;
  wire               _writeQueue_fifo_27_empty;
  wire               _writeQueue_fifo_27_full;
  wire               _writeQueue_fifo_27_error;
  wire [49:0]        _writeQueue_fifo_27_data_out;
  wire               _writeQueue_fifo_26_empty;
  wire               _writeQueue_fifo_26_full;
  wire               _writeQueue_fifo_26_error;
  wire [49:0]        _writeQueue_fifo_26_data_out;
  wire               _writeQueue_fifo_25_empty;
  wire               _writeQueue_fifo_25_full;
  wire               _writeQueue_fifo_25_error;
  wire [49:0]        _writeQueue_fifo_25_data_out;
  wire               _writeQueue_fifo_24_empty;
  wire               _writeQueue_fifo_24_full;
  wire               _writeQueue_fifo_24_error;
  wire [49:0]        _writeQueue_fifo_24_data_out;
  wire               _writeQueue_fifo_23_empty;
  wire               _writeQueue_fifo_23_full;
  wire               _writeQueue_fifo_23_error;
  wire [49:0]        _writeQueue_fifo_23_data_out;
  wire               _writeQueue_fifo_22_empty;
  wire               _writeQueue_fifo_22_full;
  wire               _writeQueue_fifo_22_error;
  wire [49:0]        _writeQueue_fifo_22_data_out;
  wire               _writeQueue_fifo_21_empty;
  wire               _writeQueue_fifo_21_full;
  wire               _writeQueue_fifo_21_error;
  wire [49:0]        _writeQueue_fifo_21_data_out;
  wire               _writeQueue_fifo_20_empty;
  wire               _writeQueue_fifo_20_full;
  wire               _writeQueue_fifo_20_error;
  wire [49:0]        _writeQueue_fifo_20_data_out;
  wire               _writeQueue_fifo_19_empty;
  wire               _writeQueue_fifo_19_full;
  wire               _writeQueue_fifo_19_error;
  wire [49:0]        _writeQueue_fifo_19_data_out;
  wire               _writeQueue_fifo_18_empty;
  wire               _writeQueue_fifo_18_full;
  wire               _writeQueue_fifo_18_error;
  wire [49:0]        _writeQueue_fifo_18_data_out;
  wire               _writeQueue_fifo_17_empty;
  wire               _writeQueue_fifo_17_full;
  wire               _writeQueue_fifo_17_error;
  wire [49:0]        _writeQueue_fifo_17_data_out;
  wire               _writeQueue_fifo_16_empty;
  wire               _writeQueue_fifo_16_full;
  wire               _writeQueue_fifo_16_error;
  wire [49:0]        _writeQueue_fifo_16_data_out;
  wire               _writeQueue_fifo_15_empty;
  wire               _writeQueue_fifo_15_full;
  wire               _writeQueue_fifo_15_error;
  wire [49:0]        _writeQueue_fifo_15_data_out;
  wire               _writeQueue_fifo_14_empty;
  wire               _writeQueue_fifo_14_full;
  wire               _writeQueue_fifo_14_error;
  wire [49:0]        _writeQueue_fifo_14_data_out;
  wire               _writeQueue_fifo_13_empty;
  wire               _writeQueue_fifo_13_full;
  wire               _writeQueue_fifo_13_error;
  wire [49:0]        _writeQueue_fifo_13_data_out;
  wire               _writeQueue_fifo_12_empty;
  wire               _writeQueue_fifo_12_full;
  wire               _writeQueue_fifo_12_error;
  wire [49:0]        _writeQueue_fifo_12_data_out;
  wire               _writeQueue_fifo_11_empty;
  wire               _writeQueue_fifo_11_full;
  wire               _writeQueue_fifo_11_error;
  wire [49:0]        _writeQueue_fifo_11_data_out;
  wire               _writeQueue_fifo_10_empty;
  wire               _writeQueue_fifo_10_full;
  wire               _writeQueue_fifo_10_error;
  wire [49:0]        _writeQueue_fifo_10_data_out;
  wire               _writeQueue_fifo_9_empty;
  wire               _writeQueue_fifo_9_full;
  wire               _writeQueue_fifo_9_error;
  wire [49:0]        _writeQueue_fifo_9_data_out;
  wire               _writeQueue_fifo_8_empty;
  wire               _writeQueue_fifo_8_full;
  wire               _writeQueue_fifo_8_error;
  wire [49:0]        _writeQueue_fifo_8_data_out;
  wire               _writeQueue_fifo_7_empty;
  wire               _writeQueue_fifo_7_full;
  wire               _writeQueue_fifo_7_error;
  wire [49:0]        _writeQueue_fifo_7_data_out;
  wire               _writeQueue_fifo_6_empty;
  wire               _writeQueue_fifo_6_full;
  wire               _writeQueue_fifo_6_error;
  wire [49:0]        _writeQueue_fifo_6_data_out;
  wire               _writeQueue_fifo_5_empty;
  wire               _writeQueue_fifo_5_full;
  wire               _writeQueue_fifo_5_error;
  wire [49:0]        _writeQueue_fifo_5_data_out;
  wire               _writeQueue_fifo_4_empty;
  wire               _writeQueue_fifo_4_full;
  wire               _writeQueue_fifo_4_error;
  wire [49:0]        _writeQueue_fifo_4_data_out;
  wire               _writeQueue_fifo_3_empty;
  wire               _writeQueue_fifo_3_full;
  wire               _writeQueue_fifo_3_error;
  wire [49:0]        _writeQueue_fifo_3_data_out;
  wire               _writeQueue_fifo_2_empty;
  wire               _writeQueue_fifo_2_full;
  wire               _writeQueue_fifo_2_error;
  wire [49:0]        _writeQueue_fifo_2_data_out;
  wire               _writeQueue_fifo_1_empty;
  wire               _writeQueue_fifo_1_full;
  wire               _writeQueue_fifo_1_error;
  wire [49:0]        _writeQueue_fifo_1_data_out;
  wire               _writeQueue_fifo_empty;
  wire               _writeQueue_fifo_full;
  wire               _writeQueue_fifo_error;
  wire [49:0]        _writeQueue_fifo_data_out;
  wire [1023:0]      _extendUnit_out;
  wire               _reduceUnit_in_ready;
  wire               _reduceUnit_out_valid;
  wire [31:0]        _reduceUnit_out_bits_data;
  wire [3:0]         _reduceUnit_out_bits_mask;
  wire               _compressUnit_out_compressValid;
  wire [31:0]        _compressUnit_writeData;
  wire               _compressUnit_stageValid;
  wire               _readData_readDataQueue_fifo_31_empty;
  wire               _readData_readDataQueue_fifo_31_full;
  wire               _readData_readDataQueue_fifo_31_error;
  wire [31:0]        _readData_readDataQueue_fifo_31_data_out;
  wire               _readData_readDataQueue_fifo_30_empty;
  wire               _readData_readDataQueue_fifo_30_full;
  wire               _readData_readDataQueue_fifo_30_error;
  wire [31:0]        _readData_readDataQueue_fifo_30_data_out;
  wire               _readData_readDataQueue_fifo_29_empty;
  wire               _readData_readDataQueue_fifo_29_full;
  wire               _readData_readDataQueue_fifo_29_error;
  wire [31:0]        _readData_readDataQueue_fifo_29_data_out;
  wire               _readData_readDataQueue_fifo_28_empty;
  wire               _readData_readDataQueue_fifo_28_full;
  wire               _readData_readDataQueue_fifo_28_error;
  wire [31:0]        _readData_readDataQueue_fifo_28_data_out;
  wire               _readData_readDataQueue_fifo_27_empty;
  wire               _readData_readDataQueue_fifo_27_full;
  wire               _readData_readDataQueue_fifo_27_error;
  wire [31:0]        _readData_readDataQueue_fifo_27_data_out;
  wire               _readData_readDataQueue_fifo_26_empty;
  wire               _readData_readDataQueue_fifo_26_full;
  wire               _readData_readDataQueue_fifo_26_error;
  wire [31:0]        _readData_readDataQueue_fifo_26_data_out;
  wire               _readData_readDataQueue_fifo_25_empty;
  wire               _readData_readDataQueue_fifo_25_full;
  wire               _readData_readDataQueue_fifo_25_error;
  wire [31:0]        _readData_readDataQueue_fifo_25_data_out;
  wire               _readData_readDataQueue_fifo_24_empty;
  wire               _readData_readDataQueue_fifo_24_full;
  wire               _readData_readDataQueue_fifo_24_error;
  wire [31:0]        _readData_readDataQueue_fifo_24_data_out;
  wire               _readData_readDataQueue_fifo_23_empty;
  wire               _readData_readDataQueue_fifo_23_full;
  wire               _readData_readDataQueue_fifo_23_error;
  wire [31:0]        _readData_readDataQueue_fifo_23_data_out;
  wire               _readData_readDataQueue_fifo_22_empty;
  wire               _readData_readDataQueue_fifo_22_full;
  wire               _readData_readDataQueue_fifo_22_error;
  wire [31:0]        _readData_readDataQueue_fifo_22_data_out;
  wire               _readData_readDataQueue_fifo_21_empty;
  wire               _readData_readDataQueue_fifo_21_full;
  wire               _readData_readDataQueue_fifo_21_error;
  wire [31:0]        _readData_readDataQueue_fifo_21_data_out;
  wire               _readData_readDataQueue_fifo_20_empty;
  wire               _readData_readDataQueue_fifo_20_full;
  wire               _readData_readDataQueue_fifo_20_error;
  wire [31:0]        _readData_readDataQueue_fifo_20_data_out;
  wire               _readData_readDataQueue_fifo_19_empty;
  wire               _readData_readDataQueue_fifo_19_full;
  wire               _readData_readDataQueue_fifo_19_error;
  wire [31:0]        _readData_readDataQueue_fifo_19_data_out;
  wire               _readData_readDataQueue_fifo_18_empty;
  wire               _readData_readDataQueue_fifo_18_full;
  wire               _readData_readDataQueue_fifo_18_error;
  wire [31:0]        _readData_readDataQueue_fifo_18_data_out;
  wire               _readData_readDataQueue_fifo_17_empty;
  wire               _readData_readDataQueue_fifo_17_full;
  wire               _readData_readDataQueue_fifo_17_error;
  wire [31:0]        _readData_readDataQueue_fifo_17_data_out;
  wire               _readData_readDataQueue_fifo_16_empty;
  wire               _readData_readDataQueue_fifo_16_full;
  wire               _readData_readDataQueue_fifo_16_error;
  wire [31:0]        _readData_readDataQueue_fifo_16_data_out;
  wire               _readData_readDataQueue_fifo_15_empty;
  wire               _readData_readDataQueue_fifo_15_full;
  wire               _readData_readDataQueue_fifo_15_error;
  wire [31:0]        _readData_readDataQueue_fifo_15_data_out;
  wire               _readData_readDataQueue_fifo_14_empty;
  wire               _readData_readDataQueue_fifo_14_full;
  wire               _readData_readDataQueue_fifo_14_error;
  wire [31:0]        _readData_readDataQueue_fifo_14_data_out;
  wire               _readData_readDataQueue_fifo_13_empty;
  wire               _readData_readDataQueue_fifo_13_full;
  wire               _readData_readDataQueue_fifo_13_error;
  wire [31:0]        _readData_readDataQueue_fifo_13_data_out;
  wire               _readData_readDataQueue_fifo_12_empty;
  wire               _readData_readDataQueue_fifo_12_full;
  wire               _readData_readDataQueue_fifo_12_error;
  wire [31:0]        _readData_readDataQueue_fifo_12_data_out;
  wire               _readData_readDataQueue_fifo_11_empty;
  wire               _readData_readDataQueue_fifo_11_full;
  wire               _readData_readDataQueue_fifo_11_error;
  wire [31:0]        _readData_readDataQueue_fifo_11_data_out;
  wire               _readData_readDataQueue_fifo_10_empty;
  wire               _readData_readDataQueue_fifo_10_full;
  wire               _readData_readDataQueue_fifo_10_error;
  wire [31:0]        _readData_readDataQueue_fifo_10_data_out;
  wire               _readData_readDataQueue_fifo_9_empty;
  wire               _readData_readDataQueue_fifo_9_full;
  wire               _readData_readDataQueue_fifo_9_error;
  wire [31:0]        _readData_readDataQueue_fifo_9_data_out;
  wire               _readData_readDataQueue_fifo_8_empty;
  wire               _readData_readDataQueue_fifo_8_full;
  wire               _readData_readDataQueue_fifo_8_error;
  wire [31:0]        _readData_readDataQueue_fifo_8_data_out;
  wire               _readData_readDataQueue_fifo_7_empty;
  wire               _readData_readDataQueue_fifo_7_full;
  wire               _readData_readDataQueue_fifo_7_error;
  wire [31:0]        _readData_readDataQueue_fifo_7_data_out;
  wire               _readData_readDataQueue_fifo_6_empty;
  wire               _readData_readDataQueue_fifo_6_full;
  wire               _readData_readDataQueue_fifo_6_error;
  wire [31:0]        _readData_readDataQueue_fifo_6_data_out;
  wire               _readData_readDataQueue_fifo_5_empty;
  wire               _readData_readDataQueue_fifo_5_full;
  wire               _readData_readDataQueue_fifo_5_error;
  wire [31:0]        _readData_readDataQueue_fifo_5_data_out;
  wire               _readData_readDataQueue_fifo_4_empty;
  wire               _readData_readDataQueue_fifo_4_full;
  wire               _readData_readDataQueue_fifo_4_error;
  wire [31:0]        _readData_readDataQueue_fifo_4_data_out;
  wire               _readData_readDataQueue_fifo_3_empty;
  wire               _readData_readDataQueue_fifo_3_full;
  wire               _readData_readDataQueue_fifo_3_error;
  wire [31:0]        _readData_readDataQueue_fifo_3_data_out;
  wire               _readData_readDataQueue_fifo_2_empty;
  wire               _readData_readDataQueue_fifo_2_full;
  wire               _readData_readDataQueue_fifo_2_error;
  wire [31:0]        _readData_readDataQueue_fifo_2_data_out;
  wire               _readData_readDataQueue_fifo_1_empty;
  wire               _readData_readDataQueue_fifo_1_full;
  wire               _readData_readDataQueue_fifo_1_error;
  wire [31:0]        _readData_readDataQueue_fifo_1_data_out;
  wire               _readData_readDataQueue_fifo_empty;
  wire               _readData_readDataQueue_fifo_full;
  wire               _readData_readDataQueue_fifo_error;
  wire [31:0]        _readData_readDataQueue_fifo_data_out;
  wire               _readMessageQueue_fifo_31_empty;
  wire               _readMessageQueue_fifo_31_full;
  wire               _readMessageQueue_fifo_31_error;
  wire [33:0]        _readMessageQueue_fifo_31_data_out;
  wire               _readMessageQueue_fifo_30_empty;
  wire               _readMessageQueue_fifo_30_full;
  wire               _readMessageQueue_fifo_30_error;
  wire [33:0]        _readMessageQueue_fifo_30_data_out;
  wire               _readMessageQueue_fifo_29_empty;
  wire               _readMessageQueue_fifo_29_full;
  wire               _readMessageQueue_fifo_29_error;
  wire [33:0]        _readMessageQueue_fifo_29_data_out;
  wire               _readMessageQueue_fifo_28_empty;
  wire               _readMessageQueue_fifo_28_full;
  wire               _readMessageQueue_fifo_28_error;
  wire [33:0]        _readMessageQueue_fifo_28_data_out;
  wire               _readMessageQueue_fifo_27_empty;
  wire               _readMessageQueue_fifo_27_full;
  wire               _readMessageQueue_fifo_27_error;
  wire [33:0]        _readMessageQueue_fifo_27_data_out;
  wire               _readMessageQueue_fifo_26_empty;
  wire               _readMessageQueue_fifo_26_full;
  wire               _readMessageQueue_fifo_26_error;
  wire [33:0]        _readMessageQueue_fifo_26_data_out;
  wire               _readMessageQueue_fifo_25_empty;
  wire               _readMessageQueue_fifo_25_full;
  wire               _readMessageQueue_fifo_25_error;
  wire [33:0]        _readMessageQueue_fifo_25_data_out;
  wire               _readMessageQueue_fifo_24_empty;
  wire               _readMessageQueue_fifo_24_full;
  wire               _readMessageQueue_fifo_24_error;
  wire [33:0]        _readMessageQueue_fifo_24_data_out;
  wire               _readMessageQueue_fifo_23_empty;
  wire               _readMessageQueue_fifo_23_full;
  wire               _readMessageQueue_fifo_23_error;
  wire [33:0]        _readMessageQueue_fifo_23_data_out;
  wire               _readMessageQueue_fifo_22_empty;
  wire               _readMessageQueue_fifo_22_full;
  wire               _readMessageQueue_fifo_22_error;
  wire [33:0]        _readMessageQueue_fifo_22_data_out;
  wire               _readMessageQueue_fifo_21_empty;
  wire               _readMessageQueue_fifo_21_full;
  wire               _readMessageQueue_fifo_21_error;
  wire [33:0]        _readMessageQueue_fifo_21_data_out;
  wire               _readMessageQueue_fifo_20_empty;
  wire               _readMessageQueue_fifo_20_full;
  wire               _readMessageQueue_fifo_20_error;
  wire [33:0]        _readMessageQueue_fifo_20_data_out;
  wire               _readMessageQueue_fifo_19_empty;
  wire               _readMessageQueue_fifo_19_full;
  wire               _readMessageQueue_fifo_19_error;
  wire [33:0]        _readMessageQueue_fifo_19_data_out;
  wire               _readMessageQueue_fifo_18_empty;
  wire               _readMessageQueue_fifo_18_full;
  wire               _readMessageQueue_fifo_18_error;
  wire [33:0]        _readMessageQueue_fifo_18_data_out;
  wire               _readMessageQueue_fifo_17_empty;
  wire               _readMessageQueue_fifo_17_full;
  wire               _readMessageQueue_fifo_17_error;
  wire [33:0]        _readMessageQueue_fifo_17_data_out;
  wire               _readMessageQueue_fifo_16_empty;
  wire               _readMessageQueue_fifo_16_full;
  wire               _readMessageQueue_fifo_16_error;
  wire [33:0]        _readMessageQueue_fifo_16_data_out;
  wire               _readMessageQueue_fifo_15_empty;
  wire               _readMessageQueue_fifo_15_full;
  wire               _readMessageQueue_fifo_15_error;
  wire [33:0]        _readMessageQueue_fifo_15_data_out;
  wire               _readMessageQueue_fifo_14_empty;
  wire               _readMessageQueue_fifo_14_full;
  wire               _readMessageQueue_fifo_14_error;
  wire [33:0]        _readMessageQueue_fifo_14_data_out;
  wire               _readMessageQueue_fifo_13_empty;
  wire               _readMessageQueue_fifo_13_full;
  wire               _readMessageQueue_fifo_13_error;
  wire [33:0]        _readMessageQueue_fifo_13_data_out;
  wire               _readMessageQueue_fifo_12_empty;
  wire               _readMessageQueue_fifo_12_full;
  wire               _readMessageQueue_fifo_12_error;
  wire [33:0]        _readMessageQueue_fifo_12_data_out;
  wire               _readMessageQueue_fifo_11_empty;
  wire               _readMessageQueue_fifo_11_full;
  wire               _readMessageQueue_fifo_11_error;
  wire [33:0]        _readMessageQueue_fifo_11_data_out;
  wire               _readMessageQueue_fifo_10_empty;
  wire               _readMessageQueue_fifo_10_full;
  wire               _readMessageQueue_fifo_10_error;
  wire [33:0]        _readMessageQueue_fifo_10_data_out;
  wire               _readMessageQueue_fifo_9_empty;
  wire               _readMessageQueue_fifo_9_full;
  wire               _readMessageQueue_fifo_9_error;
  wire [33:0]        _readMessageQueue_fifo_9_data_out;
  wire               _readMessageQueue_fifo_8_empty;
  wire               _readMessageQueue_fifo_8_full;
  wire               _readMessageQueue_fifo_8_error;
  wire [33:0]        _readMessageQueue_fifo_8_data_out;
  wire               _readMessageQueue_fifo_7_empty;
  wire               _readMessageQueue_fifo_7_full;
  wire               _readMessageQueue_fifo_7_error;
  wire [33:0]        _readMessageQueue_fifo_7_data_out;
  wire               _readMessageQueue_fifo_6_empty;
  wire               _readMessageQueue_fifo_6_full;
  wire               _readMessageQueue_fifo_6_error;
  wire [33:0]        _readMessageQueue_fifo_6_data_out;
  wire               _readMessageQueue_fifo_5_empty;
  wire               _readMessageQueue_fifo_5_full;
  wire               _readMessageQueue_fifo_5_error;
  wire [33:0]        _readMessageQueue_fifo_5_data_out;
  wire               _readMessageQueue_fifo_4_empty;
  wire               _readMessageQueue_fifo_4_full;
  wire               _readMessageQueue_fifo_4_error;
  wire [33:0]        _readMessageQueue_fifo_4_data_out;
  wire               _readMessageQueue_fifo_3_empty;
  wire               _readMessageQueue_fifo_3_full;
  wire               _readMessageQueue_fifo_3_error;
  wire [33:0]        _readMessageQueue_fifo_3_data_out;
  wire               _readMessageQueue_fifo_2_empty;
  wire               _readMessageQueue_fifo_2_full;
  wire               _readMessageQueue_fifo_2_error;
  wire [33:0]        _readMessageQueue_fifo_2_data_out;
  wire               _readMessageQueue_fifo_1_empty;
  wire               _readMessageQueue_fifo_1_full;
  wire               _readMessageQueue_fifo_1_error;
  wire [33:0]        _readMessageQueue_fifo_1_data_out;
  wire               _readMessageQueue_fifo_empty;
  wire               _readMessageQueue_fifo_full;
  wire               _readMessageQueue_fifo_error;
  wire [33:0]        _readMessageQueue_fifo_data_out;
  wire               _reorderQueueVec_fifo_31_empty;
  wire               _reorderQueueVec_fifo_31_full;
  wire               _reorderQueueVec_fifo_31_error;
  wire [63:0]        _reorderQueueVec_fifo_31_data_out;
  wire               _reorderQueueVec_fifo_30_empty;
  wire               _reorderQueueVec_fifo_30_full;
  wire               _reorderQueueVec_fifo_30_error;
  wire [63:0]        _reorderQueueVec_fifo_30_data_out;
  wire               _reorderQueueVec_fifo_29_empty;
  wire               _reorderQueueVec_fifo_29_full;
  wire               _reorderQueueVec_fifo_29_error;
  wire [63:0]        _reorderQueueVec_fifo_29_data_out;
  wire               _reorderQueueVec_fifo_28_empty;
  wire               _reorderQueueVec_fifo_28_full;
  wire               _reorderQueueVec_fifo_28_error;
  wire [63:0]        _reorderQueueVec_fifo_28_data_out;
  wire               _reorderQueueVec_fifo_27_empty;
  wire               _reorderQueueVec_fifo_27_full;
  wire               _reorderQueueVec_fifo_27_error;
  wire [63:0]        _reorderQueueVec_fifo_27_data_out;
  wire               _reorderQueueVec_fifo_26_empty;
  wire               _reorderQueueVec_fifo_26_full;
  wire               _reorderQueueVec_fifo_26_error;
  wire [63:0]        _reorderQueueVec_fifo_26_data_out;
  wire               _reorderQueueVec_fifo_25_empty;
  wire               _reorderQueueVec_fifo_25_full;
  wire               _reorderQueueVec_fifo_25_error;
  wire [63:0]        _reorderQueueVec_fifo_25_data_out;
  wire               _reorderQueueVec_fifo_24_empty;
  wire               _reorderQueueVec_fifo_24_full;
  wire               _reorderQueueVec_fifo_24_error;
  wire [63:0]        _reorderQueueVec_fifo_24_data_out;
  wire               _reorderQueueVec_fifo_23_empty;
  wire               _reorderQueueVec_fifo_23_full;
  wire               _reorderQueueVec_fifo_23_error;
  wire [63:0]        _reorderQueueVec_fifo_23_data_out;
  wire               _reorderQueueVec_fifo_22_empty;
  wire               _reorderQueueVec_fifo_22_full;
  wire               _reorderQueueVec_fifo_22_error;
  wire [63:0]        _reorderQueueVec_fifo_22_data_out;
  wire               _reorderQueueVec_fifo_21_empty;
  wire               _reorderQueueVec_fifo_21_full;
  wire               _reorderQueueVec_fifo_21_error;
  wire [63:0]        _reorderQueueVec_fifo_21_data_out;
  wire               _reorderQueueVec_fifo_20_empty;
  wire               _reorderQueueVec_fifo_20_full;
  wire               _reorderQueueVec_fifo_20_error;
  wire [63:0]        _reorderQueueVec_fifo_20_data_out;
  wire               _reorderQueueVec_fifo_19_empty;
  wire               _reorderQueueVec_fifo_19_full;
  wire               _reorderQueueVec_fifo_19_error;
  wire [63:0]        _reorderQueueVec_fifo_19_data_out;
  wire               _reorderQueueVec_fifo_18_empty;
  wire               _reorderQueueVec_fifo_18_full;
  wire               _reorderQueueVec_fifo_18_error;
  wire [63:0]        _reorderQueueVec_fifo_18_data_out;
  wire               _reorderQueueVec_fifo_17_empty;
  wire               _reorderQueueVec_fifo_17_full;
  wire               _reorderQueueVec_fifo_17_error;
  wire [63:0]        _reorderQueueVec_fifo_17_data_out;
  wire               _reorderQueueVec_fifo_16_empty;
  wire               _reorderQueueVec_fifo_16_full;
  wire               _reorderQueueVec_fifo_16_error;
  wire [63:0]        _reorderQueueVec_fifo_16_data_out;
  wire               _reorderQueueVec_fifo_15_empty;
  wire               _reorderQueueVec_fifo_15_full;
  wire               _reorderQueueVec_fifo_15_error;
  wire [63:0]        _reorderQueueVec_fifo_15_data_out;
  wire               _reorderQueueVec_fifo_14_empty;
  wire               _reorderQueueVec_fifo_14_full;
  wire               _reorderQueueVec_fifo_14_error;
  wire [63:0]        _reorderQueueVec_fifo_14_data_out;
  wire               _reorderQueueVec_fifo_13_empty;
  wire               _reorderQueueVec_fifo_13_full;
  wire               _reorderQueueVec_fifo_13_error;
  wire [63:0]        _reorderQueueVec_fifo_13_data_out;
  wire               _reorderQueueVec_fifo_12_empty;
  wire               _reorderQueueVec_fifo_12_full;
  wire               _reorderQueueVec_fifo_12_error;
  wire [63:0]        _reorderQueueVec_fifo_12_data_out;
  wire               _reorderQueueVec_fifo_11_empty;
  wire               _reorderQueueVec_fifo_11_full;
  wire               _reorderQueueVec_fifo_11_error;
  wire [63:0]        _reorderQueueVec_fifo_11_data_out;
  wire               _reorderQueueVec_fifo_10_empty;
  wire               _reorderQueueVec_fifo_10_full;
  wire               _reorderQueueVec_fifo_10_error;
  wire [63:0]        _reorderQueueVec_fifo_10_data_out;
  wire               _reorderQueueVec_fifo_9_empty;
  wire               _reorderQueueVec_fifo_9_full;
  wire               _reorderQueueVec_fifo_9_error;
  wire [63:0]        _reorderQueueVec_fifo_9_data_out;
  wire               _reorderQueueVec_fifo_8_empty;
  wire               _reorderQueueVec_fifo_8_full;
  wire               _reorderQueueVec_fifo_8_error;
  wire [63:0]        _reorderQueueVec_fifo_8_data_out;
  wire               _reorderQueueVec_fifo_7_empty;
  wire               _reorderQueueVec_fifo_7_full;
  wire               _reorderQueueVec_fifo_7_error;
  wire [63:0]        _reorderQueueVec_fifo_7_data_out;
  wire               _reorderQueueVec_fifo_6_empty;
  wire               _reorderQueueVec_fifo_6_full;
  wire               _reorderQueueVec_fifo_6_error;
  wire [63:0]        _reorderQueueVec_fifo_6_data_out;
  wire               _reorderQueueVec_fifo_5_empty;
  wire               _reorderQueueVec_fifo_5_full;
  wire               _reorderQueueVec_fifo_5_error;
  wire [63:0]        _reorderQueueVec_fifo_5_data_out;
  wire               _reorderQueueVec_fifo_4_empty;
  wire               _reorderQueueVec_fifo_4_full;
  wire               _reorderQueueVec_fifo_4_error;
  wire [63:0]        _reorderQueueVec_fifo_4_data_out;
  wire               _reorderQueueVec_fifo_3_empty;
  wire               _reorderQueueVec_fifo_3_full;
  wire               _reorderQueueVec_fifo_3_error;
  wire [63:0]        _reorderQueueVec_fifo_3_data_out;
  wire               _reorderQueueVec_fifo_2_empty;
  wire               _reorderQueueVec_fifo_2_full;
  wire               _reorderQueueVec_fifo_2_error;
  wire [63:0]        _reorderQueueVec_fifo_2_data_out;
  wire               _reorderQueueVec_fifo_1_empty;
  wire               _reorderQueueVec_fifo_1_full;
  wire               _reorderQueueVec_fifo_1_error;
  wire [63:0]        _reorderQueueVec_fifo_1_data_out;
  wire               _reorderQueueVec_fifo_empty;
  wire               _reorderQueueVec_fifo_full;
  wire               _reorderQueueVec_fifo_error;
  wire [63:0]        _reorderQueueVec_fifo_data_out;
  wire               _compressUnitResultQueue_fifo_empty;
  wire               _compressUnitResultQueue_fifo_full;
  wire               _compressUnitResultQueue_fifo_error;
  wire [1189:0]      _compressUnitResultQueue_fifo_data_out;
  wire               _readWaitQueue_fifo_empty;
  wire               _readWaitQueue_fifo_full;
  wire               _readWaitQueue_fifo_error;
  wire [103:0]       _readWaitQueue_fifo_data_out;
  wire               _readCrossBar_input_0_ready;
  wire               _readCrossBar_input_1_ready;
  wire               _readCrossBar_input_2_ready;
  wire               _readCrossBar_input_3_ready;
  wire               _readCrossBar_input_4_ready;
  wire               _readCrossBar_input_5_ready;
  wire               _readCrossBar_input_6_ready;
  wire               _readCrossBar_input_7_ready;
  wire               _readCrossBar_input_8_ready;
  wire               _readCrossBar_input_9_ready;
  wire               _readCrossBar_input_10_ready;
  wire               _readCrossBar_input_11_ready;
  wire               _readCrossBar_input_12_ready;
  wire               _readCrossBar_input_13_ready;
  wire               _readCrossBar_input_14_ready;
  wire               _readCrossBar_input_15_ready;
  wire               _readCrossBar_input_16_ready;
  wire               _readCrossBar_input_17_ready;
  wire               _readCrossBar_input_18_ready;
  wire               _readCrossBar_input_19_ready;
  wire               _readCrossBar_input_20_ready;
  wire               _readCrossBar_input_21_ready;
  wire               _readCrossBar_input_22_ready;
  wire               _readCrossBar_input_23_ready;
  wire               _readCrossBar_input_24_ready;
  wire               _readCrossBar_input_25_ready;
  wire               _readCrossBar_input_26_ready;
  wire               _readCrossBar_input_27_ready;
  wire               _readCrossBar_input_28_ready;
  wire               _readCrossBar_input_29_ready;
  wire               _readCrossBar_input_30_ready;
  wire               _readCrossBar_input_31_ready;
  wire               _readCrossBar_output_0_valid;
  wire [4:0]         _readCrossBar_output_0_bits_vs;
  wire               _readCrossBar_output_0_bits_offset;
  wire [4:0]         _readCrossBar_output_0_bits_writeIndex;
  wire               _readCrossBar_output_1_valid;
  wire [4:0]         _readCrossBar_output_1_bits_vs;
  wire               _readCrossBar_output_1_bits_offset;
  wire [4:0]         _readCrossBar_output_1_bits_writeIndex;
  wire               _readCrossBar_output_2_valid;
  wire [4:0]         _readCrossBar_output_2_bits_vs;
  wire               _readCrossBar_output_2_bits_offset;
  wire [4:0]         _readCrossBar_output_2_bits_writeIndex;
  wire               _readCrossBar_output_3_valid;
  wire [4:0]         _readCrossBar_output_3_bits_vs;
  wire               _readCrossBar_output_3_bits_offset;
  wire [4:0]         _readCrossBar_output_3_bits_writeIndex;
  wire               _readCrossBar_output_4_valid;
  wire [4:0]         _readCrossBar_output_4_bits_vs;
  wire               _readCrossBar_output_4_bits_offset;
  wire [4:0]         _readCrossBar_output_4_bits_writeIndex;
  wire               _readCrossBar_output_5_valid;
  wire [4:0]         _readCrossBar_output_5_bits_vs;
  wire               _readCrossBar_output_5_bits_offset;
  wire [4:0]         _readCrossBar_output_5_bits_writeIndex;
  wire               _readCrossBar_output_6_valid;
  wire [4:0]         _readCrossBar_output_6_bits_vs;
  wire               _readCrossBar_output_6_bits_offset;
  wire [4:0]         _readCrossBar_output_6_bits_writeIndex;
  wire               _readCrossBar_output_7_valid;
  wire [4:0]         _readCrossBar_output_7_bits_vs;
  wire               _readCrossBar_output_7_bits_offset;
  wire [4:0]         _readCrossBar_output_7_bits_writeIndex;
  wire               _readCrossBar_output_8_valid;
  wire [4:0]         _readCrossBar_output_8_bits_vs;
  wire               _readCrossBar_output_8_bits_offset;
  wire [4:0]         _readCrossBar_output_8_bits_writeIndex;
  wire               _readCrossBar_output_9_valid;
  wire [4:0]         _readCrossBar_output_9_bits_vs;
  wire               _readCrossBar_output_9_bits_offset;
  wire [4:0]         _readCrossBar_output_9_bits_writeIndex;
  wire               _readCrossBar_output_10_valid;
  wire [4:0]         _readCrossBar_output_10_bits_vs;
  wire               _readCrossBar_output_10_bits_offset;
  wire [4:0]         _readCrossBar_output_10_bits_writeIndex;
  wire               _readCrossBar_output_11_valid;
  wire [4:0]         _readCrossBar_output_11_bits_vs;
  wire               _readCrossBar_output_11_bits_offset;
  wire [4:0]         _readCrossBar_output_11_bits_writeIndex;
  wire               _readCrossBar_output_12_valid;
  wire [4:0]         _readCrossBar_output_12_bits_vs;
  wire               _readCrossBar_output_12_bits_offset;
  wire [4:0]         _readCrossBar_output_12_bits_writeIndex;
  wire               _readCrossBar_output_13_valid;
  wire [4:0]         _readCrossBar_output_13_bits_vs;
  wire               _readCrossBar_output_13_bits_offset;
  wire [4:0]         _readCrossBar_output_13_bits_writeIndex;
  wire               _readCrossBar_output_14_valid;
  wire [4:0]         _readCrossBar_output_14_bits_vs;
  wire               _readCrossBar_output_14_bits_offset;
  wire [4:0]         _readCrossBar_output_14_bits_writeIndex;
  wire               _readCrossBar_output_15_valid;
  wire [4:0]         _readCrossBar_output_15_bits_vs;
  wire               _readCrossBar_output_15_bits_offset;
  wire [4:0]         _readCrossBar_output_15_bits_writeIndex;
  wire               _readCrossBar_output_16_valid;
  wire [4:0]         _readCrossBar_output_16_bits_vs;
  wire               _readCrossBar_output_16_bits_offset;
  wire [4:0]         _readCrossBar_output_16_bits_writeIndex;
  wire               _readCrossBar_output_17_valid;
  wire [4:0]         _readCrossBar_output_17_bits_vs;
  wire               _readCrossBar_output_17_bits_offset;
  wire [4:0]         _readCrossBar_output_17_bits_writeIndex;
  wire               _readCrossBar_output_18_valid;
  wire [4:0]         _readCrossBar_output_18_bits_vs;
  wire               _readCrossBar_output_18_bits_offset;
  wire [4:0]         _readCrossBar_output_18_bits_writeIndex;
  wire               _readCrossBar_output_19_valid;
  wire [4:0]         _readCrossBar_output_19_bits_vs;
  wire               _readCrossBar_output_19_bits_offset;
  wire [4:0]         _readCrossBar_output_19_bits_writeIndex;
  wire               _readCrossBar_output_20_valid;
  wire [4:0]         _readCrossBar_output_20_bits_vs;
  wire               _readCrossBar_output_20_bits_offset;
  wire [4:0]         _readCrossBar_output_20_bits_writeIndex;
  wire               _readCrossBar_output_21_valid;
  wire [4:0]         _readCrossBar_output_21_bits_vs;
  wire               _readCrossBar_output_21_bits_offset;
  wire [4:0]         _readCrossBar_output_21_bits_writeIndex;
  wire               _readCrossBar_output_22_valid;
  wire [4:0]         _readCrossBar_output_22_bits_vs;
  wire               _readCrossBar_output_22_bits_offset;
  wire [4:0]         _readCrossBar_output_22_bits_writeIndex;
  wire               _readCrossBar_output_23_valid;
  wire [4:0]         _readCrossBar_output_23_bits_vs;
  wire               _readCrossBar_output_23_bits_offset;
  wire [4:0]         _readCrossBar_output_23_bits_writeIndex;
  wire               _readCrossBar_output_24_valid;
  wire [4:0]         _readCrossBar_output_24_bits_vs;
  wire               _readCrossBar_output_24_bits_offset;
  wire [4:0]         _readCrossBar_output_24_bits_writeIndex;
  wire               _readCrossBar_output_25_valid;
  wire [4:0]         _readCrossBar_output_25_bits_vs;
  wire               _readCrossBar_output_25_bits_offset;
  wire [4:0]         _readCrossBar_output_25_bits_writeIndex;
  wire               _readCrossBar_output_26_valid;
  wire [4:0]         _readCrossBar_output_26_bits_vs;
  wire               _readCrossBar_output_26_bits_offset;
  wire [4:0]         _readCrossBar_output_26_bits_writeIndex;
  wire               _readCrossBar_output_27_valid;
  wire [4:0]         _readCrossBar_output_27_bits_vs;
  wire               _readCrossBar_output_27_bits_offset;
  wire [4:0]         _readCrossBar_output_27_bits_writeIndex;
  wire               _readCrossBar_output_28_valid;
  wire [4:0]         _readCrossBar_output_28_bits_vs;
  wire               _readCrossBar_output_28_bits_offset;
  wire [4:0]         _readCrossBar_output_28_bits_writeIndex;
  wire               _readCrossBar_output_29_valid;
  wire [4:0]         _readCrossBar_output_29_bits_vs;
  wire               _readCrossBar_output_29_bits_offset;
  wire [4:0]         _readCrossBar_output_29_bits_writeIndex;
  wire               _readCrossBar_output_30_valid;
  wire [4:0]         _readCrossBar_output_30_bits_vs;
  wire               _readCrossBar_output_30_bits_offset;
  wire [4:0]         _readCrossBar_output_30_bits_writeIndex;
  wire               _readCrossBar_output_31_valid;
  wire [4:0]         _readCrossBar_output_31_bits_vs;
  wire               _readCrossBar_output_31_bits_offset;
  wire [4:0]         _readCrossBar_output_31_bits_writeIndex;
  wire               _accessCountQueue_fifo_empty;
  wire               _accessCountQueue_fifo_full;
  wire               _accessCountQueue_fifo_error;
  wire [191:0]       _accessCountQueue_fifo_data_out;
  wire               _slideAddressGen_indexDeq_valid;
  wire [31:0]        _slideAddressGen_indexDeq_bits_needRead;
  wire [31:0]        _slideAddressGen_indexDeq_bits_elementValid;
  wire [31:0]        _slideAddressGen_indexDeq_bits_replaceVs1;
  wire [31:0]        _slideAddressGen_indexDeq_bits_readOffset;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_0;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_1;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_2;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_3;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_4;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_5;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_6;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_7;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_8;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_9;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_10;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_11;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_12;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_13;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_14;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_15;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_16;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_17;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_18;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_19;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_20;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_21;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_22;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_23;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_24;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_25;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_26;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_27;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_28;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_29;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_30;
  wire [4:0]         _slideAddressGen_indexDeq_bits_accessLane_31;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_0;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_1;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_2;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_3;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_4;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_5;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_6;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_7;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_8;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_9;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_10;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_11;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_12;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_13;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_14;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_15;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_16;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_17;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_18;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_19;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_20;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_21;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_22;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_23;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_24;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_25;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_26;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_27;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_28;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_29;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_30;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_31;
  wire [6:0]         _slideAddressGen_indexDeq_bits_executeGroup;
  wire [63:0]        _slideAddressGen_indexDeq_bits_readDataOffset;
  wire               _slideAddressGen_indexDeq_bits_last;
  wire [6:0]         _slideAddressGen_slideGroupOut;
  wire               _exeRequestQueue_queue_fifo_31_empty;
  wire               _exeRequestQueue_queue_fifo_31_full;
  wire               _exeRequestQueue_queue_fifo_31_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_31_data_out;
  wire               _exeRequestQueue_queue_fifo_30_empty;
  wire               _exeRequestQueue_queue_fifo_30_full;
  wire               _exeRequestQueue_queue_fifo_30_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_30_data_out;
  wire               _exeRequestQueue_queue_fifo_29_empty;
  wire               _exeRequestQueue_queue_fifo_29_full;
  wire               _exeRequestQueue_queue_fifo_29_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_29_data_out;
  wire               _exeRequestQueue_queue_fifo_28_empty;
  wire               _exeRequestQueue_queue_fifo_28_full;
  wire               _exeRequestQueue_queue_fifo_28_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_28_data_out;
  wire               _exeRequestQueue_queue_fifo_27_empty;
  wire               _exeRequestQueue_queue_fifo_27_full;
  wire               _exeRequestQueue_queue_fifo_27_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_27_data_out;
  wire               _exeRequestQueue_queue_fifo_26_empty;
  wire               _exeRequestQueue_queue_fifo_26_full;
  wire               _exeRequestQueue_queue_fifo_26_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_26_data_out;
  wire               _exeRequestQueue_queue_fifo_25_empty;
  wire               _exeRequestQueue_queue_fifo_25_full;
  wire               _exeRequestQueue_queue_fifo_25_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_25_data_out;
  wire               _exeRequestQueue_queue_fifo_24_empty;
  wire               _exeRequestQueue_queue_fifo_24_full;
  wire               _exeRequestQueue_queue_fifo_24_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_24_data_out;
  wire               _exeRequestQueue_queue_fifo_23_empty;
  wire               _exeRequestQueue_queue_fifo_23_full;
  wire               _exeRequestQueue_queue_fifo_23_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_23_data_out;
  wire               _exeRequestQueue_queue_fifo_22_empty;
  wire               _exeRequestQueue_queue_fifo_22_full;
  wire               _exeRequestQueue_queue_fifo_22_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_22_data_out;
  wire               _exeRequestQueue_queue_fifo_21_empty;
  wire               _exeRequestQueue_queue_fifo_21_full;
  wire               _exeRequestQueue_queue_fifo_21_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_21_data_out;
  wire               _exeRequestQueue_queue_fifo_20_empty;
  wire               _exeRequestQueue_queue_fifo_20_full;
  wire               _exeRequestQueue_queue_fifo_20_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_20_data_out;
  wire               _exeRequestQueue_queue_fifo_19_empty;
  wire               _exeRequestQueue_queue_fifo_19_full;
  wire               _exeRequestQueue_queue_fifo_19_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_19_data_out;
  wire               _exeRequestQueue_queue_fifo_18_empty;
  wire               _exeRequestQueue_queue_fifo_18_full;
  wire               _exeRequestQueue_queue_fifo_18_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_18_data_out;
  wire               _exeRequestQueue_queue_fifo_17_empty;
  wire               _exeRequestQueue_queue_fifo_17_full;
  wire               _exeRequestQueue_queue_fifo_17_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_17_data_out;
  wire               _exeRequestQueue_queue_fifo_16_empty;
  wire               _exeRequestQueue_queue_fifo_16_full;
  wire               _exeRequestQueue_queue_fifo_16_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_16_data_out;
  wire               _exeRequestQueue_queue_fifo_15_empty;
  wire               _exeRequestQueue_queue_fifo_15_full;
  wire               _exeRequestQueue_queue_fifo_15_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_15_data_out;
  wire               _exeRequestQueue_queue_fifo_14_empty;
  wire               _exeRequestQueue_queue_fifo_14_full;
  wire               _exeRequestQueue_queue_fifo_14_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_14_data_out;
  wire               _exeRequestQueue_queue_fifo_13_empty;
  wire               _exeRequestQueue_queue_fifo_13_full;
  wire               _exeRequestQueue_queue_fifo_13_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_13_data_out;
  wire               _exeRequestQueue_queue_fifo_12_empty;
  wire               _exeRequestQueue_queue_fifo_12_full;
  wire               _exeRequestQueue_queue_fifo_12_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_12_data_out;
  wire               _exeRequestQueue_queue_fifo_11_empty;
  wire               _exeRequestQueue_queue_fifo_11_full;
  wire               _exeRequestQueue_queue_fifo_11_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_11_data_out;
  wire               _exeRequestQueue_queue_fifo_10_empty;
  wire               _exeRequestQueue_queue_fifo_10_full;
  wire               _exeRequestQueue_queue_fifo_10_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_10_data_out;
  wire               _exeRequestQueue_queue_fifo_9_empty;
  wire               _exeRequestQueue_queue_fifo_9_full;
  wire               _exeRequestQueue_queue_fifo_9_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_9_data_out;
  wire               _exeRequestQueue_queue_fifo_8_empty;
  wire               _exeRequestQueue_queue_fifo_8_full;
  wire               _exeRequestQueue_queue_fifo_8_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_8_data_out;
  wire               _exeRequestQueue_queue_fifo_7_empty;
  wire               _exeRequestQueue_queue_fifo_7_full;
  wire               _exeRequestQueue_queue_fifo_7_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_7_data_out;
  wire               _exeRequestQueue_queue_fifo_6_empty;
  wire               _exeRequestQueue_queue_fifo_6_full;
  wire               _exeRequestQueue_queue_fifo_6_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_6_data_out;
  wire               _exeRequestQueue_queue_fifo_5_empty;
  wire               _exeRequestQueue_queue_fifo_5_full;
  wire               _exeRequestQueue_queue_fifo_5_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_5_data_out;
  wire               _exeRequestQueue_queue_fifo_4_empty;
  wire               _exeRequestQueue_queue_fifo_4_full;
  wire               _exeRequestQueue_queue_fifo_4_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_4_data_out;
  wire               _exeRequestQueue_queue_fifo_3_empty;
  wire               _exeRequestQueue_queue_fifo_3_full;
  wire               _exeRequestQueue_queue_fifo_3_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_3_data_out;
  wire               _exeRequestQueue_queue_fifo_2_empty;
  wire               _exeRequestQueue_queue_fifo_2_full;
  wire               _exeRequestQueue_queue_fifo_2_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_2_data_out;
  wire               _exeRequestQueue_queue_fifo_1_empty;
  wire               _exeRequestQueue_queue_fifo_1_full;
  wire               _exeRequestQueue_queue_fifo_1_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_1_data_out;
  wire               _exeRequestQueue_queue_fifo_empty;
  wire               _exeRequestQueue_queue_fifo_full;
  wire               _exeRequestQueue_queue_fifo_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_data_out;
  wire               _maskedWrite_in_0_ready;
  wire               _maskedWrite_in_1_ready;
  wire               _maskedWrite_in_2_ready;
  wire               _maskedWrite_in_3_ready;
  wire               _maskedWrite_in_4_ready;
  wire               _maskedWrite_in_5_ready;
  wire               _maskedWrite_in_6_ready;
  wire               _maskedWrite_in_7_ready;
  wire               _maskedWrite_in_8_ready;
  wire               _maskedWrite_in_9_ready;
  wire               _maskedWrite_in_10_ready;
  wire               _maskedWrite_in_11_ready;
  wire               _maskedWrite_in_12_ready;
  wire               _maskedWrite_in_13_ready;
  wire               _maskedWrite_in_14_ready;
  wire               _maskedWrite_in_15_ready;
  wire               _maskedWrite_in_16_ready;
  wire               _maskedWrite_in_17_ready;
  wire               _maskedWrite_in_18_ready;
  wire               _maskedWrite_in_19_ready;
  wire               _maskedWrite_in_20_ready;
  wire               _maskedWrite_in_21_ready;
  wire               _maskedWrite_in_22_ready;
  wire               _maskedWrite_in_23_ready;
  wire               _maskedWrite_in_24_ready;
  wire               _maskedWrite_in_25_ready;
  wire               _maskedWrite_in_26_ready;
  wire               _maskedWrite_in_27_ready;
  wire               _maskedWrite_in_28_ready;
  wire               _maskedWrite_in_29_ready;
  wire               _maskedWrite_in_30_ready;
  wire               _maskedWrite_in_31_ready;
  wire               _maskedWrite_out_0_valid;
  wire               _maskedWrite_out_0_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_0_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_0_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_0_bits_writeData_groupCounter;
  wire               _maskedWrite_out_1_valid;
  wire               _maskedWrite_out_1_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_1_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_1_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_1_bits_writeData_groupCounter;
  wire               _maskedWrite_out_2_valid;
  wire               _maskedWrite_out_2_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_2_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_2_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_2_bits_writeData_groupCounter;
  wire               _maskedWrite_out_3_valid;
  wire               _maskedWrite_out_3_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_3_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_3_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_3_bits_writeData_groupCounter;
  wire               _maskedWrite_out_4_valid;
  wire               _maskedWrite_out_4_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_4_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_4_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_4_bits_writeData_groupCounter;
  wire               _maskedWrite_out_5_valid;
  wire               _maskedWrite_out_5_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_5_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_5_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_5_bits_writeData_groupCounter;
  wire               _maskedWrite_out_6_valid;
  wire               _maskedWrite_out_6_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_6_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_6_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_6_bits_writeData_groupCounter;
  wire               _maskedWrite_out_7_valid;
  wire               _maskedWrite_out_7_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_7_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_7_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_7_bits_writeData_groupCounter;
  wire               _maskedWrite_out_8_valid;
  wire               _maskedWrite_out_8_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_8_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_8_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_8_bits_writeData_groupCounter;
  wire               _maskedWrite_out_9_valid;
  wire               _maskedWrite_out_9_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_9_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_9_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_9_bits_writeData_groupCounter;
  wire               _maskedWrite_out_10_valid;
  wire               _maskedWrite_out_10_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_10_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_10_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_10_bits_writeData_groupCounter;
  wire               _maskedWrite_out_11_valid;
  wire               _maskedWrite_out_11_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_11_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_11_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_11_bits_writeData_groupCounter;
  wire               _maskedWrite_out_12_valid;
  wire               _maskedWrite_out_12_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_12_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_12_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_12_bits_writeData_groupCounter;
  wire               _maskedWrite_out_13_valid;
  wire               _maskedWrite_out_13_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_13_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_13_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_13_bits_writeData_groupCounter;
  wire               _maskedWrite_out_14_valid;
  wire               _maskedWrite_out_14_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_14_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_14_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_14_bits_writeData_groupCounter;
  wire               _maskedWrite_out_15_valid;
  wire               _maskedWrite_out_15_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_15_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_15_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_15_bits_writeData_groupCounter;
  wire               _maskedWrite_out_16_valid;
  wire               _maskedWrite_out_16_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_16_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_16_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_16_bits_writeData_groupCounter;
  wire               _maskedWrite_out_17_valid;
  wire               _maskedWrite_out_17_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_17_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_17_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_17_bits_writeData_groupCounter;
  wire               _maskedWrite_out_18_valid;
  wire               _maskedWrite_out_18_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_18_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_18_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_18_bits_writeData_groupCounter;
  wire               _maskedWrite_out_19_valid;
  wire               _maskedWrite_out_19_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_19_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_19_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_19_bits_writeData_groupCounter;
  wire               _maskedWrite_out_20_valid;
  wire               _maskedWrite_out_20_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_20_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_20_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_20_bits_writeData_groupCounter;
  wire               _maskedWrite_out_21_valid;
  wire               _maskedWrite_out_21_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_21_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_21_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_21_bits_writeData_groupCounter;
  wire               _maskedWrite_out_22_valid;
  wire               _maskedWrite_out_22_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_22_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_22_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_22_bits_writeData_groupCounter;
  wire               _maskedWrite_out_23_valid;
  wire               _maskedWrite_out_23_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_23_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_23_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_23_bits_writeData_groupCounter;
  wire               _maskedWrite_out_24_valid;
  wire               _maskedWrite_out_24_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_24_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_24_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_24_bits_writeData_groupCounter;
  wire               _maskedWrite_out_25_valid;
  wire               _maskedWrite_out_25_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_25_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_25_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_25_bits_writeData_groupCounter;
  wire               _maskedWrite_out_26_valid;
  wire               _maskedWrite_out_26_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_26_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_26_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_26_bits_writeData_groupCounter;
  wire               _maskedWrite_out_27_valid;
  wire               _maskedWrite_out_27_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_27_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_27_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_27_bits_writeData_groupCounter;
  wire               _maskedWrite_out_28_valid;
  wire               _maskedWrite_out_28_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_28_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_28_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_28_bits_writeData_groupCounter;
  wire               _maskedWrite_out_29_valid;
  wire               _maskedWrite_out_29_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_29_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_29_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_29_bits_writeData_groupCounter;
  wire               _maskedWrite_out_30_valid;
  wire               _maskedWrite_out_30_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_30_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_30_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_30_bits_writeData_groupCounter;
  wire               _maskedWrite_out_31_valid;
  wire               _maskedWrite_out_31_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_31_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_31_bits_writeData_mask;
  wire [4:0]         _maskedWrite_out_31_bits_writeData_groupCounter;
  wire               _maskedWrite_readChannel_0_valid;
  wire [4:0]         _maskedWrite_readChannel_0_bits_vs;
  wire               _maskedWrite_readChannel_0_bits_offset;
  wire               _maskedWrite_readChannel_1_valid;
  wire [4:0]         _maskedWrite_readChannel_1_bits_vs;
  wire               _maskedWrite_readChannel_1_bits_offset;
  wire               _maskedWrite_readChannel_2_valid;
  wire [4:0]         _maskedWrite_readChannel_2_bits_vs;
  wire               _maskedWrite_readChannel_2_bits_offset;
  wire               _maskedWrite_readChannel_3_valid;
  wire [4:0]         _maskedWrite_readChannel_3_bits_vs;
  wire               _maskedWrite_readChannel_3_bits_offset;
  wire               _maskedWrite_readChannel_4_valid;
  wire [4:0]         _maskedWrite_readChannel_4_bits_vs;
  wire               _maskedWrite_readChannel_4_bits_offset;
  wire               _maskedWrite_readChannel_5_valid;
  wire [4:0]         _maskedWrite_readChannel_5_bits_vs;
  wire               _maskedWrite_readChannel_5_bits_offset;
  wire               _maskedWrite_readChannel_6_valid;
  wire [4:0]         _maskedWrite_readChannel_6_bits_vs;
  wire               _maskedWrite_readChannel_6_bits_offset;
  wire               _maskedWrite_readChannel_7_valid;
  wire [4:0]         _maskedWrite_readChannel_7_bits_vs;
  wire               _maskedWrite_readChannel_7_bits_offset;
  wire               _maskedWrite_readChannel_8_valid;
  wire [4:0]         _maskedWrite_readChannel_8_bits_vs;
  wire               _maskedWrite_readChannel_8_bits_offset;
  wire               _maskedWrite_readChannel_9_valid;
  wire [4:0]         _maskedWrite_readChannel_9_bits_vs;
  wire               _maskedWrite_readChannel_9_bits_offset;
  wire               _maskedWrite_readChannel_10_valid;
  wire [4:0]         _maskedWrite_readChannel_10_bits_vs;
  wire               _maskedWrite_readChannel_10_bits_offset;
  wire               _maskedWrite_readChannel_11_valid;
  wire [4:0]         _maskedWrite_readChannel_11_bits_vs;
  wire               _maskedWrite_readChannel_11_bits_offset;
  wire               _maskedWrite_readChannel_12_valid;
  wire [4:0]         _maskedWrite_readChannel_12_bits_vs;
  wire               _maskedWrite_readChannel_12_bits_offset;
  wire               _maskedWrite_readChannel_13_valid;
  wire [4:0]         _maskedWrite_readChannel_13_bits_vs;
  wire               _maskedWrite_readChannel_13_bits_offset;
  wire               _maskedWrite_readChannel_14_valid;
  wire [4:0]         _maskedWrite_readChannel_14_bits_vs;
  wire               _maskedWrite_readChannel_14_bits_offset;
  wire               _maskedWrite_readChannel_15_valid;
  wire [4:0]         _maskedWrite_readChannel_15_bits_vs;
  wire               _maskedWrite_readChannel_15_bits_offset;
  wire               _maskedWrite_readChannel_16_valid;
  wire [4:0]         _maskedWrite_readChannel_16_bits_vs;
  wire               _maskedWrite_readChannel_16_bits_offset;
  wire               _maskedWrite_readChannel_17_valid;
  wire [4:0]         _maskedWrite_readChannel_17_bits_vs;
  wire               _maskedWrite_readChannel_17_bits_offset;
  wire               _maskedWrite_readChannel_18_valid;
  wire [4:0]         _maskedWrite_readChannel_18_bits_vs;
  wire               _maskedWrite_readChannel_18_bits_offset;
  wire               _maskedWrite_readChannel_19_valid;
  wire [4:0]         _maskedWrite_readChannel_19_bits_vs;
  wire               _maskedWrite_readChannel_19_bits_offset;
  wire               _maskedWrite_readChannel_20_valid;
  wire [4:0]         _maskedWrite_readChannel_20_bits_vs;
  wire               _maskedWrite_readChannel_20_bits_offset;
  wire               _maskedWrite_readChannel_21_valid;
  wire [4:0]         _maskedWrite_readChannel_21_bits_vs;
  wire               _maskedWrite_readChannel_21_bits_offset;
  wire               _maskedWrite_readChannel_22_valid;
  wire [4:0]         _maskedWrite_readChannel_22_bits_vs;
  wire               _maskedWrite_readChannel_22_bits_offset;
  wire               _maskedWrite_readChannel_23_valid;
  wire [4:0]         _maskedWrite_readChannel_23_bits_vs;
  wire               _maskedWrite_readChannel_23_bits_offset;
  wire               _maskedWrite_readChannel_24_valid;
  wire [4:0]         _maskedWrite_readChannel_24_bits_vs;
  wire               _maskedWrite_readChannel_24_bits_offset;
  wire               _maskedWrite_readChannel_25_valid;
  wire [4:0]         _maskedWrite_readChannel_25_bits_vs;
  wire               _maskedWrite_readChannel_25_bits_offset;
  wire               _maskedWrite_readChannel_26_valid;
  wire [4:0]         _maskedWrite_readChannel_26_bits_vs;
  wire               _maskedWrite_readChannel_26_bits_offset;
  wire               _maskedWrite_readChannel_27_valid;
  wire [4:0]         _maskedWrite_readChannel_27_bits_vs;
  wire               _maskedWrite_readChannel_27_bits_offset;
  wire               _maskedWrite_readChannel_28_valid;
  wire [4:0]         _maskedWrite_readChannel_28_bits_vs;
  wire               _maskedWrite_readChannel_28_bits_offset;
  wire               _maskedWrite_readChannel_29_valid;
  wire [4:0]         _maskedWrite_readChannel_29_bits_vs;
  wire               _maskedWrite_readChannel_29_bits_offset;
  wire               _maskedWrite_readChannel_30_valid;
  wire [4:0]         _maskedWrite_readChannel_30_bits_vs;
  wire               _maskedWrite_readChannel_30_bits_offset;
  wire               _maskedWrite_readChannel_31_valid;
  wire [4:0]         _maskedWrite_readChannel_31_bits_vs;
  wire               _maskedWrite_readChannel_31_bits_offset;
  wire               _maskedWrite_stageClear;
  wire               writeQueue_31_almostFull;
  wire               writeQueue_31_almostEmpty;
  wire               writeQueue_30_almostFull;
  wire               writeQueue_30_almostEmpty;
  wire               writeQueue_29_almostFull;
  wire               writeQueue_29_almostEmpty;
  wire               writeQueue_28_almostFull;
  wire               writeQueue_28_almostEmpty;
  wire               writeQueue_27_almostFull;
  wire               writeQueue_27_almostEmpty;
  wire               writeQueue_26_almostFull;
  wire               writeQueue_26_almostEmpty;
  wire               writeQueue_25_almostFull;
  wire               writeQueue_25_almostEmpty;
  wire               writeQueue_24_almostFull;
  wire               writeQueue_24_almostEmpty;
  wire               writeQueue_23_almostFull;
  wire               writeQueue_23_almostEmpty;
  wire               writeQueue_22_almostFull;
  wire               writeQueue_22_almostEmpty;
  wire               writeQueue_21_almostFull;
  wire               writeQueue_21_almostEmpty;
  wire               writeQueue_20_almostFull;
  wire               writeQueue_20_almostEmpty;
  wire               writeQueue_19_almostFull;
  wire               writeQueue_19_almostEmpty;
  wire               writeQueue_18_almostFull;
  wire               writeQueue_18_almostEmpty;
  wire               writeQueue_17_almostFull;
  wire               writeQueue_17_almostEmpty;
  wire               writeQueue_16_almostFull;
  wire               writeQueue_16_almostEmpty;
  wire               writeQueue_15_almostFull;
  wire               writeQueue_15_almostEmpty;
  wire               writeQueue_14_almostFull;
  wire               writeQueue_14_almostEmpty;
  wire               writeQueue_13_almostFull;
  wire               writeQueue_13_almostEmpty;
  wire               writeQueue_12_almostFull;
  wire               writeQueue_12_almostEmpty;
  wire               writeQueue_11_almostFull;
  wire               writeQueue_11_almostEmpty;
  wire               writeQueue_10_almostFull;
  wire               writeQueue_10_almostEmpty;
  wire               writeQueue_9_almostFull;
  wire               writeQueue_9_almostEmpty;
  wire               writeQueue_8_almostFull;
  wire               writeQueue_8_almostEmpty;
  wire               writeQueue_7_almostFull;
  wire               writeQueue_7_almostEmpty;
  wire               writeQueue_6_almostFull;
  wire               writeQueue_6_almostEmpty;
  wire               writeQueue_5_almostFull;
  wire               writeQueue_5_almostEmpty;
  wire               writeQueue_4_almostFull;
  wire               writeQueue_4_almostEmpty;
  wire               writeQueue_3_almostFull;
  wire               writeQueue_3_almostEmpty;
  wire               writeQueue_2_almostFull;
  wire               writeQueue_2_almostEmpty;
  wire               writeQueue_1_almostFull;
  wire               writeQueue_1_almostEmpty;
  wire               writeQueue_0_almostFull;
  wire               writeQueue_0_almostEmpty;
  wire               readData_readDataQueue_31_almostFull;
  wire               readData_readDataQueue_31_almostEmpty;
  wire               readData_readDataQueue_30_almostFull;
  wire               readData_readDataQueue_30_almostEmpty;
  wire               readData_readDataQueue_29_almostFull;
  wire               readData_readDataQueue_29_almostEmpty;
  wire               readData_readDataQueue_28_almostFull;
  wire               readData_readDataQueue_28_almostEmpty;
  wire               readData_readDataQueue_27_almostFull;
  wire               readData_readDataQueue_27_almostEmpty;
  wire               readData_readDataQueue_26_almostFull;
  wire               readData_readDataQueue_26_almostEmpty;
  wire               readData_readDataQueue_25_almostFull;
  wire               readData_readDataQueue_25_almostEmpty;
  wire               readData_readDataQueue_24_almostFull;
  wire               readData_readDataQueue_24_almostEmpty;
  wire               readData_readDataQueue_23_almostFull;
  wire               readData_readDataQueue_23_almostEmpty;
  wire               readData_readDataQueue_22_almostFull;
  wire               readData_readDataQueue_22_almostEmpty;
  wire               readData_readDataQueue_21_almostFull;
  wire               readData_readDataQueue_21_almostEmpty;
  wire               readData_readDataQueue_20_almostFull;
  wire               readData_readDataQueue_20_almostEmpty;
  wire               readData_readDataQueue_19_almostFull;
  wire               readData_readDataQueue_19_almostEmpty;
  wire               readData_readDataQueue_18_almostFull;
  wire               readData_readDataQueue_18_almostEmpty;
  wire               readData_readDataQueue_17_almostFull;
  wire               readData_readDataQueue_17_almostEmpty;
  wire               readData_readDataQueue_16_almostFull;
  wire               readData_readDataQueue_16_almostEmpty;
  wire               readData_readDataQueue_15_almostFull;
  wire               readData_readDataQueue_15_almostEmpty;
  wire               readData_readDataQueue_14_almostFull;
  wire               readData_readDataQueue_14_almostEmpty;
  wire               readData_readDataQueue_13_almostFull;
  wire               readData_readDataQueue_13_almostEmpty;
  wire               readData_readDataQueue_12_almostFull;
  wire               readData_readDataQueue_12_almostEmpty;
  wire               readData_readDataQueue_11_almostFull;
  wire               readData_readDataQueue_11_almostEmpty;
  wire               readData_readDataQueue_10_almostFull;
  wire               readData_readDataQueue_10_almostEmpty;
  wire               readData_readDataQueue_9_almostFull;
  wire               readData_readDataQueue_9_almostEmpty;
  wire               readData_readDataQueue_8_almostFull;
  wire               readData_readDataQueue_8_almostEmpty;
  wire               readData_readDataQueue_7_almostFull;
  wire               readData_readDataQueue_7_almostEmpty;
  wire               readData_readDataQueue_6_almostFull;
  wire               readData_readDataQueue_6_almostEmpty;
  wire               readData_readDataQueue_5_almostFull;
  wire               readData_readDataQueue_5_almostEmpty;
  wire               readData_readDataQueue_4_almostFull;
  wire               readData_readDataQueue_4_almostEmpty;
  wire               readData_readDataQueue_3_almostFull;
  wire               readData_readDataQueue_3_almostEmpty;
  wire               readData_readDataQueue_2_almostFull;
  wire               readData_readDataQueue_2_almostEmpty;
  wire               readData_readDataQueue_1_almostFull;
  wire               readData_readDataQueue_1_almostEmpty;
  wire               readData_readDataQueue_almostFull;
  wire               readData_readDataQueue_almostEmpty;
  wire               readMessageQueue_31_almostFull;
  wire               readMessageQueue_31_almostEmpty;
  wire               readMessageQueue_30_almostFull;
  wire               readMessageQueue_30_almostEmpty;
  wire               readMessageQueue_29_almostFull;
  wire               readMessageQueue_29_almostEmpty;
  wire               readMessageQueue_28_almostFull;
  wire               readMessageQueue_28_almostEmpty;
  wire               readMessageQueue_27_almostFull;
  wire               readMessageQueue_27_almostEmpty;
  wire               readMessageQueue_26_almostFull;
  wire               readMessageQueue_26_almostEmpty;
  wire               readMessageQueue_25_almostFull;
  wire               readMessageQueue_25_almostEmpty;
  wire               readMessageQueue_24_almostFull;
  wire               readMessageQueue_24_almostEmpty;
  wire               readMessageQueue_23_almostFull;
  wire               readMessageQueue_23_almostEmpty;
  wire               readMessageQueue_22_almostFull;
  wire               readMessageQueue_22_almostEmpty;
  wire               readMessageQueue_21_almostFull;
  wire               readMessageQueue_21_almostEmpty;
  wire               readMessageQueue_20_almostFull;
  wire               readMessageQueue_20_almostEmpty;
  wire               readMessageQueue_19_almostFull;
  wire               readMessageQueue_19_almostEmpty;
  wire               readMessageQueue_18_almostFull;
  wire               readMessageQueue_18_almostEmpty;
  wire               readMessageQueue_17_almostFull;
  wire               readMessageQueue_17_almostEmpty;
  wire               readMessageQueue_16_almostFull;
  wire               readMessageQueue_16_almostEmpty;
  wire               readMessageQueue_15_almostFull;
  wire               readMessageQueue_15_almostEmpty;
  wire               readMessageQueue_14_almostFull;
  wire               readMessageQueue_14_almostEmpty;
  wire               readMessageQueue_13_almostFull;
  wire               readMessageQueue_13_almostEmpty;
  wire               readMessageQueue_12_almostFull;
  wire               readMessageQueue_12_almostEmpty;
  wire               readMessageQueue_11_almostFull;
  wire               readMessageQueue_11_almostEmpty;
  wire               readMessageQueue_10_almostFull;
  wire               readMessageQueue_10_almostEmpty;
  wire               readMessageQueue_9_almostFull;
  wire               readMessageQueue_9_almostEmpty;
  wire               readMessageQueue_8_almostFull;
  wire               readMessageQueue_8_almostEmpty;
  wire               readMessageQueue_7_almostFull;
  wire               readMessageQueue_7_almostEmpty;
  wire               readMessageQueue_6_almostFull;
  wire               readMessageQueue_6_almostEmpty;
  wire               readMessageQueue_5_almostFull;
  wire               readMessageQueue_5_almostEmpty;
  wire               readMessageQueue_4_almostFull;
  wire               readMessageQueue_4_almostEmpty;
  wire               readMessageQueue_3_almostFull;
  wire               readMessageQueue_3_almostEmpty;
  wire               readMessageQueue_2_almostFull;
  wire               readMessageQueue_2_almostEmpty;
  wire               readMessageQueue_1_almostFull;
  wire               readMessageQueue_1_almostEmpty;
  wire               readMessageQueue_almostFull;
  wire               readMessageQueue_almostEmpty;
  wire               reorderQueueVec_31_almostFull;
  wire               reorderQueueVec_31_almostEmpty;
  wire               reorderQueueVec_30_almostFull;
  wire               reorderQueueVec_30_almostEmpty;
  wire               reorderQueueVec_29_almostFull;
  wire               reorderQueueVec_29_almostEmpty;
  wire               reorderQueueVec_28_almostFull;
  wire               reorderQueueVec_28_almostEmpty;
  wire               reorderQueueVec_27_almostFull;
  wire               reorderQueueVec_27_almostEmpty;
  wire               reorderQueueVec_26_almostFull;
  wire               reorderQueueVec_26_almostEmpty;
  wire               reorderQueueVec_25_almostFull;
  wire               reorderQueueVec_25_almostEmpty;
  wire               reorderQueueVec_24_almostFull;
  wire               reorderQueueVec_24_almostEmpty;
  wire               reorderQueueVec_23_almostFull;
  wire               reorderQueueVec_23_almostEmpty;
  wire               reorderQueueVec_22_almostFull;
  wire               reorderQueueVec_22_almostEmpty;
  wire               reorderQueueVec_21_almostFull;
  wire               reorderQueueVec_21_almostEmpty;
  wire               reorderQueueVec_20_almostFull;
  wire               reorderQueueVec_20_almostEmpty;
  wire               reorderQueueVec_19_almostFull;
  wire               reorderQueueVec_19_almostEmpty;
  wire               reorderQueueVec_18_almostFull;
  wire               reorderQueueVec_18_almostEmpty;
  wire               reorderQueueVec_17_almostFull;
  wire               reorderQueueVec_17_almostEmpty;
  wire               reorderQueueVec_16_almostFull;
  wire               reorderQueueVec_16_almostEmpty;
  wire               reorderQueueVec_15_almostFull;
  wire               reorderQueueVec_15_almostEmpty;
  wire               reorderQueueVec_14_almostFull;
  wire               reorderQueueVec_14_almostEmpty;
  wire               reorderQueueVec_13_almostFull;
  wire               reorderQueueVec_13_almostEmpty;
  wire               reorderQueueVec_12_almostFull;
  wire               reorderQueueVec_12_almostEmpty;
  wire               reorderQueueVec_11_almostFull;
  wire               reorderQueueVec_11_almostEmpty;
  wire               reorderQueueVec_10_almostFull;
  wire               reorderQueueVec_10_almostEmpty;
  wire               reorderQueueVec_9_almostFull;
  wire               reorderQueueVec_9_almostEmpty;
  wire               reorderQueueVec_8_almostFull;
  wire               reorderQueueVec_8_almostEmpty;
  wire               reorderQueueVec_7_almostFull;
  wire               reorderQueueVec_7_almostEmpty;
  wire               reorderQueueVec_6_almostFull;
  wire               reorderQueueVec_6_almostEmpty;
  wire               reorderQueueVec_5_almostFull;
  wire               reorderQueueVec_5_almostEmpty;
  wire               reorderQueueVec_4_almostFull;
  wire               reorderQueueVec_4_almostEmpty;
  wire               reorderQueueVec_3_almostFull;
  wire               reorderQueueVec_3_almostEmpty;
  wire               reorderQueueVec_2_almostFull;
  wire               reorderQueueVec_2_almostEmpty;
  wire               reorderQueueVec_1_almostFull;
  wire               reorderQueueVec_1_almostEmpty;
  wire               reorderQueueVec_0_almostFull;
  wire               reorderQueueVec_0_almostEmpty;
  wire               compressUnitResultQueue_almostFull;
  wire               compressUnitResultQueue_almostEmpty;
  wire               readWaitQueue_almostFull;
  wire               readWaitQueue_almostEmpty;
  wire               accessCountQueue_almostFull;
  wire               accessCountQueue_almostEmpty;
  wire               exeRequestQueue_31_almostFull;
  wire               exeRequestQueue_31_almostEmpty;
  wire               exeRequestQueue_30_almostFull;
  wire               exeRequestQueue_30_almostEmpty;
  wire               exeRequestQueue_29_almostFull;
  wire               exeRequestQueue_29_almostEmpty;
  wire               exeRequestQueue_28_almostFull;
  wire               exeRequestQueue_28_almostEmpty;
  wire               exeRequestQueue_27_almostFull;
  wire               exeRequestQueue_27_almostEmpty;
  wire               exeRequestQueue_26_almostFull;
  wire               exeRequestQueue_26_almostEmpty;
  wire               exeRequestQueue_25_almostFull;
  wire               exeRequestQueue_25_almostEmpty;
  wire               exeRequestQueue_24_almostFull;
  wire               exeRequestQueue_24_almostEmpty;
  wire               exeRequestQueue_23_almostFull;
  wire               exeRequestQueue_23_almostEmpty;
  wire               exeRequestQueue_22_almostFull;
  wire               exeRequestQueue_22_almostEmpty;
  wire               exeRequestQueue_21_almostFull;
  wire               exeRequestQueue_21_almostEmpty;
  wire               exeRequestQueue_20_almostFull;
  wire               exeRequestQueue_20_almostEmpty;
  wire               exeRequestQueue_19_almostFull;
  wire               exeRequestQueue_19_almostEmpty;
  wire               exeRequestQueue_18_almostFull;
  wire               exeRequestQueue_18_almostEmpty;
  wire               exeRequestQueue_17_almostFull;
  wire               exeRequestQueue_17_almostEmpty;
  wire               exeRequestQueue_16_almostFull;
  wire               exeRequestQueue_16_almostEmpty;
  wire               exeRequestQueue_15_almostFull;
  wire               exeRequestQueue_15_almostEmpty;
  wire               exeRequestQueue_14_almostFull;
  wire               exeRequestQueue_14_almostEmpty;
  wire               exeRequestQueue_13_almostFull;
  wire               exeRequestQueue_13_almostEmpty;
  wire               exeRequestQueue_12_almostFull;
  wire               exeRequestQueue_12_almostEmpty;
  wire               exeRequestQueue_11_almostFull;
  wire               exeRequestQueue_11_almostEmpty;
  wire               exeRequestQueue_10_almostFull;
  wire               exeRequestQueue_10_almostEmpty;
  wire               exeRequestQueue_9_almostFull;
  wire               exeRequestQueue_9_almostEmpty;
  wire               exeRequestQueue_8_almostFull;
  wire               exeRequestQueue_8_almostEmpty;
  wire               exeRequestQueue_7_almostFull;
  wire               exeRequestQueue_7_almostEmpty;
  wire               exeRequestQueue_6_almostFull;
  wire               exeRequestQueue_6_almostEmpty;
  wire               exeRequestQueue_5_almostFull;
  wire               exeRequestQueue_5_almostEmpty;
  wire               exeRequestQueue_4_almostFull;
  wire               exeRequestQueue_4_almostEmpty;
  wire               exeRequestQueue_3_almostFull;
  wire               exeRequestQueue_3_almostEmpty;
  wire               exeRequestQueue_2_almostFull;
  wire               exeRequestQueue_2_almostEmpty;
  wire               exeRequestQueue_1_almostFull;
  wire               exeRequestQueue_1_almostEmpty;
  wire               exeRequestQueue_0_almostFull;
  wire               exeRequestQueue_0_almostEmpty;
  wire [31:0]        reorderQueueVec_31_deq_bits_data;
  wire [31:0]        reorderQueueVec_30_deq_bits_data;
  wire [31:0]        reorderQueueVec_29_deq_bits_data;
  wire [31:0]        reorderQueueVec_28_deq_bits_data;
  wire [31:0]        reorderQueueVec_27_deq_bits_data;
  wire [31:0]        reorderQueueVec_26_deq_bits_data;
  wire [31:0]        reorderQueueVec_25_deq_bits_data;
  wire [31:0]        reorderQueueVec_24_deq_bits_data;
  wire [31:0]        reorderQueueVec_23_deq_bits_data;
  wire [31:0]        reorderQueueVec_22_deq_bits_data;
  wire [31:0]        reorderQueueVec_21_deq_bits_data;
  wire [31:0]        reorderQueueVec_20_deq_bits_data;
  wire [31:0]        reorderQueueVec_19_deq_bits_data;
  wire [31:0]        reorderQueueVec_18_deq_bits_data;
  wire [31:0]        reorderQueueVec_17_deq_bits_data;
  wire [31:0]        reorderQueueVec_16_deq_bits_data;
  wire [31:0]        reorderQueueVec_15_deq_bits_data;
  wire [31:0]        reorderQueueVec_14_deq_bits_data;
  wire [31:0]        reorderQueueVec_13_deq_bits_data;
  wire [31:0]        reorderQueueVec_12_deq_bits_data;
  wire [31:0]        reorderQueueVec_11_deq_bits_data;
  wire [31:0]        reorderQueueVec_10_deq_bits_data;
  wire [31:0]        reorderQueueVec_9_deq_bits_data;
  wire [31:0]        reorderQueueVec_8_deq_bits_data;
  wire [31:0]        reorderQueueVec_7_deq_bits_data;
  wire [31:0]        reorderQueueVec_6_deq_bits_data;
  wire [31:0]        reorderQueueVec_5_deq_bits_data;
  wire [31:0]        reorderQueueVec_4_deq_bits_data;
  wire [31:0]        reorderQueueVec_3_deq_bits_data;
  wire [31:0]        reorderQueueVec_2_deq_bits_data;
  wire [31:0]        reorderQueueVec_1_deq_bits_data;
  wire [31:0]        reorderQueueVec_0_deq_bits_data;
  wire [5:0]         accessCountEnq_31;
  wire [5:0]         accessCountEnq_30;
  wire [5:0]         accessCountEnq_29;
  wire [5:0]         accessCountEnq_28;
  wire [5:0]         accessCountEnq_27;
  wire [5:0]         accessCountEnq_26;
  wire [5:0]         accessCountEnq_25;
  wire [5:0]         accessCountEnq_24;
  wire [5:0]         accessCountEnq_23;
  wire [5:0]         accessCountEnq_22;
  wire [5:0]         accessCountEnq_21;
  wire [5:0]         accessCountEnq_20;
  wire [5:0]         accessCountEnq_19;
  wire [5:0]         accessCountEnq_18;
  wire [5:0]         accessCountEnq_17;
  wire [5:0]         accessCountEnq_16;
  wire [5:0]         accessCountEnq_15;
  wire [5:0]         accessCountEnq_14;
  wire [5:0]         accessCountEnq_13;
  wire [5:0]         accessCountEnq_12;
  wire [5:0]         accessCountEnq_11;
  wire [5:0]         accessCountEnq_10;
  wire [5:0]         accessCountEnq_9;
  wire [5:0]         accessCountEnq_8;
  wire [5:0]         accessCountEnq_7;
  wire [5:0]         accessCountEnq_6;
  wire [5:0]         accessCountEnq_5;
  wire [5:0]         accessCountEnq_4;
  wire [5:0]         accessCountEnq_3;
  wire [5:0]         accessCountEnq_2;
  wire [5:0]         accessCountEnq_1;
  wire [5:0]         accessCountEnq_0;
  wire               exeResp_0_ready_0 = exeResp_0_ready;
  wire               exeResp_1_ready_0 = exeResp_1_ready;
  wire               exeResp_2_ready_0 = exeResp_2_ready;
  wire               exeResp_3_ready_0 = exeResp_3_ready;
  wire               exeResp_4_ready_0 = exeResp_4_ready;
  wire               exeResp_5_ready_0 = exeResp_5_ready;
  wire               exeResp_6_ready_0 = exeResp_6_ready;
  wire               exeResp_7_ready_0 = exeResp_7_ready;
  wire               exeResp_8_ready_0 = exeResp_8_ready;
  wire               exeResp_9_ready_0 = exeResp_9_ready;
  wire               exeResp_10_ready_0 = exeResp_10_ready;
  wire               exeResp_11_ready_0 = exeResp_11_ready;
  wire               exeResp_12_ready_0 = exeResp_12_ready;
  wire               exeResp_13_ready_0 = exeResp_13_ready;
  wire               exeResp_14_ready_0 = exeResp_14_ready;
  wire               exeResp_15_ready_0 = exeResp_15_ready;
  wire               exeResp_16_ready_0 = exeResp_16_ready;
  wire               exeResp_17_ready_0 = exeResp_17_ready;
  wire               exeResp_18_ready_0 = exeResp_18_ready;
  wire               exeResp_19_ready_0 = exeResp_19_ready;
  wire               exeResp_20_ready_0 = exeResp_20_ready;
  wire               exeResp_21_ready_0 = exeResp_21_ready;
  wire               exeResp_22_ready_0 = exeResp_22_ready;
  wire               exeResp_23_ready_0 = exeResp_23_ready;
  wire               exeResp_24_ready_0 = exeResp_24_ready;
  wire               exeResp_25_ready_0 = exeResp_25_ready;
  wire               exeResp_26_ready_0 = exeResp_26_ready;
  wire               exeResp_27_ready_0 = exeResp_27_ready;
  wire               exeResp_28_ready_0 = exeResp_28_ready;
  wire               exeResp_29_ready_0 = exeResp_29_ready;
  wire               exeResp_30_ready_0 = exeResp_30_ready;
  wire               exeResp_31_ready_0 = exeResp_31_ready;
  wire               readChannel_0_ready_0 = readChannel_0_ready;
  wire               readChannel_1_ready_0 = readChannel_1_ready;
  wire               readChannel_2_ready_0 = readChannel_2_ready;
  wire               readChannel_3_ready_0 = readChannel_3_ready;
  wire               readChannel_4_ready_0 = readChannel_4_ready;
  wire               readChannel_5_ready_0 = readChannel_5_ready;
  wire               readChannel_6_ready_0 = readChannel_6_ready;
  wire               readChannel_7_ready_0 = readChannel_7_ready;
  wire               readChannel_8_ready_0 = readChannel_8_ready;
  wire               readChannel_9_ready_0 = readChannel_9_ready;
  wire               readChannel_10_ready_0 = readChannel_10_ready;
  wire               readChannel_11_ready_0 = readChannel_11_ready;
  wire               readChannel_12_ready_0 = readChannel_12_ready;
  wire               readChannel_13_ready_0 = readChannel_13_ready;
  wire               readChannel_14_ready_0 = readChannel_14_ready;
  wire               readChannel_15_ready_0 = readChannel_15_ready;
  wire               readChannel_16_ready_0 = readChannel_16_ready;
  wire               readChannel_17_ready_0 = readChannel_17_ready;
  wire               readChannel_18_ready_0 = readChannel_18_ready;
  wire               readChannel_19_ready_0 = readChannel_19_ready;
  wire               readChannel_20_ready_0 = readChannel_20_ready;
  wire               readChannel_21_ready_0 = readChannel_21_ready;
  wire               readChannel_22_ready_0 = readChannel_22_ready;
  wire               readChannel_23_ready_0 = readChannel_23_ready;
  wire               readChannel_24_ready_0 = readChannel_24_ready;
  wire               readChannel_25_ready_0 = readChannel_25_ready;
  wire               readChannel_26_ready_0 = readChannel_26_ready;
  wire               readChannel_27_ready_0 = readChannel_27_ready;
  wire               readChannel_28_ready_0 = readChannel_28_ready;
  wire               readChannel_29_ready_0 = readChannel_29_ready;
  wire               readChannel_30_ready_0 = readChannel_30_ready;
  wire               readChannel_31_ready_0 = readChannel_31_ready;
  wire               gatherData_ready_0 = gatherData_ready;
  wire               exeRequestQueue_0_enq_valid = exeReq_0_valid;
  wire [31:0]        exeRequestQueue_0_enq_bits_source1 = exeReq_0_bits_source1;
  wire [31:0]        exeRequestQueue_0_enq_bits_source2 = exeReq_0_bits_source2;
  wire [2:0]         exeRequestQueue_0_enq_bits_index = exeReq_0_bits_index;
  wire               exeRequestQueue_0_enq_bits_ffo = exeReq_0_bits_ffo;
  wire               exeRequestQueue_1_enq_valid = exeReq_1_valid;
  wire [31:0]        exeRequestQueue_1_enq_bits_source1 = exeReq_1_bits_source1;
  wire [31:0]        exeRequestQueue_1_enq_bits_source2 = exeReq_1_bits_source2;
  wire [2:0]         exeRequestQueue_1_enq_bits_index = exeReq_1_bits_index;
  wire               exeRequestQueue_1_enq_bits_ffo = exeReq_1_bits_ffo;
  wire               exeRequestQueue_2_enq_valid = exeReq_2_valid;
  wire [31:0]        exeRequestQueue_2_enq_bits_source1 = exeReq_2_bits_source1;
  wire [31:0]        exeRequestQueue_2_enq_bits_source2 = exeReq_2_bits_source2;
  wire [2:0]         exeRequestQueue_2_enq_bits_index = exeReq_2_bits_index;
  wire               exeRequestQueue_2_enq_bits_ffo = exeReq_2_bits_ffo;
  wire               exeRequestQueue_3_enq_valid = exeReq_3_valid;
  wire [31:0]        exeRequestQueue_3_enq_bits_source1 = exeReq_3_bits_source1;
  wire [31:0]        exeRequestQueue_3_enq_bits_source2 = exeReq_3_bits_source2;
  wire [2:0]         exeRequestQueue_3_enq_bits_index = exeReq_3_bits_index;
  wire               exeRequestQueue_3_enq_bits_ffo = exeReq_3_bits_ffo;
  wire               exeRequestQueue_4_enq_valid = exeReq_4_valid;
  wire [31:0]        exeRequestQueue_4_enq_bits_source1 = exeReq_4_bits_source1;
  wire [31:0]        exeRequestQueue_4_enq_bits_source2 = exeReq_4_bits_source2;
  wire [2:0]         exeRequestQueue_4_enq_bits_index = exeReq_4_bits_index;
  wire               exeRequestQueue_4_enq_bits_ffo = exeReq_4_bits_ffo;
  wire               exeRequestQueue_5_enq_valid = exeReq_5_valid;
  wire [31:0]        exeRequestQueue_5_enq_bits_source1 = exeReq_5_bits_source1;
  wire [31:0]        exeRequestQueue_5_enq_bits_source2 = exeReq_5_bits_source2;
  wire [2:0]         exeRequestQueue_5_enq_bits_index = exeReq_5_bits_index;
  wire               exeRequestQueue_5_enq_bits_ffo = exeReq_5_bits_ffo;
  wire               exeRequestQueue_6_enq_valid = exeReq_6_valid;
  wire [31:0]        exeRequestQueue_6_enq_bits_source1 = exeReq_6_bits_source1;
  wire [31:0]        exeRequestQueue_6_enq_bits_source2 = exeReq_6_bits_source2;
  wire [2:0]         exeRequestQueue_6_enq_bits_index = exeReq_6_bits_index;
  wire               exeRequestQueue_6_enq_bits_ffo = exeReq_6_bits_ffo;
  wire               exeRequestQueue_7_enq_valid = exeReq_7_valid;
  wire [31:0]        exeRequestQueue_7_enq_bits_source1 = exeReq_7_bits_source1;
  wire [31:0]        exeRequestQueue_7_enq_bits_source2 = exeReq_7_bits_source2;
  wire [2:0]         exeRequestQueue_7_enq_bits_index = exeReq_7_bits_index;
  wire               exeRequestQueue_7_enq_bits_ffo = exeReq_7_bits_ffo;
  wire               exeRequestQueue_8_enq_valid = exeReq_8_valid;
  wire [31:0]        exeRequestQueue_8_enq_bits_source1 = exeReq_8_bits_source1;
  wire [31:0]        exeRequestQueue_8_enq_bits_source2 = exeReq_8_bits_source2;
  wire [2:0]         exeRequestQueue_8_enq_bits_index = exeReq_8_bits_index;
  wire               exeRequestQueue_8_enq_bits_ffo = exeReq_8_bits_ffo;
  wire               exeRequestQueue_9_enq_valid = exeReq_9_valid;
  wire [31:0]        exeRequestQueue_9_enq_bits_source1 = exeReq_9_bits_source1;
  wire [31:0]        exeRequestQueue_9_enq_bits_source2 = exeReq_9_bits_source2;
  wire [2:0]         exeRequestQueue_9_enq_bits_index = exeReq_9_bits_index;
  wire               exeRequestQueue_9_enq_bits_ffo = exeReq_9_bits_ffo;
  wire               exeRequestQueue_10_enq_valid = exeReq_10_valid;
  wire [31:0]        exeRequestQueue_10_enq_bits_source1 = exeReq_10_bits_source1;
  wire [31:0]        exeRequestQueue_10_enq_bits_source2 = exeReq_10_bits_source2;
  wire [2:0]         exeRequestQueue_10_enq_bits_index = exeReq_10_bits_index;
  wire               exeRequestQueue_10_enq_bits_ffo = exeReq_10_bits_ffo;
  wire               exeRequestQueue_11_enq_valid = exeReq_11_valid;
  wire [31:0]        exeRequestQueue_11_enq_bits_source1 = exeReq_11_bits_source1;
  wire [31:0]        exeRequestQueue_11_enq_bits_source2 = exeReq_11_bits_source2;
  wire [2:0]         exeRequestQueue_11_enq_bits_index = exeReq_11_bits_index;
  wire               exeRequestQueue_11_enq_bits_ffo = exeReq_11_bits_ffo;
  wire               exeRequestQueue_12_enq_valid = exeReq_12_valid;
  wire [31:0]        exeRequestQueue_12_enq_bits_source1 = exeReq_12_bits_source1;
  wire [31:0]        exeRequestQueue_12_enq_bits_source2 = exeReq_12_bits_source2;
  wire [2:0]         exeRequestQueue_12_enq_bits_index = exeReq_12_bits_index;
  wire               exeRequestQueue_12_enq_bits_ffo = exeReq_12_bits_ffo;
  wire               exeRequestQueue_13_enq_valid = exeReq_13_valid;
  wire [31:0]        exeRequestQueue_13_enq_bits_source1 = exeReq_13_bits_source1;
  wire [31:0]        exeRequestQueue_13_enq_bits_source2 = exeReq_13_bits_source2;
  wire [2:0]         exeRequestQueue_13_enq_bits_index = exeReq_13_bits_index;
  wire               exeRequestQueue_13_enq_bits_ffo = exeReq_13_bits_ffo;
  wire               exeRequestQueue_14_enq_valid = exeReq_14_valid;
  wire [31:0]        exeRequestQueue_14_enq_bits_source1 = exeReq_14_bits_source1;
  wire [31:0]        exeRequestQueue_14_enq_bits_source2 = exeReq_14_bits_source2;
  wire [2:0]         exeRequestQueue_14_enq_bits_index = exeReq_14_bits_index;
  wire               exeRequestQueue_14_enq_bits_ffo = exeReq_14_bits_ffo;
  wire               exeRequestQueue_15_enq_valid = exeReq_15_valid;
  wire [31:0]        exeRequestQueue_15_enq_bits_source1 = exeReq_15_bits_source1;
  wire [31:0]        exeRequestQueue_15_enq_bits_source2 = exeReq_15_bits_source2;
  wire [2:0]         exeRequestQueue_15_enq_bits_index = exeReq_15_bits_index;
  wire               exeRequestQueue_15_enq_bits_ffo = exeReq_15_bits_ffo;
  wire               exeRequestQueue_16_enq_valid = exeReq_16_valid;
  wire [31:0]        exeRequestQueue_16_enq_bits_source1 = exeReq_16_bits_source1;
  wire [31:0]        exeRequestQueue_16_enq_bits_source2 = exeReq_16_bits_source2;
  wire [2:0]         exeRequestQueue_16_enq_bits_index = exeReq_16_bits_index;
  wire               exeRequestQueue_16_enq_bits_ffo = exeReq_16_bits_ffo;
  wire               exeRequestQueue_17_enq_valid = exeReq_17_valid;
  wire [31:0]        exeRequestQueue_17_enq_bits_source1 = exeReq_17_bits_source1;
  wire [31:0]        exeRequestQueue_17_enq_bits_source2 = exeReq_17_bits_source2;
  wire [2:0]         exeRequestQueue_17_enq_bits_index = exeReq_17_bits_index;
  wire               exeRequestQueue_17_enq_bits_ffo = exeReq_17_bits_ffo;
  wire               exeRequestQueue_18_enq_valid = exeReq_18_valid;
  wire [31:0]        exeRequestQueue_18_enq_bits_source1 = exeReq_18_bits_source1;
  wire [31:0]        exeRequestQueue_18_enq_bits_source2 = exeReq_18_bits_source2;
  wire [2:0]         exeRequestQueue_18_enq_bits_index = exeReq_18_bits_index;
  wire               exeRequestQueue_18_enq_bits_ffo = exeReq_18_bits_ffo;
  wire               exeRequestQueue_19_enq_valid = exeReq_19_valid;
  wire [31:0]        exeRequestQueue_19_enq_bits_source1 = exeReq_19_bits_source1;
  wire [31:0]        exeRequestQueue_19_enq_bits_source2 = exeReq_19_bits_source2;
  wire [2:0]         exeRequestQueue_19_enq_bits_index = exeReq_19_bits_index;
  wire               exeRequestQueue_19_enq_bits_ffo = exeReq_19_bits_ffo;
  wire               exeRequestQueue_20_enq_valid = exeReq_20_valid;
  wire [31:0]        exeRequestQueue_20_enq_bits_source1 = exeReq_20_bits_source1;
  wire [31:0]        exeRequestQueue_20_enq_bits_source2 = exeReq_20_bits_source2;
  wire [2:0]         exeRequestQueue_20_enq_bits_index = exeReq_20_bits_index;
  wire               exeRequestQueue_20_enq_bits_ffo = exeReq_20_bits_ffo;
  wire               exeRequestQueue_21_enq_valid = exeReq_21_valid;
  wire [31:0]        exeRequestQueue_21_enq_bits_source1 = exeReq_21_bits_source1;
  wire [31:0]        exeRequestQueue_21_enq_bits_source2 = exeReq_21_bits_source2;
  wire [2:0]         exeRequestQueue_21_enq_bits_index = exeReq_21_bits_index;
  wire               exeRequestQueue_21_enq_bits_ffo = exeReq_21_bits_ffo;
  wire               exeRequestQueue_22_enq_valid = exeReq_22_valid;
  wire [31:0]        exeRequestQueue_22_enq_bits_source1 = exeReq_22_bits_source1;
  wire [31:0]        exeRequestQueue_22_enq_bits_source2 = exeReq_22_bits_source2;
  wire [2:0]         exeRequestQueue_22_enq_bits_index = exeReq_22_bits_index;
  wire               exeRequestQueue_22_enq_bits_ffo = exeReq_22_bits_ffo;
  wire               exeRequestQueue_23_enq_valid = exeReq_23_valid;
  wire [31:0]        exeRequestQueue_23_enq_bits_source1 = exeReq_23_bits_source1;
  wire [31:0]        exeRequestQueue_23_enq_bits_source2 = exeReq_23_bits_source2;
  wire [2:0]         exeRequestQueue_23_enq_bits_index = exeReq_23_bits_index;
  wire               exeRequestQueue_23_enq_bits_ffo = exeReq_23_bits_ffo;
  wire               exeRequestQueue_24_enq_valid = exeReq_24_valid;
  wire [31:0]        exeRequestQueue_24_enq_bits_source1 = exeReq_24_bits_source1;
  wire [31:0]        exeRequestQueue_24_enq_bits_source2 = exeReq_24_bits_source2;
  wire [2:0]         exeRequestQueue_24_enq_bits_index = exeReq_24_bits_index;
  wire               exeRequestQueue_24_enq_bits_ffo = exeReq_24_bits_ffo;
  wire               exeRequestQueue_25_enq_valid = exeReq_25_valid;
  wire [31:0]        exeRequestQueue_25_enq_bits_source1 = exeReq_25_bits_source1;
  wire [31:0]        exeRequestQueue_25_enq_bits_source2 = exeReq_25_bits_source2;
  wire [2:0]         exeRequestQueue_25_enq_bits_index = exeReq_25_bits_index;
  wire               exeRequestQueue_25_enq_bits_ffo = exeReq_25_bits_ffo;
  wire               exeRequestQueue_26_enq_valid = exeReq_26_valid;
  wire [31:0]        exeRequestQueue_26_enq_bits_source1 = exeReq_26_bits_source1;
  wire [31:0]        exeRequestQueue_26_enq_bits_source2 = exeReq_26_bits_source2;
  wire [2:0]         exeRequestQueue_26_enq_bits_index = exeReq_26_bits_index;
  wire               exeRequestQueue_26_enq_bits_ffo = exeReq_26_bits_ffo;
  wire               exeRequestQueue_27_enq_valid = exeReq_27_valid;
  wire [31:0]        exeRequestQueue_27_enq_bits_source1 = exeReq_27_bits_source1;
  wire [31:0]        exeRequestQueue_27_enq_bits_source2 = exeReq_27_bits_source2;
  wire [2:0]         exeRequestQueue_27_enq_bits_index = exeReq_27_bits_index;
  wire               exeRequestQueue_27_enq_bits_ffo = exeReq_27_bits_ffo;
  wire               exeRequestQueue_28_enq_valid = exeReq_28_valid;
  wire [31:0]        exeRequestQueue_28_enq_bits_source1 = exeReq_28_bits_source1;
  wire [31:0]        exeRequestQueue_28_enq_bits_source2 = exeReq_28_bits_source2;
  wire [2:0]         exeRequestQueue_28_enq_bits_index = exeReq_28_bits_index;
  wire               exeRequestQueue_28_enq_bits_ffo = exeReq_28_bits_ffo;
  wire               exeRequestQueue_29_enq_valid = exeReq_29_valid;
  wire [31:0]        exeRequestQueue_29_enq_bits_source1 = exeReq_29_bits_source1;
  wire [31:0]        exeRequestQueue_29_enq_bits_source2 = exeReq_29_bits_source2;
  wire [2:0]         exeRequestQueue_29_enq_bits_index = exeReq_29_bits_index;
  wire               exeRequestQueue_29_enq_bits_ffo = exeReq_29_bits_ffo;
  wire               exeRequestQueue_30_enq_valid = exeReq_30_valid;
  wire [31:0]        exeRequestQueue_30_enq_bits_source1 = exeReq_30_bits_source1;
  wire [31:0]        exeRequestQueue_30_enq_bits_source2 = exeReq_30_bits_source2;
  wire [2:0]         exeRequestQueue_30_enq_bits_index = exeReq_30_bits_index;
  wire               exeRequestQueue_30_enq_bits_ffo = exeReq_30_bits_ffo;
  wire               exeRequestQueue_31_enq_valid = exeReq_31_valid;
  wire [31:0]        exeRequestQueue_31_enq_bits_source1 = exeReq_31_bits_source1;
  wire [31:0]        exeRequestQueue_31_enq_bits_source2 = exeReq_31_bits_source2;
  wire [2:0]         exeRequestQueue_31_enq_bits_index = exeReq_31_bits_index;
  wire               exeRequestQueue_31_enq_bits_ffo = exeReq_31_bits_ffo;
  wire               reorderQueueVec_0_enq_valid = readResult_0_valid;
  wire               reorderQueueVec_1_enq_valid = readResult_1_valid;
  wire               reorderQueueVec_2_enq_valid = readResult_2_valid;
  wire               reorderQueueVec_3_enq_valid = readResult_3_valid;
  wire               reorderQueueVec_4_enq_valid = readResult_4_valid;
  wire               reorderQueueVec_5_enq_valid = readResult_5_valid;
  wire               reorderQueueVec_6_enq_valid = readResult_6_valid;
  wire               reorderQueueVec_7_enq_valid = readResult_7_valid;
  wire               reorderQueueVec_8_enq_valid = readResult_8_valid;
  wire               reorderQueueVec_9_enq_valid = readResult_9_valid;
  wire               reorderQueueVec_10_enq_valid = readResult_10_valid;
  wire               reorderQueueVec_11_enq_valid = readResult_11_valid;
  wire               reorderQueueVec_12_enq_valid = readResult_12_valid;
  wire               reorderQueueVec_13_enq_valid = readResult_13_valid;
  wire               reorderQueueVec_14_enq_valid = readResult_14_valid;
  wire               reorderQueueVec_15_enq_valid = readResult_15_valid;
  wire               reorderQueueVec_16_enq_valid = readResult_16_valid;
  wire               reorderQueueVec_17_enq_valid = readResult_17_valid;
  wire               reorderQueueVec_18_enq_valid = readResult_18_valid;
  wire               reorderQueueVec_19_enq_valid = readResult_19_valid;
  wire               reorderQueueVec_20_enq_valid = readResult_20_valid;
  wire               reorderQueueVec_21_enq_valid = readResult_21_valid;
  wire               reorderQueueVec_22_enq_valid = readResult_22_valid;
  wire               reorderQueueVec_23_enq_valid = readResult_23_valid;
  wire               reorderQueueVec_24_enq_valid = readResult_24_valid;
  wire               reorderQueueVec_25_enq_valid = readResult_25_valid;
  wire               reorderQueueVec_26_enq_valid = readResult_26_valid;
  wire               reorderQueueVec_27_enq_valid = readResult_27_valid;
  wire               reorderQueueVec_28_enq_valid = readResult_28_valid;
  wire               reorderQueueVec_29_enq_valid = readResult_29_valid;
  wire               reorderQueueVec_30_enq_valid = readResult_30_valid;
  wire               reorderQueueVec_31_enq_valid = readResult_31_valid;
  wire               readMessageQueue_deq_ready = readResult_0_valid;
  wire               readMessageQueue_1_deq_ready = readResult_1_valid;
  wire               readMessageQueue_2_deq_ready = readResult_2_valid;
  wire               readMessageQueue_3_deq_ready = readResult_3_valid;
  wire               readMessageQueue_4_deq_ready = readResult_4_valid;
  wire               readMessageQueue_5_deq_ready = readResult_5_valid;
  wire               readMessageQueue_6_deq_ready = readResult_6_valid;
  wire               readMessageQueue_7_deq_ready = readResult_7_valid;
  wire               readMessageQueue_8_deq_ready = readResult_8_valid;
  wire               readMessageQueue_9_deq_ready = readResult_9_valid;
  wire               readMessageQueue_10_deq_ready = readResult_10_valid;
  wire               readMessageQueue_11_deq_ready = readResult_11_valid;
  wire               readMessageQueue_12_deq_ready = readResult_12_valid;
  wire               readMessageQueue_13_deq_ready = readResult_13_valid;
  wire               readMessageQueue_14_deq_ready = readResult_14_valid;
  wire               readMessageQueue_15_deq_ready = readResult_15_valid;
  wire               readMessageQueue_16_deq_ready = readResult_16_valid;
  wire               readMessageQueue_17_deq_ready = readResult_17_valid;
  wire               readMessageQueue_18_deq_ready = readResult_18_valid;
  wire               readMessageQueue_19_deq_ready = readResult_19_valid;
  wire               readMessageQueue_20_deq_ready = readResult_20_valid;
  wire               readMessageQueue_21_deq_ready = readResult_21_valid;
  wire               readMessageQueue_22_deq_ready = readResult_22_valid;
  wire               readMessageQueue_23_deq_ready = readResult_23_valid;
  wire               readMessageQueue_24_deq_ready = readResult_24_valid;
  wire               readMessageQueue_25_deq_ready = readResult_25_valid;
  wire               readMessageQueue_26_deq_ready = readResult_26_valid;
  wire               readMessageQueue_27_deq_ready = readResult_27_valid;
  wire               readMessageQueue_28_deq_ready = readResult_28_valid;
  wire               readMessageQueue_29_deq_ready = readResult_29_valid;
  wire               readMessageQueue_30_deq_ready = readResult_30_valid;
  wire               readMessageQueue_31_deq_ready = readResult_31_valid;
  wire [7:0]         checkVec_checkResult_lo_lo_lo_15 = 8'h0;
  wire [7:0]         checkVec_checkResult_lo_lo_hi_15 = 8'h0;
  wire [7:0]         checkVec_checkResult_lo_hi_lo_15 = 8'h0;
  wire [7:0]         checkVec_checkResult_lo_hi_hi_15 = 8'h0;
  wire [7:0]         checkVec_checkResult_hi_lo_lo_15 = 8'h0;
  wire [7:0]         checkVec_checkResult_hi_lo_hi_15 = 8'h0;
  wire [7:0]         checkVec_checkResult_hi_hi_lo_15 = 8'h0;
  wire [7:0]         checkVec_checkResult_hi_hi_hi_15 = 8'h0;
  wire [7:0]         checkVec_checkResult_lo_lo_lo_lo_14 = 8'hFF;
  wire [7:0]         checkVec_checkResult_lo_lo_lo_hi_14 = 8'hFF;
  wire [7:0]         checkVec_checkResult_lo_lo_hi_lo_14 = 8'hFF;
  wire [7:0]         checkVec_checkResult_lo_lo_hi_hi_14 = 8'hFF;
  wire [7:0]         checkVec_checkResult_lo_hi_lo_lo_14 = 8'hFF;
  wire [7:0]         checkVec_checkResult_lo_hi_lo_hi_14 = 8'hFF;
  wire [7:0]         checkVec_checkResult_lo_hi_hi_lo_14 = 8'hFF;
  wire [7:0]         checkVec_checkResult_lo_hi_hi_hi_14 = 8'hFF;
  wire [7:0]         checkVec_checkResult_hi_lo_lo_lo_14 = 8'hFF;
  wire [7:0]         checkVec_checkResult_hi_lo_lo_hi_14 = 8'hFF;
  wire [7:0]         checkVec_checkResult_hi_lo_hi_lo_14 = 8'hFF;
  wire [7:0]         checkVec_checkResult_hi_lo_hi_hi_14 = 8'hFF;
  wire [7:0]         checkVec_checkResult_hi_hi_lo_lo_14 = 8'hFF;
  wire [7:0]         checkVec_checkResult_hi_hi_lo_hi_14 = 8'hFF;
  wire [7:0]         checkVec_checkResult_hi_hi_hi_lo_14 = 8'hFF;
  wire [7:0]         checkVec_checkResult_hi_hi_hi_hi_14 = 8'hFF;
  wire [1:0]         checkVec_checkResultVec_0_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_1_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_2_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_3_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_4_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_5_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_6_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_7_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_8_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_9_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_10_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_11_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_12_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_13_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_14_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_15_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_16_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_17_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_18_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_19_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_20_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_21_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_22_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_23_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_24_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_25_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_26_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_27_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_28_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_29_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_30_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_31_1_2 = 2'h0;
  wire [15:0]        checkVec_checkResult_lo_lo_lo_14 = 16'hFFFF;
  wire [15:0]        checkVec_checkResult_lo_lo_hi_14 = 16'hFFFF;
  wire [15:0]        checkVec_checkResult_lo_hi_lo_14 = 16'hFFFF;
  wire [15:0]        checkVec_checkResult_lo_hi_hi_14 = 16'hFFFF;
  wire [15:0]        checkVec_checkResult_hi_lo_lo_14 = 16'hFFFF;
  wire [15:0]        checkVec_checkResult_hi_lo_hi_14 = 16'hFFFF;
  wire [15:0]        checkVec_checkResult_hi_hi_lo_14 = 16'hFFFF;
  wire [15:0]        checkVec_checkResult_hi_hi_hi_14 = 16'hFFFF;
  wire [31:0]        checkVec_checkResult_lo_lo_14 = 32'hFFFFFFFF;
  wire [31:0]        checkVec_checkResult_lo_hi_14 = 32'hFFFFFFFF;
  wire [31:0]        checkVec_checkResult_hi_lo_14 = 32'hFFFFFFFF;
  wire [31:0]        checkVec_checkResult_hi_hi_14 = 32'hFFFFFFFF;
  wire [63:0]        checkVec_checkResult_lo_14 = 64'hFFFFFFFFFFFFFFFF;
  wire [63:0]        checkVec_checkResult_hi_14 = 64'hFFFFFFFFFFFFFFFF;
  wire [127:0]       checkVec_2_0 = 128'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
  wire [3:0]         checkVec_checkResult_lo_lo_lo_lo_15 = 4'h0;
  wire [3:0]         checkVec_checkResult_lo_lo_lo_hi_15 = 4'h0;
  wire [3:0]         checkVec_checkResult_lo_lo_hi_lo_15 = 4'h0;
  wire [3:0]         checkVec_checkResult_lo_lo_hi_hi_15 = 4'h0;
  wire [3:0]         checkVec_checkResult_lo_hi_lo_lo_15 = 4'h0;
  wire [3:0]         checkVec_checkResult_lo_hi_lo_hi_15 = 4'h0;
  wire [3:0]         checkVec_checkResult_lo_hi_hi_lo_15 = 4'h0;
  wire [3:0]         checkVec_checkResult_lo_hi_hi_hi_15 = 4'h0;
  wire [3:0]         checkVec_checkResult_hi_lo_lo_lo_15 = 4'h0;
  wire [3:0]         checkVec_checkResult_hi_lo_lo_hi_15 = 4'h0;
  wire [3:0]         checkVec_checkResult_hi_lo_hi_lo_15 = 4'h0;
  wire [3:0]         checkVec_checkResult_hi_lo_hi_hi_15 = 4'h0;
  wire [3:0]         checkVec_checkResult_hi_hi_lo_lo_15 = 4'h0;
  wire [3:0]         checkVec_checkResult_hi_hi_lo_hi_15 = 4'h0;
  wire [3:0]         checkVec_checkResult_hi_hi_hi_lo_15 = 4'h0;
  wire [3:0]         checkVec_checkResult_hi_hi_hi_hi_15 = 4'h0;
  wire [15:0]        checkVec_checkResult_lo_lo_15 = 16'h0;
  wire [15:0]        checkVec_checkResult_lo_hi_15 = 16'h0;
  wire [15:0]        checkVec_checkResult_hi_lo_15 = 16'h0;
  wire [15:0]        checkVec_checkResult_hi_hi_15 = 16'h0;
  wire [63:0]        checkVec_2_1 = 64'h0;
  wire [4:0]         readVS1Req_requestIndex = 5'h0;
  wire [4:0]         selectExecuteReq_0_bits_requestIndex = 5'h0;
  wire [4:0]         selectExecuteReq_1_bits_requestIndex = 5'h1;
  wire [4:0]         selectExecuteReq_2_bits_requestIndex = 5'h2;
  wire [4:0]         selectExecuteReq_3_bits_requestIndex = 5'h3;
  wire [4:0]         selectExecuteReq_4_bits_requestIndex = 5'h4;
  wire [4:0]         selectExecuteReq_5_bits_requestIndex = 5'h5;
  wire [4:0]         selectExecuteReq_6_bits_requestIndex = 5'h6;
  wire [4:0]         selectExecuteReq_7_bits_requestIndex = 5'h7;
  wire [4:0]         selectExecuteReq_8_bits_requestIndex = 5'h8;
  wire [4:0]         selectExecuteReq_9_bits_requestIndex = 5'h9;
  wire [4:0]         selectExecuteReq_10_bits_requestIndex = 5'hA;
  wire [4:0]         selectExecuteReq_11_bits_requestIndex = 5'hB;
  wire [4:0]         selectExecuteReq_12_bits_requestIndex = 5'hC;
  wire [4:0]         selectExecuteReq_13_bits_requestIndex = 5'hD;
  wire [4:0]         selectExecuteReq_14_bits_requestIndex = 5'hE;
  wire [4:0]         selectExecuteReq_15_bits_requestIndex = 5'hF;
  wire [4:0]         selectExecuteReq_16_bits_requestIndex = 5'h10;
  wire [4:0]         selectExecuteReq_17_bits_requestIndex = 5'h11;
  wire [4:0]         selectExecuteReq_18_bits_requestIndex = 5'h12;
  wire [4:0]         selectExecuteReq_19_bits_requestIndex = 5'h13;
  wire [4:0]         selectExecuteReq_20_bits_requestIndex = 5'h14;
  wire [4:0]         selectExecuteReq_21_bits_requestIndex = 5'h15;
  wire [4:0]         selectExecuteReq_22_bits_requestIndex = 5'h16;
  wire [4:0]         selectExecuteReq_23_bits_requestIndex = 5'h17;
  wire [4:0]         selectExecuteReq_24_bits_requestIndex = 5'h18;
  wire [4:0]         selectExecuteReq_25_bits_requestIndex = 5'h19;
  wire [4:0]         selectExecuteReq_26_bits_requestIndex = 5'h1A;
  wire [4:0]         selectExecuteReq_27_bits_requestIndex = 5'h1B;
  wire [4:0]         selectExecuteReq_28_bits_requestIndex = 5'h1C;
  wire [4:0]         selectExecuteReq_29_bits_requestIndex = 5'h1D;
  wire [4:0]         selectExecuteReq_30_bits_requestIndex = 5'h1E;
  wire [4:0]         selectExecuteReq_31_bits_requestIndex = 5'h1F;
  wire               vs1Split_0_2 = 1'h1;
  wire               vs1Split_1_2 = 1'h1;
  wire               vs1Split_2_2 = 1'h1;
  wire [31:0]        checkVec_checkResult_lo_15 = 32'h0;
  wire [31:0]        checkVec_checkResult_hi_15 = 32'h0;
  wire [1:0]         readChannel_0_bits_readSource = 2'h2;
  wire [1:0]         readChannel_1_bits_readSource = 2'h2;
  wire [1:0]         readChannel_2_bits_readSource = 2'h2;
  wire [1:0]         readChannel_3_bits_readSource = 2'h2;
  wire [1:0]         readChannel_4_bits_readSource = 2'h2;
  wire [1:0]         readChannel_5_bits_readSource = 2'h2;
  wire [1:0]         readChannel_6_bits_readSource = 2'h2;
  wire [1:0]         readChannel_7_bits_readSource = 2'h2;
  wire [1:0]         readChannel_8_bits_readSource = 2'h2;
  wire [1:0]         readChannel_9_bits_readSource = 2'h2;
  wire [1:0]         readChannel_10_bits_readSource = 2'h2;
  wire [1:0]         readChannel_11_bits_readSource = 2'h2;
  wire [1:0]         readChannel_12_bits_readSource = 2'h2;
  wire [1:0]         readChannel_13_bits_readSource = 2'h2;
  wire [1:0]         readChannel_14_bits_readSource = 2'h2;
  wire [1:0]         readChannel_15_bits_readSource = 2'h2;
  wire [1:0]         readChannel_16_bits_readSource = 2'h2;
  wire [1:0]         readChannel_17_bits_readSource = 2'h2;
  wire [1:0]         readChannel_18_bits_readSource = 2'h2;
  wire [1:0]         readChannel_19_bits_readSource = 2'h2;
  wire [1:0]         readChannel_20_bits_readSource = 2'h2;
  wire [1:0]         readChannel_21_bits_readSource = 2'h2;
  wire [1:0]         readChannel_22_bits_readSource = 2'h2;
  wire [1:0]         readChannel_23_bits_readSource = 2'h2;
  wire [1:0]         readChannel_24_bits_readSource = 2'h2;
  wire [1:0]         readChannel_25_bits_readSource = 2'h2;
  wire [1:0]         readChannel_26_bits_readSource = 2'h2;
  wire [1:0]         readChannel_27_bits_readSource = 2'h2;
  wire [1:0]         readChannel_28_bits_readSource = 2'h2;
  wire [1:0]         readChannel_29_bits_readSource = 2'h2;
  wire [1:0]         readChannel_30_bits_readSource = 2'h2;
  wire [1:0]         readChannel_31_bits_readSource = 2'h2;
  wire               exeResp_0_bits_last = 1'h0;
  wire               exeResp_1_bits_last = 1'h0;
  wire               exeResp_2_bits_last = 1'h0;
  wire               exeResp_3_bits_last = 1'h0;
  wire               exeResp_4_bits_last = 1'h0;
  wire               exeResp_5_bits_last = 1'h0;
  wire               exeResp_6_bits_last = 1'h0;
  wire               exeResp_7_bits_last = 1'h0;
  wire               exeResp_8_bits_last = 1'h0;
  wire               exeResp_9_bits_last = 1'h0;
  wire               exeResp_10_bits_last = 1'h0;
  wire               exeResp_11_bits_last = 1'h0;
  wire               exeResp_12_bits_last = 1'h0;
  wire               exeResp_13_bits_last = 1'h0;
  wire               exeResp_14_bits_last = 1'h0;
  wire               exeResp_15_bits_last = 1'h0;
  wire               exeResp_16_bits_last = 1'h0;
  wire               exeResp_17_bits_last = 1'h0;
  wire               exeResp_18_bits_last = 1'h0;
  wire               exeResp_19_bits_last = 1'h0;
  wire               exeResp_20_bits_last = 1'h0;
  wire               exeResp_21_bits_last = 1'h0;
  wire               exeResp_22_bits_last = 1'h0;
  wire               exeResp_23_bits_last = 1'h0;
  wire               exeResp_24_bits_last = 1'h0;
  wire               exeResp_25_bits_last = 1'h0;
  wire               exeResp_26_bits_last = 1'h0;
  wire               exeResp_27_bits_last = 1'h0;
  wire               exeResp_28_bits_last = 1'h0;
  wire               exeResp_29_bits_last = 1'h0;
  wire               exeResp_30_bits_last = 1'h0;
  wire               exeResp_31_bits_last = 1'h0;
  wire               writeRequest_0_ffoByOther = 1'h0;
  wire               writeRequest_1_ffoByOther = 1'h0;
  wire               writeRequest_2_ffoByOther = 1'h0;
  wire               writeRequest_3_ffoByOther = 1'h0;
  wire               writeRequest_4_ffoByOther = 1'h0;
  wire               writeRequest_5_ffoByOther = 1'h0;
  wire               writeRequest_6_ffoByOther = 1'h0;
  wire               writeRequest_7_ffoByOther = 1'h0;
  wire               writeRequest_8_ffoByOther = 1'h0;
  wire               writeRequest_9_ffoByOther = 1'h0;
  wire               writeRequest_10_ffoByOther = 1'h0;
  wire               writeRequest_11_ffoByOther = 1'h0;
  wire               writeRequest_12_ffoByOther = 1'h0;
  wire               writeRequest_13_ffoByOther = 1'h0;
  wire               writeRequest_14_ffoByOther = 1'h0;
  wire               writeRequest_15_ffoByOther = 1'h0;
  wire               writeRequest_16_ffoByOther = 1'h0;
  wire               writeRequest_17_ffoByOther = 1'h0;
  wire               writeRequest_18_ffoByOther = 1'h0;
  wire               writeRequest_19_ffoByOther = 1'h0;
  wire               writeRequest_20_ffoByOther = 1'h0;
  wire               writeRequest_21_ffoByOther = 1'h0;
  wire               writeRequest_22_ffoByOther = 1'h0;
  wire               writeRequest_23_ffoByOther = 1'h0;
  wire               writeRequest_24_ffoByOther = 1'h0;
  wire               writeRequest_25_ffoByOther = 1'h0;
  wire               writeRequest_26_ffoByOther = 1'h0;
  wire               writeRequest_27_ffoByOther = 1'h0;
  wire               writeRequest_28_ffoByOther = 1'h0;
  wire               writeRequest_29_ffoByOther = 1'h0;
  wire               writeRequest_30_ffoByOther = 1'h0;
  wire               writeRequest_31_ffoByOther = 1'h0;
  wire               writeQueue_0_deq_ready = exeResp_0_ready_0;
  wire               writeQueue_0_deq_valid;
  wire [3:0]         writeQueue_0_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_0_deq_bits_writeData_data;
  wire               writeQueue_1_deq_ready = exeResp_1_ready_0;
  wire               writeQueue_1_deq_valid;
  wire [3:0]         writeQueue_1_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_1_deq_bits_writeData_data;
  wire               writeQueue_2_deq_ready = exeResp_2_ready_0;
  wire               writeQueue_2_deq_valid;
  wire [3:0]         writeQueue_2_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_2_deq_bits_writeData_data;
  wire               writeQueue_3_deq_ready = exeResp_3_ready_0;
  wire               writeQueue_3_deq_valid;
  wire [3:0]         writeQueue_3_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_3_deq_bits_writeData_data;
  wire               writeQueue_4_deq_ready = exeResp_4_ready_0;
  wire               writeQueue_4_deq_valid;
  wire [3:0]         writeQueue_4_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_4_deq_bits_writeData_data;
  wire               writeQueue_5_deq_ready = exeResp_5_ready_0;
  wire               writeQueue_5_deq_valid;
  wire [3:0]         writeQueue_5_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_5_deq_bits_writeData_data;
  wire               writeQueue_6_deq_ready = exeResp_6_ready_0;
  wire               writeQueue_6_deq_valid;
  wire [3:0]         writeQueue_6_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_6_deq_bits_writeData_data;
  wire               writeQueue_7_deq_ready = exeResp_7_ready_0;
  wire               writeQueue_7_deq_valid;
  wire [3:0]         writeQueue_7_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_7_deq_bits_writeData_data;
  wire               writeQueue_8_deq_ready = exeResp_8_ready_0;
  wire               writeQueue_8_deq_valid;
  wire [3:0]         writeQueue_8_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_8_deq_bits_writeData_data;
  wire               writeQueue_9_deq_ready = exeResp_9_ready_0;
  wire               writeQueue_9_deq_valid;
  wire [3:0]         writeQueue_9_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_9_deq_bits_writeData_data;
  wire               writeQueue_10_deq_ready = exeResp_10_ready_0;
  wire               writeQueue_10_deq_valid;
  wire [3:0]         writeQueue_10_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_10_deq_bits_writeData_data;
  wire               writeQueue_11_deq_ready = exeResp_11_ready_0;
  wire               writeQueue_11_deq_valid;
  wire [3:0]         writeQueue_11_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_11_deq_bits_writeData_data;
  wire               writeQueue_12_deq_ready = exeResp_12_ready_0;
  wire               writeQueue_12_deq_valid;
  wire [3:0]         writeQueue_12_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_12_deq_bits_writeData_data;
  wire               writeQueue_13_deq_ready = exeResp_13_ready_0;
  wire               writeQueue_13_deq_valid;
  wire [3:0]         writeQueue_13_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_13_deq_bits_writeData_data;
  wire               writeQueue_14_deq_ready = exeResp_14_ready_0;
  wire               writeQueue_14_deq_valid;
  wire [3:0]         writeQueue_14_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_14_deq_bits_writeData_data;
  wire               writeQueue_15_deq_ready = exeResp_15_ready_0;
  wire               writeQueue_15_deq_valid;
  wire [3:0]         writeQueue_15_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_15_deq_bits_writeData_data;
  wire               writeQueue_16_deq_ready = exeResp_16_ready_0;
  wire               writeQueue_16_deq_valid;
  wire [3:0]         writeQueue_16_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_16_deq_bits_writeData_data;
  wire               writeQueue_17_deq_ready = exeResp_17_ready_0;
  wire               writeQueue_17_deq_valid;
  wire [3:0]         writeQueue_17_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_17_deq_bits_writeData_data;
  wire               writeQueue_18_deq_ready = exeResp_18_ready_0;
  wire               writeQueue_18_deq_valid;
  wire [3:0]         writeQueue_18_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_18_deq_bits_writeData_data;
  wire               writeQueue_19_deq_ready = exeResp_19_ready_0;
  wire               writeQueue_19_deq_valid;
  wire [3:0]         writeQueue_19_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_19_deq_bits_writeData_data;
  wire               writeQueue_20_deq_ready = exeResp_20_ready_0;
  wire               writeQueue_20_deq_valid;
  wire [3:0]         writeQueue_20_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_20_deq_bits_writeData_data;
  wire               writeQueue_21_deq_ready = exeResp_21_ready_0;
  wire               writeQueue_21_deq_valid;
  wire [3:0]         writeQueue_21_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_21_deq_bits_writeData_data;
  wire               writeQueue_22_deq_ready = exeResp_22_ready_0;
  wire               writeQueue_22_deq_valid;
  wire [3:0]         writeQueue_22_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_22_deq_bits_writeData_data;
  wire               writeQueue_23_deq_ready = exeResp_23_ready_0;
  wire               writeQueue_23_deq_valid;
  wire [3:0]         writeQueue_23_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_23_deq_bits_writeData_data;
  wire               writeQueue_24_deq_ready = exeResp_24_ready_0;
  wire               writeQueue_24_deq_valid;
  wire [3:0]         writeQueue_24_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_24_deq_bits_writeData_data;
  wire               writeQueue_25_deq_ready = exeResp_25_ready_0;
  wire               writeQueue_25_deq_valid;
  wire [3:0]         writeQueue_25_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_25_deq_bits_writeData_data;
  wire               writeQueue_26_deq_ready = exeResp_26_ready_0;
  wire               writeQueue_26_deq_valid;
  wire [3:0]         writeQueue_26_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_26_deq_bits_writeData_data;
  wire               writeQueue_27_deq_ready = exeResp_27_ready_0;
  wire               writeQueue_27_deq_valid;
  wire [3:0]         writeQueue_27_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_27_deq_bits_writeData_data;
  wire               writeQueue_28_deq_ready = exeResp_28_ready_0;
  wire               writeQueue_28_deq_valid;
  wire [3:0]         writeQueue_28_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_28_deq_bits_writeData_data;
  wire               writeQueue_29_deq_ready = exeResp_29_ready_0;
  wire               writeQueue_29_deq_valid;
  wire [3:0]         writeQueue_29_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_29_deq_bits_writeData_data;
  wire               writeQueue_30_deq_ready = exeResp_30_ready_0;
  wire               writeQueue_30_deq_valid;
  wire [3:0]         writeQueue_30_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_30_deq_bits_writeData_data;
  wire               writeQueue_31_deq_ready = exeResp_31_ready_0;
  wire               writeQueue_31_deq_valid;
  wire [3:0]         writeQueue_31_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_31_deq_bits_writeData_data;
  wire               gatherResponse;
  reg  [31:0]        v0_0;
  reg  [31:0]        v0_1;
  reg  [31:0]        v0_2;
  reg  [31:0]        v0_3;
  reg  [31:0]        v0_4;
  reg  [31:0]        v0_5;
  reg  [31:0]        v0_6;
  reg  [31:0]        v0_7;
  reg  [31:0]        v0_8;
  reg  [31:0]        v0_9;
  reg  [31:0]        v0_10;
  reg  [31:0]        v0_11;
  reg  [31:0]        v0_12;
  reg  [31:0]        v0_13;
  reg  [31:0]        v0_14;
  reg  [31:0]        v0_15;
  reg  [31:0]        v0_16;
  reg  [31:0]        v0_17;
  reg  [31:0]        v0_18;
  reg  [31:0]        v0_19;
  reg  [31:0]        v0_20;
  reg  [31:0]        v0_21;
  reg  [31:0]        v0_22;
  reg  [31:0]        v0_23;
  reg  [31:0]        v0_24;
  reg  [31:0]        v0_25;
  reg  [31:0]        v0_26;
  reg  [31:0]        v0_27;
  reg  [31:0]        v0_28;
  reg  [31:0]        v0_29;
  reg  [31:0]        v0_30;
  reg  [31:0]        v0_31;
  reg  [31:0]        v0_32;
  reg  [31:0]        v0_33;
  reg  [31:0]        v0_34;
  reg  [31:0]        v0_35;
  reg  [31:0]        v0_36;
  reg  [31:0]        v0_37;
  reg  [31:0]        v0_38;
  reg  [31:0]        v0_39;
  reg  [31:0]        v0_40;
  reg  [31:0]        v0_41;
  reg  [31:0]        v0_42;
  reg  [31:0]        v0_43;
  reg  [31:0]        v0_44;
  reg  [31:0]        v0_45;
  reg  [31:0]        v0_46;
  reg  [31:0]        v0_47;
  reg  [31:0]        v0_48;
  reg  [31:0]        v0_49;
  reg  [31:0]        v0_50;
  reg  [31:0]        v0_51;
  reg  [31:0]        v0_52;
  reg  [31:0]        v0_53;
  reg  [31:0]        v0_54;
  reg  [31:0]        v0_55;
  reg  [31:0]        v0_56;
  reg  [31:0]        v0_57;
  reg  [31:0]        v0_58;
  reg  [31:0]        v0_59;
  reg  [31:0]        v0_60;
  reg  [31:0]        v0_61;
  reg  [31:0]        v0_62;
  reg  [31:0]        v0_63;
  wire [15:0]        maskExt_lo = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt = {maskExt_hi, maskExt_lo};
  wire [15:0]        maskExt_lo_1 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_1 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_1 = {maskExt_hi_1, maskExt_lo_1};
  wire [15:0]        maskExt_lo_2 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_2 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_2 = {maskExt_hi_2, maskExt_lo_2};
  wire [15:0]        maskExt_lo_3 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_3 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_3 = {maskExt_hi_3, maskExt_lo_3};
  wire [15:0]        maskExt_lo_4 = {{8{v0UpdateVec_4_bits_mask[1]}}, {8{v0UpdateVec_4_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_4 = {{8{v0UpdateVec_4_bits_mask[3]}}, {8{v0UpdateVec_4_bits_mask[2]}}};
  wire [31:0]        maskExt_4 = {maskExt_hi_4, maskExt_lo_4};
  wire [15:0]        maskExt_lo_5 = {{8{v0UpdateVec_5_bits_mask[1]}}, {8{v0UpdateVec_5_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_5 = {{8{v0UpdateVec_5_bits_mask[3]}}, {8{v0UpdateVec_5_bits_mask[2]}}};
  wire [31:0]        maskExt_5 = {maskExt_hi_5, maskExt_lo_5};
  wire [15:0]        maskExt_lo_6 = {{8{v0UpdateVec_6_bits_mask[1]}}, {8{v0UpdateVec_6_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_6 = {{8{v0UpdateVec_6_bits_mask[3]}}, {8{v0UpdateVec_6_bits_mask[2]}}};
  wire [31:0]        maskExt_6 = {maskExt_hi_6, maskExt_lo_6};
  wire [15:0]        maskExt_lo_7 = {{8{v0UpdateVec_7_bits_mask[1]}}, {8{v0UpdateVec_7_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_7 = {{8{v0UpdateVec_7_bits_mask[3]}}, {8{v0UpdateVec_7_bits_mask[2]}}};
  wire [31:0]        maskExt_7 = {maskExt_hi_7, maskExt_lo_7};
  wire [15:0]        maskExt_lo_8 = {{8{v0UpdateVec_8_bits_mask[1]}}, {8{v0UpdateVec_8_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_8 = {{8{v0UpdateVec_8_bits_mask[3]}}, {8{v0UpdateVec_8_bits_mask[2]}}};
  wire [31:0]        maskExt_8 = {maskExt_hi_8, maskExt_lo_8};
  wire [15:0]        maskExt_lo_9 = {{8{v0UpdateVec_9_bits_mask[1]}}, {8{v0UpdateVec_9_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_9 = {{8{v0UpdateVec_9_bits_mask[3]}}, {8{v0UpdateVec_9_bits_mask[2]}}};
  wire [31:0]        maskExt_9 = {maskExt_hi_9, maskExt_lo_9};
  wire [15:0]        maskExt_lo_10 = {{8{v0UpdateVec_10_bits_mask[1]}}, {8{v0UpdateVec_10_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_10 = {{8{v0UpdateVec_10_bits_mask[3]}}, {8{v0UpdateVec_10_bits_mask[2]}}};
  wire [31:0]        maskExt_10 = {maskExt_hi_10, maskExt_lo_10};
  wire [15:0]        maskExt_lo_11 = {{8{v0UpdateVec_11_bits_mask[1]}}, {8{v0UpdateVec_11_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_11 = {{8{v0UpdateVec_11_bits_mask[3]}}, {8{v0UpdateVec_11_bits_mask[2]}}};
  wire [31:0]        maskExt_11 = {maskExt_hi_11, maskExt_lo_11};
  wire [15:0]        maskExt_lo_12 = {{8{v0UpdateVec_12_bits_mask[1]}}, {8{v0UpdateVec_12_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_12 = {{8{v0UpdateVec_12_bits_mask[3]}}, {8{v0UpdateVec_12_bits_mask[2]}}};
  wire [31:0]        maskExt_12 = {maskExt_hi_12, maskExt_lo_12};
  wire [15:0]        maskExt_lo_13 = {{8{v0UpdateVec_13_bits_mask[1]}}, {8{v0UpdateVec_13_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_13 = {{8{v0UpdateVec_13_bits_mask[3]}}, {8{v0UpdateVec_13_bits_mask[2]}}};
  wire [31:0]        maskExt_13 = {maskExt_hi_13, maskExt_lo_13};
  wire [15:0]        maskExt_lo_14 = {{8{v0UpdateVec_14_bits_mask[1]}}, {8{v0UpdateVec_14_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_14 = {{8{v0UpdateVec_14_bits_mask[3]}}, {8{v0UpdateVec_14_bits_mask[2]}}};
  wire [31:0]        maskExt_14 = {maskExt_hi_14, maskExt_lo_14};
  wire [15:0]        maskExt_lo_15 = {{8{v0UpdateVec_15_bits_mask[1]}}, {8{v0UpdateVec_15_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_15 = {{8{v0UpdateVec_15_bits_mask[3]}}, {8{v0UpdateVec_15_bits_mask[2]}}};
  wire [31:0]        maskExt_15 = {maskExt_hi_15, maskExt_lo_15};
  wire [15:0]        maskExt_lo_16 = {{8{v0UpdateVec_16_bits_mask[1]}}, {8{v0UpdateVec_16_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_16 = {{8{v0UpdateVec_16_bits_mask[3]}}, {8{v0UpdateVec_16_bits_mask[2]}}};
  wire [31:0]        maskExt_16 = {maskExt_hi_16, maskExt_lo_16};
  wire [15:0]        maskExt_lo_17 = {{8{v0UpdateVec_17_bits_mask[1]}}, {8{v0UpdateVec_17_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_17 = {{8{v0UpdateVec_17_bits_mask[3]}}, {8{v0UpdateVec_17_bits_mask[2]}}};
  wire [31:0]        maskExt_17 = {maskExt_hi_17, maskExt_lo_17};
  wire [15:0]        maskExt_lo_18 = {{8{v0UpdateVec_18_bits_mask[1]}}, {8{v0UpdateVec_18_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_18 = {{8{v0UpdateVec_18_bits_mask[3]}}, {8{v0UpdateVec_18_bits_mask[2]}}};
  wire [31:0]        maskExt_18 = {maskExt_hi_18, maskExt_lo_18};
  wire [15:0]        maskExt_lo_19 = {{8{v0UpdateVec_19_bits_mask[1]}}, {8{v0UpdateVec_19_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_19 = {{8{v0UpdateVec_19_bits_mask[3]}}, {8{v0UpdateVec_19_bits_mask[2]}}};
  wire [31:0]        maskExt_19 = {maskExt_hi_19, maskExt_lo_19};
  wire [15:0]        maskExt_lo_20 = {{8{v0UpdateVec_20_bits_mask[1]}}, {8{v0UpdateVec_20_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_20 = {{8{v0UpdateVec_20_bits_mask[3]}}, {8{v0UpdateVec_20_bits_mask[2]}}};
  wire [31:0]        maskExt_20 = {maskExt_hi_20, maskExt_lo_20};
  wire [15:0]        maskExt_lo_21 = {{8{v0UpdateVec_21_bits_mask[1]}}, {8{v0UpdateVec_21_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_21 = {{8{v0UpdateVec_21_bits_mask[3]}}, {8{v0UpdateVec_21_bits_mask[2]}}};
  wire [31:0]        maskExt_21 = {maskExt_hi_21, maskExt_lo_21};
  wire [15:0]        maskExt_lo_22 = {{8{v0UpdateVec_22_bits_mask[1]}}, {8{v0UpdateVec_22_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_22 = {{8{v0UpdateVec_22_bits_mask[3]}}, {8{v0UpdateVec_22_bits_mask[2]}}};
  wire [31:0]        maskExt_22 = {maskExt_hi_22, maskExt_lo_22};
  wire [15:0]        maskExt_lo_23 = {{8{v0UpdateVec_23_bits_mask[1]}}, {8{v0UpdateVec_23_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_23 = {{8{v0UpdateVec_23_bits_mask[3]}}, {8{v0UpdateVec_23_bits_mask[2]}}};
  wire [31:0]        maskExt_23 = {maskExt_hi_23, maskExt_lo_23};
  wire [15:0]        maskExt_lo_24 = {{8{v0UpdateVec_24_bits_mask[1]}}, {8{v0UpdateVec_24_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_24 = {{8{v0UpdateVec_24_bits_mask[3]}}, {8{v0UpdateVec_24_bits_mask[2]}}};
  wire [31:0]        maskExt_24 = {maskExt_hi_24, maskExt_lo_24};
  wire [15:0]        maskExt_lo_25 = {{8{v0UpdateVec_25_bits_mask[1]}}, {8{v0UpdateVec_25_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_25 = {{8{v0UpdateVec_25_bits_mask[3]}}, {8{v0UpdateVec_25_bits_mask[2]}}};
  wire [31:0]        maskExt_25 = {maskExt_hi_25, maskExt_lo_25};
  wire [15:0]        maskExt_lo_26 = {{8{v0UpdateVec_26_bits_mask[1]}}, {8{v0UpdateVec_26_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_26 = {{8{v0UpdateVec_26_bits_mask[3]}}, {8{v0UpdateVec_26_bits_mask[2]}}};
  wire [31:0]        maskExt_26 = {maskExt_hi_26, maskExt_lo_26};
  wire [15:0]        maskExt_lo_27 = {{8{v0UpdateVec_27_bits_mask[1]}}, {8{v0UpdateVec_27_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_27 = {{8{v0UpdateVec_27_bits_mask[3]}}, {8{v0UpdateVec_27_bits_mask[2]}}};
  wire [31:0]        maskExt_27 = {maskExt_hi_27, maskExt_lo_27};
  wire [15:0]        maskExt_lo_28 = {{8{v0UpdateVec_28_bits_mask[1]}}, {8{v0UpdateVec_28_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_28 = {{8{v0UpdateVec_28_bits_mask[3]}}, {8{v0UpdateVec_28_bits_mask[2]}}};
  wire [31:0]        maskExt_28 = {maskExt_hi_28, maskExt_lo_28};
  wire [15:0]        maskExt_lo_29 = {{8{v0UpdateVec_29_bits_mask[1]}}, {8{v0UpdateVec_29_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_29 = {{8{v0UpdateVec_29_bits_mask[3]}}, {8{v0UpdateVec_29_bits_mask[2]}}};
  wire [31:0]        maskExt_29 = {maskExt_hi_29, maskExt_lo_29};
  wire [15:0]        maskExt_lo_30 = {{8{v0UpdateVec_30_bits_mask[1]}}, {8{v0UpdateVec_30_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_30 = {{8{v0UpdateVec_30_bits_mask[3]}}, {8{v0UpdateVec_30_bits_mask[2]}}};
  wire [31:0]        maskExt_30 = {maskExt_hi_30, maskExt_lo_30};
  wire [15:0]        maskExt_lo_31 = {{8{v0UpdateVec_31_bits_mask[1]}}, {8{v0UpdateVec_31_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_31 = {{8{v0UpdateVec_31_bits_mask[3]}}, {8{v0UpdateVec_31_bits_mask[2]}}};
  wire [31:0]        maskExt_31 = {maskExt_hi_31, maskExt_lo_31};
  wire [15:0]        maskExt_lo_32 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_32 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_32 = {maskExt_hi_32, maskExt_lo_32};
  wire [15:0]        maskExt_lo_33 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_33 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_33 = {maskExt_hi_33, maskExt_lo_33};
  wire [15:0]        maskExt_lo_34 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_34 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_34 = {maskExt_hi_34, maskExt_lo_34};
  wire [15:0]        maskExt_lo_35 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_35 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_35 = {maskExt_hi_35, maskExt_lo_35};
  wire [15:0]        maskExt_lo_36 = {{8{v0UpdateVec_4_bits_mask[1]}}, {8{v0UpdateVec_4_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_36 = {{8{v0UpdateVec_4_bits_mask[3]}}, {8{v0UpdateVec_4_bits_mask[2]}}};
  wire [31:0]        maskExt_36 = {maskExt_hi_36, maskExt_lo_36};
  wire [15:0]        maskExt_lo_37 = {{8{v0UpdateVec_5_bits_mask[1]}}, {8{v0UpdateVec_5_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_37 = {{8{v0UpdateVec_5_bits_mask[3]}}, {8{v0UpdateVec_5_bits_mask[2]}}};
  wire [31:0]        maskExt_37 = {maskExt_hi_37, maskExt_lo_37};
  wire [15:0]        maskExt_lo_38 = {{8{v0UpdateVec_6_bits_mask[1]}}, {8{v0UpdateVec_6_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_38 = {{8{v0UpdateVec_6_bits_mask[3]}}, {8{v0UpdateVec_6_bits_mask[2]}}};
  wire [31:0]        maskExt_38 = {maskExt_hi_38, maskExt_lo_38};
  wire [15:0]        maskExt_lo_39 = {{8{v0UpdateVec_7_bits_mask[1]}}, {8{v0UpdateVec_7_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_39 = {{8{v0UpdateVec_7_bits_mask[3]}}, {8{v0UpdateVec_7_bits_mask[2]}}};
  wire [31:0]        maskExt_39 = {maskExt_hi_39, maskExt_lo_39};
  wire [15:0]        maskExt_lo_40 = {{8{v0UpdateVec_8_bits_mask[1]}}, {8{v0UpdateVec_8_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_40 = {{8{v0UpdateVec_8_bits_mask[3]}}, {8{v0UpdateVec_8_bits_mask[2]}}};
  wire [31:0]        maskExt_40 = {maskExt_hi_40, maskExt_lo_40};
  wire [15:0]        maskExt_lo_41 = {{8{v0UpdateVec_9_bits_mask[1]}}, {8{v0UpdateVec_9_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_41 = {{8{v0UpdateVec_9_bits_mask[3]}}, {8{v0UpdateVec_9_bits_mask[2]}}};
  wire [31:0]        maskExt_41 = {maskExt_hi_41, maskExt_lo_41};
  wire [15:0]        maskExt_lo_42 = {{8{v0UpdateVec_10_bits_mask[1]}}, {8{v0UpdateVec_10_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_42 = {{8{v0UpdateVec_10_bits_mask[3]}}, {8{v0UpdateVec_10_bits_mask[2]}}};
  wire [31:0]        maskExt_42 = {maskExt_hi_42, maskExt_lo_42};
  wire [15:0]        maskExt_lo_43 = {{8{v0UpdateVec_11_bits_mask[1]}}, {8{v0UpdateVec_11_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_43 = {{8{v0UpdateVec_11_bits_mask[3]}}, {8{v0UpdateVec_11_bits_mask[2]}}};
  wire [31:0]        maskExt_43 = {maskExt_hi_43, maskExt_lo_43};
  wire [15:0]        maskExt_lo_44 = {{8{v0UpdateVec_12_bits_mask[1]}}, {8{v0UpdateVec_12_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_44 = {{8{v0UpdateVec_12_bits_mask[3]}}, {8{v0UpdateVec_12_bits_mask[2]}}};
  wire [31:0]        maskExt_44 = {maskExt_hi_44, maskExt_lo_44};
  wire [15:0]        maskExt_lo_45 = {{8{v0UpdateVec_13_bits_mask[1]}}, {8{v0UpdateVec_13_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_45 = {{8{v0UpdateVec_13_bits_mask[3]}}, {8{v0UpdateVec_13_bits_mask[2]}}};
  wire [31:0]        maskExt_45 = {maskExt_hi_45, maskExt_lo_45};
  wire [15:0]        maskExt_lo_46 = {{8{v0UpdateVec_14_bits_mask[1]}}, {8{v0UpdateVec_14_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_46 = {{8{v0UpdateVec_14_bits_mask[3]}}, {8{v0UpdateVec_14_bits_mask[2]}}};
  wire [31:0]        maskExt_46 = {maskExt_hi_46, maskExt_lo_46};
  wire [15:0]        maskExt_lo_47 = {{8{v0UpdateVec_15_bits_mask[1]}}, {8{v0UpdateVec_15_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_47 = {{8{v0UpdateVec_15_bits_mask[3]}}, {8{v0UpdateVec_15_bits_mask[2]}}};
  wire [31:0]        maskExt_47 = {maskExt_hi_47, maskExt_lo_47};
  wire [15:0]        maskExt_lo_48 = {{8{v0UpdateVec_16_bits_mask[1]}}, {8{v0UpdateVec_16_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_48 = {{8{v0UpdateVec_16_bits_mask[3]}}, {8{v0UpdateVec_16_bits_mask[2]}}};
  wire [31:0]        maskExt_48 = {maskExt_hi_48, maskExt_lo_48};
  wire [15:0]        maskExt_lo_49 = {{8{v0UpdateVec_17_bits_mask[1]}}, {8{v0UpdateVec_17_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_49 = {{8{v0UpdateVec_17_bits_mask[3]}}, {8{v0UpdateVec_17_bits_mask[2]}}};
  wire [31:0]        maskExt_49 = {maskExt_hi_49, maskExt_lo_49};
  wire [15:0]        maskExt_lo_50 = {{8{v0UpdateVec_18_bits_mask[1]}}, {8{v0UpdateVec_18_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_50 = {{8{v0UpdateVec_18_bits_mask[3]}}, {8{v0UpdateVec_18_bits_mask[2]}}};
  wire [31:0]        maskExt_50 = {maskExt_hi_50, maskExt_lo_50};
  wire [15:0]        maskExt_lo_51 = {{8{v0UpdateVec_19_bits_mask[1]}}, {8{v0UpdateVec_19_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_51 = {{8{v0UpdateVec_19_bits_mask[3]}}, {8{v0UpdateVec_19_bits_mask[2]}}};
  wire [31:0]        maskExt_51 = {maskExt_hi_51, maskExt_lo_51};
  wire [15:0]        maskExt_lo_52 = {{8{v0UpdateVec_20_bits_mask[1]}}, {8{v0UpdateVec_20_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_52 = {{8{v0UpdateVec_20_bits_mask[3]}}, {8{v0UpdateVec_20_bits_mask[2]}}};
  wire [31:0]        maskExt_52 = {maskExt_hi_52, maskExt_lo_52};
  wire [15:0]        maskExt_lo_53 = {{8{v0UpdateVec_21_bits_mask[1]}}, {8{v0UpdateVec_21_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_53 = {{8{v0UpdateVec_21_bits_mask[3]}}, {8{v0UpdateVec_21_bits_mask[2]}}};
  wire [31:0]        maskExt_53 = {maskExt_hi_53, maskExt_lo_53};
  wire [15:0]        maskExt_lo_54 = {{8{v0UpdateVec_22_bits_mask[1]}}, {8{v0UpdateVec_22_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_54 = {{8{v0UpdateVec_22_bits_mask[3]}}, {8{v0UpdateVec_22_bits_mask[2]}}};
  wire [31:0]        maskExt_54 = {maskExt_hi_54, maskExt_lo_54};
  wire [15:0]        maskExt_lo_55 = {{8{v0UpdateVec_23_bits_mask[1]}}, {8{v0UpdateVec_23_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_55 = {{8{v0UpdateVec_23_bits_mask[3]}}, {8{v0UpdateVec_23_bits_mask[2]}}};
  wire [31:0]        maskExt_55 = {maskExt_hi_55, maskExt_lo_55};
  wire [15:0]        maskExt_lo_56 = {{8{v0UpdateVec_24_bits_mask[1]}}, {8{v0UpdateVec_24_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_56 = {{8{v0UpdateVec_24_bits_mask[3]}}, {8{v0UpdateVec_24_bits_mask[2]}}};
  wire [31:0]        maskExt_56 = {maskExt_hi_56, maskExt_lo_56};
  wire [15:0]        maskExt_lo_57 = {{8{v0UpdateVec_25_bits_mask[1]}}, {8{v0UpdateVec_25_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_57 = {{8{v0UpdateVec_25_bits_mask[3]}}, {8{v0UpdateVec_25_bits_mask[2]}}};
  wire [31:0]        maskExt_57 = {maskExt_hi_57, maskExt_lo_57};
  wire [15:0]        maskExt_lo_58 = {{8{v0UpdateVec_26_bits_mask[1]}}, {8{v0UpdateVec_26_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_58 = {{8{v0UpdateVec_26_bits_mask[3]}}, {8{v0UpdateVec_26_bits_mask[2]}}};
  wire [31:0]        maskExt_58 = {maskExt_hi_58, maskExt_lo_58};
  wire [15:0]        maskExt_lo_59 = {{8{v0UpdateVec_27_bits_mask[1]}}, {8{v0UpdateVec_27_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_59 = {{8{v0UpdateVec_27_bits_mask[3]}}, {8{v0UpdateVec_27_bits_mask[2]}}};
  wire [31:0]        maskExt_59 = {maskExt_hi_59, maskExt_lo_59};
  wire [15:0]        maskExt_lo_60 = {{8{v0UpdateVec_28_bits_mask[1]}}, {8{v0UpdateVec_28_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_60 = {{8{v0UpdateVec_28_bits_mask[3]}}, {8{v0UpdateVec_28_bits_mask[2]}}};
  wire [31:0]        maskExt_60 = {maskExt_hi_60, maskExt_lo_60};
  wire [15:0]        maskExt_lo_61 = {{8{v0UpdateVec_29_bits_mask[1]}}, {8{v0UpdateVec_29_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_61 = {{8{v0UpdateVec_29_bits_mask[3]}}, {8{v0UpdateVec_29_bits_mask[2]}}};
  wire [31:0]        maskExt_61 = {maskExt_hi_61, maskExt_lo_61};
  wire [15:0]        maskExt_lo_62 = {{8{v0UpdateVec_30_bits_mask[1]}}, {8{v0UpdateVec_30_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_62 = {{8{v0UpdateVec_30_bits_mask[3]}}, {8{v0UpdateVec_30_bits_mask[2]}}};
  wire [31:0]        maskExt_62 = {maskExt_hi_62, maskExt_lo_62};
  wire [15:0]        maskExt_lo_63 = {{8{v0UpdateVec_31_bits_mask[1]}}, {8{v0UpdateVec_31_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_63 = {{8{v0UpdateVec_31_bits_mask[3]}}, {8{v0UpdateVec_31_bits_mask[2]}}};
  wire [31:0]        maskExt_63 = {maskExt_hi_63, maskExt_lo_63};
  wire [63:0]        _GEN = {v0_1, v0_0};
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo;
  assign regroupV0_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_1;
  assign regroupV0_lo_lo_lo_lo_lo_1 = _GEN;
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_2;
  assign regroupV0_lo_lo_lo_lo_lo_2 = _GEN;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]        selectReadStageMask_lo_lo_lo_lo_lo;
  assign selectReadStageMask_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_lo;
  assign maskSplit_maskSelect_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_lo_1;
  assign maskSplit_maskSelect_lo_lo_lo_lo_lo_1 = _GEN;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_lo_2;
  assign maskSplit_maskSelect_lo_lo_lo_lo_lo_2 = _GEN;
  wire [63:0]        maskForDestination_lo_lo_lo_lo_lo;
  assign maskForDestination_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]        _GEN_0 = {v0_3, v0_2};
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi;
  assign regroupV0_lo_lo_lo_lo_hi = _GEN_0;
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_1;
  assign regroupV0_lo_lo_lo_lo_hi_1 = _GEN_0;
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_2;
  assign regroupV0_lo_lo_lo_lo_hi_2 = _GEN_0;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi = _GEN_0;
  wire [63:0]        selectReadStageMask_lo_lo_lo_lo_hi;
  assign selectReadStageMask_lo_lo_lo_lo_hi = _GEN_0;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_hi;
  assign maskSplit_maskSelect_lo_lo_lo_lo_hi = _GEN_0;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_hi_1;
  assign maskSplit_maskSelect_lo_lo_lo_lo_hi_1 = _GEN_0;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_hi_2;
  assign maskSplit_maskSelect_lo_lo_lo_lo_hi_2 = _GEN_0;
  wire [63:0]        maskForDestination_lo_lo_lo_lo_hi;
  assign maskForDestination_lo_lo_lo_lo_hi = _GEN_0;
  wire [127:0]       regroupV0_lo_lo_lo_lo = {regroupV0_lo_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo_lo};
  wire [63:0]        _GEN_1 = {v0_5, v0_4};
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo;
  assign regroupV0_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_1;
  assign regroupV0_lo_lo_lo_hi_lo_1 = _GEN_1;
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_2;
  assign regroupV0_lo_lo_lo_hi_lo_2 = _GEN_1;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]        selectReadStageMask_lo_lo_lo_hi_lo;
  assign selectReadStageMask_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_lo;
  assign maskSplit_maskSelect_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_lo_1;
  assign maskSplit_maskSelect_lo_lo_lo_hi_lo_1 = _GEN_1;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_lo_2;
  assign maskSplit_maskSelect_lo_lo_lo_hi_lo_2 = _GEN_1;
  wire [63:0]        maskForDestination_lo_lo_lo_hi_lo;
  assign maskForDestination_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]        _GEN_2 = {v0_7, v0_6};
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi;
  assign regroupV0_lo_lo_lo_hi_hi = _GEN_2;
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_1;
  assign regroupV0_lo_lo_lo_hi_hi_1 = _GEN_2;
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_2;
  assign regroupV0_lo_lo_lo_hi_hi_2 = _GEN_2;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi = _GEN_2;
  wire [63:0]        selectReadStageMask_lo_lo_lo_hi_hi;
  assign selectReadStageMask_lo_lo_lo_hi_hi = _GEN_2;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_hi;
  assign maskSplit_maskSelect_lo_lo_lo_hi_hi = _GEN_2;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_hi_1;
  assign maskSplit_maskSelect_lo_lo_lo_hi_hi_1 = _GEN_2;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_hi_2;
  assign maskSplit_maskSelect_lo_lo_lo_hi_hi_2 = _GEN_2;
  wire [63:0]        maskForDestination_lo_lo_lo_hi_hi;
  assign maskForDestination_lo_lo_lo_hi_hi = _GEN_2;
  wire [127:0]       regroupV0_lo_lo_lo_hi = {regroupV0_lo_lo_lo_hi_hi, regroupV0_lo_lo_lo_hi_lo};
  wire [255:0]       regroupV0_lo_lo_lo = {regroupV0_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo};
  wire [63:0]        _GEN_3 = {v0_9, v0_8};
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo;
  assign regroupV0_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_1;
  assign regroupV0_lo_lo_hi_lo_lo_1 = _GEN_3;
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_2;
  assign regroupV0_lo_lo_hi_lo_lo_2 = _GEN_3;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]        selectReadStageMask_lo_lo_hi_lo_lo;
  assign selectReadStageMask_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_lo;
  assign maskSplit_maskSelect_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_lo_1;
  assign maskSplit_maskSelect_lo_lo_hi_lo_lo_1 = _GEN_3;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_lo_2;
  assign maskSplit_maskSelect_lo_lo_hi_lo_lo_2 = _GEN_3;
  wire [63:0]        maskForDestination_lo_lo_hi_lo_lo;
  assign maskForDestination_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]        _GEN_4 = {v0_11, v0_10};
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi;
  assign regroupV0_lo_lo_hi_lo_hi = _GEN_4;
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_1;
  assign regroupV0_lo_lo_hi_lo_hi_1 = _GEN_4;
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_2;
  assign regroupV0_lo_lo_hi_lo_hi_2 = _GEN_4;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi = _GEN_4;
  wire [63:0]        selectReadStageMask_lo_lo_hi_lo_hi;
  assign selectReadStageMask_lo_lo_hi_lo_hi = _GEN_4;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_hi;
  assign maskSplit_maskSelect_lo_lo_hi_lo_hi = _GEN_4;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_hi_1;
  assign maskSplit_maskSelect_lo_lo_hi_lo_hi_1 = _GEN_4;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_hi_2;
  assign maskSplit_maskSelect_lo_lo_hi_lo_hi_2 = _GEN_4;
  wire [63:0]        maskForDestination_lo_lo_hi_lo_hi;
  assign maskForDestination_lo_lo_hi_lo_hi = _GEN_4;
  wire [127:0]       regroupV0_lo_lo_hi_lo = {regroupV0_lo_lo_hi_lo_hi, regroupV0_lo_lo_hi_lo_lo};
  wire [63:0]        _GEN_5 = {v0_13, v0_12};
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo;
  assign regroupV0_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_1;
  assign regroupV0_lo_lo_hi_hi_lo_1 = _GEN_5;
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_2;
  assign regroupV0_lo_lo_hi_hi_lo_2 = _GEN_5;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]        selectReadStageMask_lo_lo_hi_hi_lo;
  assign selectReadStageMask_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_lo;
  assign maskSplit_maskSelect_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_lo_1;
  assign maskSplit_maskSelect_lo_lo_hi_hi_lo_1 = _GEN_5;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_lo_2;
  assign maskSplit_maskSelect_lo_lo_hi_hi_lo_2 = _GEN_5;
  wire [63:0]        maskForDestination_lo_lo_hi_hi_lo;
  assign maskForDestination_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]        _GEN_6 = {v0_15, v0_14};
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi;
  assign regroupV0_lo_lo_hi_hi_hi = _GEN_6;
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_1;
  assign regroupV0_lo_lo_hi_hi_hi_1 = _GEN_6;
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_2;
  assign regroupV0_lo_lo_hi_hi_hi_2 = _GEN_6;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi = _GEN_6;
  wire [63:0]        selectReadStageMask_lo_lo_hi_hi_hi;
  assign selectReadStageMask_lo_lo_hi_hi_hi = _GEN_6;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_hi;
  assign maskSplit_maskSelect_lo_lo_hi_hi_hi = _GEN_6;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_hi_1;
  assign maskSplit_maskSelect_lo_lo_hi_hi_hi_1 = _GEN_6;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_hi_2;
  assign maskSplit_maskSelect_lo_lo_hi_hi_hi_2 = _GEN_6;
  wire [63:0]        maskForDestination_lo_lo_hi_hi_hi;
  assign maskForDestination_lo_lo_hi_hi_hi = _GEN_6;
  wire [127:0]       regroupV0_lo_lo_hi_hi = {regroupV0_lo_lo_hi_hi_hi, regroupV0_lo_lo_hi_hi_lo};
  wire [255:0]       regroupV0_lo_lo_hi = {regroupV0_lo_lo_hi_hi, regroupV0_lo_lo_hi_lo};
  wire [511:0]       regroupV0_lo_lo = {regroupV0_lo_lo_hi, regroupV0_lo_lo_lo};
  wire [63:0]        _GEN_7 = {v0_17, v0_16};
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo;
  assign regroupV0_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_1;
  assign regroupV0_lo_hi_lo_lo_lo_1 = _GEN_7;
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_2;
  assign regroupV0_lo_hi_lo_lo_lo_2 = _GEN_7;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]        selectReadStageMask_lo_hi_lo_lo_lo;
  assign selectReadStageMask_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_lo;
  assign maskSplit_maskSelect_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_lo_1;
  assign maskSplit_maskSelect_lo_hi_lo_lo_lo_1 = _GEN_7;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_lo_2;
  assign maskSplit_maskSelect_lo_hi_lo_lo_lo_2 = _GEN_7;
  wire [63:0]        maskForDestination_lo_hi_lo_lo_lo;
  assign maskForDestination_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]        _GEN_8 = {v0_19, v0_18};
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi;
  assign regroupV0_lo_hi_lo_lo_hi = _GEN_8;
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_1;
  assign regroupV0_lo_hi_lo_lo_hi_1 = _GEN_8;
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_2;
  assign regroupV0_lo_hi_lo_lo_hi_2 = _GEN_8;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi = _GEN_8;
  wire [63:0]        selectReadStageMask_lo_hi_lo_lo_hi;
  assign selectReadStageMask_lo_hi_lo_lo_hi = _GEN_8;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_hi;
  assign maskSplit_maskSelect_lo_hi_lo_lo_hi = _GEN_8;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_hi_1;
  assign maskSplit_maskSelect_lo_hi_lo_lo_hi_1 = _GEN_8;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_hi_2;
  assign maskSplit_maskSelect_lo_hi_lo_lo_hi_2 = _GEN_8;
  wire [63:0]        maskForDestination_lo_hi_lo_lo_hi;
  assign maskForDestination_lo_hi_lo_lo_hi = _GEN_8;
  wire [127:0]       regroupV0_lo_hi_lo_lo = {regroupV0_lo_hi_lo_lo_hi, regroupV0_lo_hi_lo_lo_lo};
  wire [63:0]        _GEN_9 = {v0_21, v0_20};
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo;
  assign regroupV0_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_1;
  assign regroupV0_lo_hi_lo_hi_lo_1 = _GEN_9;
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_2;
  assign regroupV0_lo_hi_lo_hi_lo_2 = _GEN_9;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]        selectReadStageMask_lo_hi_lo_hi_lo;
  assign selectReadStageMask_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_lo;
  assign maskSplit_maskSelect_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_lo_1;
  assign maskSplit_maskSelect_lo_hi_lo_hi_lo_1 = _GEN_9;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_lo_2;
  assign maskSplit_maskSelect_lo_hi_lo_hi_lo_2 = _GEN_9;
  wire [63:0]        maskForDestination_lo_hi_lo_hi_lo;
  assign maskForDestination_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]        _GEN_10 = {v0_23, v0_22};
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi;
  assign regroupV0_lo_hi_lo_hi_hi = _GEN_10;
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_1;
  assign regroupV0_lo_hi_lo_hi_hi_1 = _GEN_10;
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_2;
  assign regroupV0_lo_hi_lo_hi_hi_2 = _GEN_10;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi = _GEN_10;
  wire [63:0]        selectReadStageMask_lo_hi_lo_hi_hi;
  assign selectReadStageMask_lo_hi_lo_hi_hi = _GEN_10;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_hi;
  assign maskSplit_maskSelect_lo_hi_lo_hi_hi = _GEN_10;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_hi_1;
  assign maskSplit_maskSelect_lo_hi_lo_hi_hi_1 = _GEN_10;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_hi_2;
  assign maskSplit_maskSelect_lo_hi_lo_hi_hi_2 = _GEN_10;
  wire [63:0]        maskForDestination_lo_hi_lo_hi_hi;
  assign maskForDestination_lo_hi_lo_hi_hi = _GEN_10;
  wire [127:0]       regroupV0_lo_hi_lo_hi = {regroupV0_lo_hi_lo_hi_hi, regroupV0_lo_hi_lo_hi_lo};
  wire [255:0]       regroupV0_lo_hi_lo = {regroupV0_lo_hi_lo_hi, regroupV0_lo_hi_lo_lo};
  wire [63:0]        _GEN_11 = {v0_25, v0_24};
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo;
  assign regroupV0_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_1;
  assign regroupV0_lo_hi_hi_lo_lo_1 = _GEN_11;
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_2;
  assign regroupV0_lo_hi_hi_lo_lo_2 = _GEN_11;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]        selectReadStageMask_lo_hi_hi_lo_lo;
  assign selectReadStageMask_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_lo;
  assign maskSplit_maskSelect_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_lo_1;
  assign maskSplit_maskSelect_lo_hi_hi_lo_lo_1 = _GEN_11;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_lo_2;
  assign maskSplit_maskSelect_lo_hi_hi_lo_lo_2 = _GEN_11;
  wire [63:0]        maskForDestination_lo_hi_hi_lo_lo;
  assign maskForDestination_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]        _GEN_12 = {v0_27, v0_26};
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi;
  assign regroupV0_lo_hi_hi_lo_hi = _GEN_12;
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_1;
  assign regroupV0_lo_hi_hi_lo_hi_1 = _GEN_12;
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_2;
  assign regroupV0_lo_hi_hi_lo_hi_2 = _GEN_12;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi = _GEN_12;
  wire [63:0]        selectReadStageMask_lo_hi_hi_lo_hi;
  assign selectReadStageMask_lo_hi_hi_lo_hi = _GEN_12;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_hi;
  assign maskSplit_maskSelect_lo_hi_hi_lo_hi = _GEN_12;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_hi_1;
  assign maskSplit_maskSelect_lo_hi_hi_lo_hi_1 = _GEN_12;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_hi_2;
  assign maskSplit_maskSelect_lo_hi_hi_lo_hi_2 = _GEN_12;
  wire [63:0]        maskForDestination_lo_hi_hi_lo_hi;
  assign maskForDestination_lo_hi_hi_lo_hi = _GEN_12;
  wire [127:0]       regroupV0_lo_hi_hi_lo = {regroupV0_lo_hi_hi_lo_hi, regroupV0_lo_hi_hi_lo_lo};
  wire [63:0]        _GEN_13 = {v0_29, v0_28};
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo;
  assign regroupV0_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_1;
  assign regroupV0_lo_hi_hi_hi_lo_1 = _GEN_13;
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_2;
  assign regroupV0_lo_hi_hi_hi_lo_2 = _GEN_13;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]        selectReadStageMask_lo_hi_hi_hi_lo;
  assign selectReadStageMask_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_lo;
  assign maskSplit_maskSelect_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_lo_1;
  assign maskSplit_maskSelect_lo_hi_hi_hi_lo_1 = _GEN_13;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_lo_2;
  assign maskSplit_maskSelect_lo_hi_hi_hi_lo_2 = _GEN_13;
  wire [63:0]        maskForDestination_lo_hi_hi_hi_lo;
  assign maskForDestination_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]        _GEN_14 = {v0_31, v0_30};
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi;
  assign regroupV0_lo_hi_hi_hi_hi = _GEN_14;
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_1;
  assign regroupV0_lo_hi_hi_hi_hi_1 = _GEN_14;
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_2;
  assign regroupV0_lo_hi_hi_hi_hi_2 = _GEN_14;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi = _GEN_14;
  wire [63:0]        selectReadStageMask_lo_hi_hi_hi_hi;
  assign selectReadStageMask_lo_hi_hi_hi_hi = _GEN_14;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_hi;
  assign maskSplit_maskSelect_lo_hi_hi_hi_hi = _GEN_14;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_hi_1;
  assign maskSplit_maskSelect_lo_hi_hi_hi_hi_1 = _GEN_14;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_hi_2;
  assign maskSplit_maskSelect_lo_hi_hi_hi_hi_2 = _GEN_14;
  wire [63:0]        maskForDestination_lo_hi_hi_hi_hi;
  assign maskForDestination_lo_hi_hi_hi_hi = _GEN_14;
  wire [127:0]       regroupV0_lo_hi_hi_hi = {regroupV0_lo_hi_hi_hi_hi, regroupV0_lo_hi_hi_hi_lo};
  wire [255:0]       regroupV0_lo_hi_hi = {regroupV0_lo_hi_hi_hi, regroupV0_lo_hi_hi_lo};
  wire [511:0]       regroupV0_lo_hi = {regroupV0_lo_hi_hi, regroupV0_lo_hi_lo};
  wire [1023:0]      regroupV0_lo = {regroupV0_lo_hi, regroupV0_lo_lo};
  wire [63:0]        _GEN_15 = {v0_33, v0_32};
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo;
  assign regroupV0_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_1;
  assign regroupV0_hi_lo_lo_lo_lo_1 = _GEN_15;
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_2;
  assign regroupV0_hi_lo_lo_lo_lo_2 = _GEN_15;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]        selectReadStageMask_hi_lo_lo_lo_lo;
  assign selectReadStageMask_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_lo;
  assign maskSplit_maskSelect_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_lo_1;
  assign maskSplit_maskSelect_hi_lo_lo_lo_lo_1 = _GEN_15;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_lo_2;
  assign maskSplit_maskSelect_hi_lo_lo_lo_lo_2 = _GEN_15;
  wire [63:0]        maskForDestination_hi_lo_lo_lo_lo;
  assign maskForDestination_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]        _GEN_16 = {v0_35, v0_34};
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi;
  assign regroupV0_hi_lo_lo_lo_hi = _GEN_16;
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_1;
  assign regroupV0_hi_lo_lo_lo_hi_1 = _GEN_16;
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_2;
  assign regroupV0_hi_lo_lo_lo_hi_2 = _GEN_16;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi = _GEN_16;
  wire [63:0]        selectReadStageMask_hi_lo_lo_lo_hi;
  assign selectReadStageMask_hi_lo_lo_lo_hi = _GEN_16;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_hi;
  assign maskSplit_maskSelect_hi_lo_lo_lo_hi = _GEN_16;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_hi_1;
  assign maskSplit_maskSelect_hi_lo_lo_lo_hi_1 = _GEN_16;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_hi_2;
  assign maskSplit_maskSelect_hi_lo_lo_lo_hi_2 = _GEN_16;
  wire [63:0]        maskForDestination_hi_lo_lo_lo_hi;
  assign maskForDestination_hi_lo_lo_lo_hi = _GEN_16;
  wire [127:0]       regroupV0_hi_lo_lo_lo = {regroupV0_hi_lo_lo_lo_hi, regroupV0_hi_lo_lo_lo_lo};
  wire [63:0]        _GEN_17 = {v0_37, v0_36};
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo;
  assign regroupV0_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_1;
  assign regroupV0_hi_lo_lo_hi_lo_1 = _GEN_17;
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_2;
  assign regroupV0_hi_lo_lo_hi_lo_2 = _GEN_17;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]        selectReadStageMask_hi_lo_lo_hi_lo;
  assign selectReadStageMask_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_lo;
  assign maskSplit_maskSelect_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_lo_1;
  assign maskSplit_maskSelect_hi_lo_lo_hi_lo_1 = _GEN_17;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_lo_2;
  assign maskSplit_maskSelect_hi_lo_lo_hi_lo_2 = _GEN_17;
  wire [63:0]        maskForDestination_hi_lo_lo_hi_lo;
  assign maskForDestination_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]        _GEN_18 = {v0_39, v0_38};
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi;
  assign regroupV0_hi_lo_lo_hi_hi = _GEN_18;
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_1;
  assign regroupV0_hi_lo_lo_hi_hi_1 = _GEN_18;
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_2;
  assign regroupV0_hi_lo_lo_hi_hi_2 = _GEN_18;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi = _GEN_18;
  wire [63:0]        selectReadStageMask_hi_lo_lo_hi_hi;
  assign selectReadStageMask_hi_lo_lo_hi_hi = _GEN_18;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_hi;
  assign maskSplit_maskSelect_hi_lo_lo_hi_hi = _GEN_18;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_hi_1;
  assign maskSplit_maskSelect_hi_lo_lo_hi_hi_1 = _GEN_18;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_hi_2;
  assign maskSplit_maskSelect_hi_lo_lo_hi_hi_2 = _GEN_18;
  wire [63:0]        maskForDestination_hi_lo_lo_hi_hi;
  assign maskForDestination_hi_lo_lo_hi_hi = _GEN_18;
  wire [127:0]       regroupV0_hi_lo_lo_hi = {regroupV0_hi_lo_lo_hi_hi, regroupV0_hi_lo_lo_hi_lo};
  wire [255:0]       regroupV0_hi_lo_lo = {regroupV0_hi_lo_lo_hi, regroupV0_hi_lo_lo_lo};
  wire [63:0]        _GEN_19 = {v0_41, v0_40};
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo;
  assign regroupV0_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_1;
  assign regroupV0_hi_lo_hi_lo_lo_1 = _GEN_19;
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_2;
  assign regroupV0_hi_lo_hi_lo_lo_2 = _GEN_19;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]        selectReadStageMask_hi_lo_hi_lo_lo;
  assign selectReadStageMask_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_lo;
  assign maskSplit_maskSelect_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_lo_1;
  assign maskSplit_maskSelect_hi_lo_hi_lo_lo_1 = _GEN_19;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_lo_2;
  assign maskSplit_maskSelect_hi_lo_hi_lo_lo_2 = _GEN_19;
  wire [63:0]        maskForDestination_hi_lo_hi_lo_lo;
  assign maskForDestination_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]        _GEN_20 = {v0_43, v0_42};
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi;
  assign regroupV0_hi_lo_hi_lo_hi = _GEN_20;
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_1;
  assign regroupV0_hi_lo_hi_lo_hi_1 = _GEN_20;
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_2;
  assign regroupV0_hi_lo_hi_lo_hi_2 = _GEN_20;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi = _GEN_20;
  wire [63:0]        selectReadStageMask_hi_lo_hi_lo_hi;
  assign selectReadStageMask_hi_lo_hi_lo_hi = _GEN_20;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_hi;
  assign maskSplit_maskSelect_hi_lo_hi_lo_hi = _GEN_20;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_hi_1;
  assign maskSplit_maskSelect_hi_lo_hi_lo_hi_1 = _GEN_20;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_hi_2;
  assign maskSplit_maskSelect_hi_lo_hi_lo_hi_2 = _GEN_20;
  wire [63:0]        maskForDestination_hi_lo_hi_lo_hi;
  assign maskForDestination_hi_lo_hi_lo_hi = _GEN_20;
  wire [127:0]       regroupV0_hi_lo_hi_lo = {regroupV0_hi_lo_hi_lo_hi, regroupV0_hi_lo_hi_lo_lo};
  wire [63:0]        _GEN_21 = {v0_45, v0_44};
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo;
  assign regroupV0_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_1;
  assign regroupV0_hi_lo_hi_hi_lo_1 = _GEN_21;
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_2;
  assign regroupV0_hi_lo_hi_hi_lo_2 = _GEN_21;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]        selectReadStageMask_hi_lo_hi_hi_lo;
  assign selectReadStageMask_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_lo;
  assign maskSplit_maskSelect_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_lo_1;
  assign maskSplit_maskSelect_hi_lo_hi_hi_lo_1 = _GEN_21;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_lo_2;
  assign maskSplit_maskSelect_hi_lo_hi_hi_lo_2 = _GEN_21;
  wire [63:0]        maskForDestination_hi_lo_hi_hi_lo;
  assign maskForDestination_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]        _GEN_22 = {v0_47, v0_46};
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi;
  assign regroupV0_hi_lo_hi_hi_hi = _GEN_22;
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_1;
  assign regroupV0_hi_lo_hi_hi_hi_1 = _GEN_22;
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_2;
  assign regroupV0_hi_lo_hi_hi_hi_2 = _GEN_22;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi = _GEN_22;
  wire [63:0]        selectReadStageMask_hi_lo_hi_hi_hi;
  assign selectReadStageMask_hi_lo_hi_hi_hi = _GEN_22;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_hi;
  assign maskSplit_maskSelect_hi_lo_hi_hi_hi = _GEN_22;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_hi_1;
  assign maskSplit_maskSelect_hi_lo_hi_hi_hi_1 = _GEN_22;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_hi_2;
  assign maskSplit_maskSelect_hi_lo_hi_hi_hi_2 = _GEN_22;
  wire [63:0]        maskForDestination_hi_lo_hi_hi_hi;
  assign maskForDestination_hi_lo_hi_hi_hi = _GEN_22;
  wire [127:0]       regroupV0_hi_lo_hi_hi = {regroupV0_hi_lo_hi_hi_hi, regroupV0_hi_lo_hi_hi_lo};
  wire [255:0]       regroupV0_hi_lo_hi = {regroupV0_hi_lo_hi_hi, regroupV0_hi_lo_hi_lo};
  wire [511:0]       regroupV0_hi_lo = {regroupV0_hi_lo_hi, regroupV0_hi_lo_lo};
  wire [63:0]        _GEN_23 = {v0_49, v0_48};
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo;
  assign regroupV0_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_1;
  assign regroupV0_hi_hi_lo_lo_lo_1 = _GEN_23;
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_2;
  assign regroupV0_hi_hi_lo_lo_lo_2 = _GEN_23;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]        selectReadStageMask_hi_hi_lo_lo_lo;
  assign selectReadStageMask_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_lo;
  assign maskSplit_maskSelect_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_lo_1;
  assign maskSplit_maskSelect_hi_hi_lo_lo_lo_1 = _GEN_23;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_lo_2;
  assign maskSplit_maskSelect_hi_hi_lo_lo_lo_2 = _GEN_23;
  wire [63:0]        maskForDestination_hi_hi_lo_lo_lo;
  assign maskForDestination_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]        _GEN_24 = {v0_51, v0_50};
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi;
  assign regroupV0_hi_hi_lo_lo_hi = _GEN_24;
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_1;
  assign regroupV0_hi_hi_lo_lo_hi_1 = _GEN_24;
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_2;
  assign regroupV0_hi_hi_lo_lo_hi_2 = _GEN_24;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi = _GEN_24;
  wire [63:0]        selectReadStageMask_hi_hi_lo_lo_hi;
  assign selectReadStageMask_hi_hi_lo_lo_hi = _GEN_24;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_hi;
  assign maskSplit_maskSelect_hi_hi_lo_lo_hi = _GEN_24;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_hi_1;
  assign maskSplit_maskSelect_hi_hi_lo_lo_hi_1 = _GEN_24;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_hi_2;
  assign maskSplit_maskSelect_hi_hi_lo_lo_hi_2 = _GEN_24;
  wire [63:0]        maskForDestination_hi_hi_lo_lo_hi;
  assign maskForDestination_hi_hi_lo_lo_hi = _GEN_24;
  wire [127:0]       regroupV0_hi_hi_lo_lo = {regroupV0_hi_hi_lo_lo_hi, regroupV0_hi_hi_lo_lo_lo};
  wire [63:0]        _GEN_25 = {v0_53, v0_52};
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo;
  assign regroupV0_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_1;
  assign regroupV0_hi_hi_lo_hi_lo_1 = _GEN_25;
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_2;
  assign regroupV0_hi_hi_lo_hi_lo_2 = _GEN_25;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]        selectReadStageMask_hi_hi_lo_hi_lo;
  assign selectReadStageMask_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_lo;
  assign maskSplit_maskSelect_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_lo_1;
  assign maskSplit_maskSelect_hi_hi_lo_hi_lo_1 = _GEN_25;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_lo_2;
  assign maskSplit_maskSelect_hi_hi_lo_hi_lo_2 = _GEN_25;
  wire [63:0]        maskForDestination_hi_hi_lo_hi_lo;
  assign maskForDestination_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]        _GEN_26 = {v0_55, v0_54};
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi;
  assign regroupV0_hi_hi_lo_hi_hi = _GEN_26;
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_1;
  assign regroupV0_hi_hi_lo_hi_hi_1 = _GEN_26;
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_2;
  assign regroupV0_hi_hi_lo_hi_hi_2 = _GEN_26;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi = _GEN_26;
  wire [63:0]        selectReadStageMask_hi_hi_lo_hi_hi;
  assign selectReadStageMask_hi_hi_lo_hi_hi = _GEN_26;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_hi;
  assign maskSplit_maskSelect_hi_hi_lo_hi_hi = _GEN_26;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_hi_1;
  assign maskSplit_maskSelect_hi_hi_lo_hi_hi_1 = _GEN_26;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_hi_2;
  assign maskSplit_maskSelect_hi_hi_lo_hi_hi_2 = _GEN_26;
  wire [63:0]        maskForDestination_hi_hi_lo_hi_hi;
  assign maskForDestination_hi_hi_lo_hi_hi = _GEN_26;
  wire [127:0]       regroupV0_hi_hi_lo_hi = {regroupV0_hi_hi_lo_hi_hi, regroupV0_hi_hi_lo_hi_lo};
  wire [255:0]       regroupV0_hi_hi_lo = {regroupV0_hi_hi_lo_hi, regroupV0_hi_hi_lo_lo};
  wire [63:0]        _GEN_27 = {v0_57, v0_56};
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo;
  assign regroupV0_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_1;
  assign regroupV0_hi_hi_hi_lo_lo_1 = _GEN_27;
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_2;
  assign regroupV0_hi_hi_hi_lo_lo_2 = _GEN_27;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]        selectReadStageMask_hi_hi_hi_lo_lo;
  assign selectReadStageMask_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_lo;
  assign maskSplit_maskSelect_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_lo_1;
  assign maskSplit_maskSelect_hi_hi_hi_lo_lo_1 = _GEN_27;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_lo_2;
  assign maskSplit_maskSelect_hi_hi_hi_lo_lo_2 = _GEN_27;
  wire [63:0]        maskForDestination_hi_hi_hi_lo_lo;
  assign maskForDestination_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]        _GEN_28 = {v0_59, v0_58};
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi;
  assign regroupV0_hi_hi_hi_lo_hi = _GEN_28;
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_1;
  assign regroupV0_hi_hi_hi_lo_hi_1 = _GEN_28;
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_2;
  assign regroupV0_hi_hi_hi_lo_hi_2 = _GEN_28;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi = _GEN_28;
  wire [63:0]        selectReadStageMask_hi_hi_hi_lo_hi;
  assign selectReadStageMask_hi_hi_hi_lo_hi = _GEN_28;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_hi;
  assign maskSplit_maskSelect_hi_hi_hi_lo_hi = _GEN_28;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_hi_1;
  assign maskSplit_maskSelect_hi_hi_hi_lo_hi_1 = _GEN_28;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_hi_2;
  assign maskSplit_maskSelect_hi_hi_hi_lo_hi_2 = _GEN_28;
  wire [63:0]        maskForDestination_hi_hi_hi_lo_hi;
  assign maskForDestination_hi_hi_hi_lo_hi = _GEN_28;
  wire [127:0]       regroupV0_hi_hi_hi_lo = {regroupV0_hi_hi_hi_lo_hi, regroupV0_hi_hi_hi_lo_lo};
  wire [63:0]        _GEN_29 = {v0_61, v0_60};
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo;
  assign regroupV0_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_1;
  assign regroupV0_hi_hi_hi_hi_lo_1 = _GEN_29;
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_2;
  assign regroupV0_hi_hi_hi_hi_lo_2 = _GEN_29;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]        selectReadStageMask_hi_hi_hi_hi_lo;
  assign selectReadStageMask_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_lo;
  assign maskSplit_maskSelect_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_lo_1;
  assign maskSplit_maskSelect_hi_hi_hi_hi_lo_1 = _GEN_29;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_lo_2;
  assign maskSplit_maskSelect_hi_hi_hi_hi_lo_2 = _GEN_29;
  wire [63:0]        maskForDestination_hi_hi_hi_hi_lo;
  assign maskForDestination_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]        _GEN_30 = {v0_63, v0_62};
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi;
  assign regroupV0_hi_hi_hi_hi_hi = _GEN_30;
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_1;
  assign regroupV0_hi_hi_hi_hi_hi_1 = _GEN_30;
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_2;
  assign regroupV0_hi_hi_hi_hi_hi_2 = _GEN_30;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi = _GEN_30;
  wire [63:0]        selectReadStageMask_hi_hi_hi_hi_hi;
  assign selectReadStageMask_hi_hi_hi_hi_hi = _GEN_30;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_hi;
  assign maskSplit_maskSelect_hi_hi_hi_hi_hi = _GEN_30;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_hi_1;
  assign maskSplit_maskSelect_hi_hi_hi_hi_hi_1 = _GEN_30;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_hi_2;
  assign maskSplit_maskSelect_hi_hi_hi_hi_hi_2 = _GEN_30;
  wire [63:0]        maskForDestination_hi_hi_hi_hi_hi;
  assign maskForDestination_hi_hi_hi_hi_hi = _GEN_30;
  wire [127:0]       regroupV0_hi_hi_hi_hi = {regroupV0_hi_hi_hi_hi_hi, regroupV0_hi_hi_hi_hi_lo};
  wire [255:0]       regroupV0_hi_hi_hi = {regroupV0_hi_hi_hi_hi, regroupV0_hi_hi_hi_lo};
  wire [511:0]       regroupV0_hi_hi = {regroupV0_hi_hi_hi, regroupV0_hi_hi_lo};
  wire [1023:0]      regroupV0_hi = {regroupV0_hi_hi, regroupV0_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_1 = {regroupV0_lo[131:128], regroupV0_lo[3:0]};
  wire [7:0]         regroupV0_lo_lo_hi_1 = {regroupV0_lo[387:384], regroupV0_lo[259:256]};
  wire [15:0]        regroupV0_lo_lo_1 = {regroupV0_lo_lo_hi_1, regroupV0_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_1 = {regroupV0_lo[643:640], regroupV0_lo[515:512]};
  wire [7:0]         regroupV0_lo_hi_hi_1 = {regroupV0_lo[899:896], regroupV0_lo[771:768]};
  wire [15:0]        regroupV0_lo_hi_1 = {regroupV0_lo_hi_hi_1, regroupV0_lo_hi_lo_1};
  wire [31:0]        regroupV0_lo_1 = {regroupV0_lo_hi_1, regroupV0_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_1 = {regroupV0_hi[131:128], regroupV0_hi[3:0]};
  wire [7:0]         regroupV0_hi_lo_hi_1 = {regroupV0_hi[387:384], regroupV0_hi[259:256]};
  wire [15:0]        regroupV0_hi_lo_1 = {regroupV0_hi_lo_hi_1, regroupV0_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_1 = {regroupV0_hi[643:640], regroupV0_hi[515:512]};
  wire [7:0]         regroupV0_hi_hi_hi_1 = {regroupV0_hi[899:896], regroupV0_hi[771:768]};
  wire [15:0]        regroupV0_hi_hi_1 = {regroupV0_hi_hi_hi_1, regroupV0_hi_hi_lo_1};
  wire [31:0]        regroupV0_hi_1 = {regroupV0_hi_hi_1, regroupV0_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_2 = {regroupV0_lo[135:132], regroupV0_lo[7:4]};
  wire [7:0]         regroupV0_lo_lo_hi_2 = {regroupV0_lo[391:388], regroupV0_lo[263:260]};
  wire [15:0]        regroupV0_lo_lo_2 = {regroupV0_lo_lo_hi_2, regroupV0_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_2 = {regroupV0_lo[647:644], regroupV0_lo[519:516]};
  wire [7:0]         regroupV0_lo_hi_hi_2 = {regroupV0_lo[903:900], regroupV0_lo[775:772]};
  wire [15:0]        regroupV0_lo_hi_2 = {regroupV0_lo_hi_hi_2, regroupV0_lo_hi_lo_2};
  wire [31:0]        regroupV0_lo_2 = {regroupV0_lo_hi_2, regroupV0_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_2 = {regroupV0_hi[135:132], regroupV0_hi[7:4]};
  wire [7:0]         regroupV0_hi_lo_hi_2 = {regroupV0_hi[391:388], regroupV0_hi[263:260]};
  wire [15:0]        regroupV0_hi_lo_2 = {regroupV0_hi_lo_hi_2, regroupV0_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_2 = {regroupV0_hi[647:644], regroupV0_hi[519:516]};
  wire [7:0]         regroupV0_hi_hi_hi_2 = {regroupV0_hi[903:900], regroupV0_hi[775:772]};
  wire [15:0]        regroupV0_hi_hi_2 = {regroupV0_hi_hi_hi_2, regroupV0_hi_hi_lo_2};
  wire [31:0]        regroupV0_hi_2 = {regroupV0_hi_hi_2, regroupV0_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_3 = {regroupV0_lo[139:136], regroupV0_lo[11:8]};
  wire [7:0]         regroupV0_lo_lo_hi_3 = {regroupV0_lo[395:392], regroupV0_lo[267:264]};
  wire [15:0]        regroupV0_lo_lo_3 = {regroupV0_lo_lo_hi_3, regroupV0_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_3 = {regroupV0_lo[651:648], regroupV0_lo[523:520]};
  wire [7:0]         regroupV0_lo_hi_hi_3 = {regroupV0_lo[907:904], regroupV0_lo[779:776]};
  wire [15:0]        regroupV0_lo_hi_3 = {regroupV0_lo_hi_hi_3, regroupV0_lo_hi_lo_3};
  wire [31:0]        regroupV0_lo_3 = {regroupV0_lo_hi_3, regroupV0_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_3 = {regroupV0_hi[139:136], regroupV0_hi[11:8]};
  wire [7:0]         regroupV0_hi_lo_hi_3 = {regroupV0_hi[395:392], regroupV0_hi[267:264]};
  wire [15:0]        regroupV0_hi_lo_3 = {regroupV0_hi_lo_hi_3, regroupV0_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_3 = {regroupV0_hi[651:648], regroupV0_hi[523:520]};
  wire [7:0]         regroupV0_hi_hi_hi_3 = {regroupV0_hi[907:904], regroupV0_hi[779:776]};
  wire [15:0]        regroupV0_hi_hi_3 = {regroupV0_hi_hi_hi_3, regroupV0_hi_hi_lo_3};
  wire [31:0]        regroupV0_hi_3 = {regroupV0_hi_hi_3, regroupV0_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_4 = {regroupV0_lo[143:140], regroupV0_lo[15:12]};
  wire [7:0]         regroupV0_lo_lo_hi_4 = {regroupV0_lo[399:396], regroupV0_lo[271:268]};
  wire [15:0]        regroupV0_lo_lo_4 = {regroupV0_lo_lo_hi_4, regroupV0_lo_lo_lo_4};
  wire [7:0]         regroupV0_lo_hi_lo_4 = {regroupV0_lo[655:652], regroupV0_lo[527:524]};
  wire [7:0]         regroupV0_lo_hi_hi_4 = {regroupV0_lo[911:908], regroupV0_lo[783:780]};
  wire [15:0]        regroupV0_lo_hi_4 = {regroupV0_lo_hi_hi_4, regroupV0_lo_hi_lo_4};
  wire [31:0]        regroupV0_lo_4 = {regroupV0_lo_hi_4, regroupV0_lo_lo_4};
  wire [7:0]         regroupV0_hi_lo_lo_4 = {regroupV0_hi[143:140], regroupV0_hi[15:12]};
  wire [7:0]         regroupV0_hi_lo_hi_4 = {regroupV0_hi[399:396], regroupV0_hi[271:268]};
  wire [15:0]        regroupV0_hi_lo_4 = {regroupV0_hi_lo_hi_4, regroupV0_hi_lo_lo_4};
  wire [7:0]         regroupV0_hi_hi_lo_4 = {regroupV0_hi[655:652], regroupV0_hi[527:524]};
  wire [7:0]         regroupV0_hi_hi_hi_4 = {regroupV0_hi[911:908], regroupV0_hi[783:780]};
  wire [15:0]        regroupV0_hi_hi_4 = {regroupV0_hi_hi_hi_4, regroupV0_hi_hi_lo_4};
  wire [31:0]        regroupV0_hi_4 = {regroupV0_hi_hi_4, regroupV0_hi_lo_4};
  wire [7:0]         regroupV0_lo_lo_lo_5 = {regroupV0_lo[147:144], regroupV0_lo[19:16]};
  wire [7:0]         regroupV0_lo_lo_hi_5 = {regroupV0_lo[403:400], regroupV0_lo[275:272]};
  wire [15:0]        regroupV0_lo_lo_5 = {regroupV0_lo_lo_hi_5, regroupV0_lo_lo_lo_5};
  wire [7:0]         regroupV0_lo_hi_lo_5 = {regroupV0_lo[659:656], regroupV0_lo[531:528]};
  wire [7:0]         regroupV0_lo_hi_hi_5 = {regroupV0_lo[915:912], regroupV0_lo[787:784]};
  wire [15:0]        regroupV0_lo_hi_5 = {regroupV0_lo_hi_hi_5, regroupV0_lo_hi_lo_5};
  wire [31:0]        regroupV0_lo_5 = {regroupV0_lo_hi_5, regroupV0_lo_lo_5};
  wire [7:0]         regroupV0_hi_lo_lo_5 = {regroupV0_hi[147:144], regroupV0_hi[19:16]};
  wire [7:0]         regroupV0_hi_lo_hi_5 = {regroupV0_hi[403:400], regroupV0_hi[275:272]};
  wire [15:0]        regroupV0_hi_lo_5 = {regroupV0_hi_lo_hi_5, regroupV0_hi_lo_lo_5};
  wire [7:0]         regroupV0_hi_hi_lo_5 = {regroupV0_hi[659:656], regroupV0_hi[531:528]};
  wire [7:0]         regroupV0_hi_hi_hi_5 = {regroupV0_hi[915:912], regroupV0_hi[787:784]};
  wire [15:0]        regroupV0_hi_hi_5 = {regroupV0_hi_hi_hi_5, regroupV0_hi_hi_lo_5};
  wire [31:0]        regroupV0_hi_5 = {regroupV0_hi_hi_5, regroupV0_hi_lo_5};
  wire [7:0]         regroupV0_lo_lo_lo_6 = {regroupV0_lo[151:148], regroupV0_lo[23:20]};
  wire [7:0]         regroupV0_lo_lo_hi_6 = {regroupV0_lo[407:404], regroupV0_lo[279:276]};
  wire [15:0]        regroupV0_lo_lo_6 = {regroupV0_lo_lo_hi_6, regroupV0_lo_lo_lo_6};
  wire [7:0]         regroupV0_lo_hi_lo_6 = {regroupV0_lo[663:660], regroupV0_lo[535:532]};
  wire [7:0]         regroupV0_lo_hi_hi_6 = {regroupV0_lo[919:916], regroupV0_lo[791:788]};
  wire [15:0]        regroupV0_lo_hi_6 = {regroupV0_lo_hi_hi_6, regroupV0_lo_hi_lo_6};
  wire [31:0]        regroupV0_lo_6 = {regroupV0_lo_hi_6, regroupV0_lo_lo_6};
  wire [7:0]         regroupV0_hi_lo_lo_6 = {regroupV0_hi[151:148], regroupV0_hi[23:20]};
  wire [7:0]         regroupV0_hi_lo_hi_6 = {regroupV0_hi[407:404], regroupV0_hi[279:276]};
  wire [15:0]        regroupV0_hi_lo_6 = {regroupV0_hi_lo_hi_6, regroupV0_hi_lo_lo_6};
  wire [7:0]         regroupV0_hi_hi_lo_6 = {regroupV0_hi[663:660], regroupV0_hi[535:532]};
  wire [7:0]         regroupV0_hi_hi_hi_6 = {regroupV0_hi[919:916], regroupV0_hi[791:788]};
  wire [15:0]        regroupV0_hi_hi_6 = {regroupV0_hi_hi_hi_6, regroupV0_hi_hi_lo_6};
  wire [31:0]        regroupV0_hi_6 = {regroupV0_hi_hi_6, regroupV0_hi_lo_6};
  wire [7:0]         regroupV0_lo_lo_lo_7 = {regroupV0_lo[155:152], regroupV0_lo[27:24]};
  wire [7:0]         regroupV0_lo_lo_hi_7 = {regroupV0_lo[411:408], regroupV0_lo[283:280]};
  wire [15:0]        regroupV0_lo_lo_7 = {regroupV0_lo_lo_hi_7, regroupV0_lo_lo_lo_7};
  wire [7:0]         regroupV0_lo_hi_lo_7 = {regroupV0_lo[667:664], regroupV0_lo[539:536]};
  wire [7:0]         regroupV0_lo_hi_hi_7 = {regroupV0_lo[923:920], regroupV0_lo[795:792]};
  wire [15:0]        regroupV0_lo_hi_7 = {regroupV0_lo_hi_hi_7, regroupV0_lo_hi_lo_7};
  wire [31:0]        regroupV0_lo_7 = {regroupV0_lo_hi_7, regroupV0_lo_lo_7};
  wire [7:0]         regroupV0_hi_lo_lo_7 = {regroupV0_hi[155:152], regroupV0_hi[27:24]};
  wire [7:0]         regroupV0_hi_lo_hi_7 = {regroupV0_hi[411:408], regroupV0_hi[283:280]};
  wire [15:0]        regroupV0_hi_lo_7 = {regroupV0_hi_lo_hi_7, regroupV0_hi_lo_lo_7};
  wire [7:0]         regroupV0_hi_hi_lo_7 = {regroupV0_hi[667:664], regroupV0_hi[539:536]};
  wire [7:0]         regroupV0_hi_hi_hi_7 = {regroupV0_hi[923:920], regroupV0_hi[795:792]};
  wire [15:0]        regroupV0_hi_hi_7 = {regroupV0_hi_hi_hi_7, regroupV0_hi_hi_lo_7};
  wire [31:0]        regroupV0_hi_7 = {regroupV0_hi_hi_7, regroupV0_hi_lo_7};
  wire [7:0]         regroupV0_lo_lo_lo_8 = {regroupV0_lo[159:156], regroupV0_lo[31:28]};
  wire [7:0]         regroupV0_lo_lo_hi_8 = {regroupV0_lo[415:412], regroupV0_lo[287:284]};
  wire [15:0]        regroupV0_lo_lo_8 = {regroupV0_lo_lo_hi_8, regroupV0_lo_lo_lo_8};
  wire [7:0]         regroupV0_lo_hi_lo_8 = {regroupV0_lo[671:668], regroupV0_lo[543:540]};
  wire [7:0]         regroupV0_lo_hi_hi_8 = {regroupV0_lo[927:924], regroupV0_lo[799:796]};
  wire [15:0]        regroupV0_lo_hi_8 = {regroupV0_lo_hi_hi_8, regroupV0_lo_hi_lo_8};
  wire [31:0]        regroupV0_lo_8 = {regroupV0_lo_hi_8, regroupV0_lo_lo_8};
  wire [7:0]         regroupV0_hi_lo_lo_8 = {regroupV0_hi[159:156], regroupV0_hi[31:28]};
  wire [7:0]         regroupV0_hi_lo_hi_8 = {regroupV0_hi[415:412], regroupV0_hi[287:284]};
  wire [15:0]        regroupV0_hi_lo_8 = {regroupV0_hi_lo_hi_8, regroupV0_hi_lo_lo_8};
  wire [7:0]         regroupV0_hi_hi_lo_8 = {regroupV0_hi[671:668], regroupV0_hi[543:540]};
  wire [7:0]         regroupV0_hi_hi_hi_8 = {regroupV0_hi[927:924], regroupV0_hi[799:796]};
  wire [15:0]        regroupV0_hi_hi_8 = {regroupV0_hi_hi_hi_8, regroupV0_hi_hi_lo_8};
  wire [31:0]        regroupV0_hi_8 = {regroupV0_hi_hi_8, regroupV0_hi_lo_8};
  wire [7:0]         regroupV0_lo_lo_lo_9 = {regroupV0_lo[163:160], regroupV0_lo[35:32]};
  wire [7:0]         regroupV0_lo_lo_hi_9 = {regroupV0_lo[419:416], regroupV0_lo[291:288]};
  wire [15:0]        regroupV0_lo_lo_9 = {regroupV0_lo_lo_hi_9, regroupV0_lo_lo_lo_9};
  wire [7:0]         regroupV0_lo_hi_lo_9 = {regroupV0_lo[675:672], regroupV0_lo[547:544]};
  wire [7:0]         regroupV0_lo_hi_hi_9 = {regroupV0_lo[931:928], regroupV0_lo[803:800]};
  wire [15:0]        regroupV0_lo_hi_9 = {regroupV0_lo_hi_hi_9, regroupV0_lo_hi_lo_9};
  wire [31:0]        regroupV0_lo_9 = {regroupV0_lo_hi_9, regroupV0_lo_lo_9};
  wire [7:0]         regroupV0_hi_lo_lo_9 = {regroupV0_hi[163:160], regroupV0_hi[35:32]};
  wire [7:0]         regroupV0_hi_lo_hi_9 = {regroupV0_hi[419:416], regroupV0_hi[291:288]};
  wire [15:0]        regroupV0_hi_lo_9 = {regroupV0_hi_lo_hi_9, regroupV0_hi_lo_lo_9};
  wire [7:0]         regroupV0_hi_hi_lo_9 = {regroupV0_hi[675:672], regroupV0_hi[547:544]};
  wire [7:0]         regroupV0_hi_hi_hi_9 = {regroupV0_hi[931:928], regroupV0_hi[803:800]};
  wire [15:0]        regroupV0_hi_hi_9 = {regroupV0_hi_hi_hi_9, regroupV0_hi_hi_lo_9};
  wire [31:0]        regroupV0_hi_9 = {regroupV0_hi_hi_9, regroupV0_hi_lo_9};
  wire [7:0]         regroupV0_lo_lo_lo_10 = {regroupV0_lo[167:164], regroupV0_lo[39:36]};
  wire [7:0]         regroupV0_lo_lo_hi_10 = {regroupV0_lo[423:420], regroupV0_lo[295:292]};
  wire [15:0]        regroupV0_lo_lo_10 = {regroupV0_lo_lo_hi_10, regroupV0_lo_lo_lo_10};
  wire [7:0]         regroupV0_lo_hi_lo_10 = {regroupV0_lo[679:676], regroupV0_lo[551:548]};
  wire [7:0]         regroupV0_lo_hi_hi_10 = {regroupV0_lo[935:932], regroupV0_lo[807:804]};
  wire [15:0]        regroupV0_lo_hi_10 = {regroupV0_lo_hi_hi_10, regroupV0_lo_hi_lo_10};
  wire [31:0]        regroupV0_lo_10 = {regroupV0_lo_hi_10, regroupV0_lo_lo_10};
  wire [7:0]         regroupV0_hi_lo_lo_10 = {regroupV0_hi[167:164], regroupV0_hi[39:36]};
  wire [7:0]         regroupV0_hi_lo_hi_10 = {regroupV0_hi[423:420], regroupV0_hi[295:292]};
  wire [15:0]        regroupV0_hi_lo_10 = {regroupV0_hi_lo_hi_10, regroupV0_hi_lo_lo_10};
  wire [7:0]         regroupV0_hi_hi_lo_10 = {regroupV0_hi[679:676], regroupV0_hi[551:548]};
  wire [7:0]         regroupV0_hi_hi_hi_10 = {regroupV0_hi[935:932], regroupV0_hi[807:804]};
  wire [15:0]        regroupV0_hi_hi_10 = {regroupV0_hi_hi_hi_10, regroupV0_hi_hi_lo_10};
  wire [31:0]        regroupV0_hi_10 = {regroupV0_hi_hi_10, regroupV0_hi_lo_10};
  wire [7:0]         regroupV0_lo_lo_lo_11 = {regroupV0_lo[171:168], regroupV0_lo[43:40]};
  wire [7:0]         regroupV0_lo_lo_hi_11 = {regroupV0_lo[427:424], regroupV0_lo[299:296]};
  wire [15:0]        regroupV0_lo_lo_11 = {regroupV0_lo_lo_hi_11, regroupV0_lo_lo_lo_11};
  wire [7:0]         regroupV0_lo_hi_lo_11 = {regroupV0_lo[683:680], regroupV0_lo[555:552]};
  wire [7:0]         regroupV0_lo_hi_hi_11 = {regroupV0_lo[939:936], regroupV0_lo[811:808]};
  wire [15:0]        regroupV0_lo_hi_11 = {regroupV0_lo_hi_hi_11, regroupV0_lo_hi_lo_11};
  wire [31:0]        regroupV0_lo_11 = {regroupV0_lo_hi_11, regroupV0_lo_lo_11};
  wire [7:0]         regroupV0_hi_lo_lo_11 = {regroupV0_hi[171:168], regroupV0_hi[43:40]};
  wire [7:0]         regroupV0_hi_lo_hi_11 = {regroupV0_hi[427:424], regroupV0_hi[299:296]};
  wire [15:0]        regroupV0_hi_lo_11 = {regroupV0_hi_lo_hi_11, regroupV0_hi_lo_lo_11};
  wire [7:0]         regroupV0_hi_hi_lo_11 = {regroupV0_hi[683:680], regroupV0_hi[555:552]};
  wire [7:0]         regroupV0_hi_hi_hi_11 = {regroupV0_hi[939:936], regroupV0_hi[811:808]};
  wire [15:0]        regroupV0_hi_hi_11 = {regroupV0_hi_hi_hi_11, regroupV0_hi_hi_lo_11};
  wire [31:0]        regroupV0_hi_11 = {regroupV0_hi_hi_11, regroupV0_hi_lo_11};
  wire [7:0]         regroupV0_lo_lo_lo_12 = {regroupV0_lo[175:172], regroupV0_lo[47:44]};
  wire [7:0]         regroupV0_lo_lo_hi_12 = {regroupV0_lo[431:428], regroupV0_lo[303:300]};
  wire [15:0]        regroupV0_lo_lo_12 = {regroupV0_lo_lo_hi_12, regroupV0_lo_lo_lo_12};
  wire [7:0]         regroupV0_lo_hi_lo_12 = {regroupV0_lo[687:684], regroupV0_lo[559:556]};
  wire [7:0]         regroupV0_lo_hi_hi_12 = {regroupV0_lo[943:940], regroupV0_lo[815:812]};
  wire [15:0]        regroupV0_lo_hi_12 = {regroupV0_lo_hi_hi_12, regroupV0_lo_hi_lo_12};
  wire [31:0]        regroupV0_lo_12 = {regroupV0_lo_hi_12, regroupV0_lo_lo_12};
  wire [7:0]         regroupV0_hi_lo_lo_12 = {regroupV0_hi[175:172], regroupV0_hi[47:44]};
  wire [7:0]         regroupV0_hi_lo_hi_12 = {regroupV0_hi[431:428], regroupV0_hi[303:300]};
  wire [15:0]        regroupV0_hi_lo_12 = {regroupV0_hi_lo_hi_12, regroupV0_hi_lo_lo_12};
  wire [7:0]         regroupV0_hi_hi_lo_12 = {regroupV0_hi[687:684], regroupV0_hi[559:556]};
  wire [7:0]         regroupV0_hi_hi_hi_12 = {regroupV0_hi[943:940], regroupV0_hi[815:812]};
  wire [15:0]        regroupV0_hi_hi_12 = {regroupV0_hi_hi_hi_12, regroupV0_hi_hi_lo_12};
  wire [31:0]        regroupV0_hi_12 = {regroupV0_hi_hi_12, regroupV0_hi_lo_12};
  wire [7:0]         regroupV0_lo_lo_lo_13 = {regroupV0_lo[179:176], regroupV0_lo[51:48]};
  wire [7:0]         regroupV0_lo_lo_hi_13 = {regroupV0_lo[435:432], regroupV0_lo[307:304]};
  wire [15:0]        regroupV0_lo_lo_13 = {regroupV0_lo_lo_hi_13, regroupV0_lo_lo_lo_13};
  wire [7:0]         regroupV0_lo_hi_lo_13 = {regroupV0_lo[691:688], regroupV0_lo[563:560]};
  wire [7:0]         regroupV0_lo_hi_hi_13 = {regroupV0_lo[947:944], regroupV0_lo[819:816]};
  wire [15:0]        regroupV0_lo_hi_13 = {regroupV0_lo_hi_hi_13, regroupV0_lo_hi_lo_13};
  wire [31:0]        regroupV0_lo_13 = {regroupV0_lo_hi_13, regroupV0_lo_lo_13};
  wire [7:0]         regroupV0_hi_lo_lo_13 = {regroupV0_hi[179:176], regroupV0_hi[51:48]};
  wire [7:0]         regroupV0_hi_lo_hi_13 = {regroupV0_hi[435:432], regroupV0_hi[307:304]};
  wire [15:0]        regroupV0_hi_lo_13 = {regroupV0_hi_lo_hi_13, regroupV0_hi_lo_lo_13};
  wire [7:0]         regroupV0_hi_hi_lo_13 = {regroupV0_hi[691:688], regroupV0_hi[563:560]};
  wire [7:0]         regroupV0_hi_hi_hi_13 = {regroupV0_hi[947:944], regroupV0_hi[819:816]};
  wire [15:0]        regroupV0_hi_hi_13 = {regroupV0_hi_hi_hi_13, regroupV0_hi_hi_lo_13};
  wire [31:0]        regroupV0_hi_13 = {regroupV0_hi_hi_13, regroupV0_hi_lo_13};
  wire [7:0]         regroupV0_lo_lo_lo_14 = {regroupV0_lo[183:180], regroupV0_lo[55:52]};
  wire [7:0]         regroupV0_lo_lo_hi_14 = {regroupV0_lo[439:436], regroupV0_lo[311:308]};
  wire [15:0]        regroupV0_lo_lo_14 = {regroupV0_lo_lo_hi_14, regroupV0_lo_lo_lo_14};
  wire [7:0]         regroupV0_lo_hi_lo_14 = {regroupV0_lo[695:692], regroupV0_lo[567:564]};
  wire [7:0]         regroupV0_lo_hi_hi_14 = {regroupV0_lo[951:948], regroupV0_lo[823:820]};
  wire [15:0]        regroupV0_lo_hi_14 = {regroupV0_lo_hi_hi_14, regroupV0_lo_hi_lo_14};
  wire [31:0]        regroupV0_lo_14 = {regroupV0_lo_hi_14, regroupV0_lo_lo_14};
  wire [7:0]         regroupV0_hi_lo_lo_14 = {regroupV0_hi[183:180], regroupV0_hi[55:52]};
  wire [7:0]         regroupV0_hi_lo_hi_14 = {regroupV0_hi[439:436], regroupV0_hi[311:308]};
  wire [15:0]        regroupV0_hi_lo_14 = {regroupV0_hi_lo_hi_14, regroupV0_hi_lo_lo_14};
  wire [7:0]         regroupV0_hi_hi_lo_14 = {regroupV0_hi[695:692], regroupV0_hi[567:564]};
  wire [7:0]         regroupV0_hi_hi_hi_14 = {regroupV0_hi[951:948], regroupV0_hi[823:820]};
  wire [15:0]        regroupV0_hi_hi_14 = {regroupV0_hi_hi_hi_14, regroupV0_hi_hi_lo_14};
  wire [31:0]        regroupV0_hi_14 = {regroupV0_hi_hi_14, regroupV0_hi_lo_14};
  wire [7:0]         regroupV0_lo_lo_lo_15 = {regroupV0_lo[187:184], regroupV0_lo[59:56]};
  wire [7:0]         regroupV0_lo_lo_hi_15 = {regroupV0_lo[443:440], regroupV0_lo[315:312]};
  wire [15:0]        regroupV0_lo_lo_15 = {regroupV0_lo_lo_hi_15, regroupV0_lo_lo_lo_15};
  wire [7:0]         regroupV0_lo_hi_lo_15 = {regroupV0_lo[699:696], regroupV0_lo[571:568]};
  wire [7:0]         regroupV0_lo_hi_hi_15 = {regroupV0_lo[955:952], regroupV0_lo[827:824]};
  wire [15:0]        regroupV0_lo_hi_15 = {regroupV0_lo_hi_hi_15, regroupV0_lo_hi_lo_15};
  wire [31:0]        regroupV0_lo_15 = {regroupV0_lo_hi_15, regroupV0_lo_lo_15};
  wire [7:0]         regroupV0_hi_lo_lo_15 = {regroupV0_hi[187:184], regroupV0_hi[59:56]};
  wire [7:0]         regroupV0_hi_lo_hi_15 = {regroupV0_hi[443:440], regroupV0_hi[315:312]};
  wire [15:0]        regroupV0_hi_lo_15 = {regroupV0_hi_lo_hi_15, regroupV0_hi_lo_lo_15};
  wire [7:0]         regroupV0_hi_hi_lo_15 = {regroupV0_hi[699:696], regroupV0_hi[571:568]};
  wire [7:0]         regroupV0_hi_hi_hi_15 = {regroupV0_hi[955:952], regroupV0_hi[827:824]};
  wire [15:0]        regroupV0_hi_hi_15 = {regroupV0_hi_hi_hi_15, regroupV0_hi_hi_lo_15};
  wire [31:0]        regroupV0_hi_15 = {regroupV0_hi_hi_15, regroupV0_hi_lo_15};
  wire [7:0]         regroupV0_lo_lo_lo_16 = {regroupV0_lo[191:188], regroupV0_lo[63:60]};
  wire [7:0]         regroupV0_lo_lo_hi_16 = {regroupV0_lo[447:444], regroupV0_lo[319:316]};
  wire [15:0]        regroupV0_lo_lo_16 = {regroupV0_lo_lo_hi_16, regroupV0_lo_lo_lo_16};
  wire [7:0]         regroupV0_lo_hi_lo_16 = {regroupV0_lo[703:700], regroupV0_lo[575:572]};
  wire [7:0]         regroupV0_lo_hi_hi_16 = {regroupV0_lo[959:956], regroupV0_lo[831:828]};
  wire [15:0]        regroupV0_lo_hi_16 = {regroupV0_lo_hi_hi_16, regroupV0_lo_hi_lo_16};
  wire [31:0]        regroupV0_lo_16 = {regroupV0_lo_hi_16, regroupV0_lo_lo_16};
  wire [7:0]         regroupV0_hi_lo_lo_16 = {regroupV0_hi[191:188], regroupV0_hi[63:60]};
  wire [7:0]         regroupV0_hi_lo_hi_16 = {regroupV0_hi[447:444], regroupV0_hi[319:316]};
  wire [15:0]        regroupV0_hi_lo_16 = {regroupV0_hi_lo_hi_16, regroupV0_hi_lo_lo_16};
  wire [7:0]         regroupV0_hi_hi_lo_16 = {regroupV0_hi[703:700], regroupV0_hi[575:572]};
  wire [7:0]         regroupV0_hi_hi_hi_16 = {regroupV0_hi[959:956], regroupV0_hi[831:828]};
  wire [15:0]        regroupV0_hi_hi_16 = {regroupV0_hi_hi_hi_16, regroupV0_hi_hi_lo_16};
  wire [31:0]        regroupV0_hi_16 = {regroupV0_hi_hi_16, regroupV0_hi_lo_16};
  wire [7:0]         regroupV0_lo_lo_lo_17 = {regroupV0_lo[195:192], regroupV0_lo[67:64]};
  wire [7:0]         regroupV0_lo_lo_hi_17 = {regroupV0_lo[451:448], regroupV0_lo[323:320]};
  wire [15:0]        regroupV0_lo_lo_17 = {regroupV0_lo_lo_hi_17, regroupV0_lo_lo_lo_17};
  wire [7:0]         regroupV0_lo_hi_lo_17 = {regroupV0_lo[707:704], regroupV0_lo[579:576]};
  wire [7:0]         regroupV0_lo_hi_hi_17 = {regroupV0_lo[963:960], regroupV0_lo[835:832]};
  wire [15:0]        regroupV0_lo_hi_17 = {regroupV0_lo_hi_hi_17, regroupV0_lo_hi_lo_17};
  wire [31:0]        regroupV0_lo_17 = {regroupV0_lo_hi_17, regroupV0_lo_lo_17};
  wire [7:0]         regroupV0_hi_lo_lo_17 = {regroupV0_hi[195:192], regroupV0_hi[67:64]};
  wire [7:0]         regroupV0_hi_lo_hi_17 = {regroupV0_hi[451:448], regroupV0_hi[323:320]};
  wire [15:0]        regroupV0_hi_lo_17 = {regroupV0_hi_lo_hi_17, regroupV0_hi_lo_lo_17};
  wire [7:0]         regroupV0_hi_hi_lo_17 = {regroupV0_hi[707:704], regroupV0_hi[579:576]};
  wire [7:0]         regroupV0_hi_hi_hi_17 = {regroupV0_hi[963:960], regroupV0_hi[835:832]};
  wire [15:0]        regroupV0_hi_hi_17 = {regroupV0_hi_hi_hi_17, regroupV0_hi_hi_lo_17};
  wire [31:0]        regroupV0_hi_17 = {regroupV0_hi_hi_17, regroupV0_hi_lo_17};
  wire [7:0]         regroupV0_lo_lo_lo_18 = {regroupV0_lo[199:196], regroupV0_lo[71:68]};
  wire [7:0]         regroupV0_lo_lo_hi_18 = {regroupV0_lo[455:452], regroupV0_lo[327:324]};
  wire [15:0]        regroupV0_lo_lo_18 = {regroupV0_lo_lo_hi_18, regroupV0_lo_lo_lo_18};
  wire [7:0]         regroupV0_lo_hi_lo_18 = {regroupV0_lo[711:708], regroupV0_lo[583:580]};
  wire [7:0]         regroupV0_lo_hi_hi_18 = {regroupV0_lo[967:964], regroupV0_lo[839:836]};
  wire [15:0]        regroupV0_lo_hi_18 = {regroupV0_lo_hi_hi_18, regroupV0_lo_hi_lo_18};
  wire [31:0]        regroupV0_lo_18 = {regroupV0_lo_hi_18, regroupV0_lo_lo_18};
  wire [7:0]         regroupV0_hi_lo_lo_18 = {regroupV0_hi[199:196], regroupV0_hi[71:68]};
  wire [7:0]         regroupV0_hi_lo_hi_18 = {regroupV0_hi[455:452], regroupV0_hi[327:324]};
  wire [15:0]        regroupV0_hi_lo_18 = {regroupV0_hi_lo_hi_18, regroupV0_hi_lo_lo_18};
  wire [7:0]         regroupV0_hi_hi_lo_18 = {regroupV0_hi[711:708], regroupV0_hi[583:580]};
  wire [7:0]         regroupV0_hi_hi_hi_18 = {regroupV0_hi[967:964], regroupV0_hi[839:836]};
  wire [15:0]        regroupV0_hi_hi_18 = {regroupV0_hi_hi_hi_18, regroupV0_hi_hi_lo_18};
  wire [31:0]        regroupV0_hi_18 = {regroupV0_hi_hi_18, regroupV0_hi_lo_18};
  wire [7:0]         regroupV0_lo_lo_lo_19 = {regroupV0_lo[203:200], regroupV0_lo[75:72]};
  wire [7:0]         regroupV0_lo_lo_hi_19 = {regroupV0_lo[459:456], regroupV0_lo[331:328]};
  wire [15:0]        regroupV0_lo_lo_19 = {regroupV0_lo_lo_hi_19, regroupV0_lo_lo_lo_19};
  wire [7:0]         regroupV0_lo_hi_lo_19 = {regroupV0_lo[715:712], regroupV0_lo[587:584]};
  wire [7:0]         regroupV0_lo_hi_hi_19 = {regroupV0_lo[971:968], regroupV0_lo[843:840]};
  wire [15:0]        regroupV0_lo_hi_19 = {regroupV0_lo_hi_hi_19, regroupV0_lo_hi_lo_19};
  wire [31:0]        regroupV0_lo_19 = {regroupV0_lo_hi_19, regroupV0_lo_lo_19};
  wire [7:0]         regroupV0_hi_lo_lo_19 = {regroupV0_hi[203:200], regroupV0_hi[75:72]};
  wire [7:0]         regroupV0_hi_lo_hi_19 = {regroupV0_hi[459:456], regroupV0_hi[331:328]};
  wire [15:0]        regroupV0_hi_lo_19 = {regroupV0_hi_lo_hi_19, regroupV0_hi_lo_lo_19};
  wire [7:0]         regroupV0_hi_hi_lo_19 = {regroupV0_hi[715:712], regroupV0_hi[587:584]};
  wire [7:0]         regroupV0_hi_hi_hi_19 = {regroupV0_hi[971:968], regroupV0_hi[843:840]};
  wire [15:0]        regroupV0_hi_hi_19 = {regroupV0_hi_hi_hi_19, regroupV0_hi_hi_lo_19};
  wire [31:0]        regroupV0_hi_19 = {regroupV0_hi_hi_19, regroupV0_hi_lo_19};
  wire [7:0]         regroupV0_lo_lo_lo_20 = {regroupV0_lo[207:204], regroupV0_lo[79:76]};
  wire [7:0]         regroupV0_lo_lo_hi_20 = {regroupV0_lo[463:460], regroupV0_lo[335:332]};
  wire [15:0]        regroupV0_lo_lo_20 = {regroupV0_lo_lo_hi_20, regroupV0_lo_lo_lo_20};
  wire [7:0]         regroupV0_lo_hi_lo_20 = {regroupV0_lo[719:716], regroupV0_lo[591:588]};
  wire [7:0]         regroupV0_lo_hi_hi_20 = {regroupV0_lo[975:972], regroupV0_lo[847:844]};
  wire [15:0]        regroupV0_lo_hi_20 = {regroupV0_lo_hi_hi_20, regroupV0_lo_hi_lo_20};
  wire [31:0]        regroupV0_lo_20 = {regroupV0_lo_hi_20, regroupV0_lo_lo_20};
  wire [7:0]         regroupV0_hi_lo_lo_20 = {regroupV0_hi[207:204], regroupV0_hi[79:76]};
  wire [7:0]         regroupV0_hi_lo_hi_20 = {regroupV0_hi[463:460], regroupV0_hi[335:332]};
  wire [15:0]        regroupV0_hi_lo_20 = {regroupV0_hi_lo_hi_20, regroupV0_hi_lo_lo_20};
  wire [7:0]         regroupV0_hi_hi_lo_20 = {regroupV0_hi[719:716], regroupV0_hi[591:588]};
  wire [7:0]         regroupV0_hi_hi_hi_20 = {regroupV0_hi[975:972], regroupV0_hi[847:844]};
  wire [15:0]        regroupV0_hi_hi_20 = {regroupV0_hi_hi_hi_20, regroupV0_hi_hi_lo_20};
  wire [31:0]        regroupV0_hi_20 = {regroupV0_hi_hi_20, regroupV0_hi_lo_20};
  wire [7:0]         regroupV0_lo_lo_lo_21 = {regroupV0_lo[211:208], regroupV0_lo[83:80]};
  wire [7:0]         regroupV0_lo_lo_hi_21 = {regroupV0_lo[467:464], regroupV0_lo[339:336]};
  wire [15:0]        regroupV0_lo_lo_21 = {regroupV0_lo_lo_hi_21, regroupV0_lo_lo_lo_21};
  wire [7:0]         regroupV0_lo_hi_lo_21 = {regroupV0_lo[723:720], regroupV0_lo[595:592]};
  wire [7:0]         regroupV0_lo_hi_hi_21 = {regroupV0_lo[979:976], regroupV0_lo[851:848]};
  wire [15:0]        regroupV0_lo_hi_21 = {regroupV0_lo_hi_hi_21, regroupV0_lo_hi_lo_21};
  wire [31:0]        regroupV0_lo_21 = {regroupV0_lo_hi_21, regroupV0_lo_lo_21};
  wire [7:0]         regroupV0_hi_lo_lo_21 = {regroupV0_hi[211:208], regroupV0_hi[83:80]};
  wire [7:0]         regroupV0_hi_lo_hi_21 = {regroupV0_hi[467:464], regroupV0_hi[339:336]};
  wire [15:0]        regroupV0_hi_lo_21 = {regroupV0_hi_lo_hi_21, regroupV0_hi_lo_lo_21};
  wire [7:0]         regroupV0_hi_hi_lo_21 = {regroupV0_hi[723:720], regroupV0_hi[595:592]};
  wire [7:0]         regroupV0_hi_hi_hi_21 = {regroupV0_hi[979:976], regroupV0_hi[851:848]};
  wire [15:0]        regroupV0_hi_hi_21 = {regroupV0_hi_hi_hi_21, regroupV0_hi_hi_lo_21};
  wire [31:0]        regroupV0_hi_21 = {regroupV0_hi_hi_21, regroupV0_hi_lo_21};
  wire [7:0]         regroupV0_lo_lo_lo_22 = {regroupV0_lo[215:212], regroupV0_lo[87:84]};
  wire [7:0]         regroupV0_lo_lo_hi_22 = {regroupV0_lo[471:468], regroupV0_lo[343:340]};
  wire [15:0]        regroupV0_lo_lo_22 = {regroupV0_lo_lo_hi_22, regroupV0_lo_lo_lo_22};
  wire [7:0]         regroupV0_lo_hi_lo_22 = {regroupV0_lo[727:724], regroupV0_lo[599:596]};
  wire [7:0]         regroupV0_lo_hi_hi_22 = {regroupV0_lo[983:980], regroupV0_lo[855:852]};
  wire [15:0]        regroupV0_lo_hi_22 = {regroupV0_lo_hi_hi_22, regroupV0_lo_hi_lo_22};
  wire [31:0]        regroupV0_lo_22 = {regroupV0_lo_hi_22, regroupV0_lo_lo_22};
  wire [7:0]         regroupV0_hi_lo_lo_22 = {regroupV0_hi[215:212], regroupV0_hi[87:84]};
  wire [7:0]         regroupV0_hi_lo_hi_22 = {regroupV0_hi[471:468], regroupV0_hi[343:340]};
  wire [15:0]        regroupV0_hi_lo_22 = {regroupV0_hi_lo_hi_22, regroupV0_hi_lo_lo_22};
  wire [7:0]         regroupV0_hi_hi_lo_22 = {regroupV0_hi[727:724], regroupV0_hi[599:596]};
  wire [7:0]         regroupV0_hi_hi_hi_22 = {regroupV0_hi[983:980], regroupV0_hi[855:852]};
  wire [15:0]        regroupV0_hi_hi_22 = {regroupV0_hi_hi_hi_22, regroupV0_hi_hi_lo_22};
  wire [31:0]        regroupV0_hi_22 = {regroupV0_hi_hi_22, regroupV0_hi_lo_22};
  wire [7:0]         regroupV0_lo_lo_lo_23 = {regroupV0_lo[219:216], regroupV0_lo[91:88]};
  wire [7:0]         regroupV0_lo_lo_hi_23 = {regroupV0_lo[475:472], regroupV0_lo[347:344]};
  wire [15:0]        regroupV0_lo_lo_23 = {regroupV0_lo_lo_hi_23, regroupV0_lo_lo_lo_23};
  wire [7:0]         regroupV0_lo_hi_lo_23 = {regroupV0_lo[731:728], regroupV0_lo[603:600]};
  wire [7:0]         regroupV0_lo_hi_hi_23 = {regroupV0_lo[987:984], regroupV0_lo[859:856]};
  wire [15:0]        regroupV0_lo_hi_23 = {regroupV0_lo_hi_hi_23, regroupV0_lo_hi_lo_23};
  wire [31:0]        regroupV0_lo_23 = {regroupV0_lo_hi_23, regroupV0_lo_lo_23};
  wire [7:0]         regroupV0_hi_lo_lo_23 = {regroupV0_hi[219:216], regroupV0_hi[91:88]};
  wire [7:0]         regroupV0_hi_lo_hi_23 = {regroupV0_hi[475:472], regroupV0_hi[347:344]};
  wire [15:0]        regroupV0_hi_lo_23 = {regroupV0_hi_lo_hi_23, regroupV0_hi_lo_lo_23};
  wire [7:0]         regroupV0_hi_hi_lo_23 = {regroupV0_hi[731:728], regroupV0_hi[603:600]};
  wire [7:0]         regroupV0_hi_hi_hi_23 = {regroupV0_hi[987:984], regroupV0_hi[859:856]};
  wire [15:0]        regroupV0_hi_hi_23 = {regroupV0_hi_hi_hi_23, regroupV0_hi_hi_lo_23};
  wire [31:0]        regroupV0_hi_23 = {regroupV0_hi_hi_23, regroupV0_hi_lo_23};
  wire [7:0]         regroupV0_lo_lo_lo_24 = {regroupV0_lo[223:220], regroupV0_lo[95:92]};
  wire [7:0]         regroupV0_lo_lo_hi_24 = {regroupV0_lo[479:476], regroupV0_lo[351:348]};
  wire [15:0]        regroupV0_lo_lo_24 = {regroupV0_lo_lo_hi_24, regroupV0_lo_lo_lo_24};
  wire [7:0]         regroupV0_lo_hi_lo_24 = {regroupV0_lo[735:732], regroupV0_lo[607:604]};
  wire [7:0]         regroupV0_lo_hi_hi_24 = {regroupV0_lo[991:988], regroupV0_lo[863:860]};
  wire [15:0]        regroupV0_lo_hi_24 = {regroupV0_lo_hi_hi_24, regroupV0_lo_hi_lo_24};
  wire [31:0]        regroupV0_lo_24 = {regroupV0_lo_hi_24, regroupV0_lo_lo_24};
  wire [7:0]         regroupV0_hi_lo_lo_24 = {regroupV0_hi[223:220], regroupV0_hi[95:92]};
  wire [7:0]         regroupV0_hi_lo_hi_24 = {regroupV0_hi[479:476], regroupV0_hi[351:348]};
  wire [15:0]        regroupV0_hi_lo_24 = {regroupV0_hi_lo_hi_24, regroupV0_hi_lo_lo_24};
  wire [7:0]         regroupV0_hi_hi_lo_24 = {regroupV0_hi[735:732], regroupV0_hi[607:604]};
  wire [7:0]         regroupV0_hi_hi_hi_24 = {regroupV0_hi[991:988], regroupV0_hi[863:860]};
  wire [15:0]        regroupV0_hi_hi_24 = {regroupV0_hi_hi_hi_24, regroupV0_hi_hi_lo_24};
  wire [31:0]        regroupV0_hi_24 = {regroupV0_hi_hi_24, regroupV0_hi_lo_24};
  wire [7:0]         regroupV0_lo_lo_lo_25 = {regroupV0_lo[227:224], regroupV0_lo[99:96]};
  wire [7:0]         regroupV0_lo_lo_hi_25 = {regroupV0_lo[483:480], regroupV0_lo[355:352]};
  wire [15:0]        regroupV0_lo_lo_25 = {regroupV0_lo_lo_hi_25, regroupV0_lo_lo_lo_25};
  wire [7:0]         regroupV0_lo_hi_lo_25 = {regroupV0_lo[739:736], regroupV0_lo[611:608]};
  wire [7:0]         regroupV0_lo_hi_hi_25 = {regroupV0_lo[995:992], regroupV0_lo[867:864]};
  wire [15:0]        regroupV0_lo_hi_25 = {regroupV0_lo_hi_hi_25, regroupV0_lo_hi_lo_25};
  wire [31:0]        regroupV0_lo_25 = {regroupV0_lo_hi_25, regroupV0_lo_lo_25};
  wire [7:0]         regroupV0_hi_lo_lo_25 = {regroupV0_hi[227:224], regroupV0_hi[99:96]};
  wire [7:0]         regroupV0_hi_lo_hi_25 = {regroupV0_hi[483:480], regroupV0_hi[355:352]};
  wire [15:0]        regroupV0_hi_lo_25 = {regroupV0_hi_lo_hi_25, regroupV0_hi_lo_lo_25};
  wire [7:0]         regroupV0_hi_hi_lo_25 = {regroupV0_hi[739:736], regroupV0_hi[611:608]};
  wire [7:0]         regroupV0_hi_hi_hi_25 = {regroupV0_hi[995:992], regroupV0_hi[867:864]};
  wire [15:0]        regroupV0_hi_hi_25 = {regroupV0_hi_hi_hi_25, regroupV0_hi_hi_lo_25};
  wire [31:0]        regroupV0_hi_25 = {regroupV0_hi_hi_25, regroupV0_hi_lo_25};
  wire [7:0]         regroupV0_lo_lo_lo_26 = {regroupV0_lo[231:228], regroupV0_lo[103:100]};
  wire [7:0]         regroupV0_lo_lo_hi_26 = {regroupV0_lo[487:484], regroupV0_lo[359:356]};
  wire [15:0]        regroupV0_lo_lo_26 = {regroupV0_lo_lo_hi_26, regroupV0_lo_lo_lo_26};
  wire [7:0]         regroupV0_lo_hi_lo_26 = {regroupV0_lo[743:740], regroupV0_lo[615:612]};
  wire [7:0]         regroupV0_lo_hi_hi_26 = {regroupV0_lo[999:996], regroupV0_lo[871:868]};
  wire [15:0]        regroupV0_lo_hi_26 = {regroupV0_lo_hi_hi_26, regroupV0_lo_hi_lo_26};
  wire [31:0]        regroupV0_lo_26 = {regroupV0_lo_hi_26, regroupV0_lo_lo_26};
  wire [7:0]         regroupV0_hi_lo_lo_26 = {regroupV0_hi[231:228], regroupV0_hi[103:100]};
  wire [7:0]         regroupV0_hi_lo_hi_26 = {regroupV0_hi[487:484], regroupV0_hi[359:356]};
  wire [15:0]        regroupV0_hi_lo_26 = {regroupV0_hi_lo_hi_26, regroupV0_hi_lo_lo_26};
  wire [7:0]         regroupV0_hi_hi_lo_26 = {regroupV0_hi[743:740], regroupV0_hi[615:612]};
  wire [7:0]         regroupV0_hi_hi_hi_26 = {regroupV0_hi[999:996], regroupV0_hi[871:868]};
  wire [15:0]        regroupV0_hi_hi_26 = {regroupV0_hi_hi_hi_26, regroupV0_hi_hi_lo_26};
  wire [31:0]        regroupV0_hi_26 = {regroupV0_hi_hi_26, regroupV0_hi_lo_26};
  wire [7:0]         regroupV0_lo_lo_lo_27 = {regroupV0_lo[235:232], regroupV0_lo[107:104]};
  wire [7:0]         regroupV0_lo_lo_hi_27 = {regroupV0_lo[491:488], regroupV0_lo[363:360]};
  wire [15:0]        regroupV0_lo_lo_27 = {regroupV0_lo_lo_hi_27, regroupV0_lo_lo_lo_27};
  wire [7:0]         regroupV0_lo_hi_lo_27 = {regroupV0_lo[747:744], regroupV0_lo[619:616]};
  wire [7:0]         regroupV0_lo_hi_hi_27 = {regroupV0_lo[1003:1000], regroupV0_lo[875:872]};
  wire [15:0]        regroupV0_lo_hi_27 = {regroupV0_lo_hi_hi_27, regroupV0_lo_hi_lo_27};
  wire [31:0]        regroupV0_lo_27 = {regroupV0_lo_hi_27, regroupV0_lo_lo_27};
  wire [7:0]         regroupV0_hi_lo_lo_27 = {regroupV0_hi[235:232], regroupV0_hi[107:104]};
  wire [7:0]         regroupV0_hi_lo_hi_27 = {regroupV0_hi[491:488], regroupV0_hi[363:360]};
  wire [15:0]        regroupV0_hi_lo_27 = {regroupV0_hi_lo_hi_27, regroupV0_hi_lo_lo_27};
  wire [7:0]         regroupV0_hi_hi_lo_27 = {regroupV0_hi[747:744], regroupV0_hi[619:616]};
  wire [7:0]         regroupV0_hi_hi_hi_27 = {regroupV0_hi[1003:1000], regroupV0_hi[875:872]};
  wire [15:0]        regroupV0_hi_hi_27 = {regroupV0_hi_hi_hi_27, regroupV0_hi_hi_lo_27};
  wire [31:0]        regroupV0_hi_27 = {regroupV0_hi_hi_27, regroupV0_hi_lo_27};
  wire [7:0]         regroupV0_lo_lo_lo_28 = {regroupV0_lo[239:236], regroupV0_lo[111:108]};
  wire [7:0]         regroupV0_lo_lo_hi_28 = {regroupV0_lo[495:492], regroupV0_lo[367:364]};
  wire [15:0]        regroupV0_lo_lo_28 = {regroupV0_lo_lo_hi_28, regroupV0_lo_lo_lo_28};
  wire [7:0]         regroupV0_lo_hi_lo_28 = {regroupV0_lo[751:748], regroupV0_lo[623:620]};
  wire [7:0]         regroupV0_lo_hi_hi_28 = {regroupV0_lo[1007:1004], regroupV0_lo[879:876]};
  wire [15:0]        regroupV0_lo_hi_28 = {regroupV0_lo_hi_hi_28, regroupV0_lo_hi_lo_28};
  wire [31:0]        regroupV0_lo_28 = {regroupV0_lo_hi_28, regroupV0_lo_lo_28};
  wire [7:0]         regroupV0_hi_lo_lo_28 = {regroupV0_hi[239:236], regroupV0_hi[111:108]};
  wire [7:0]         regroupV0_hi_lo_hi_28 = {regroupV0_hi[495:492], regroupV0_hi[367:364]};
  wire [15:0]        regroupV0_hi_lo_28 = {regroupV0_hi_lo_hi_28, regroupV0_hi_lo_lo_28};
  wire [7:0]         regroupV0_hi_hi_lo_28 = {regroupV0_hi[751:748], regroupV0_hi[623:620]};
  wire [7:0]         regroupV0_hi_hi_hi_28 = {regroupV0_hi[1007:1004], regroupV0_hi[879:876]};
  wire [15:0]        regroupV0_hi_hi_28 = {regroupV0_hi_hi_hi_28, regroupV0_hi_hi_lo_28};
  wire [31:0]        regroupV0_hi_28 = {regroupV0_hi_hi_28, regroupV0_hi_lo_28};
  wire [7:0]         regroupV0_lo_lo_lo_29 = {regroupV0_lo[243:240], regroupV0_lo[115:112]};
  wire [7:0]         regroupV0_lo_lo_hi_29 = {regroupV0_lo[499:496], regroupV0_lo[371:368]};
  wire [15:0]        regroupV0_lo_lo_29 = {regroupV0_lo_lo_hi_29, regroupV0_lo_lo_lo_29};
  wire [7:0]         regroupV0_lo_hi_lo_29 = {regroupV0_lo[755:752], regroupV0_lo[627:624]};
  wire [7:0]         regroupV0_lo_hi_hi_29 = {regroupV0_lo[1011:1008], regroupV0_lo[883:880]};
  wire [15:0]        regroupV0_lo_hi_29 = {regroupV0_lo_hi_hi_29, regroupV0_lo_hi_lo_29};
  wire [31:0]        regroupV0_lo_29 = {regroupV0_lo_hi_29, regroupV0_lo_lo_29};
  wire [7:0]         regroupV0_hi_lo_lo_29 = {regroupV0_hi[243:240], regroupV0_hi[115:112]};
  wire [7:0]         regroupV0_hi_lo_hi_29 = {regroupV0_hi[499:496], regroupV0_hi[371:368]};
  wire [15:0]        regroupV0_hi_lo_29 = {regroupV0_hi_lo_hi_29, regroupV0_hi_lo_lo_29};
  wire [7:0]         regroupV0_hi_hi_lo_29 = {regroupV0_hi[755:752], regroupV0_hi[627:624]};
  wire [7:0]         regroupV0_hi_hi_hi_29 = {regroupV0_hi[1011:1008], regroupV0_hi[883:880]};
  wire [15:0]        regroupV0_hi_hi_29 = {regroupV0_hi_hi_hi_29, regroupV0_hi_hi_lo_29};
  wire [31:0]        regroupV0_hi_29 = {regroupV0_hi_hi_29, regroupV0_hi_lo_29};
  wire [7:0]         regroupV0_lo_lo_lo_30 = {regroupV0_lo[247:244], regroupV0_lo[119:116]};
  wire [7:0]         regroupV0_lo_lo_hi_30 = {regroupV0_lo[503:500], regroupV0_lo[375:372]};
  wire [15:0]        regroupV0_lo_lo_30 = {regroupV0_lo_lo_hi_30, regroupV0_lo_lo_lo_30};
  wire [7:0]         regroupV0_lo_hi_lo_30 = {regroupV0_lo[759:756], regroupV0_lo[631:628]};
  wire [7:0]         regroupV0_lo_hi_hi_30 = {regroupV0_lo[1015:1012], regroupV0_lo[887:884]};
  wire [15:0]        regroupV0_lo_hi_30 = {regroupV0_lo_hi_hi_30, regroupV0_lo_hi_lo_30};
  wire [31:0]        regroupV0_lo_30 = {regroupV0_lo_hi_30, regroupV0_lo_lo_30};
  wire [7:0]         regroupV0_hi_lo_lo_30 = {regroupV0_hi[247:244], regroupV0_hi[119:116]};
  wire [7:0]         regroupV0_hi_lo_hi_30 = {regroupV0_hi[503:500], regroupV0_hi[375:372]};
  wire [15:0]        regroupV0_hi_lo_30 = {regroupV0_hi_lo_hi_30, regroupV0_hi_lo_lo_30};
  wire [7:0]         regroupV0_hi_hi_lo_30 = {regroupV0_hi[759:756], regroupV0_hi[631:628]};
  wire [7:0]         regroupV0_hi_hi_hi_30 = {regroupV0_hi[1015:1012], regroupV0_hi[887:884]};
  wire [15:0]        regroupV0_hi_hi_30 = {regroupV0_hi_hi_hi_30, regroupV0_hi_hi_lo_30};
  wire [31:0]        regroupV0_hi_30 = {regroupV0_hi_hi_30, regroupV0_hi_lo_30};
  wire [7:0]         regroupV0_lo_lo_lo_31 = {regroupV0_lo[251:248], regroupV0_lo[123:120]};
  wire [7:0]         regroupV0_lo_lo_hi_31 = {regroupV0_lo[507:504], regroupV0_lo[379:376]};
  wire [15:0]        regroupV0_lo_lo_31 = {regroupV0_lo_lo_hi_31, regroupV0_lo_lo_lo_31};
  wire [7:0]         regroupV0_lo_hi_lo_31 = {regroupV0_lo[763:760], regroupV0_lo[635:632]};
  wire [7:0]         regroupV0_lo_hi_hi_31 = {regroupV0_lo[1019:1016], regroupV0_lo[891:888]};
  wire [15:0]        regroupV0_lo_hi_31 = {regroupV0_lo_hi_hi_31, regroupV0_lo_hi_lo_31};
  wire [31:0]        regroupV0_lo_31 = {regroupV0_lo_hi_31, regroupV0_lo_lo_31};
  wire [7:0]         regroupV0_hi_lo_lo_31 = {regroupV0_hi[251:248], regroupV0_hi[123:120]};
  wire [7:0]         regroupV0_hi_lo_hi_31 = {regroupV0_hi[507:504], regroupV0_hi[379:376]};
  wire [15:0]        regroupV0_hi_lo_31 = {regroupV0_hi_lo_hi_31, regroupV0_hi_lo_lo_31};
  wire [7:0]         regroupV0_hi_hi_lo_31 = {regroupV0_hi[763:760], regroupV0_hi[635:632]};
  wire [7:0]         regroupV0_hi_hi_hi_31 = {regroupV0_hi[1019:1016], regroupV0_hi[891:888]};
  wire [15:0]        regroupV0_hi_hi_31 = {regroupV0_hi_hi_hi_31, regroupV0_hi_hi_lo_31};
  wire [31:0]        regroupV0_hi_31 = {regroupV0_hi_hi_31, regroupV0_hi_lo_31};
  wire [7:0]         regroupV0_lo_lo_lo_32 = {regroupV0_lo[255:252], regroupV0_lo[127:124]};
  wire [7:0]         regroupV0_lo_lo_hi_32 = {regroupV0_lo[511:508], regroupV0_lo[383:380]};
  wire [15:0]        regroupV0_lo_lo_32 = {regroupV0_lo_lo_hi_32, regroupV0_lo_lo_lo_32};
  wire [7:0]         regroupV0_lo_hi_lo_32 = {regroupV0_lo[767:764], regroupV0_lo[639:636]};
  wire [7:0]         regroupV0_lo_hi_hi_32 = {regroupV0_lo[1023:1020], regroupV0_lo[895:892]};
  wire [15:0]        regroupV0_lo_hi_32 = {regroupV0_lo_hi_hi_32, regroupV0_lo_hi_lo_32};
  wire [31:0]        regroupV0_lo_32 = {regroupV0_lo_hi_32, regroupV0_lo_lo_32};
  wire [7:0]         regroupV0_hi_lo_lo_32 = {regroupV0_hi[255:252], regroupV0_hi[127:124]};
  wire [7:0]         regroupV0_hi_lo_hi_32 = {regroupV0_hi[511:508], regroupV0_hi[383:380]};
  wire [15:0]        regroupV0_hi_lo_32 = {regroupV0_hi_lo_hi_32, regroupV0_hi_lo_lo_32};
  wire [7:0]         regroupV0_hi_hi_lo_32 = {regroupV0_hi[767:764], regroupV0_hi[639:636]};
  wire [7:0]         regroupV0_hi_hi_hi_32 = {regroupV0_hi[1023:1020], regroupV0_hi[895:892]};
  wire [15:0]        regroupV0_hi_hi_32 = {regroupV0_hi_hi_hi_32, regroupV0_hi_hi_lo_32};
  wire [31:0]        regroupV0_hi_32 = {regroupV0_hi_hi_32, regroupV0_hi_lo_32};
  wire [127:0]       regroupV0_lo_lo_lo_lo_1 = {regroupV0_hi_2, regroupV0_lo_2, regroupV0_hi_1, regroupV0_lo_1};
  wire [127:0]       regroupV0_lo_lo_lo_hi_1 = {regroupV0_hi_4, regroupV0_lo_4, regroupV0_hi_3, regroupV0_lo_3};
  wire [255:0]       regroupV0_lo_lo_lo_33 = {regroupV0_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_1};
  wire [127:0]       regroupV0_lo_lo_hi_lo_1 = {regroupV0_hi_6, regroupV0_lo_6, regroupV0_hi_5, regroupV0_lo_5};
  wire [127:0]       regroupV0_lo_lo_hi_hi_1 = {regroupV0_hi_8, regroupV0_lo_8, regroupV0_hi_7, regroupV0_lo_7};
  wire [255:0]       regroupV0_lo_lo_hi_33 = {regroupV0_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_1};
  wire [511:0]       regroupV0_lo_lo_33 = {regroupV0_lo_lo_hi_33, regroupV0_lo_lo_lo_33};
  wire [127:0]       regroupV0_lo_hi_lo_lo_1 = {regroupV0_hi_10, regroupV0_lo_10, regroupV0_hi_9, regroupV0_lo_9};
  wire [127:0]       regroupV0_lo_hi_lo_hi_1 = {regroupV0_hi_12, regroupV0_lo_12, regroupV0_hi_11, regroupV0_lo_11};
  wire [255:0]       regroupV0_lo_hi_lo_33 = {regroupV0_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_1};
  wire [127:0]       regroupV0_lo_hi_hi_lo_1 = {regroupV0_hi_14, regroupV0_lo_14, regroupV0_hi_13, regroupV0_lo_13};
  wire [127:0]       regroupV0_lo_hi_hi_hi_1 = {regroupV0_hi_16, regroupV0_lo_16, regroupV0_hi_15, regroupV0_lo_15};
  wire [255:0]       regroupV0_lo_hi_hi_33 = {regroupV0_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_1};
  wire [511:0]       regroupV0_lo_hi_33 = {regroupV0_lo_hi_hi_33, regroupV0_lo_hi_lo_33};
  wire [1023:0]      regroupV0_lo_33 = {regroupV0_lo_hi_33, regroupV0_lo_lo_33};
  wire [127:0]       regroupV0_hi_lo_lo_lo_1 = {regroupV0_hi_18, regroupV0_lo_18, regroupV0_hi_17, regroupV0_lo_17};
  wire [127:0]       regroupV0_hi_lo_lo_hi_1 = {regroupV0_hi_20, regroupV0_lo_20, regroupV0_hi_19, regroupV0_lo_19};
  wire [255:0]       regroupV0_hi_lo_lo_33 = {regroupV0_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_1};
  wire [127:0]       regroupV0_hi_lo_hi_lo_1 = {regroupV0_hi_22, regroupV0_lo_22, regroupV0_hi_21, regroupV0_lo_21};
  wire [127:0]       regroupV0_hi_lo_hi_hi_1 = {regroupV0_hi_24, regroupV0_lo_24, regroupV0_hi_23, regroupV0_lo_23};
  wire [255:0]       regroupV0_hi_lo_hi_33 = {regroupV0_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_1};
  wire [511:0]       regroupV0_hi_lo_33 = {regroupV0_hi_lo_hi_33, regroupV0_hi_lo_lo_33};
  wire [127:0]       regroupV0_hi_hi_lo_lo_1 = {regroupV0_hi_26, regroupV0_lo_26, regroupV0_hi_25, regroupV0_lo_25};
  wire [127:0]       regroupV0_hi_hi_lo_hi_1 = {regroupV0_hi_28, regroupV0_lo_28, regroupV0_hi_27, regroupV0_lo_27};
  wire [255:0]       regroupV0_hi_hi_lo_33 = {regroupV0_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_1};
  wire [127:0]       regroupV0_hi_hi_hi_lo_1 = {regroupV0_hi_30, regroupV0_lo_30, regroupV0_hi_29, regroupV0_lo_29};
  wire [127:0]       regroupV0_hi_hi_hi_hi_1 = {regroupV0_hi_32, regroupV0_lo_32, regroupV0_hi_31, regroupV0_lo_31};
  wire [255:0]       regroupV0_hi_hi_hi_33 = {regroupV0_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_1};
  wire [511:0]       regroupV0_hi_hi_33 = {regroupV0_hi_hi_hi_33, regroupV0_hi_hi_lo_33};
  wire [1023:0]      regroupV0_hi_33 = {regroupV0_hi_hi_33, regroupV0_hi_lo_33};
  wire [2047:0]      regroupV0_0 = {regroupV0_hi_33, regroupV0_lo_33};
  wire [127:0]       regroupV0_lo_lo_lo_lo_2 = {regroupV0_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_1};
  wire [127:0]       regroupV0_lo_lo_lo_hi_2 = {regroupV0_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_1};
  wire [255:0]       regroupV0_lo_lo_lo_34 = {regroupV0_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_2};
  wire [127:0]       regroupV0_lo_lo_hi_lo_2 = {regroupV0_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_1};
  wire [127:0]       regroupV0_lo_lo_hi_hi_2 = {regroupV0_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_1};
  wire [255:0]       regroupV0_lo_lo_hi_34 = {regroupV0_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_2};
  wire [511:0]       regroupV0_lo_lo_34 = {regroupV0_lo_lo_hi_34, regroupV0_lo_lo_lo_34};
  wire [127:0]       regroupV0_lo_hi_lo_lo_2 = {regroupV0_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_1};
  wire [127:0]       regroupV0_lo_hi_lo_hi_2 = {regroupV0_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_1};
  wire [255:0]       regroupV0_lo_hi_lo_34 = {regroupV0_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_2};
  wire [127:0]       regroupV0_lo_hi_hi_lo_2 = {regroupV0_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_1};
  wire [127:0]       regroupV0_lo_hi_hi_hi_2 = {regroupV0_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_1};
  wire [255:0]       regroupV0_lo_hi_hi_34 = {regroupV0_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_2};
  wire [511:0]       regroupV0_lo_hi_34 = {regroupV0_lo_hi_hi_34, regroupV0_lo_hi_lo_34};
  wire [1023:0]      regroupV0_lo_34 = {regroupV0_lo_hi_34, regroupV0_lo_lo_34};
  wire [127:0]       regroupV0_hi_lo_lo_lo_2 = {regroupV0_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_1};
  wire [127:0]       regroupV0_hi_lo_lo_hi_2 = {regroupV0_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_1};
  wire [255:0]       regroupV0_hi_lo_lo_34 = {regroupV0_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_2};
  wire [127:0]       regroupV0_hi_lo_hi_lo_2 = {regroupV0_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_1};
  wire [127:0]       regroupV0_hi_lo_hi_hi_2 = {regroupV0_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_1};
  wire [255:0]       regroupV0_hi_lo_hi_34 = {regroupV0_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_2};
  wire [511:0]       regroupV0_hi_lo_34 = {regroupV0_hi_lo_hi_34, regroupV0_hi_lo_lo_34};
  wire [127:0]       regroupV0_hi_hi_lo_lo_2 = {regroupV0_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_1};
  wire [127:0]       regroupV0_hi_hi_lo_hi_2 = {regroupV0_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_1};
  wire [255:0]       regroupV0_hi_hi_lo_34 = {regroupV0_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_2};
  wire [127:0]       regroupV0_hi_hi_hi_lo_2 = {regroupV0_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_1};
  wire [127:0]       regroupV0_hi_hi_hi_hi_2 = {regroupV0_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_1};
  wire [255:0]       regroupV0_hi_hi_hi_34 = {regroupV0_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_2};
  wire [511:0]       regroupV0_hi_hi_34 = {regroupV0_hi_hi_hi_34, regroupV0_hi_hi_lo_34};
  wire [1023:0]      regroupV0_hi_34 = {regroupV0_hi_hi_34, regroupV0_hi_lo_34};
  wire [3:0]         regroupV0_lo_lo_lo_lo_3 = {regroupV0_lo_34[65:64], regroupV0_lo_34[1:0]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_3 = {regroupV0_lo_34[193:192], regroupV0_lo_34[129:128]};
  wire [7:0]         regroupV0_lo_lo_lo_35 = {regroupV0_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_hi_lo_3 = {regroupV0_lo_34[321:320], regroupV0_lo_34[257:256]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_3 = {regroupV0_lo_34[449:448], regroupV0_lo_34[385:384]};
  wire [7:0]         regroupV0_lo_lo_hi_35 = {regroupV0_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_35 = {regroupV0_lo_lo_hi_35, regroupV0_lo_lo_lo_35};
  wire [3:0]         regroupV0_lo_hi_lo_lo_3 = {regroupV0_lo_34[577:576], regroupV0_lo_34[513:512]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_3 = {regroupV0_lo_34[705:704], regroupV0_lo_34[641:640]};
  wire [7:0]         regroupV0_lo_hi_lo_35 = {regroupV0_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_hi_lo_3 = {regroupV0_lo_34[833:832], regroupV0_lo_34[769:768]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_3 = {regroupV0_lo_34[961:960], regroupV0_lo_34[897:896]};
  wire [7:0]         regroupV0_lo_hi_hi_35 = {regroupV0_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_35 = {regroupV0_lo_hi_hi_35, regroupV0_lo_hi_lo_35};
  wire [31:0]        regroupV0_lo_35 = {regroupV0_lo_hi_35, regroupV0_lo_lo_35};
  wire [3:0]         regroupV0_hi_lo_lo_lo_3 = {regroupV0_hi_34[65:64], regroupV0_hi_34[1:0]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_3 = {regroupV0_hi_34[193:192], regroupV0_hi_34[129:128]};
  wire [7:0]         regroupV0_hi_lo_lo_35 = {regroupV0_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_hi_lo_3 = {regroupV0_hi_34[321:320], regroupV0_hi_34[257:256]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_3 = {regroupV0_hi_34[449:448], regroupV0_hi_34[385:384]};
  wire [7:0]         regroupV0_hi_lo_hi_35 = {regroupV0_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_35 = {regroupV0_hi_lo_hi_35, regroupV0_hi_lo_lo_35};
  wire [3:0]         regroupV0_hi_hi_lo_lo_3 = {regroupV0_hi_34[577:576], regroupV0_hi_34[513:512]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_3 = {regroupV0_hi_34[705:704], regroupV0_hi_34[641:640]};
  wire [7:0]         regroupV0_hi_hi_lo_35 = {regroupV0_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_hi_lo_3 = {regroupV0_hi_34[833:832], regroupV0_hi_34[769:768]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_3 = {regroupV0_hi_34[961:960], regroupV0_hi_34[897:896]};
  wire [7:0]         regroupV0_hi_hi_hi_35 = {regroupV0_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_35 = {regroupV0_hi_hi_hi_35, regroupV0_hi_hi_lo_35};
  wire [31:0]        regroupV0_hi_35 = {regroupV0_hi_hi_35, regroupV0_hi_lo_35};
  wire [3:0]         regroupV0_lo_lo_lo_lo_4 = {regroupV0_lo_34[67:66], regroupV0_lo_34[3:2]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_4 = {regroupV0_lo_34[195:194], regroupV0_lo_34[131:130]};
  wire [7:0]         regroupV0_lo_lo_lo_36 = {regroupV0_lo_lo_lo_hi_4, regroupV0_lo_lo_lo_lo_4};
  wire [3:0]         regroupV0_lo_lo_hi_lo_4 = {regroupV0_lo_34[323:322], regroupV0_lo_34[259:258]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_4 = {regroupV0_lo_34[451:450], regroupV0_lo_34[387:386]};
  wire [7:0]         regroupV0_lo_lo_hi_36 = {regroupV0_lo_lo_hi_hi_4, regroupV0_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_36 = {regroupV0_lo_lo_hi_36, regroupV0_lo_lo_lo_36};
  wire [3:0]         regroupV0_lo_hi_lo_lo_4 = {regroupV0_lo_34[579:578], regroupV0_lo_34[515:514]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_4 = {regroupV0_lo_34[707:706], regroupV0_lo_34[643:642]};
  wire [7:0]         regroupV0_lo_hi_lo_36 = {regroupV0_lo_hi_lo_hi_4, regroupV0_lo_hi_lo_lo_4};
  wire [3:0]         regroupV0_lo_hi_hi_lo_4 = {regroupV0_lo_34[835:834], regroupV0_lo_34[771:770]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_4 = {regroupV0_lo_34[963:962], regroupV0_lo_34[899:898]};
  wire [7:0]         regroupV0_lo_hi_hi_36 = {regroupV0_lo_hi_hi_hi_4, regroupV0_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_36 = {regroupV0_lo_hi_hi_36, regroupV0_lo_hi_lo_36};
  wire [31:0]        regroupV0_lo_36 = {regroupV0_lo_hi_36, regroupV0_lo_lo_36};
  wire [3:0]         regroupV0_hi_lo_lo_lo_4 = {regroupV0_hi_34[67:66], regroupV0_hi_34[3:2]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_4 = {regroupV0_hi_34[195:194], regroupV0_hi_34[131:130]};
  wire [7:0]         regroupV0_hi_lo_lo_36 = {regroupV0_hi_lo_lo_hi_4, regroupV0_hi_lo_lo_lo_4};
  wire [3:0]         regroupV0_hi_lo_hi_lo_4 = {regroupV0_hi_34[323:322], regroupV0_hi_34[259:258]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_4 = {regroupV0_hi_34[451:450], regroupV0_hi_34[387:386]};
  wire [7:0]         regroupV0_hi_lo_hi_36 = {regroupV0_hi_lo_hi_hi_4, regroupV0_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_36 = {regroupV0_hi_lo_hi_36, regroupV0_hi_lo_lo_36};
  wire [3:0]         regroupV0_hi_hi_lo_lo_4 = {regroupV0_hi_34[579:578], regroupV0_hi_34[515:514]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_4 = {regroupV0_hi_34[707:706], regroupV0_hi_34[643:642]};
  wire [7:0]         regroupV0_hi_hi_lo_36 = {regroupV0_hi_hi_lo_hi_4, regroupV0_hi_hi_lo_lo_4};
  wire [3:0]         regroupV0_hi_hi_hi_lo_4 = {regroupV0_hi_34[835:834], regroupV0_hi_34[771:770]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_4 = {regroupV0_hi_34[963:962], regroupV0_hi_34[899:898]};
  wire [7:0]         regroupV0_hi_hi_hi_36 = {regroupV0_hi_hi_hi_hi_4, regroupV0_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_36 = {regroupV0_hi_hi_hi_36, regroupV0_hi_hi_lo_36};
  wire [31:0]        regroupV0_hi_36 = {regroupV0_hi_hi_36, regroupV0_hi_lo_36};
  wire [3:0]         regroupV0_lo_lo_lo_lo_5 = {regroupV0_lo_34[69:68], regroupV0_lo_34[5:4]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_5 = {regroupV0_lo_34[197:196], regroupV0_lo_34[133:132]};
  wire [7:0]         regroupV0_lo_lo_lo_37 = {regroupV0_lo_lo_lo_hi_5, regroupV0_lo_lo_lo_lo_5};
  wire [3:0]         regroupV0_lo_lo_hi_lo_5 = {regroupV0_lo_34[325:324], regroupV0_lo_34[261:260]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_5 = {regroupV0_lo_34[453:452], regroupV0_lo_34[389:388]};
  wire [7:0]         regroupV0_lo_lo_hi_37 = {regroupV0_lo_lo_hi_hi_5, regroupV0_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_37 = {regroupV0_lo_lo_hi_37, regroupV0_lo_lo_lo_37};
  wire [3:0]         regroupV0_lo_hi_lo_lo_5 = {regroupV0_lo_34[581:580], regroupV0_lo_34[517:516]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_5 = {regroupV0_lo_34[709:708], regroupV0_lo_34[645:644]};
  wire [7:0]         regroupV0_lo_hi_lo_37 = {regroupV0_lo_hi_lo_hi_5, regroupV0_lo_hi_lo_lo_5};
  wire [3:0]         regroupV0_lo_hi_hi_lo_5 = {regroupV0_lo_34[837:836], regroupV0_lo_34[773:772]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_5 = {regroupV0_lo_34[965:964], regroupV0_lo_34[901:900]};
  wire [7:0]         regroupV0_lo_hi_hi_37 = {regroupV0_lo_hi_hi_hi_5, regroupV0_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_37 = {regroupV0_lo_hi_hi_37, regroupV0_lo_hi_lo_37};
  wire [31:0]        regroupV0_lo_37 = {regroupV0_lo_hi_37, regroupV0_lo_lo_37};
  wire [3:0]         regroupV0_hi_lo_lo_lo_5 = {regroupV0_hi_34[69:68], regroupV0_hi_34[5:4]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_5 = {regroupV0_hi_34[197:196], regroupV0_hi_34[133:132]};
  wire [7:0]         regroupV0_hi_lo_lo_37 = {regroupV0_hi_lo_lo_hi_5, regroupV0_hi_lo_lo_lo_5};
  wire [3:0]         regroupV0_hi_lo_hi_lo_5 = {regroupV0_hi_34[325:324], regroupV0_hi_34[261:260]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_5 = {regroupV0_hi_34[453:452], regroupV0_hi_34[389:388]};
  wire [7:0]         regroupV0_hi_lo_hi_37 = {regroupV0_hi_lo_hi_hi_5, regroupV0_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_37 = {regroupV0_hi_lo_hi_37, regroupV0_hi_lo_lo_37};
  wire [3:0]         regroupV0_hi_hi_lo_lo_5 = {regroupV0_hi_34[581:580], regroupV0_hi_34[517:516]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_5 = {regroupV0_hi_34[709:708], regroupV0_hi_34[645:644]};
  wire [7:0]         regroupV0_hi_hi_lo_37 = {regroupV0_hi_hi_lo_hi_5, regroupV0_hi_hi_lo_lo_5};
  wire [3:0]         regroupV0_hi_hi_hi_lo_5 = {regroupV0_hi_34[837:836], regroupV0_hi_34[773:772]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_5 = {regroupV0_hi_34[965:964], regroupV0_hi_34[901:900]};
  wire [7:0]         regroupV0_hi_hi_hi_37 = {regroupV0_hi_hi_hi_hi_5, regroupV0_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_37 = {regroupV0_hi_hi_hi_37, regroupV0_hi_hi_lo_37};
  wire [31:0]        regroupV0_hi_37 = {regroupV0_hi_hi_37, regroupV0_hi_lo_37};
  wire [3:0]         regroupV0_lo_lo_lo_lo_6 = {regroupV0_lo_34[71:70], regroupV0_lo_34[7:6]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_6 = {regroupV0_lo_34[199:198], regroupV0_lo_34[135:134]};
  wire [7:0]         regroupV0_lo_lo_lo_38 = {regroupV0_lo_lo_lo_hi_6, regroupV0_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_hi_lo_6 = {regroupV0_lo_34[327:326], regroupV0_lo_34[263:262]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_6 = {regroupV0_lo_34[455:454], regroupV0_lo_34[391:390]};
  wire [7:0]         regroupV0_lo_lo_hi_38 = {regroupV0_lo_lo_hi_hi_6, regroupV0_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_38 = {regroupV0_lo_lo_hi_38, regroupV0_lo_lo_lo_38};
  wire [3:0]         regroupV0_lo_hi_lo_lo_6 = {regroupV0_lo_34[583:582], regroupV0_lo_34[519:518]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_6 = {regroupV0_lo_34[711:710], regroupV0_lo_34[647:646]};
  wire [7:0]         regroupV0_lo_hi_lo_38 = {regroupV0_lo_hi_lo_hi_6, regroupV0_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_hi_lo_6 = {regroupV0_lo_34[839:838], regroupV0_lo_34[775:774]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_6 = {regroupV0_lo_34[967:966], regroupV0_lo_34[903:902]};
  wire [7:0]         regroupV0_lo_hi_hi_38 = {regroupV0_lo_hi_hi_hi_6, regroupV0_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_38 = {regroupV0_lo_hi_hi_38, regroupV0_lo_hi_lo_38};
  wire [31:0]        regroupV0_lo_38 = {regroupV0_lo_hi_38, regroupV0_lo_lo_38};
  wire [3:0]         regroupV0_hi_lo_lo_lo_6 = {regroupV0_hi_34[71:70], regroupV0_hi_34[7:6]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_6 = {regroupV0_hi_34[199:198], regroupV0_hi_34[135:134]};
  wire [7:0]         regroupV0_hi_lo_lo_38 = {regroupV0_hi_lo_lo_hi_6, regroupV0_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_hi_lo_6 = {regroupV0_hi_34[327:326], regroupV0_hi_34[263:262]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_6 = {regroupV0_hi_34[455:454], regroupV0_hi_34[391:390]};
  wire [7:0]         regroupV0_hi_lo_hi_38 = {regroupV0_hi_lo_hi_hi_6, regroupV0_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_38 = {regroupV0_hi_lo_hi_38, regroupV0_hi_lo_lo_38};
  wire [3:0]         regroupV0_hi_hi_lo_lo_6 = {regroupV0_hi_34[583:582], regroupV0_hi_34[519:518]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_6 = {regroupV0_hi_34[711:710], regroupV0_hi_34[647:646]};
  wire [7:0]         regroupV0_hi_hi_lo_38 = {regroupV0_hi_hi_lo_hi_6, regroupV0_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_hi_lo_6 = {regroupV0_hi_34[839:838], regroupV0_hi_34[775:774]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_6 = {regroupV0_hi_34[967:966], regroupV0_hi_34[903:902]};
  wire [7:0]         regroupV0_hi_hi_hi_38 = {regroupV0_hi_hi_hi_hi_6, regroupV0_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_38 = {regroupV0_hi_hi_hi_38, regroupV0_hi_hi_lo_38};
  wire [31:0]        regroupV0_hi_38 = {regroupV0_hi_hi_38, regroupV0_hi_lo_38};
  wire [3:0]         regroupV0_lo_lo_lo_lo_7 = {regroupV0_lo_34[73:72], regroupV0_lo_34[9:8]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_7 = {regroupV0_lo_34[201:200], regroupV0_lo_34[137:136]};
  wire [7:0]         regroupV0_lo_lo_lo_39 = {regroupV0_lo_lo_lo_hi_7, regroupV0_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_hi_lo_7 = {regroupV0_lo_34[329:328], regroupV0_lo_34[265:264]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_7 = {regroupV0_lo_34[457:456], regroupV0_lo_34[393:392]};
  wire [7:0]         regroupV0_lo_lo_hi_39 = {regroupV0_lo_lo_hi_hi_7, regroupV0_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_39 = {regroupV0_lo_lo_hi_39, regroupV0_lo_lo_lo_39};
  wire [3:0]         regroupV0_lo_hi_lo_lo_7 = {regroupV0_lo_34[585:584], regroupV0_lo_34[521:520]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_7 = {regroupV0_lo_34[713:712], regroupV0_lo_34[649:648]};
  wire [7:0]         regroupV0_lo_hi_lo_39 = {regroupV0_lo_hi_lo_hi_7, regroupV0_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_hi_lo_7 = {regroupV0_lo_34[841:840], regroupV0_lo_34[777:776]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_7 = {regroupV0_lo_34[969:968], regroupV0_lo_34[905:904]};
  wire [7:0]         regroupV0_lo_hi_hi_39 = {regroupV0_lo_hi_hi_hi_7, regroupV0_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_39 = {regroupV0_lo_hi_hi_39, regroupV0_lo_hi_lo_39};
  wire [31:0]        regroupV0_lo_39 = {regroupV0_lo_hi_39, regroupV0_lo_lo_39};
  wire [3:0]         regroupV0_hi_lo_lo_lo_7 = {regroupV0_hi_34[73:72], regroupV0_hi_34[9:8]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_7 = {regroupV0_hi_34[201:200], regroupV0_hi_34[137:136]};
  wire [7:0]         regroupV0_hi_lo_lo_39 = {regroupV0_hi_lo_lo_hi_7, regroupV0_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_hi_lo_7 = {regroupV0_hi_34[329:328], regroupV0_hi_34[265:264]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_7 = {regroupV0_hi_34[457:456], regroupV0_hi_34[393:392]};
  wire [7:0]         regroupV0_hi_lo_hi_39 = {regroupV0_hi_lo_hi_hi_7, regroupV0_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_39 = {regroupV0_hi_lo_hi_39, regroupV0_hi_lo_lo_39};
  wire [3:0]         regroupV0_hi_hi_lo_lo_7 = {regroupV0_hi_34[585:584], regroupV0_hi_34[521:520]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_7 = {regroupV0_hi_34[713:712], regroupV0_hi_34[649:648]};
  wire [7:0]         regroupV0_hi_hi_lo_39 = {regroupV0_hi_hi_lo_hi_7, regroupV0_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_hi_lo_7 = {regroupV0_hi_34[841:840], regroupV0_hi_34[777:776]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_7 = {regroupV0_hi_34[969:968], regroupV0_hi_34[905:904]};
  wire [7:0]         regroupV0_hi_hi_hi_39 = {regroupV0_hi_hi_hi_hi_7, regroupV0_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_39 = {regroupV0_hi_hi_hi_39, regroupV0_hi_hi_lo_39};
  wire [31:0]        regroupV0_hi_39 = {regroupV0_hi_hi_39, regroupV0_hi_lo_39};
  wire [3:0]         regroupV0_lo_lo_lo_lo_8 = {regroupV0_lo_34[75:74], regroupV0_lo_34[11:10]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_8 = {regroupV0_lo_34[203:202], regroupV0_lo_34[139:138]};
  wire [7:0]         regroupV0_lo_lo_lo_40 = {regroupV0_lo_lo_lo_hi_8, regroupV0_lo_lo_lo_lo_8};
  wire [3:0]         regroupV0_lo_lo_hi_lo_8 = {regroupV0_lo_34[331:330], regroupV0_lo_34[267:266]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_8 = {regroupV0_lo_34[459:458], regroupV0_lo_34[395:394]};
  wire [7:0]         regroupV0_lo_lo_hi_40 = {regroupV0_lo_lo_hi_hi_8, regroupV0_lo_lo_hi_lo_8};
  wire [15:0]        regroupV0_lo_lo_40 = {regroupV0_lo_lo_hi_40, regroupV0_lo_lo_lo_40};
  wire [3:0]         regroupV0_lo_hi_lo_lo_8 = {regroupV0_lo_34[587:586], regroupV0_lo_34[523:522]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_8 = {regroupV0_lo_34[715:714], regroupV0_lo_34[651:650]};
  wire [7:0]         regroupV0_lo_hi_lo_40 = {regroupV0_lo_hi_lo_hi_8, regroupV0_lo_hi_lo_lo_8};
  wire [3:0]         regroupV0_lo_hi_hi_lo_8 = {regroupV0_lo_34[843:842], regroupV0_lo_34[779:778]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_8 = {regroupV0_lo_34[971:970], regroupV0_lo_34[907:906]};
  wire [7:0]         regroupV0_lo_hi_hi_40 = {regroupV0_lo_hi_hi_hi_8, regroupV0_lo_hi_hi_lo_8};
  wire [15:0]        regroupV0_lo_hi_40 = {regroupV0_lo_hi_hi_40, regroupV0_lo_hi_lo_40};
  wire [31:0]        regroupV0_lo_40 = {regroupV0_lo_hi_40, regroupV0_lo_lo_40};
  wire [3:0]         regroupV0_hi_lo_lo_lo_8 = {regroupV0_hi_34[75:74], regroupV0_hi_34[11:10]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_8 = {regroupV0_hi_34[203:202], regroupV0_hi_34[139:138]};
  wire [7:0]         regroupV0_hi_lo_lo_40 = {regroupV0_hi_lo_lo_hi_8, regroupV0_hi_lo_lo_lo_8};
  wire [3:0]         regroupV0_hi_lo_hi_lo_8 = {regroupV0_hi_34[331:330], regroupV0_hi_34[267:266]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_8 = {regroupV0_hi_34[459:458], regroupV0_hi_34[395:394]};
  wire [7:0]         regroupV0_hi_lo_hi_40 = {regroupV0_hi_lo_hi_hi_8, regroupV0_hi_lo_hi_lo_8};
  wire [15:0]        regroupV0_hi_lo_40 = {regroupV0_hi_lo_hi_40, regroupV0_hi_lo_lo_40};
  wire [3:0]         regroupV0_hi_hi_lo_lo_8 = {regroupV0_hi_34[587:586], regroupV0_hi_34[523:522]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_8 = {regroupV0_hi_34[715:714], regroupV0_hi_34[651:650]};
  wire [7:0]         regroupV0_hi_hi_lo_40 = {regroupV0_hi_hi_lo_hi_8, regroupV0_hi_hi_lo_lo_8};
  wire [3:0]         regroupV0_hi_hi_hi_lo_8 = {regroupV0_hi_34[843:842], regroupV0_hi_34[779:778]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_8 = {regroupV0_hi_34[971:970], regroupV0_hi_34[907:906]};
  wire [7:0]         regroupV0_hi_hi_hi_40 = {regroupV0_hi_hi_hi_hi_8, regroupV0_hi_hi_hi_lo_8};
  wire [15:0]        regroupV0_hi_hi_40 = {regroupV0_hi_hi_hi_40, regroupV0_hi_hi_lo_40};
  wire [31:0]        regroupV0_hi_40 = {regroupV0_hi_hi_40, regroupV0_hi_lo_40};
  wire [3:0]         regroupV0_lo_lo_lo_lo_9 = {regroupV0_lo_34[77:76], regroupV0_lo_34[13:12]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_9 = {regroupV0_lo_34[205:204], regroupV0_lo_34[141:140]};
  wire [7:0]         regroupV0_lo_lo_lo_41 = {regroupV0_lo_lo_lo_hi_9, regroupV0_lo_lo_lo_lo_9};
  wire [3:0]         regroupV0_lo_lo_hi_lo_9 = {regroupV0_lo_34[333:332], regroupV0_lo_34[269:268]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_9 = {regroupV0_lo_34[461:460], regroupV0_lo_34[397:396]};
  wire [7:0]         regroupV0_lo_lo_hi_41 = {regroupV0_lo_lo_hi_hi_9, regroupV0_lo_lo_hi_lo_9};
  wire [15:0]        regroupV0_lo_lo_41 = {regroupV0_lo_lo_hi_41, regroupV0_lo_lo_lo_41};
  wire [3:0]         regroupV0_lo_hi_lo_lo_9 = {regroupV0_lo_34[589:588], regroupV0_lo_34[525:524]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_9 = {regroupV0_lo_34[717:716], regroupV0_lo_34[653:652]};
  wire [7:0]         regroupV0_lo_hi_lo_41 = {regroupV0_lo_hi_lo_hi_9, regroupV0_lo_hi_lo_lo_9};
  wire [3:0]         regroupV0_lo_hi_hi_lo_9 = {regroupV0_lo_34[845:844], regroupV0_lo_34[781:780]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_9 = {regroupV0_lo_34[973:972], regroupV0_lo_34[909:908]};
  wire [7:0]         regroupV0_lo_hi_hi_41 = {regroupV0_lo_hi_hi_hi_9, regroupV0_lo_hi_hi_lo_9};
  wire [15:0]        regroupV0_lo_hi_41 = {regroupV0_lo_hi_hi_41, regroupV0_lo_hi_lo_41};
  wire [31:0]        regroupV0_lo_41 = {regroupV0_lo_hi_41, regroupV0_lo_lo_41};
  wire [3:0]         regroupV0_hi_lo_lo_lo_9 = {regroupV0_hi_34[77:76], regroupV0_hi_34[13:12]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_9 = {regroupV0_hi_34[205:204], regroupV0_hi_34[141:140]};
  wire [7:0]         regroupV0_hi_lo_lo_41 = {regroupV0_hi_lo_lo_hi_9, regroupV0_hi_lo_lo_lo_9};
  wire [3:0]         regroupV0_hi_lo_hi_lo_9 = {regroupV0_hi_34[333:332], regroupV0_hi_34[269:268]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_9 = {regroupV0_hi_34[461:460], regroupV0_hi_34[397:396]};
  wire [7:0]         regroupV0_hi_lo_hi_41 = {regroupV0_hi_lo_hi_hi_9, regroupV0_hi_lo_hi_lo_9};
  wire [15:0]        regroupV0_hi_lo_41 = {regroupV0_hi_lo_hi_41, regroupV0_hi_lo_lo_41};
  wire [3:0]         regroupV0_hi_hi_lo_lo_9 = {regroupV0_hi_34[589:588], regroupV0_hi_34[525:524]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_9 = {regroupV0_hi_34[717:716], regroupV0_hi_34[653:652]};
  wire [7:0]         regroupV0_hi_hi_lo_41 = {regroupV0_hi_hi_lo_hi_9, regroupV0_hi_hi_lo_lo_9};
  wire [3:0]         regroupV0_hi_hi_hi_lo_9 = {regroupV0_hi_34[845:844], regroupV0_hi_34[781:780]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_9 = {regroupV0_hi_34[973:972], regroupV0_hi_34[909:908]};
  wire [7:0]         regroupV0_hi_hi_hi_41 = {regroupV0_hi_hi_hi_hi_9, regroupV0_hi_hi_hi_lo_9};
  wire [15:0]        regroupV0_hi_hi_41 = {regroupV0_hi_hi_hi_41, regroupV0_hi_hi_lo_41};
  wire [31:0]        regroupV0_hi_41 = {regroupV0_hi_hi_41, regroupV0_hi_lo_41};
  wire [3:0]         regroupV0_lo_lo_lo_lo_10 = {regroupV0_lo_34[79:78], regroupV0_lo_34[15:14]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_10 = {regroupV0_lo_34[207:206], regroupV0_lo_34[143:142]};
  wire [7:0]         regroupV0_lo_lo_lo_42 = {regroupV0_lo_lo_lo_hi_10, regroupV0_lo_lo_lo_lo_10};
  wire [3:0]         regroupV0_lo_lo_hi_lo_10 = {regroupV0_lo_34[335:334], regroupV0_lo_34[271:270]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_10 = {regroupV0_lo_34[463:462], regroupV0_lo_34[399:398]};
  wire [7:0]         regroupV0_lo_lo_hi_42 = {regroupV0_lo_lo_hi_hi_10, regroupV0_lo_lo_hi_lo_10};
  wire [15:0]        regroupV0_lo_lo_42 = {regroupV0_lo_lo_hi_42, regroupV0_lo_lo_lo_42};
  wire [3:0]         regroupV0_lo_hi_lo_lo_10 = {regroupV0_lo_34[591:590], regroupV0_lo_34[527:526]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_10 = {regroupV0_lo_34[719:718], regroupV0_lo_34[655:654]};
  wire [7:0]         regroupV0_lo_hi_lo_42 = {regroupV0_lo_hi_lo_hi_10, regroupV0_lo_hi_lo_lo_10};
  wire [3:0]         regroupV0_lo_hi_hi_lo_10 = {regroupV0_lo_34[847:846], regroupV0_lo_34[783:782]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_10 = {regroupV0_lo_34[975:974], regroupV0_lo_34[911:910]};
  wire [7:0]         regroupV0_lo_hi_hi_42 = {regroupV0_lo_hi_hi_hi_10, regroupV0_lo_hi_hi_lo_10};
  wire [15:0]        regroupV0_lo_hi_42 = {regroupV0_lo_hi_hi_42, regroupV0_lo_hi_lo_42};
  wire [31:0]        regroupV0_lo_42 = {regroupV0_lo_hi_42, regroupV0_lo_lo_42};
  wire [3:0]         regroupV0_hi_lo_lo_lo_10 = {regroupV0_hi_34[79:78], regroupV0_hi_34[15:14]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_10 = {regroupV0_hi_34[207:206], regroupV0_hi_34[143:142]};
  wire [7:0]         regroupV0_hi_lo_lo_42 = {regroupV0_hi_lo_lo_hi_10, regroupV0_hi_lo_lo_lo_10};
  wire [3:0]         regroupV0_hi_lo_hi_lo_10 = {regroupV0_hi_34[335:334], regroupV0_hi_34[271:270]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_10 = {regroupV0_hi_34[463:462], regroupV0_hi_34[399:398]};
  wire [7:0]         regroupV0_hi_lo_hi_42 = {regroupV0_hi_lo_hi_hi_10, regroupV0_hi_lo_hi_lo_10};
  wire [15:0]        regroupV0_hi_lo_42 = {regroupV0_hi_lo_hi_42, regroupV0_hi_lo_lo_42};
  wire [3:0]         regroupV0_hi_hi_lo_lo_10 = {regroupV0_hi_34[591:590], regroupV0_hi_34[527:526]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_10 = {regroupV0_hi_34[719:718], regroupV0_hi_34[655:654]};
  wire [7:0]         regroupV0_hi_hi_lo_42 = {regroupV0_hi_hi_lo_hi_10, regroupV0_hi_hi_lo_lo_10};
  wire [3:0]         regroupV0_hi_hi_hi_lo_10 = {regroupV0_hi_34[847:846], regroupV0_hi_34[783:782]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_10 = {regroupV0_hi_34[975:974], regroupV0_hi_34[911:910]};
  wire [7:0]         regroupV0_hi_hi_hi_42 = {regroupV0_hi_hi_hi_hi_10, regroupV0_hi_hi_hi_lo_10};
  wire [15:0]        regroupV0_hi_hi_42 = {regroupV0_hi_hi_hi_42, regroupV0_hi_hi_lo_42};
  wire [31:0]        regroupV0_hi_42 = {regroupV0_hi_hi_42, regroupV0_hi_lo_42};
  wire [3:0]         regroupV0_lo_lo_lo_lo_11 = {regroupV0_lo_34[81:80], regroupV0_lo_34[17:16]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_11 = {regroupV0_lo_34[209:208], regroupV0_lo_34[145:144]};
  wire [7:0]         regroupV0_lo_lo_lo_43 = {regroupV0_lo_lo_lo_hi_11, regroupV0_lo_lo_lo_lo_11};
  wire [3:0]         regroupV0_lo_lo_hi_lo_11 = {regroupV0_lo_34[337:336], regroupV0_lo_34[273:272]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_11 = {regroupV0_lo_34[465:464], regroupV0_lo_34[401:400]};
  wire [7:0]         regroupV0_lo_lo_hi_43 = {regroupV0_lo_lo_hi_hi_11, regroupV0_lo_lo_hi_lo_11};
  wire [15:0]        regroupV0_lo_lo_43 = {regroupV0_lo_lo_hi_43, regroupV0_lo_lo_lo_43};
  wire [3:0]         regroupV0_lo_hi_lo_lo_11 = {regroupV0_lo_34[593:592], regroupV0_lo_34[529:528]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_11 = {regroupV0_lo_34[721:720], regroupV0_lo_34[657:656]};
  wire [7:0]         regroupV0_lo_hi_lo_43 = {regroupV0_lo_hi_lo_hi_11, regroupV0_lo_hi_lo_lo_11};
  wire [3:0]         regroupV0_lo_hi_hi_lo_11 = {regroupV0_lo_34[849:848], regroupV0_lo_34[785:784]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_11 = {regroupV0_lo_34[977:976], regroupV0_lo_34[913:912]};
  wire [7:0]         regroupV0_lo_hi_hi_43 = {regroupV0_lo_hi_hi_hi_11, regroupV0_lo_hi_hi_lo_11};
  wire [15:0]        regroupV0_lo_hi_43 = {regroupV0_lo_hi_hi_43, regroupV0_lo_hi_lo_43};
  wire [31:0]        regroupV0_lo_43 = {regroupV0_lo_hi_43, regroupV0_lo_lo_43};
  wire [3:0]         regroupV0_hi_lo_lo_lo_11 = {regroupV0_hi_34[81:80], regroupV0_hi_34[17:16]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_11 = {regroupV0_hi_34[209:208], regroupV0_hi_34[145:144]};
  wire [7:0]         regroupV0_hi_lo_lo_43 = {regroupV0_hi_lo_lo_hi_11, regroupV0_hi_lo_lo_lo_11};
  wire [3:0]         regroupV0_hi_lo_hi_lo_11 = {regroupV0_hi_34[337:336], regroupV0_hi_34[273:272]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_11 = {regroupV0_hi_34[465:464], regroupV0_hi_34[401:400]};
  wire [7:0]         regroupV0_hi_lo_hi_43 = {regroupV0_hi_lo_hi_hi_11, regroupV0_hi_lo_hi_lo_11};
  wire [15:0]        regroupV0_hi_lo_43 = {regroupV0_hi_lo_hi_43, regroupV0_hi_lo_lo_43};
  wire [3:0]         regroupV0_hi_hi_lo_lo_11 = {regroupV0_hi_34[593:592], regroupV0_hi_34[529:528]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_11 = {regroupV0_hi_34[721:720], regroupV0_hi_34[657:656]};
  wire [7:0]         regroupV0_hi_hi_lo_43 = {regroupV0_hi_hi_lo_hi_11, regroupV0_hi_hi_lo_lo_11};
  wire [3:0]         regroupV0_hi_hi_hi_lo_11 = {regroupV0_hi_34[849:848], regroupV0_hi_34[785:784]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_11 = {regroupV0_hi_34[977:976], regroupV0_hi_34[913:912]};
  wire [7:0]         regroupV0_hi_hi_hi_43 = {regroupV0_hi_hi_hi_hi_11, regroupV0_hi_hi_hi_lo_11};
  wire [15:0]        regroupV0_hi_hi_43 = {regroupV0_hi_hi_hi_43, regroupV0_hi_hi_lo_43};
  wire [31:0]        regroupV0_hi_43 = {regroupV0_hi_hi_43, regroupV0_hi_lo_43};
  wire [3:0]         regroupV0_lo_lo_lo_lo_12 = {regroupV0_lo_34[83:82], regroupV0_lo_34[19:18]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_12 = {regroupV0_lo_34[211:210], regroupV0_lo_34[147:146]};
  wire [7:0]         regroupV0_lo_lo_lo_44 = {regroupV0_lo_lo_lo_hi_12, regroupV0_lo_lo_lo_lo_12};
  wire [3:0]         regroupV0_lo_lo_hi_lo_12 = {regroupV0_lo_34[339:338], regroupV0_lo_34[275:274]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_12 = {regroupV0_lo_34[467:466], regroupV0_lo_34[403:402]};
  wire [7:0]         regroupV0_lo_lo_hi_44 = {regroupV0_lo_lo_hi_hi_12, regroupV0_lo_lo_hi_lo_12};
  wire [15:0]        regroupV0_lo_lo_44 = {regroupV0_lo_lo_hi_44, regroupV0_lo_lo_lo_44};
  wire [3:0]         regroupV0_lo_hi_lo_lo_12 = {regroupV0_lo_34[595:594], regroupV0_lo_34[531:530]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_12 = {regroupV0_lo_34[723:722], regroupV0_lo_34[659:658]};
  wire [7:0]         regroupV0_lo_hi_lo_44 = {regroupV0_lo_hi_lo_hi_12, regroupV0_lo_hi_lo_lo_12};
  wire [3:0]         regroupV0_lo_hi_hi_lo_12 = {regroupV0_lo_34[851:850], regroupV0_lo_34[787:786]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_12 = {regroupV0_lo_34[979:978], regroupV0_lo_34[915:914]};
  wire [7:0]         regroupV0_lo_hi_hi_44 = {regroupV0_lo_hi_hi_hi_12, regroupV0_lo_hi_hi_lo_12};
  wire [15:0]        regroupV0_lo_hi_44 = {regroupV0_lo_hi_hi_44, regroupV0_lo_hi_lo_44};
  wire [31:0]        regroupV0_lo_44 = {regroupV0_lo_hi_44, regroupV0_lo_lo_44};
  wire [3:0]         regroupV0_hi_lo_lo_lo_12 = {regroupV0_hi_34[83:82], regroupV0_hi_34[19:18]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_12 = {regroupV0_hi_34[211:210], regroupV0_hi_34[147:146]};
  wire [7:0]         regroupV0_hi_lo_lo_44 = {regroupV0_hi_lo_lo_hi_12, regroupV0_hi_lo_lo_lo_12};
  wire [3:0]         regroupV0_hi_lo_hi_lo_12 = {regroupV0_hi_34[339:338], regroupV0_hi_34[275:274]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_12 = {regroupV0_hi_34[467:466], regroupV0_hi_34[403:402]};
  wire [7:0]         regroupV0_hi_lo_hi_44 = {regroupV0_hi_lo_hi_hi_12, regroupV0_hi_lo_hi_lo_12};
  wire [15:0]        regroupV0_hi_lo_44 = {regroupV0_hi_lo_hi_44, regroupV0_hi_lo_lo_44};
  wire [3:0]         regroupV0_hi_hi_lo_lo_12 = {regroupV0_hi_34[595:594], regroupV0_hi_34[531:530]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_12 = {regroupV0_hi_34[723:722], regroupV0_hi_34[659:658]};
  wire [7:0]         regroupV0_hi_hi_lo_44 = {regroupV0_hi_hi_lo_hi_12, regroupV0_hi_hi_lo_lo_12};
  wire [3:0]         regroupV0_hi_hi_hi_lo_12 = {regroupV0_hi_34[851:850], regroupV0_hi_34[787:786]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_12 = {regroupV0_hi_34[979:978], regroupV0_hi_34[915:914]};
  wire [7:0]         regroupV0_hi_hi_hi_44 = {regroupV0_hi_hi_hi_hi_12, regroupV0_hi_hi_hi_lo_12};
  wire [15:0]        regroupV0_hi_hi_44 = {regroupV0_hi_hi_hi_44, regroupV0_hi_hi_lo_44};
  wire [31:0]        regroupV0_hi_44 = {regroupV0_hi_hi_44, regroupV0_hi_lo_44};
  wire [3:0]         regroupV0_lo_lo_lo_lo_13 = {regroupV0_lo_34[85:84], regroupV0_lo_34[21:20]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_13 = {regroupV0_lo_34[213:212], regroupV0_lo_34[149:148]};
  wire [7:0]         regroupV0_lo_lo_lo_45 = {regroupV0_lo_lo_lo_hi_13, regroupV0_lo_lo_lo_lo_13};
  wire [3:0]         regroupV0_lo_lo_hi_lo_13 = {regroupV0_lo_34[341:340], regroupV0_lo_34[277:276]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_13 = {regroupV0_lo_34[469:468], regroupV0_lo_34[405:404]};
  wire [7:0]         regroupV0_lo_lo_hi_45 = {regroupV0_lo_lo_hi_hi_13, regroupV0_lo_lo_hi_lo_13};
  wire [15:0]        regroupV0_lo_lo_45 = {regroupV0_lo_lo_hi_45, regroupV0_lo_lo_lo_45};
  wire [3:0]         regroupV0_lo_hi_lo_lo_13 = {regroupV0_lo_34[597:596], regroupV0_lo_34[533:532]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_13 = {regroupV0_lo_34[725:724], regroupV0_lo_34[661:660]};
  wire [7:0]         regroupV0_lo_hi_lo_45 = {regroupV0_lo_hi_lo_hi_13, regroupV0_lo_hi_lo_lo_13};
  wire [3:0]         regroupV0_lo_hi_hi_lo_13 = {regroupV0_lo_34[853:852], regroupV0_lo_34[789:788]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_13 = {regroupV0_lo_34[981:980], regroupV0_lo_34[917:916]};
  wire [7:0]         regroupV0_lo_hi_hi_45 = {regroupV0_lo_hi_hi_hi_13, regroupV0_lo_hi_hi_lo_13};
  wire [15:0]        regroupV0_lo_hi_45 = {regroupV0_lo_hi_hi_45, regroupV0_lo_hi_lo_45};
  wire [31:0]        regroupV0_lo_45 = {regroupV0_lo_hi_45, regroupV0_lo_lo_45};
  wire [3:0]         regroupV0_hi_lo_lo_lo_13 = {regroupV0_hi_34[85:84], regroupV0_hi_34[21:20]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_13 = {regroupV0_hi_34[213:212], regroupV0_hi_34[149:148]};
  wire [7:0]         regroupV0_hi_lo_lo_45 = {regroupV0_hi_lo_lo_hi_13, regroupV0_hi_lo_lo_lo_13};
  wire [3:0]         regroupV0_hi_lo_hi_lo_13 = {regroupV0_hi_34[341:340], regroupV0_hi_34[277:276]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_13 = {regroupV0_hi_34[469:468], regroupV0_hi_34[405:404]};
  wire [7:0]         regroupV0_hi_lo_hi_45 = {regroupV0_hi_lo_hi_hi_13, regroupV0_hi_lo_hi_lo_13};
  wire [15:0]        regroupV0_hi_lo_45 = {regroupV0_hi_lo_hi_45, regroupV0_hi_lo_lo_45};
  wire [3:0]         regroupV0_hi_hi_lo_lo_13 = {regroupV0_hi_34[597:596], regroupV0_hi_34[533:532]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_13 = {regroupV0_hi_34[725:724], regroupV0_hi_34[661:660]};
  wire [7:0]         regroupV0_hi_hi_lo_45 = {regroupV0_hi_hi_lo_hi_13, regroupV0_hi_hi_lo_lo_13};
  wire [3:0]         regroupV0_hi_hi_hi_lo_13 = {regroupV0_hi_34[853:852], regroupV0_hi_34[789:788]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_13 = {regroupV0_hi_34[981:980], regroupV0_hi_34[917:916]};
  wire [7:0]         regroupV0_hi_hi_hi_45 = {regroupV0_hi_hi_hi_hi_13, regroupV0_hi_hi_hi_lo_13};
  wire [15:0]        regroupV0_hi_hi_45 = {regroupV0_hi_hi_hi_45, regroupV0_hi_hi_lo_45};
  wire [31:0]        regroupV0_hi_45 = {regroupV0_hi_hi_45, regroupV0_hi_lo_45};
  wire [3:0]         regroupV0_lo_lo_lo_lo_14 = {regroupV0_lo_34[87:86], regroupV0_lo_34[23:22]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_14 = {regroupV0_lo_34[215:214], regroupV0_lo_34[151:150]};
  wire [7:0]         regroupV0_lo_lo_lo_46 = {regroupV0_lo_lo_lo_hi_14, regroupV0_lo_lo_lo_lo_14};
  wire [3:0]         regroupV0_lo_lo_hi_lo_14 = {regroupV0_lo_34[343:342], regroupV0_lo_34[279:278]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_14 = {regroupV0_lo_34[471:470], regroupV0_lo_34[407:406]};
  wire [7:0]         regroupV0_lo_lo_hi_46 = {regroupV0_lo_lo_hi_hi_14, regroupV0_lo_lo_hi_lo_14};
  wire [15:0]        regroupV0_lo_lo_46 = {regroupV0_lo_lo_hi_46, regroupV0_lo_lo_lo_46};
  wire [3:0]         regroupV0_lo_hi_lo_lo_14 = {regroupV0_lo_34[599:598], regroupV0_lo_34[535:534]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_14 = {regroupV0_lo_34[727:726], regroupV0_lo_34[663:662]};
  wire [7:0]         regroupV0_lo_hi_lo_46 = {regroupV0_lo_hi_lo_hi_14, regroupV0_lo_hi_lo_lo_14};
  wire [3:0]         regroupV0_lo_hi_hi_lo_14 = {regroupV0_lo_34[855:854], regroupV0_lo_34[791:790]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_14 = {regroupV0_lo_34[983:982], regroupV0_lo_34[919:918]};
  wire [7:0]         regroupV0_lo_hi_hi_46 = {regroupV0_lo_hi_hi_hi_14, regroupV0_lo_hi_hi_lo_14};
  wire [15:0]        regroupV0_lo_hi_46 = {regroupV0_lo_hi_hi_46, regroupV0_lo_hi_lo_46};
  wire [31:0]        regroupV0_lo_46 = {regroupV0_lo_hi_46, regroupV0_lo_lo_46};
  wire [3:0]         regroupV0_hi_lo_lo_lo_14 = {regroupV0_hi_34[87:86], regroupV0_hi_34[23:22]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_14 = {regroupV0_hi_34[215:214], regroupV0_hi_34[151:150]};
  wire [7:0]         regroupV0_hi_lo_lo_46 = {regroupV0_hi_lo_lo_hi_14, regroupV0_hi_lo_lo_lo_14};
  wire [3:0]         regroupV0_hi_lo_hi_lo_14 = {regroupV0_hi_34[343:342], regroupV0_hi_34[279:278]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_14 = {regroupV0_hi_34[471:470], regroupV0_hi_34[407:406]};
  wire [7:0]         regroupV0_hi_lo_hi_46 = {regroupV0_hi_lo_hi_hi_14, regroupV0_hi_lo_hi_lo_14};
  wire [15:0]        regroupV0_hi_lo_46 = {regroupV0_hi_lo_hi_46, regroupV0_hi_lo_lo_46};
  wire [3:0]         regroupV0_hi_hi_lo_lo_14 = {regroupV0_hi_34[599:598], regroupV0_hi_34[535:534]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_14 = {regroupV0_hi_34[727:726], regroupV0_hi_34[663:662]};
  wire [7:0]         regroupV0_hi_hi_lo_46 = {regroupV0_hi_hi_lo_hi_14, regroupV0_hi_hi_lo_lo_14};
  wire [3:0]         regroupV0_hi_hi_hi_lo_14 = {regroupV0_hi_34[855:854], regroupV0_hi_34[791:790]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_14 = {regroupV0_hi_34[983:982], regroupV0_hi_34[919:918]};
  wire [7:0]         regroupV0_hi_hi_hi_46 = {regroupV0_hi_hi_hi_hi_14, regroupV0_hi_hi_hi_lo_14};
  wire [15:0]        regroupV0_hi_hi_46 = {regroupV0_hi_hi_hi_46, regroupV0_hi_hi_lo_46};
  wire [31:0]        regroupV0_hi_46 = {regroupV0_hi_hi_46, regroupV0_hi_lo_46};
  wire [3:0]         regroupV0_lo_lo_lo_lo_15 = {regroupV0_lo_34[89:88], regroupV0_lo_34[25:24]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_15 = {regroupV0_lo_34[217:216], regroupV0_lo_34[153:152]};
  wire [7:0]         regroupV0_lo_lo_lo_47 = {regroupV0_lo_lo_lo_hi_15, regroupV0_lo_lo_lo_lo_15};
  wire [3:0]         regroupV0_lo_lo_hi_lo_15 = {regroupV0_lo_34[345:344], regroupV0_lo_34[281:280]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_15 = {regroupV0_lo_34[473:472], regroupV0_lo_34[409:408]};
  wire [7:0]         regroupV0_lo_lo_hi_47 = {regroupV0_lo_lo_hi_hi_15, regroupV0_lo_lo_hi_lo_15};
  wire [15:0]        regroupV0_lo_lo_47 = {regroupV0_lo_lo_hi_47, regroupV0_lo_lo_lo_47};
  wire [3:0]         regroupV0_lo_hi_lo_lo_15 = {regroupV0_lo_34[601:600], regroupV0_lo_34[537:536]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_15 = {regroupV0_lo_34[729:728], regroupV0_lo_34[665:664]};
  wire [7:0]         regroupV0_lo_hi_lo_47 = {regroupV0_lo_hi_lo_hi_15, regroupV0_lo_hi_lo_lo_15};
  wire [3:0]         regroupV0_lo_hi_hi_lo_15 = {regroupV0_lo_34[857:856], regroupV0_lo_34[793:792]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_15 = {regroupV0_lo_34[985:984], regroupV0_lo_34[921:920]};
  wire [7:0]         regroupV0_lo_hi_hi_47 = {regroupV0_lo_hi_hi_hi_15, regroupV0_lo_hi_hi_lo_15};
  wire [15:0]        regroupV0_lo_hi_47 = {regroupV0_lo_hi_hi_47, regroupV0_lo_hi_lo_47};
  wire [31:0]        regroupV0_lo_47 = {regroupV0_lo_hi_47, regroupV0_lo_lo_47};
  wire [3:0]         regroupV0_hi_lo_lo_lo_15 = {regroupV0_hi_34[89:88], regroupV0_hi_34[25:24]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_15 = {regroupV0_hi_34[217:216], regroupV0_hi_34[153:152]};
  wire [7:0]         regroupV0_hi_lo_lo_47 = {regroupV0_hi_lo_lo_hi_15, regroupV0_hi_lo_lo_lo_15};
  wire [3:0]         regroupV0_hi_lo_hi_lo_15 = {regroupV0_hi_34[345:344], regroupV0_hi_34[281:280]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_15 = {regroupV0_hi_34[473:472], regroupV0_hi_34[409:408]};
  wire [7:0]         regroupV0_hi_lo_hi_47 = {regroupV0_hi_lo_hi_hi_15, regroupV0_hi_lo_hi_lo_15};
  wire [15:0]        regroupV0_hi_lo_47 = {regroupV0_hi_lo_hi_47, regroupV0_hi_lo_lo_47};
  wire [3:0]         regroupV0_hi_hi_lo_lo_15 = {regroupV0_hi_34[601:600], regroupV0_hi_34[537:536]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_15 = {regroupV0_hi_34[729:728], regroupV0_hi_34[665:664]};
  wire [7:0]         regroupV0_hi_hi_lo_47 = {regroupV0_hi_hi_lo_hi_15, regroupV0_hi_hi_lo_lo_15};
  wire [3:0]         regroupV0_hi_hi_hi_lo_15 = {regroupV0_hi_34[857:856], regroupV0_hi_34[793:792]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_15 = {regroupV0_hi_34[985:984], regroupV0_hi_34[921:920]};
  wire [7:0]         regroupV0_hi_hi_hi_47 = {regroupV0_hi_hi_hi_hi_15, regroupV0_hi_hi_hi_lo_15};
  wire [15:0]        regroupV0_hi_hi_47 = {regroupV0_hi_hi_hi_47, regroupV0_hi_hi_lo_47};
  wire [31:0]        regroupV0_hi_47 = {regroupV0_hi_hi_47, regroupV0_hi_lo_47};
  wire [3:0]         regroupV0_lo_lo_lo_lo_16 = {regroupV0_lo_34[91:90], regroupV0_lo_34[27:26]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_16 = {regroupV0_lo_34[219:218], regroupV0_lo_34[155:154]};
  wire [7:0]         regroupV0_lo_lo_lo_48 = {regroupV0_lo_lo_lo_hi_16, regroupV0_lo_lo_lo_lo_16};
  wire [3:0]         regroupV0_lo_lo_hi_lo_16 = {regroupV0_lo_34[347:346], regroupV0_lo_34[283:282]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_16 = {regroupV0_lo_34[475:474], regroupV0_lo_34[411:410]};
  wire [7:0]         regroupV0_lo_lo_hi_48 = {regroupV0_lo_lo_hi_hi_16, regroupV0_lo_lo_hi_lo_16};
  wire [15:0]        regroupV0_lo_lo_48 = {regroupV0_lo_lo_hi_48, regroupV0_lo_lo_lo_48};
  wire [3:0]         regroupV0_lo_hi_lo_lo_16 = {regroupV0_lo_34[603:602], regroupV0_lo_34[539:538]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_16 = {regroupV0_lo_34[731:730], regroupV0_lo_34[667:666]};
  wire [7:0]         regroupV0_lo_hi_lo_48 = {regroupV0_lo_hi_lo_hi_16, regroupV0_lo_hi_lo_lo_16};
  wire [3:0]         regroupV0_lo_hi_hi_lo_16 = {regroupV0_lo_34[859:858], regroupV0_lo_34[795:794]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_16 = {regroupV0_lo_34[987:986], regroupV0_lo_34[923:922]};
  wire [7:0]         regroupV0_lo_hi_hi_48 = {regroupV0_lo_hi_hi_hi_16, regroupV0_lo_hi_hi_lo_16};
  wire [15:0]        regroupV0_lo_hi_48 = {regroupV0_lo_hi_hi_48, regroupV0_lo_hi_lo_48};
  wire [31:0]        regroupV0_lo_48 = {regroupV0_lo_hi_48, regroupV0_lo_lo_48};
  wire [3:0]         regroupV0_hi_lo_lo_lo_16 = {regroupV0_hi_34[91:90], regroupV0_hi_34[27:26]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_16 = {regroupV0_hi_34[219:218], regroupV0_hi_34[155:154]};
  wire [7:0]         regroupV0_hi_lo_lo_48 = {regroupV0_hi_lo_lo_hi_16, regroupV0_hi_lo_lo_lo_16};
  wire [3:0]         regroupV0_hi_lo_hi_lo_16 = {regroupV0_hi_34[347:346], regroupV0_hi_34[283:282]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_16 = {regroupV0_hi_34[475:474], regroupV0_hi_34[411:410]};
  wire [7:0]         regroupV0_hi_lo_hi_48 = {regroupV0_hi_lo_hi_hi_16, regroupV0_hi_lo_hi_lo_16};
  wire [15:0]        regroupV0_hi_lo_48 = {regroupV0_hi_lo_hi_48, regroupV0_hi_lo_lo_48};
  wire [3:0]         regroupV0_hi_hi_lo_lo_16 = {regroupV0_hi_34[603:602], regroupV0_hi_34[539:538]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_16 = {regroupV0_hi_34[731:730], regroupV0_hi_34[667:666]};
  wire [7:0]         regroupV0_hi_hi_lo_48 = {regroupV0_hi_hi_lo_hi_16, regroupV0_hi_hi_lo_lo_16};
  wire [3:0]         regroupV0_hi_hi_hi_lo_16 = {regroupV0_hi_34[859:858], regroupV0_hi_34[795:794]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_16 = {regroupV0_hi_34[987:986], regroupV0_hi_34[923:922]};
  wire [7:0]         regroupV0_hi_hi_hi_48 = {regroupV0_hi_hi_hi_hi_16, regroupV0_hi_hi_hi_lo_16};
  wire [15:0]        regroupV0_hi_hi_48 = {regroupV0_hi_hi_hi_48, regroupV0_hi_hi_lo_48};
  wire [31:0]        regroupV0_hi_48 = {regroupV0_hi_hi_48, regroupV0_hi_lo_48};
  wire [3:0]         regroupV0_lo_lo_lo_lo_17 = {regroupV0_lo_34[93:92], regroupV0_lo_34[29:28]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_17 = {regroupV0_lo_34[221:220], regroupV0_lo_34[157:156]};
  wire [7:0]         regroupV0_lo_lo_lo_49 = {regroupV0_lo_lo_lo_hi_17, regroupV0_lo_lo_lo_lo_17};
  wire [3:0]         regroupV0_lo_lo_hi_lo_17 = {regroupV0_lo_34[349:348], regroupV0_lo_34[285:284]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_17 = {regroupV0_lo_34[477:476], regroupV0_lo_34[413:412]};
  wire [7:0]         regroupV0_lo_lo_hi_49 = {regroupV0_lo_lo_hi_hi_17, regroupV0_lo_lo_hi_lo_17};
  wire [15:0]        regroupV0_lo_lo_49 = {regroupV0_lo_lo_hi_49, regroupV0_lo_lo_lo_49};
  wire [3:0]         regroupV0_lo_hi_lo_lo_17 = {regroupV0_lo_34[605:604], regroupV0_lo_34[541:540]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_17 = {regroupV0_lo_34[733:732], regroupV0_lo_34[669:668]};
  wire [7:0]         regroupV0_lo_hi_lo_49 = {regroupV0_lo_hi_lo_hi_17, regroupV0_lo_hi_lo_lo_17};
  wire [3:0]         regroupV0_lo_hi_hi_lo_17 = {regroupV0_lo_34[861:860], regroupV0_lo_34[797:796]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_17 = {regroupV0_lo_34[989:988], regroupV0_lo_34[925:924]};
  wire [7:0]         regroupV0_lo_hi_hi_49 = {regroupV0_lo_hi_hi_hi_17, regroupV0_lo_hi_hi_lo_17};
  wire [15:0]        regroupV0_lo_hi_49 = {regroupV0_lo_hi_hi_49, regroupV0_lo_hi_lo_49};
  wire [31:0]        regroupV0_lo_49 = {regroupV0_lo_hi_49, regroupV0_lo_lo_49};
  wire [3:0]         regroupV0_hi_lo_lo_lo_17 = {regroupV0_hi_34[93:92], regroupV0_hi_34[29:28]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_17 = {regroupV0_hi_34[221:220], regroupV0_hi_34[157:156]};
  wire [7:0]         regroupV0_hi_lo_lo_49 = {regroupV0_hi_lo_lo_hi_17, regroupV0_hi_lo_lo_lo_17};
  wire [3:0]         regroupV0_hi_lo_hi_lo_17 = {regroupV0_hi_34[349:348], regroupV0_hi_34[285:284]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_17 = {regroupV0_hi_34[477:476], regroupV0_hi_34[413:412]};
  wire [7:0]         regroupV0_hi_lo_hi_49 = {regroupV0_hi_lo_hi_hi_17, regroupV0_hi_lo_hi_lo_17};
  wire [15:0]        regroupV0_hi_lo_49 = {regroupV0_hi_lo_hi_49, regroupV0_hi_lo_lo_49};
  wire [3:0]         regroupV0_hi_hi_lo_lo_17 = {regroupV0_hi_34[605:604], regroupV0_hi_34[541:540]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_17 = {regroupV0_hi_34[733:732], regroupV0_hi_34[669:668]};
  wire [7:0]         regroupV0_hi_hi_lo_49 = {regroupV0_hi_hi_lo_hi_17, regroupV0_hi_hi_lo_lo_17};
  wire [3:0]         regroupV0_hi_hi_hi_lo_17 = {regroupV0_hi_34[861:860], regroupV0_hi_34[797:796]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_17 = {regroupV0_hi_34[989:988], regroupV0_hi_34[925:924]};
  wire [7:0]         regroupV0_hi_hi_hi_49 = {regroupV0_hi_hi_hi_hi_17, regroupV0_hi_hi_hi_lo_17};
  wire [15:0]        regroupV0_hi_hi_49 = {regroupV0_hi_hi_hi_49, regroupV0_hi_hi_lo_49};
  wire [31:0]        regroupV0_hi_49 = {regroupV0_hi_hi_49, regroupV0_hi_lo_49};
  wire [3:0]         regroupV0_lo_lo_lo_lo_18 = {regroupV0_lo_34[95:94], regroupV0_lo_34[31:30]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_18 = {regroupV0_lo_34[223:222], regroupV0_lo_34[159:158]};
  wire [7:0]         regroupV0_lo_lo_lo_50 = {regroupV0_lo_lo_lo_hi_18, regroupV0_lo_lo_lo_lo_18};
  wire [3:0]         regroupV0_lo_lo_hi_lo_18 = {regroupV0_lo_34[351:350], regroupV0_lo_34[287:286]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_18 = {regroupV0_lo_34[479:478], regroupV0_lo_34[415:414]};
  wire [7:0]         regroupV0_lo_lo_hi_50 = {regroupV0_lo_lo_hi_hi_18, regroupV0_lo_lo_hi_lo_18};
  wire [15:0]        regroupV0_lo_lo_50 = {regroupV0_lo_lo_hi_50, regroupV0_lo_lo_lo_50};
  wire [3:0]         regroupV0_lo_hi_lo_lo_18 = {regroupV0_lo_34[607:606], regroupV0_lo_34[543:542]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_18 = {regroupV0_lo_34[735:734], regroupV0_lo_34[671:670]};
  wire [7:0]         regroupV0_lo_hi_lo_50 = {regroupV0_lo_hi_lo_hi_18, regroupV0_lo_hi_lo_lo_18};
  wire [3:0]         regroupV0_lo_hi_hi_lo_18 = {regroupV0_lo_34[863:862], regroupV0_lo_34[799:798]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_18 = {regroupV0_lo_34[991:990], regroupV0_lo_34[927:926]};
  wire [7:0]         regroupV0_lo_hi_hi_50 = {regroupV0_lo_hi_hi_hi_18, regroupV0_lo_hi_hi_lo_18};
  wire [15:0]        regroupV0_lo_hi_50 = {regroupV0_lo_hi_hi_50, regroupV0_lo_hi_lo_50};
  wire [31:0]        regroupV0_lo_50 = {regroupV0_lo_hi_50, regroupV0_lo_lo_50};
  wire [3:0]         regroupV0_hi_lo_lo_lo_18 = {regroupV0_hi_34[95:94], regroupV0_hi_34[31:30]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_18 = {regroupV0_hi_34[223:222], regroupV0_hi_34[159:158]};
  wire [7:0]         regroupV0_hi_lo_lo_50 = {regroupV0_hi_lo_lo_hi_18, regroupV0_hi_lo_lo_lo_18};
  wire [3:0]         regroupV0_hi_lo_hi_lo_18 = {regroupV0_hi_34[351:350], regroupV0_hi_34[287:286]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_18 = {regroupV0_hi_34[479:478], regroupV0_hi_34[415:414]};
  wire [7:0]         regroupV0_hi_lo_hi_50 = {regroupV0_hi_lo_hi_hi_18, regroupV0_hi_lo_hi_lo_18};
  wire [15:0]        regroupV0_hi_lo_50 = {regroupV0_hi_lo_hi_50, regroupV0_hi_lo_lo_50};
  wire [3:0]         regroupV0_hi_hi_lo_lo_18 = {regroupV0_hi_34[607:606], regroupV0_hi_34[543:542]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_18 = {regroupV0_hi_34[735:734], regroupV0_hi_34[671:670]};
  wire [7:0]         regroupV0_hi_hi_lo_50 = {regroupV0_hi_hi_lo_hi_18, regroupV0_hi_hi_lo_lo_18};
  wire [3:0]         regroupV0_hi_hi_hi_lo_18 = {regroupV0_hi_34[863:862], regroupV0_hi_34[799:798]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_18 = {regroupV0_hi_34[991:990], regroupV0_hi_34[927:926]};
  wire [7:0]         regroupV0_hi_hi_hi_50 = {regroupV0_hi_hi_hi_hi_18, regroupV0_hi_hi_hi_lo_18};
  wire [15:0]        regroupV0_hi_hi_50 = {regroupV0_hi_hi_hi_50, regroupV0_hi_hi_lo_50};
  wire [31:0]        regroupV0_hi_50 = {regroupV0_hi_hi_50, regroupV0_hi_lo_50};
  wire [3:0]         regroupV0_lo_lo_lo_lo_19 = {regroupV0_lo_34[97:96], regroupV0_lo_34[33:32]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_19 = {regroupV0_lo_34[225:224], regroupV0_lo_34[161:160]};
  wire [7:0]         regroupV0_lo_lo_lo_51 = {regroupV0_lo_lo_lo_hi_19, regroupV0_lo_lo_lo_lo_19};
  wire [3:0]         regroupV0_lo_lo_hi_lo_19 = {regroupV0_lo_34[353:352], regroupV0_lo_34[289:288]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_19 = {regroupV0_lo_34[481:480], regroupV0_lo_34[417:416]};
  wire [7:0]         regroupV0_lo_lo_hi_51 = {regroupV0_lo_lo_hi_hi_19, regroupV0_lo_lo_hi_lo_19};
  wire [15:0]        regroupV0_lo_lo_51 = {regroupV0_lo_lo_hi_51, regroupV0_lo_lo_lo_51};
  wire [3:0]         regroupV0_lo_hi_lo_lo_19 = {regroupV0_lo_34[609:608], regroupV0_lo_34[545:544]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_19 = {regroupV0_lo_34[737:736], regroupV0_lo_34[673:672]};
  wire [7:0]         regroupV0_lo_hi_lo_51 = {regroupV0_lo_hi_lo_hi_19, regroupV0_lo_hi_lo_lo_19};
  wire [3:0]         regroupV0_lo_hi_hi_lo_19 = {regroupV0_lo_34[865:864], regroupV0_lo_34[801:800]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_19 = {regroupV0_lo_34[993:992], regroupV0_lo_34[929:928]};
  wire [7:0]         regroupV0_lo_hi_hi_51 = {regroupV0_lo_hi_hi_hi_19, regroupV0_lo_hi_hi_lo_19};
  wire [15:0]        regroupV0_lo_hi_51 = {regroupV0_lo_hi_hi_51, regroupV0_lo_hi_lo_51};
  wire [31:0]        regroupV0_lo_51 = {regroupV0_lo_hi_51, regroupV0_lo_lo_51};
  wire [3:0]         regroupV0_hi_lo_lo_lo_19 = {regroupV0_hi_34[97:96], regroupV0_hi_34[33:32]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_19 = {regroupV0_hi_34[225:224], regroupV0_hi_34[161:160]};
  wire [7:0]         regroupV0_hi_lo_lo_51 = {regroupV0_hi_lo_lo_hi_19, regroupV0_hi_lo_lo_lo_19};
  wire [3:0]         regroupV0_hi_lo_hi_lo_19 = {regroupV0_hi_34[353:352], regroupV0_hi_34[289:288]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_19 = {regroupV0_hi_34[481:480], regroupV0_hi_34[417:416]};
  wire [7:0]         regroupV0_hi_lo_hi_51 = {regroupV0_hi_lo_hi_hi_19, regroupV0_hi_lo_hi_lo_19};
  wire [15:0]        regroupV0_hi_lo_51 = {regroupV0_hi_lo_hi_51, regroupV0_hi_lo_lo_51};
  wire [3:0]         regroupV0_hi_hi_lo_lo_19 = {regroupV0_hi_34[609:608], regroupV0_hi_34[545:544]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_19 = {regroupV0_hi_34[737:736], regroupV0_hi_34[673:672]};
  wire [7:0]         regroupV0_hi_hi_lo_51 = {regroupV0_hi_hi_lo_hi_19, regroupV0_hi_hi_lo_lo_19};
  wire [3:0]         regroupV0_hi_hi_hi_lo_19 = {regroupV0_hi_34[865:864], regroupV0_hi_34[801:800]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_19 = {regroupV0_hi_34[993:992], regroupV0_hi_34[929:928]};
  wire [7:0]         regroupV0_hi_hi_hi_51 = {regroupV0_hi_hi_hi_hi_19, regroupV0_hi_hi_hi_lo_19};
  wire [15:0]        regroupV0_hi_hi_51 = {regroupV0_hi_hi_hi_51, regroupV0_hi_hi_lo_51};
  wire [31:0]        regroupV0_hi_51 = {regroupV0_hi_hi_51, regroupV0_hi_lo_51};
  wire [3:0]         regroupV0_lo_lo_lo_lo_20 = {regroupV0_lo_34[99:98], regroupV0_lo_34[35:34]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_20 = {regroupV0_lo_34[227:226], regroupV0_lo_34[163:162]};
  wire [7:0]         regroupV0_lo_lo_lo_52 = {regroupV0_lo_lo_lo_hi_20, regroupV0_lo_lo_lo_lo_20};
  wire [3:0]         regroupV0_lo_lo_hi_lo_20 = {regroupV0_lo_34[355:354], regroupV0_lo_34[291:290]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_20 = {regroupV0_lo_34[483:482], regroupV0_lo_34[419:418]};
  wire [7:0]         regroupV0_lo_lo_hi_52 = {regroupV0_lo_lo_hi_hi_20, regroupV0_lo_lo_hi_lo_20};
  wire [15:0]        regroupV0_lo_lo_52 = {regroupV0_lo_lo_hi_52, regroupV0_lo_lo_lo_52};
  wire [3:0]         regroupV0_lo_hi_lo_lo_20 = {regroupV0_lo_34[611:610], regroupV0_lo_34[547:546]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_20 = {regroupV0_lo_34[739:738], regroupV0_lo_34[675:674]};
  wire [7:0]         regroupV0_lo_hi_lo_52 = {regroupV0_lo_hi_lo_hi_20, regroupV0_lo_hi_lo_lo_20};
  wire [3:0]         regroupV0_lo_hi_hi_lo_20 = {regroupV0_lo_34[867:866], regroupV0_lo_34[803:802]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_20 = {regroupV0_lo_34[995:994], regroupV0_lo_34[931:930]};
  wire [7:0]         regroupV0_lo_hi_hi_52 = {regroupV0_lo_hi_hi_hi_20, regroupV0_lo_hi_hi_lo_20};
  wire [15:0]        regroupV0_lo_hi_52 = {regroupV0_lo_hi_hi_52, regroupV0_lo_hi_lo_52};
  wire [31:0]        regroupV0_lo_52 = {regroupV0_lo_hi_52, regroupV0_lo_lo_52};
  wire [3:0]         regroupV0_hi_lo_lo_lo_20 = {regroupV0_hi_34[99:98], regroupV0_hi_34[35:34]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_20 = {regroupV0_hi_34[227:226], regroupV0_hi_34[163:162]};
  wire [7:0]         regroupV0_hi_lo_lo_52 = {regroupV0_hi_lo_lo_hi_20, regroupV0_hi_lo_lo_lo_20};
  wire [3:0]         regroupV0_hi_lo_hi_lo_20 = {regroupV0_hi_34[355:354], regroupV0_hi_34[291:290]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_20 = {regroupV0_hi_34[483:482], regroupV0_hi_34[419:418]};
  wire [7:0]         regroupV0_hi_lo_hi_52 = {regroupV0_hi_lo_hi_hi_20, regroupV0_hi_lo_hi_lo_20};
  wire [15:0]        regroupV0_hi_lo_52 = {regroupV0_hi_lo_hi_52, regroupV0_hi_lo_lo_52};
  wire [3:0]         regroupV0_hi_hi_lo_lo_20 = {regroupV0_hi_34[611:610], regroupV0_hi_34[547:546]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_20 = {regroupV0_hi_34[739:738], regroupV0_hi_34[675:674]};
  wire [7:0]         regroupV0_hi_hi_lo_52 = {regroupV0_hi_hi_lo_hi_20, regroupV0_hi_hi_lo_lo_20};
  wire [3:0]         regroupV0_hi_hi_hi_lo_20 = {regroupV0_hi_34[867:866], regroupV0_hi_34[803:802]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_20 = {regroupV0_hi_34[995:994], regroupV0_hi_34[931:930]};
  wire [7:0]         regroupV0_hi_hi_hi_52 = {regroupV0_hi_hi_hi_hi_20, regroupV0_hi_hi_hi_lo_20};
  wire [15:0]        regroupV0_hi_hi_52 = {regroupV0_hi_hi_hi_52, regroupV0_hi_hi_lo_52};
  wire [31:0]        regroupV0_hi_52 = {regroupV0_hi_hi_52, regroupV0_hi_lo_52};
  wire [3:0]         regroupV0_lo_lo_lo_lo_21 = {regroupV0_lo_34[101:100], regroupV0_lo_34[37:36]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_21 = {regroupV0_lo_34[229:228], regroupV0_lo_34[165:164]};
  wire [7:0]         regroupV0_lo_lo_lo_53 = {regroupV0_lo_lo_lo_hi_21, regroupV0_lo_lo_lo_lo_21};
  wire [3:0]         regroupV0_lo_lo_hi_lo_21 = {regroupV0_lo_34[357:356], regroupV0_lo_34[293:292]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_21 = {regroupV0_lo_34[485:484], regroupV0_lo_34[421:420]};
  wire [7:0]         regroupV0_lo_lo_hi_53 = {regroupV0_lo_lo_hi_hi_21, regroupV0_lo_lo_hi_lo_21};
  wire [15:0]        regroupV0_lo_lo_53 = {regroupV0_lo_lo_hi_53, regroupV0_lo_lo_lo_53};
  wire [3:0]         regroupV0_lo_hi_lo_lo_21 = {regroupV0_lo_34[613:612], regroupV0_lo_34[549:548]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_21 = {regroupV0_lo_34[741:740], regroupV0_lo_34[677:676]};
  wire [7:0]         regroupV0_lo_hi_lo_53 = {regroupV0_lo_hi_lo_hi_21, regroupV0_lo_hi_lo_lo_21};
  wire [3:0]         regroupV0_lo_hi_hi_lo_21 = {regroupV0_lo_34[869:868], regroupV0_lo_34[805:804]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_21 = {regroupV0_lo_34[997:996], regroupV0_lo_34[933:932]};
  wire [7:0]         regroupV0_lo_hi_hi_53 = {regroupV0_lo_hi_hi_hi_21, regroupV0_lo_hi_hi_lo_21};
  wire [15:0]        regroupV0_lo_hi_53 = {regroupV0_lo_hi_hi_53, regroupV0_lo_hi_lo_53};
  wire [31:0]        regroupV0_lo_53 = {regroupV0_lo_hi_53, regroupV0_lo_lo_53};
  wire [3:0]         regroupV0_hi_lo_lo_lo_21 = {regroupV0_hi_34[101:100], regroupV0_hi_34[37:36]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_21 = {regroupV0_hi_34[229:228], regroupV0_hi_34[165:164]};
  wire [7:0]         regroupV0_hi_lo_lo_53 = {regroupV0_hi_lo_lo_hi_21, regroupV0_hi_lo_lo_lo_21};
  wire [3:0]         regroupV0_hi_lo_hi_lo_21 = {regroupV0_hi_34[357:356], regroupV0_hi_34[293:292]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_21 = {regroupV0_hi_34[485:484], regroupV0_hi_34[421:420]};
  wire [7:0]         regroupV0_hi_lo_hi_53 = {regroupV0_hi_lo_hi_hi_21, regroupV0_hi_lo_hi_lo_21};
  wire [15:0]        regroupV0_hi_lo_53 = {regroupV0_hi_lo_hi_53, regroupV0_hi_lo_lo_53};
  wire [3:0]         regroupV0_hi_hi_lo_lo_21 = {regroupV0_hi_34[613:612], regroupV0_hi_34[549:548]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_21 = {regroupV0_hi_34[741:740], regroupV0_hi_34[677:676]};
  wire [7:0]         regroupV0_hi_hi_lo_53 = {regroupV0_hi_hi_lo_hi_21, regroupV0_hi_hi_lo_lo_21};
  wire [3:0]         regroupV0_hi_hi_hi_lo_21 = {regroupV0_hi_34[869:868], regroupV0_hi_34[805:804]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_21 = {regroupV0_hi_34[997:996], regroupV0_hi_34[933:932]};
  wire [7:0]         regroupV0_hi_hi_hi_53 = {regroupV0_hi_hi_hi_hi_21, regroupV0_hi_hi_hi_lo_21};
  wire [15:0]        regroupV0_hi_hi_53 = {regroupV0_hi_hi_hi_53, regroupV0_hi_hi_lo_53};
  wire [31:0]        regroupV0_hi_53 = {regroupV0_hi_hi_53, regroupV0_hi_lo_53};
  wire [3:0]         regroupV0_lo_lo_lo_lo_22 = {regroupV0_lo_34[103:102], regroupV0_lo_34[39:38]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_22 = {regroupV0_lo_34[231:230], regroupV0_lo_34[167:166]};
  wire [7:0]         regroupV0_lo_lo_lo_54 = {regroupV0_lo_lo_lo_hi_22, regroupV0_lo_lo_lo_lo_22};
  wire [3:0]         regroupV0_lo_lo_hi_lo_22 = {regroupV0_lo_34[359:358], regroupV0_lo_34[295:294]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_22 = {regroupV0_lo_34[487:486], regroupV0_lo_34[423:422]};
  wire [7:0]         regroupV0_lo_lo_hi_54 = {regroupV0_lo_lo_hi_hi_22, regroupV0_lo_lo_hi_lo_22};
  wire [15:0]        regroupV0_lo_lo_54 = {regroupV0_lo_lo_hi_54, regroupV0_lo_lo_lo_54};
  wire [3:0]         regroupV0_lo_hi_lo_lo_22 = {regroupV0_lo_34[615:614], regroupV0_lo_34[551:550]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_22 = {regroupV0_lo_34[743:742], regroupV0_lo_34[679:678]};
  wire [7:0]         regroupV0_lo_hi_lo_54 = {regroupV0_lo_hi_lo_hi_22, regroupV0_lo_hi_lo_lo_22};
  wire [3:0]         regroupV0_lo_hi_hi_lo_22 = {regroupV0_lo_34[871:870], regroupV0_lo_34[807:806]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_22 = {regroupV0_lo_34[999:998], regroupV0_lo_34[935:934]};
  wire [7:0]         regroupV0_lo_hi_hi_54 = {regroupV0_lo_hi_hi_hi_22, regroupV0_lo_hi_hi_lo_22};
  wire [15:0]        regroupV0_lo_hi_54 = {regroupV0_lo_hi_hi_54, regroupV0_lo_hi_lo_54};
  wire [31:0]        regroupV0_lo_54 = {regroupV0_lo_hi_54, regroupV0_lo_lo_54};
  wire [3:0]         regroupV0_hi_lo_lo_lo_22 = {regroupV0_hi_34[103:102], regroupV0_hi_34[39:38]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_22 = {regroupV0_hi_34[231:230], regroupV0_hi_34[167:166]};
  wire [7:0]         regroupV0_hi_lo_lo_54 = {regroupV0_hi_lo_lo_hi_22, regroupV0_hi_lo_lo_lo_22};
  wire [3:0]         regroupV0_hi_lo_hi_lo_22 = {regroupV0_hi_34[359:358], regroupV0_hi_34[295:294]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_22 = {regroupV0_hi_34[487:486], regroupV0_hi_34[423:422]};
  wire [7:0]         regroupV0_hi_lo_hi_54 = {regroupV0_hi_lo_hi_hi_22, regroupV0_hi_lo_hi_lo_22};
  wire [15:0]        regroupV0_hi_lo_54 = {regroupV0_hi_lo_hi_54, regroupV0_hi_lo_lo_54};
  wire [3:0]         regroupV0_hi_hi_lo_lo_22 = {regroupV0_hi_34[615:614], regroupV0_hi_34[551:550]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_22 = {regroupV0_hi_34[743:742], regroupV0_hi_34[679:678]};
  wire [7:0]         regroupV0_hi_hi_lo_54 = {regroupV0_hi_hi_lo_hi_22, regroupV0_hi_hi_lo_lo_22};
  wire [3:0]         regroupV0_hi_hi_hi_lo_22 = {regroupV0_hi_34[871:870], regroupV0_hi_34[807:806]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_22 = {regroupV0_hi_34[999:998], regroupV0_hi_34[935:934]};
  wire [7:0]         regroupV0_hi_hi_hi_54 = {regroupV0_hi_hi_hi_hi_22, regroupV0_hi_hi_hi_lo_22};
  wire [15:0]        regroupV0_hi_hi_54 = {regroupV0_hi_hi_hi_54, regroupV0_hi_hi_lo_54};
  wire [31:0]        regroupV0_hi_54 = {regroupV0_hi_hi_54, regroupV0_hi_lo_54};
  wire [3:0]         regroupV0_lo_lo_lo_lo_23 = {regroupV0_lo_34[105:104], regroupV0_lo_34[41:40]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_23 = {regroupV0_lo_34[233:232], regroupV0_lo_34[169:168]};
  wire [7:0]         regroupV0_lo_lo_lo_55 = {regroupV0_lo_lo_lo_hi_23, regroupV0_lo_lo_lo_lo_23};
  wire [3:0]         regroupV0_lo_lo_hi_lo_23 = {regroupV0_lo_34[361:360], regroupV0_lo_34[297:296]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_23 = {regroupV0_lo_34[489:488], regroupV0_lo_34[425:424]};
  wire [7:0]         regroupV0_lo_lo_hi_55 = {regroupV0_lo_lo_hi_hi_23, regroupV0_lo_lo_hi_lo_23};
  wire [15:0]        regroupV0_lo_lo_55 = {regroupV0_lo_lo_hi_55, regroupV0_lo_lo_lo_55};
  wire [3:0]         regroupV0_lo_hi_lo_lo_23 = {regroupV0_lo_34[617:616], regroupV0_lo_34[553:552]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_23 = {regroupV0_lo_34[745:744], regroupV0_lo_34[681:680]};
  wire [7:0]         regroupV0_lo_hi_lo_55 = {regroupV0_lo_hi_lo_hi_23, regroupV0_lo_hi_lo_lo_23};
  wire [3:0]         regroupV0_lo_hi_hi_lo_23 = {regroupV0_lo_34[873:872], regroupV0_lo_34[809:808]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_23 = {regroupV0_lo_34[1001:1000], regroupV0_lo_34[937:936]};
  wire [7:0]         regroupV0_lo_hi_hi_55 = {regroupV0_lo_hi_hi_hi_23, regroupV0_lo_hi_hi_lo_23};
  wire [15:0]        regroupV0_lo_hi_55 = {regroupV0_lo_hi_hi_55, regroupV0_lo_hi_lo_55};
  wire [31:0]        regroupV0_lo_55 = {regroupV0_lo_hi_55, regroupV0_lo_lo_55};
  wire [3:0]         regroupV0_hi_lo_lo_lo_23 = {regroupV0_hi_34[105:104], regroupV0_hi_34[41:40]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_23 = {regroupV0_hi_34[233:232], regroupV0_hi_34[169:168]};
  wire [7:0]         regroupV0_hi_lo_lo_55 = {regroupV0_hi_lo_lo_hi_23, regroupV0_hi_lo_lo_lo_23};
  wire [3:0]         regroupV0_hi_lo_hi_lo_23 = {regroupV0_hi_34[361:360], regroupV0_hi_34[297:296]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_23 = {regroupV0_hi_34[489:488], regroupV0_hi_34[425:424]};
  wire [7:0]         regroupV0_hi_lo_hi_55 = {regroupV0_hi_lo_hi_hi_23, regroupV0_hi_lo_hi_lo_23};
  wire [15:0]        regroupV0_hi_lo_55 = {regroupV0_hi_lo_hi_55, regroupV0_hi_lo_lo_55};
  wire [3:0]         regroupV0_hi_hi_lo_lo_23 = {regroupV0_hi_34[617:616], regroupV0_hi_34[553:552]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_23 = {regroupV0_hi_34[745:744], regroupV0_hi_34[681:680]};
  wire [7:0]         regroupV0_hi_hi_lo_55 = {regroupV0_hi_hi_lo_hi_23, regroupV0_hi_hi_lo_lo_23};
  wire [3:0]         regroupV0_hi_hi_hi_lo_23 = {regroupV0_hi_34[873:872], regroupV0_hi_34[809:808]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_23 = {regroupV0_hi_34[1001:1000], regroupV0_hi_34[937:936]};
  wire [7:0]         regroupV0_hi_hi_hi_55 = {regroupV0_hi_hi_hi_hi_23, regroupV0_hi_hi_hi_lo_23};
  wire [15:0]        regroupV0_hi_hi_55 = {regroupV0_hi_hi_hi_55, regroupV0_hi_hi_lo_55};
  wire [31:0]        regroupV0_hi_55 = {regroupV0_hi_hi_55, regroupV0_hi_lo_55};
  wire [3:0]         regroupV0_lo_lo_lo_lo_24 = {regroupV0_lo_34[107:106], regroupV0_lo_34[43:42]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_24 = {regroupV0_lo_34[235:234], regroupV0_lo_34[171:170]};
  wire [7:0]         regroupV0_lo_lo_lo_56 = {regroupV0_lo_lo_lo_hi_24, regroupV0_lo_lo_lo_lo_24};
  wire [3:0]         regroupV0_lo_lo_hi_lo_24 = {regroupV0_lo_34[363:362], regroupV0_lo_34[299:298]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_24 = {regroupV0_lo_34[491:490], regroupV0_lo_34[427:426]};
  wire [7:0]         regroupV0_lo_lo_hi_56 = {regroupV0_lo_lo_hi_hi_24, regroupV0_lo_lo_hi_lo_24};
  wire [15:0]        regroupV0_lo_lo_56 = {regroupV0_lo_lo_hi_56, regroupV0_lo_lo_lo_56};
  wire [3:0]         regroupV0_lo_hi_lo_lo_24 = {regroupV0_lo_34[619:618], regroupV0_lo_34[555:554]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_24 = {regroupV0_lo_34[747:746], regroupV0_lo_34[683:682]};
  wire [7:0]         regroupV0_lo_hi_lo_56 = {regroupV0_lo_hi_lo_hi_24, regroupV0_lo_hi_lo_lo_24};
  wire [3:0]         regroupV0_lo_hi_hi_lo_24 = {regroupV0_lo_34[875:874], regroupV0_lo_34[811:810]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_24 = {regroupV0_lo_34[1003:1002], regroupV0_lo_34[939:938]};
  wire [7:0]         regroupV0_lo_hi_hi_56 = {regroupV0_lo_hi_hi_hi_24, regroupV0_lo_hi_hi_lo_24};
  wire [15:0]        regroupV0_lo_hi_56 = {regroupV0_lo_hi_hi_56, regroupV0_lo_hi_lo_56};
  wire [31:0]        regroupV0_lo_56 = {regroupV0_lo_hi_56, regroupV0_lo_lo_56};
  wire [3:0]         regroupV0_hi_lo_lo_lo_24 = {regroupV0_hi_34[107:106], regroupV0_hi_34[43:42]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_24 = {regroupV0_hi_34[235:234], regroupV0_hi_34[171:170]};
  wire [7:0]         regroupV0_hi_lo_lo_56 = {regroupV0_hi_lo_lo_hi_24, regroupV0_hi_lo_lo_lo_24};
  wire [3:0]         regroupV0_hi_lo_hi_lo_24 = {regroupV0_hi_34[363:362], regroupV0_hi_34[299:298]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_24 = {regroupV0_hi_34[491:490], regroupV0_hi_34[427:426]};
  wire [7:0]         regroupV0_hi_lo_hi_56 = {regroupV0_hi_lo_hi_hi_24, regroupV0_hi_lo_hi_lo_24};
  wire [15:0]        regroupV0_hi_lo_56 = {regroupV0_hi_lo_hi_56, regroupV0_hi_lo_lo_56};
  wire [3:0]         regroupV0_hi_hi_lo_lo_24 = {regroupV0_hi_34[619:618], regroupV0_hi_34[555:554]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_24 = {regroupV0_hi_34[747:746], regroupV0_hi_34[683:682]};
  wire [7:0]         regroupV0_hi_hi_lo_56 = {regroupV0_hi_hi_lo_hi_24, regroupV0_hi_hi_lo_lo_24};
  wire [3:0]         regroupV0_hi_hi_hi_lo_24 = {regroupV0_hi_34[875:874], regroupV0_hi_34[811:810]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_24 = {regroupV0_hi_34[1003:1002], regroupV0_hi_34[939:938]};
  wire [7:0]         regroupV0_hi_hi_hi_56 = {regroupV0_hi_hi_hi_hi_24, regroupV0_hi_hi_hi_lo_24};
  wire [15:0]        regroupV0_hi_hi_56 = {regroupV0_hi_hi_hi_56, regroupV0_hi_hi_lo_56};
  wire [31:0]        regroupV0_hi_56 = {regroupV0_hi_hi_56, regroupV0_hi_lo_56};
  wire [3:0]         regroupV0_lo_lo_lo_lo_25 = {regroupV0_lo_34[109:108], regroupV0_lo_34[45:44]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_25 = {regroupV0_lo_34[237:236], regroupV0_lo_34[173:172]};
  wire [7:0]         regroupV0_lo_lo_lo_57 = {regroupV0_lo_lo_lo_hi_25, regroupV0_lo_lo_lo_lo_25};
  wire [3:0]         regroupV0_lo_lo_hi_lo_25 = {regroupV0_lo_34[365:364], regroupV0_lo_34[301:300]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_25 = {regroupV0_lo_34[493:492], regroupV0_lo_34[429:428]};
  wire [7:0]         regroupV0_lo_lo_hi_57 = {regroupV0_lo_lo_hi_hi_25, regroupV0_lo_lo_hi_lo_25};
  wire [15:0]        regroupV0_lo_lo_57 = {regroupV0_lo_lo_hi_57, regroupV0_lo_lo_lo_57};
  wire [3:0]         regroupV0_lo_hi_lo_lo_25 = {regroupV0_lo_34[621:620], regroupV0_lo_34[557:556]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_25 = {regroupV0_lo_34[749:748], regroupV0_lo_34[685:684]};
  wire [7:0]         regroupV0_lo_hi_lo_57 = {regroupV0_lo_hi_lo_hi_25, regroupV0_lo_hi_lo_lo_25};
  wire [3:0]         regroupV0_lo_hi_hi_lo_25 = {regroupV0_lo_34[877:876], regroupV0_lo_34[813:812]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_25 = {regroupV0_lo_34[1005:1004], regroupV0_lo_34[941:940]};
  wire [7:0]         regroupV0_lo_hi_hi_57 = {regroupV0_lo_hi_hi_hi_25, regroupV0_lo_hi_hi_lo_25};
  wire [15:0]        regroupV0_lo_hi_57 = {regroupV0_lo_hi_hi_57, regroupV0_lo_hi_lo_57};
  wire [31:0]        regroupV0_lo_57 = {regroupV0_lo_hi_57, regroupV0_lo_lo_57};
  wire [3:0]         regroupV0_hi_lo_lo_lo_25 = {regroupV0_hi_34[109:108], regroupV0_hi_34[45:44]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_25 = {regroupV0_hi_34[237:236], regroupV0_hi_34[173:172]};
  wire [7:0]         regroupV0_hi_lo_lo_57 = {regroupV0_hi_lo_lo_hi_25, regroupV0_hi_lo_lo_lo_25};
  wire [3:0]         regroupV0_hi_lo_hi_lo_25 = {regroupV0_hi_34[365:364], regroupV0_hi_34[301:300]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_25 = {regroupV0_hi_34[493:492], regroupV0_hi_34[429:428]};
  wire [7:0]         regroupV0_hi_lo_hi_57 = {regroupV0_hi_lo_hi_hi_25, regroupV0_hi_lo_hi_lo_25};
  wire [15:0]        regroupV0_hi_lo_57 = {regroupV0_hi_lo_hi_57, regroupV0_hi_lo_lo_57};
  wire [3:0]         regroupV0_hi_hi_lo_lo_25 = {regroupV0_hi_34[621:620], regroupV0_hi_34[557:556]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_25 = {regroupV0_hi_34[749:748], regroupV0_hi_34[685:684]};
  wire [7:0]         regroupV0_hi_hi_lo_57 = {regroupV0_hi_hi_lo_hi_25, regroupV0_hi_hi_lo_lo_25};
  wire [3:0]         regroupV0_hi_hi_hi_lo_25 = {regroupV0_hi_34[877:876], regroupV0_hi_34[813:812]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_25 = {regroupV0_hi_34[1005:1004], regroupV0_hi_34[941:940]};
  wire [7:0]         regroupV0_hi_hi_hi_57 = {regroupV0_hi_hi_hi_hi_25, regroupV0_hi_hi_hi_lo_25};
  wire [15:0]        regroupV0_hi_hi_57 = {regroupV0_hi_hi_hi_57, regroupV0_hi_hi_lo_57};
  wire [31:0]        regroupV0_hi_57 = {regroupV0_hi_hi_57, regroupV0_hi_lo_57};
  wire [3:0]         regroupV0_lo_lo_lo_lo_26 = {regroupV0_lo_34[111:110], regroupV0_lo_34[47:46]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_26 = {regroupV0_lo_34[239:238], regroupV0_lo_34[175:174]};
  wire [7:0]         regroupV0_lo_lo_lo_58 = {regroupV0_lo_lo_lo_hi_26, regroupV0_lo_lo_lo_lo_26};
  wire [3:0]         regroupV0_lo_lo_hi_lo_26 = {regroupV0_lo_34[367:366], regroupV0_lo_34[303:302]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_26 = {regroupV0_lo_34[495:494], regroupV0_lo_34[431:430]};
  wire [7:0]         regroupV0_lo_lo_hi_58 = {regroupV0_lo_lo_hi_hi_26, regroupV0_lo_lo_hi_lo_26};
  wire [15:0]        regroupV0_lo_lo_58 = {regroupV0_lo_lo_hi_58, regroupV0_lo_lo_lo_58};
  wire [3:0]         regroupV0_lo_hi_lo_lo_26 = {regroupV0_lo_34[623:622], regroupV0_lo_34[559:558]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_26 = {regroupV0_lo_34[751:750], regroupV0_lo_34[687:686]};
  wire [7:0]         regroupV0_lo_hi_lo_58 = {regroupV0_lo_hi_lo_hi_26, regroupV0_lo_hi_lo_lo_26};
  wire [3:0]         regroupV0_lo_hi_hi_lo_26 = {regroupV0_lo_34[879:878], regroupV0_lo_34[815:814]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_26 = {regroupV0_lo_34[1007:1006], regroupV0_lo_34[943:942]};
  wire [7:0]         regroupV0_lo_hi_hi_58 = {regroupV0_lo_hi_hi_hi_26, regroupV0_lo_hi_hi_lo_26};
  wire [15:0]        regroupV0_lo_hi_58 = {regroupV0_lo_hi_hi_58, regroupV0_lo_hi_lo_58};
  wire [31:0]        regroupV0_lo_58 = {regroupV0_lo_hi_58, regroupV0_lo_lo_58};
  wire [3:0]         regroupV0_hi_lo_lo_lo_26 = {regroupV0_hi_34[111:110], regroupV0_hi_34[47:46]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_26 = {regroupV0_hi_34[239:238], regroupV0_hi_34[175:174]};
  wire [7:0]         regroupV0_hi_lo_lo_58 = {regroupV0_hi_lo_lo_hi_26, regroupV0_hi_lo_lo_lo_26};
  wire [3:0]         regroupV0_hi_lo_hi_lo_26 = {regroupV0_hi_34[367:366], regroupV0_hi_34[303:302]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_26 = {regroupV0_hi_34[495:494], regroupV0_hi_34[431:430]};
  wire [7:0]         regroupV0_hi_lo_hi_58 = {regroupV0_hi_lo_hi_hi_26, regroupV0_hi_lo_hi_lo_26};
  wire [15:0]        regroupV0_hi_lo_58 = {regroupV0_hi_lo_hi_58, regroupV0_hi_lo_lo_58};
  wire [3:0]         regroupV0_hi_hi_lo_lo_26 = {regroupV0_hi_34[623:622], regroupV0_hi_34[559:558]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_26 = {regroupV0_hi_34[751:750], regroupV0_hi_34[687:686]};
  wire [7:0]         regroupV0_hi_hi_lo_58 = {regroupV0_hi_hi_lo_hi_26, regroupV0_hi_hi_lo_lo_26};
  wire [3:0]         regroupV0_hi_hi_hi_lo_26 = {regroupV0_hi_34[879:878], regroupV0_hi_34[815:814]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_26 = {regroupV0_hi_34[1007:1006], regroupV0_hi_34[943:942]};
  wire [7:0]         regroupV0_hi_hi_hi_58 = {regroupV0_hi_hi_hi_hi_26, regroupV0_hi_hi_hi_lo_26};
  wire [15:0]        regroupV0_hi_hi_58 = {regroupV0_hi_hi_hi_58, regroupV0_hi_hi_lo_58};
  wire [31:0]        regroupV0_hi_58 = {regroupV0_hi_hi_58, regroupV0_hi_lo_58};
  wire [3:0]         regroupV0_lo_lo_lo_lo_27 = {regroupV0_lo_34[113:112], regroupV0_lo_34[49:48]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_27 = {regroupV0_lo_34[241:240], regroupV0_lo_34[177:176]};
  wire [7:0]         regroupV0_lo_lo_lo_59 = {regroupV0_lo_lo_lo_hi_27, regroupV0_lo_lo_lo_lo_27};
  wire [3:0]         regroupV0_lo_lo_hi_lo_27 = {regroupV0_lo_34[369:368], regroupV0_lo_34[305:304]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_27 = {regroupV0_lo_34[497:496], regroupV0_lo_34[433:432]};
  wire [7:0]         regroupV0_lo_lo_hi_59 = {regroupV0_lo_lo_hi_hi_27, regroupV0_lo_lo_hi_lo_27};
  wire [15:0]        regroupV0_lo_lo_59 = {regroupV0_lo_lo_hi_59, regroupV0_lo_lo_lo_59};
  wire [3:0]         regroupV0_lo_hi_lo_lo_27 = {regroupV0_lo_34[625:624], regroupV0_lo_34[561:560]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_27 = {regroupV0_lo_34[753:752], regroupV0_lo_34[689:688]};
  wire [7:0]         regroupV0_lo_hi_lo_59 = {regroupV0_lo_hi_lo_hi_27, regroupV0_lo_hi_lo_lo_27};
  wire [3:0]         regroupV0_lo_hi_hi_lo_27 = {regroupV0_lo_34[881:880], regroupV0_lo_34[817:816]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_27 = {regroupV0_lo_34[1009:1008], regroupV0_lo_34[945:944]};
  wire [7:0]         regroupV0_lo_hi_hi_59 = {regroupV0_lo_hi_hi_hi_27, regroupV0_lo_hi_hi_lo_27};
  wire [15:0]        regroupV0_lo_hi_59 = {regroupV0_lo_hi_hi_59, regroupV0_lo_hi_lo_59};
  wire [31:0]        regroupV0_lo_59 = {regroupV0_lo_hi_59, regroupV0_lo_lo_59};
  wire [3:0]         regroupV0_hi_lo_lo_lo_27 = {regroupV0_hi_34[113:112], regroupV0_hi_34[49:48]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_27 = {regroupV0_hi_34[241:240], regroupV0_hi_34[177:176]};
  wire [7:0]         regroupV0_hi_lo_lo_59 = {regroupV0_hi_lo_lo_hi_27, regroupV0_hi_lo_lo_lo_27};
  wire [3:0]         regroupV0_hi_lo_hi_lo_27 = {regroupV0_hi_34[369:368], regroupV0_hi_34[305:304]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_27 = {regroupV0_hi_34[497:496], regroupV0_hi_34[433:432]};
  wire [7:0]         regroupV0_hi_lo_hi_59 = {regroupV0_hi_lo_hi_hi_27, regroupV0_hi_lo_hi_lo_27};
  wire [15:0]        regroupV0_hi_lo_59 = {regroupV0_hi_lo_hi_59, regroupV0_hi_lo_lo_59};
  wire [3:0]         regroupV0_hi_hi_lo_lo_27 = {regroupV0_hi_34[625:624], regroupV0_hi_34[561:560]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_27 = {regroupV0_hi_34[753:752], regroupV0_hi_34[689:688]};
  wire [7:0]         regroupV0_hi_hi_lo_59 = {regroupV0_hi_hi_lo_hi_27, regroupV0_hi_hi_lo_lo_27};
  wire [3:0]         regroupV0_hi_hi_hi_lo_27 = {regroupV0_hi_34[881:880], regroupV0_hi_34[817:816]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_27 = {regroupV0_hi_34[1009:1008], regroupV0_hi_34[945:944]};
  wire [7:0]         regroupV0_hi_hi_hi_59 = {regroupV0_hi_hi_hi_hi_27, regroupV0_hi_hi_hi_lo_27};
  wire [15:0]        regroupV0_hi_hi_59 = {regroupV0_hi_hi_hi_59, regroupV0_hi_hi_lo_59};
  wire [31:0]        regroupV0_hi_59 = {regroupV0_hi_hi_59, regroupV0_hi_lo_59};
  wire [3:0]         regroupV0_lo_lo_lo_lo_28 = {regroupV0_lo_34[115:114], regroupV0_lo_34[51:50]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_28 = {regroupV0_lo_34[243:242], regroupV0_lo_34[179:178]};
  wire [7:0]         regroupV0_lo_lo_lo_60 = {regroupV0_lo_lo_lo_hi_28, regroupV0_lo_lo_lo_lo_28};
  wire [3:0]         regroupV0_lo_lo_hi_lo_28 = {regroupV0_lo_34[371:370], regroupV0_lo_34[307:306]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_28 = {regroupV0_lo_34[499:498], regroupV0_lo_34[435:434]};
  wire [7:0]         regroupV0_lo_lo_hi_60 = {regroupV0_lo_lo_hi_hi_28, regroupV0_lo_lo_hi_lo_28};
  wire [15:0]        regroupV0_lo_lo_60 = {regroupV0_lo_lo_hi_60, regroupV0_lo_lo_lo_60};
  wire [3:0]         regroupV0_lo_hi_lo_lo_28 = {regroupV0_lo_34[627:626], regroupV0_lo_34[563:562]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_28 = {regroupV0_lo_34[755:754], regroupV0_lo_34[691:690]};
  wire [7:0]         regroupV0_lo_hi_lo_60 = {regroupV0_lo_hi_lo_hi_28, regroupV0_lo_hi_lo_lo_28};
  wire [3:0]         regroupV0_lo_hi_hi_lo_28 = {regroupV0_lo_34[883:882], regroupV0_lo_34[819:818]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_28 = {regroupV0_lo_34[1011:1010], regroupV0_lo_34[947:946]};
  wire [7:0]         regroupV0_lo_hi_hi_60 = {regroupV0_lo_hi_hi_hi_28, regroupV0_lo_hi_hi_lo_28};
  wire [15:0]        regroupV0_lo_hi_60 = {regroupV0_lo_hi_hi_60, regroupV0_lo_hi_lo_60};
  wire [31:0]        regroupV0_lo_60 = {regroupV0_lo_hi_60, regroupV0_lo_lo_60};
  wire [3:0]         regroupV0_hi_lo_lo_lo_28 = {regroupV0_hi_34[115:114], regroupV0_hi_34[51:50]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_28 = {regroupV0_hi_34[243:242], regroupV0_hi_34[179:178]};
  wire [7:0]         regroupV0_hi_lo_lo_60 = {regroupV0_hi_lo_lo_hi_28, regroupV0_hi_lo_lo_lo_28};
  wire [3:0]         regroupV0_hi_lo_hi_lo_28 = {regroupV0_hi_34[371:370], regroupV0_hi_34[307:306]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_28 = {regroupV0_hi_34[499:498], regroupV0_hi_34[435:434]};
  wire [7:0]         regroupV0_hi_lo_hi_60 = {regroupV0_hi_lo_hi_hi_28, regroupV0_hi_lo_hi_lo_28};
  wire [15:0]        regroupV0_hi_lo_60 = {regroupV0_hi_lo_hi_60, regroupV0_hi_lo_lo_60};
  wire [3:0]         regroupV0_hi_hi_lo_lo_28 = {regroupV0_hi_34[627:626], regroupV0_hi_34[563:562]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_28 = {regroupV0_hi_34[755:754], regroupV0_hi_34[691:690]};
  wire [7:0]         regroupV0_hi_hi_lo_60 = {regroupV0_hi_hi_lo_hi_28, regroupV0_hi_hi_lo_lo_28};
  wire [3:0]         regroupV0_hi_hi_hi_lo_28 = {regroupV0_hi_34[883:882], regroupV0_hi_34[819:818]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_28 = {regroupV0_hi_34[1011:1010], regroupV0_hi_34[947:946]};
  wire [7:0]         regroupV0_hi_hi_hi_60 = {regroupV0_hi_hi_hi_hi_28, regroupV0_hi_hi_hi_lo_28};
  wire [15:0]        regroupV0_hi_hi_60 = {regroupV0_hi_hi_hi_60, regroupV0_hi_hi_lo_60};
  wire [31:0]        regroupV0_hi_60 = {regroupV0_hi_hi_60, regroupV0_hi_lo_60};
  wire [3:0]         regroupV0_lo_lo_lo_lo_29 = {regroupV0_lo_34[117:116], regroupV0_lo_34[53:52]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_29 = {regroupV0_lo_34[245:244], regroupV0_lo_34[181:180]};
  wire [7:0]         regroupV0_lo_lo_lo_61 = {regroupV0_lo_lo_lo_hi_29, regroupV0_lo_lo_lo_lo_29};
  wire [3:0]         regroupV0_lo_lo_hi_lo_29 = {regroupV0_lo_34[373:372], regroupV0_lo_34[309:308]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_29 = {regroupV0_lo_34[501:500], regroupV0_lo_34[437:436]};
  wire [7:0]         regroupV0_lo_lo_hi_61 = {regroupV0_lo_lo_hi_hi_29, regroupV0_lo_lo_hi_lo_29};
  wire [15:0]        regroupV0_lo_lo_61 = {regroupV0_lo_lo_hi_61, regroupV0_lo_lo_lo_61};
  wire [3:0]         regroupV0_lo_hi_lo_lo_29 = {regroupV0_lo_34[629:628], regroupV0_lo_34[565:564]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_29 = {regroupV0_lo_34[757:756], regroupV0_lo_34[693:692]};
  wire [7:0]         regroupV0_lo_hi_lo_61 = {regroupV0_lo_hi_lo_hi_29, regroupV0_lo_hi_lo_lo_29};
  wire [3:0]         regroupV0_lo_hi_hi_lo_29 = {regroupV0_lo_34[885:884], regroupV0_lo_34[821:820]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_29 = {regroupV0_lo_34[1013:1012], regroupV0_lo_34[949:948]};
  wire [7:0]         regroupV0_lo_hi_hi_61 = {regroupV0_lo_hi_hi_hi_29, regroupV0_lo_hi_hi_lo_29};
  wire [15:0]        regroupV0_lo_hi_61 = {regroupV0_lo_hi_hi_61, regroupV0_lo_hi_lo_61};
  wire [31:0]        regroupV0_lo_61 = {regroupV0_lo_hi_61, regroupV0_lo_lo_61};
  wire [3:0]         regroupV0_hi_lo_lo_lo_29 = {regroupV0_hi_34[117:116], regroupV0_hi_34[53:52]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_29 = {regroupV0_hi_34[245:244], regroupV0_hi_34[181:180]};
  wire [7:0]         regroupV0_hi_lo_lo_61 = {regroupV0_hi_lo_lo_hi_29, regroupV0_hi_lo_lo_lo_29};
  wire [3:0]         regroupV0_hi_lo_hi_lo_29 = {regroupV0_hi_34[373:372], regroupV0_hi_34[309:308]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_29 = {regroupV0_hi_34[501:500], regroupV0_hi_34[437:436]};
  wire [7:0]         regroupV0_hi_lo_hi_61 = {regroupV0_hi_lo_hi_hi_29, regroupV0_hi_lo_hi_lo_29};
  wire [15:0]        regroupV0_hi_lo_61 = {regroupV0_hi_lo_hi_61, regroupV0_hi_lo_lo_61};
  wire [3:0]         regroupV0_hi_hi_lo_lo_29 = {regroupV0_hi_34[629:628], regroupV0_hi_34[565:564]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_29 = {regroupV0_hi_34[757:756], regroupV0_hi_34[693:692]};
  wire [7:0]         regroupV0_hi_hi_lo_61 = {regroupV0_hi_hi_lo_hi_29, regroupV0_hi_hi_lo_lo_29};
  wire [3:0]         regroupV0_hi_hi_hi_lo_29 = {regroupV0_hi_34[885:884], regroupV0_hi_34[821:820]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_29 = {regroupV0_hi_34[1013:1012], regroupV0_hi_34[949:948]};
  wire [7:0]         regroupV0_hi_hi_hi_61 = {regroupV0_hi_hi_hi_hi_29, regroupV0_hi_hi_hi_lo_29};
  wire [15:0]        regroupV0_hi_hi_61 = {regroupV0_hi_hi_hi_61, regroupV0_hi_hi_lo_61};
  wire [31:0]        regroupV0_hi_61 = {regroupV0_hi_hi_61, regroupV0_hi_lo_61};
  wire [3:0]         regroupV0_lo_lo_lo_lo_30 = {regroupV0_lo_34[119:118], regroupV0_lo_34[55:54]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_30 = {regroupV0_lo_34[247:246], regroupV0_lo_34[183:182]};
  wire [7:0]         regroupV0_lo_lo_lo_62 = {regroupV0_lo_lo_lo_hi_30, regroupV0_lo_lo_lo_lo_30};
  wire [3:0]         regroupV0_lo_lo_hi_lo_30 = {regroupV0_lo_34[375:374], regroupV0_lo_34[311:310]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_30 = {regroupV0_lo_34[503:502], regroupV0_lo_34[439:438]};
  wire [7:0]         regroupV0_lo_lo_hi_62 = {regroupV0_lo_lo_hi_hi_30, regroupV0_lo_lo_hi_lo_30};
  wire [15:0]        regroupV0_lo_lo_62 = {regroupV0_lo_lo_hi_62, regroupV0_lo_lo_lo_62};
  wire [3:0]         regroupV0_lo_hi_lo_lo_30 = {regroupV0_lo_34[631:630], regroupV0_lo_34[567:566]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_30 = {regroupV0_lo_34[759:758], regroupV0_lo_34[695:694]};
  wire [7:0]         regroupV0_lo_hi_lo_62 = {regroupV0_lo_hi_lo_hi_30, regroupV0_lo_hi_lo_lo_30};
  wire [3:0]         regroupV0_lo_hi_hi_lo_30 = {regroupV0_lo_34[887:886], regroupV0_lo_34[823:822]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_30 = {regroupV0_lo_34[1015:1014], regroupV0_lo_34[951:950]};
  wire [7:0]         regroupV0_lo_hi_hi_62 = {regroupV0_lo_hi_hi_hi_30, regroupV0_lo_hi_hi_lo_30};
  wire [15:0]        regroupV0_lo_hi_62 = {regroupV0_lo_hi_hi_62, regroupV0_lo_hi_lo_62};
  wire [31:0]        regroupV0_lo_62 = {regroupV0_lo_hi_62, regroupV0_lo_lo_62};
  wire [3:0]         regroupV0_hi_lo_lo_lo_30 = {regroupV0_hi_34[119:118], regroupV0_hi_34[55:54]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_30 = {regroupV0_hi_34[247:246], regroupV0_hi_34[183:182]};
  wire [7:0]         regroupV0_hi_lo_lo_62 = {regroupV0_hi_lo_lo_hi_30, regroupV0_hi_lo_lo_lo_30};
  wire [3:0]         regroupV0_hi_lo_hi_lo_30 = {regroupV0_hi_34[375:374], regroupV0_hi_34[311:310]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_30 = {regroupV0_hi_34[503:502], regroupV0_hi_34[439:438]};
  wire [7:0]         regroupV0_hi_lo_hi_62 = {regroupV0_hi_lo_hi_hi_30, regroupV0_hi_lo_hi_lo_30};
  wire [15:0]        regroupV0_hi_lo_62 = {regroupV0_hi_lo_hi_62, regroupV0_hi_lo_lo_62};
  wire [3:0]         regroupV0_hi_hi_lo_lo_30 = {regroupV0_hi_34[631:630], regroupV0_hi_34[567:566]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_30 = {regroupV0_hi_34[759:758], regroupV0_hi_34[695:694]};
  wire [7:0]         regroupV0_hi_hi_lo_62 = {regroupV0_hi_hi_lo_hi_30, regroupV0_hi_hi_lo_lo_30};
  wire [3:0]         regroupV0_hi_hi_hi_lo_30 = {regroupV0_hi_34[887:886], regroupV0_hi_34[823:822]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_30 = {regroupV0_hi_34[1015:1014], regroupV0_hi_34[951:950]};
  wire [7:0]         regroupV0_hi_hi_hi_62 = {regroupV0_hi_hi_hi_hi_30, regroupV0_hi_hi_hi_lo_30};
  wire [15:0]        regroupV0_hi_hi_62 = {regroupV0_hi_hi_hi_62, regroupV0_hi_hi_lo_62};
  wire [31:0]        regroupV0_hi_62 = {regroupV0_hi_hi_62, regroupV0_hi_lo_62};
  wire [3:0]         regroupV0_lo_lo_lo_lo_31 = {regroupV0_lo_34[121:120], regroupV0_lo_34[57:56]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_31 = {regroupV0_lo_34[249:248], regroupV0_lo_34[185:184]};
  wire [7:0]         regroupV0_lo_lo_lo_63 = {regroupV0_lo_lo_lo_hi_31, regroupV0_lo_lo_lo_lo_31};
  wire [3:0]         regroupV0_lo_lo_hi_lo_31 = {regroupV0_lo_34[377:376], regroupV0_lo_34[313:312]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_31 = {regroupV0_lo_34[505:504], regroupV0_lo_34[441:440]};
  wire [7:0]         regroupV0_lo_lo_hi_63 = {regroupV0_lo_lo_hi_hi_31, regroupV0_lo_lo_hi_lo_31};
  wire [15:0]        regroupV0_lo_lo_63 = {regroupV0_lo_lo_hi_63, regroupV0_lo_lo_lo_63};
  wire [3:0]         regroupV0_lo_hi_lo_lo_31 = {regroupV0_lo_34[633:632], regroupV0_lo_34[569:568]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_31 = {regroupV0_lo_34[761:760], regroupV0_lo_34[697:696]};
  wire [7:0]         regroupV0_lo_hi_lo_63 = {regroupV0_lo_hi_lo_hi_31, regroupV0_lo_hi_lo_lo_31};
  wire [3:0]         regroupV0_lo_hi_hi_lo_31 = {regroupV0_lo_34[889:888], regroupV0_lo_34[825:824]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_31 = {regroupV0_lo_34[1017:1016], regroupV0_lo_34[953:952]};
  wire [7:0]         regroupV0_lo_hi_hi_63 = {regroupV0_lo_hi_hi_hi_31, regroupV0_lo_hi_hi_lo_31};
  wire [15:0]        regroupV0_lo_hi_63 = {regroupV0_lo_hi_hi_63, regroupV0_lo_hi_lo_63};
  wire [31:0]        regroupV0_lo_63 = {regroupV0_lo_hi_63, regroupV0_lo_lo_63};
  wire [3:0]         regroupV0_hi_lo_lo_lo_31 = {regroupV0_hi_34[121:120], regroupV0_hi_34[57:56]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_31 = {regroupV0_hi_34[249:248], regroupV0_hi_34[185:184]};
  wire [7:0]         regroupV0_hi_lo_lo_63 = {regroupV0_hi_lo_lo_hi_31, regroupV0_hi_lo_lo_lo_31};
  wire [3:0]         regroupV0_hi_lo_hi_lo_31 = {regroupV0_hi_34[377:376], regroupV0_hi_34[313:312]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_31 = {regroupV0_hi_34[505:504], regroupV0_hi_34[441:440]};
  wire [7:0]         regroupV0_hi_lo_hi_63 = {regroupV0_hi_lo_hi_hi_31, regroupV0_hi_lo_hi_lo_31};
  wire [15:0]        regroupV0_hi_lo_63 = {regroupV0_hi_lo_hi_63, regroupV0_hi_lo_lo_63};
  wire [3:0]         regroupV0_hi_hi_lo_lo_31 = {regroupV0_hi_34[633:632], regroupV0_hi_34[569:568]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_31 = {regroupV0_hi_34[761:760], regroupV0_hi_34[697:696]};
  wire [7:0]         regroupV0_hi_hi_lo_63 = {regroupV0_hi_hi_lo_hi_31, regroupV0_hi_hi_lo_lo_31};
  wire [3:0]         regroupV0_hi_hi_hi_lo_31 = {regroupV0_hi_34[889:888], regroupV0_hi_34[825:824]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_31 = {regroupV0_hi_34[1017:1016], regroupV0_hi_34[953:952]};
  wire [7:0]         regroupV0_hi_hi_hi_63 = {regroupV0_hi_hi_hi_hi_31, regroupV0_hi_hi_hi_lo_31};
  wire [15:0]        regroupV0_hi_hi_63 = {regroupV0_hi_hi_hi_63, regroupV0_hi_hi_lo_63};
  wire [31:0]        regroupV0_hi_63 = {regroupV0_hi_hi_63, regroupV0_hi_lo_63};
  wire [3:0]         regroupV0_lo_lo_lo_lo_32 = {regroupV0_lo_34[123:122], regroupV0_lo_34[59:58]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_32 = {regroupV0_lo_34[251:250], regroupV0_lo_34[187:186]};
  wire [7:0]         regroupV0_lo_lo_lo_64 = {regroupV0_lo_lo_lo_hi_32, regroupV0_lo_lo_lo_lo_32};
  wire [3:0]         regroupV0_lo_lo_hi_lo_32 = {regroupV0_lo_34[379:378], regroupV0_lo_34[315:314]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_32 = {regroupV0_lo_34[507:506], regroupV0_lo_34[443:442]};
  wire [7:0]         regroupV0_lo_lo_hi_64 = {regroupV0_lo_lo_hi_hi_32, regroupV0_lo_lo_hi_lo_32};
  wire [15:0]        regroupV0_lo_lo_64 = {regroupV0_lo_lo_hi_64, regroupV0_lo_lo_lo_64};
  wire [3:0]         regroupV0_lo_hi_lo_lo_32 = {regroupV0_lo_34[635:634], regroupV0_lo_34[571:570]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_32 = {regroupV0_lo_34[763:762], regroupV0_lo_34[699:698]};
  wire [7:0]         regroupV0_lo_hi_lo_64 = {regroupV0_lo_hi_lo_hi_32, regroupV0_lo_hi_lo_lo_32};
  wire [3:0]         regroupV0_lo_hi_hi_lo_32 = {regroupV0_lo_34[891:890], regroupV0_lo_34[827:826]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_32 = {regroupV0_lo_34[1019:1018], regroupV0_lo_34[955:954]};
  wire [7:0]         regroupV0_lo_hi_hi_64 = {regroupV0_lo_hi_hi_hi_32, regroupV0_lo_hi_hi_lo_32};
  wire [15:0]        regroupV0_lo_hi_64 = {regroupV0_lo_hi_hi_64, regroupV0_lo_hi_lo_64};
  wire [31:0]        regroupV0_lo_64 = {regroupV0_lo_hi_64, regroupV0_lo_lo_64};
  wire [3:0]         regroupV0_hi_lo_lo_lo_32 = {regroupV0_hi_34[123:122], regroupV0_hi_34[59:58]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_32 = {regroupV0_hi_34[251:250], regroupV0_hi_34[187:186]};
  wire [7:0]         regroupV0_hi_lo_lo_64 = {regroupV0_hi_lo_lo_hi_32, regroupV0_hi_lo_lo_lo_32};
  wire [3:0]         regroupV0_hi_lo_hi_lo_32 = {regroupV0_hi_34[379:378], regroupV0_hi_34[315:314]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_32 = {regroupV0_hi_34[507:506], regroupV0_hi_34[443:442]};
  wire [7:0]         regroupV0_hi_lo_hi_64 = {regroupV0_hi_lo_hi_hi_32, regroupV0_hi_lo_hi_lo_32};
  wire [15:0]        regroupV0_hi_lo_64 = {regroupV0_hi_lo_hi_64, regroupV0_hi_lo_lo_64};
  wire [3:0]         regroupV0_hi_hi_lo_lo_32 = {regroupV0_hi_34[635:634], regroupV0_hi_34[571:570]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_32 = {regroupV0_hi_34[763:762], regroupV0_hi_34[699:698]};
  wire [7:0]         regroupV0_hi_hi_lo_64 = {regroupV0_hi_hi_lo_hi_32, regroupV0_hi_hi_lo_lo_32};
  wire [3:0]         regroupV0_hi_hi_hi_lo_32 = {regroupV0_hi_34[891:890], regroupV0_hi_34[827:826]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_32 = {regroupV0_hi_34[1019:1018], regroupV0_hi_34[955:954]};
  wire [7:0]         regroupV0_hi_hi_hi_64 = {regroupV0_hi_hi_hi_hi_32, regroupV0_hi_hi_hi_lo_32};
  wire [15:0]        regroupV0_hi_hi_64 = {regroupV0_hi_hi_hi_64, regroupV0_hi_hi_lo_64};
  wire [31:0]        regroupV0_hi_64 = {regroupV0_hi_hi_64, regroupV0_hi_lo_64};
  wire [3:0]         regroupV0_lo_lo_lo_lo_33 = {regroupV0_lo_34[125:124], regroupV0_lo_34[61:60]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_33 = {regroupV0_lo_34[253:252], regroupV0_lo_34[189:188]};
  wire [7:0]         regroupV0_lo_lo_lo_65 = {regroupV0_lo_lo_lo_hi_33, regroupV0_lo_lo_lo_lo_33};
  wire [3:0]         regroupV0_lo_lo_hi_lo_33 = {regroupV0_lo_34[381:380], regroupV0_lo_34[317:316]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_33 = {regroupV0_lo_34[509:508], regroupV0_lo_34[445:444]};
  wire [7:0]         regroupV0_lo_lo_hi_65 = {regroupV0_lo_lo_hi_hi_33, regroupV0_lo_lo_hi_lo_33};
  wire [15:0]        regroupV0_lo_lo_65 = {regroupV0_lo_lo_hi_65, regroupV0_lo_lo_lo_65};
  wire [3:0]         regroupV0_lo_hi_lo_lo_33 = {regroupV0_lo_34[637:636], regroupV0_lo_34[573:572]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_33 = {regroupV0_lo_34[765:764], regroupV0_lo_34[701:700]};
  wire [7:0]         regroupV0_lo_hi_lo_65 = {regroupV0_lo_hi_lo_hi_33, regroupV0_lo_hi_lo_lo_33};
  wire [3:0]         regroupV0_lo_hi_hi_lo_33 = {regroupV0_lo_34[893:892], regroupV0_lo_34[829:828]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_33 = {regroupV0_lo_34[1021:1020], regroupV0_lo_34[957:956]};
  wire [7:0]         regroupV0_lo_hi_hi_65 = {regroupV0_lo_hi_hi_hi_33, regroupV0_lo_hi_hi_lo_33};
  wire [15:0]        regroupV0_lo_hi_65 = {regroupV0_lo_hi_hi_65, regroupV0_lo_hi_lo_65};
  wire [31:0]        regroupV0_lo_65 = {regroupV0_lo_hi_65, regroupV0_lo_lo_65};
  wire [3:0]         regroupV0_hi_lo_lo_lo_33 = {regroupV0_hi_34[125:124], regroupV0_hi_34[61:60]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_33 = {regroupV0_hi_34[253:252], regroupV0_hi_34[189:188]};
  wire [7:0]         regroupV0_hi_lo_lo_65 = {regroupV0_hi_lo_lo_hi_33, regroupV0_hi_lo_lo_lo_33};
  wire [3:0]         regroupV0_hi_lo_hi_lo_33 = {regroupV0_hi_34[381:380], regroupV0_hi_34[317:316]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_33 = {regroupV0_hi_34[509:508], regroupV0_hi_34[445:444]};
  wire [7:0]         regroupV0_hi_lo_hi_65 = {regroupV0_hi_lo_hi_hi_33, regroupV0_hi_lo_hi_lo_33};
  wire [15:0]        regroupV0_hi_lo_65 = {regroupV0_hi_lo_hi_65, regroupV0_hi_lo_lo_65};
  wire [3:0]         regroupV0_hi_hi_lo_lo_33 = {regroupV0_hi_34[637:636], regroupV0_hi_34[573:572]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_33 = {regroupV0_hi_34[765:764], regroupV0_hi_34[701:700]};
  wire [7:0]         regroupV0_hi_hi_lo_65 = {regroupV0_hi_hi_lo_hi_33, regroupV0_hi_hi_lo_lo_33};
  wire [3:0]         regroupV0_hi_hi_hi_lo_33 = {regroupV0_hi_34[893:892], regroupV0_hi_34[829:828]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_33 = {regroupV0_hi_34[1021:1020], regroupV0_hi_34[957:956]};
  wire [7:0]         regroupV0_hi_hi_hi_65 = {regroupV0_hi_hi_hi_hi_33, regroupV0_hi_hi_hi_lo_33};
  wire [15:0]        regroupV0_hi_hi_65 = {regroupV0_hi_hi_hi_65, regroupV0_hi_hi_lo_65};
  wire [31:0]        regroupV0_hi_65 = {regroupV0_hi_hi_65, regroupV0_hi_lo_65};
  wire [3:0]         regroupV0_lo_lo_lo_lo_34 = {regroupV0_lo_34[127:126], regroupV0_lo_34[63:62]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_34 = {regroupV0_lo_34[255:254], regroupV0_lo_34[191:190]};
  wire [7:0]         regroupV0_lo_lo_lo_66 = {regroupV0_lo_lo_lo_hi_34, regroupV0_lo_lo_lo_lo_34};
  wire [3:0]         regroupV0_lo_lo_hi_lo_34 = {regroupV0_lo_34[383:382], regroupV0_lo_34[319:318]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_34 = {regroupV0_lo_34[511:510], regroupV0_lo_34[447:446]};
  wire [7:0]         regroupV0_lo_lo_hi_66 = {regroupV0_lo_lo_hi_hi_34, regroupV0_lo_lo_hi_lo_34};
  wire [15:0]        regroupV0_lo_lo_66 = {regroupV0_lo_lo_hi_66, regroupV0_lo_lo_lo_66};
  wire [3:0]         regroupV0_lo_hi_lo_lo_34 = {regroupV0_lo_34[639:638], regroupV0_lo_34[575:574]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_34 = {regroupV0_lo_34[767:766], regroupV0_lo_34[703:702]};
  wire [7:0]         regroupV0_lo_hi_lo_66 = {regroupV0_lo_hi_lo_hi_34, regroupV0_lo_hi_lo_lo_34};
  wire [3:0]         regroupV0_lo_hi_hi_lo_34 = {regroupV0_lo_34[895:894], regroupV0_lo_34[831:830]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_34 = {regroupV0_lo_34[1023:1022], regroupV0_lo_34[959:958]};
  wire [7:0]         regroupV0_lo_hi_hi_66 = {regroupV0_lo_hi_hi_hi_34, regroupV0_lo_hi_hi_lo_34};
  wire [15:0]        regroupV0_lo_hi_66 = {regroupV0_lo_hi_hi_66, regroupV0_lo_hi_lo_66};
  wire [31:0]        regroupV0_lo_66 = {regroupV0_lo_hi_66, regroupV0_lo_lo_66};
  wire [3:0]         regroupV0_hi_lo_lo_lo_34 = {regroupV0_hi_34[127:126], regroupV0_hi_34[63:62]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_34 = {regroupV0_hi_34[255:254], regroupV0_hi_34[191:190]};
  wire [7:0]         regroupV0_hi_lo_lo_66 = {regroupV0_hi_lo_lo_hi_34, regroupV0_hi_lo_lo_lo_34};
  wire [3:0]         regroupV0_hi_lo_hi_lo_34 = {regroupV0_hi_34[383:382], regroupV0_hi_34[319:318]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_34 = {regroupV0_hi_34[511:510], regroupV0_hi_34[447:446]};
  wire [7:0]         regroupV0_hi_lo_hi_66 = {regroupV0_hi_lo_hi_hi_34, regroupV0_hi_lo_hi_lo_34};
  wire [15:0]        regroupV0_hi_lo_66 = {regroupV0_hi_lo_hi_66, regroupV0_hi_lo_lo_66};
  wire [3:0]         regroupV0_hi_hi_lo_lo_34 = {regroupV0_hi_34[639:638], regroupV0_hi_34[575:574]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_34 = {regroupV0_hi_34[767:766], regroupV0_hi_34[703:702]};
  wire [7:0]         regroupV0_hi_hi_lo_66 = {regroupV0_hi_hi_lo_hi_34, regroupV0_hi_hi_lo_lo_34};
  wire [3:0]         regroupV0_hi_hi_hi_lo_34 = {regroupV0_hi_34[895:894], regroupV0_hi_34[831:830]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_34 = {regroupV0_hi_34[1023:1022], regroupV0_hi_34[959:958]};
  wire [7:0]         regroupV0_hi_hi_hi_66 = {regroupV0_hi_hi_hi_hi_34, regroupV0_hi_hi_hi_lo_34};
  wire [15:0]        regroupV0_hi_hi_66 = {regroupV0_hi_hi_hi_66, regroupV0_hi_hi_lo_66};
  wire [31:0]        regroupV0_hi_66 = {regroupV0_hi_hi_66, regroupV0_hi_lo_66};
  wire [127:0]       regroupV0_lo_lo_lo_lo_35 = {regroupV0_hi_36, regroupV0_lo_36, regroupV0_hi_35, regroupV0_lo_35};
  wire [127:0]       regroupV0_lo_lo_lo_hi_35 = {regroupV0_hi_38, regroupV0_lo_38, regroupV0_hi_37, regroupV0_lo_37};
  wire [255:0]       regroupV0_lo_lo_lo_67 = {regroupV0_lo_lo_lo_hi_35, regroupV0_lo_lo_lo_lo_35};
  wire [127:0]       regroupV0_lo_lo_hi_lo_35 = {regroupV0_hi_40, regroupV0_lo_40, regroupV0_hi_39, regroupV0_lo_39};
  wire [127:0]       regroupV0_lo_lo_hi_hi_35 = {regroupV0_hi_42, regroupV0_lo_42, regroupV0_hi_41, regroupV0_lo_41};
  wire [255:0]       regroupV0_lo_lo_hi_67 = {regroupV0_lo_lo_hi_hi_35, regroupV0_lo_lo_hi_lo_35};
  wire [511:0]       regroupV0_lo_lo_67 = {regroupV0_lo_lo_hi_67, regroupV0_lo_lo_lo_67};
  wire [127:0]       regroupV0_lo_hi_lo_lo_35 = {regroupV0_hi_44, regroupV0_lo_44, regroupV0_hi_43, regroupV0_lo_43};
  wire [127:0]       regroupV0_lo_hi_lo_hi_35 = {regroupV0_hi_46, regroupV0_lo_46, regroupV0_hi_45, regroupV0_lo_45};
  wire [255:0]       regroupV0_lo_hi_lo_67 = {regroupV0_lo_hi_lo_hi_35, regroupV0_lo_hi_lo_lo_35};
  wire [127:0]       regroupV0_lo_hi_hi_lo_35 = {regroupV0_hi_48, regroupV0_lo_48, regroupV0_hi_47, regroupV0_lo_47};
  wire [127:0]       regroupV0_lo_hi_hi_hi_35 = {regroupV0_hi_50, regroupV0_lo_50, regroupV0_hi_49, regroupV0_lo_49};
  wire [255:0]       regroupV0_lo_hi_hi_67 = {regroupV0_lo_hi_hi_hi_35, regroupV0_lo_hi_hi_lo_35};
  wire [511:0]       regroupV0_lo_hi_67 = {regroupV0_lo_hi_hi_67, regroupV0_lo_hi_lo_67};
  wire [1023:0]      regroupV0_lo_67 = {regroupV0_lo_hi_67, regroupV0_lo_lo_67};
  wire [127:0]       regroupV0_hi_lo_lo_lo_35 = {regroupV0_hi_52, regroupV0_lo_52, regroupV0_hi_51, regroupV0_lo_51};
  wire [127:0]       regroupV0_hi_lo_lo_hi_35 = {regroupV0_hi_54, regroupV0_lo_54, regroupV0_hi_53, regroupV0_lo_53};
  wire [255:0]       regroupV0_hi_lo_lo_67 = {regroupV0_hi_lo_lo_hi_35, regroupV0_hi_lo_lo_lo_35};
  wire [127:0]       regroupV0_hi_lo_hi_lo_35 = {regroupV0_hi_56, regroupV0_lo_56, regroupV0_hi_55, regroupV0_lo_55};
  wire [127:0]       regroupV0_hi_lo_hi_hi_35 = {regroupV0_hi_58, regroupV0_lo_58, regroupV0_hi_57, regroupV0_lo_57};
  wire [255:0]       regroupV0_hi_lo_hi_67 = {regroupV0_hi_lo_hi_hi_35, regroupV0_hi_lo_hi_lo_35};
  wire [511:0]       regroupV0_hi_lo_67 = {regroupV0_hi_lo_hi_67, regroupV0_hi_lo_lo_67};
  wire [127:0]       regroupV0_hi_hi_lo_lo_35 = {regroupV0_hi_60, regroupV0_lo_60, regroupV0_hi_59, regroupV0_lo_59};
  wire [127:0]       regroupV0_hi_hi_lo_hi_35 = {regroupV0_hi_62, regroupV0_lo_62, regroupV0_hi_61, regroupV0_lo_61};
  wire [255:0]       regroupV0_hi_hi_lo_67 = {regroupV0_hi_hi_lo_hi_35, regroupV0_hi_hi_lo_lo_35};
  wire [127:0]       regroupV0_hi_hi_hi_lo_35 = {regroupV0_hi_64, regroupV0_lo_64, regroupV0_hi_63, regroupV0_lo_63};
  wire [127:0]       regroupV0_hi_hi_hi_hi_35 = {regroupV0_hi_66, regroupV0_lo_66, regroupV0_hi_65, regroupV0_lo_65};
  wire [255:0]       regroupV0_hi_hi_hi_67 = {regroupV0_hi_hi_hi_hi_35, regroupV0_hi_hi_hi_lo_35};
  wire [511:0]       regroupV0_hi_hi_67 = {regroupV0_hi_hi_hi_67, regroupV0_hi_hi_lo_67};
  wire [1023:0]      regroupV0_hi_67 = {regroupV0_hi_hi_67, regroupV0_hi_lo_67};
  wire [2047:0]      regroupV0_1 = {regroupV0_hi_67, regroupV0_lo_67};
  wire [127:0]       regroupV0_lo_lo_lo_lo_36 = {regroupV0_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_2};
  wire [127:0]       regroupV0_lo_lo_lo_hi_36 = {regroupV0_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_2};
  wire [255:0]       regroupV0_lo_lo_lo_68 = {regroupV0_lo_lo_lo_hi_36, regroupV0_lo_lo_lo_lo_36};
  wire [127:0]       regroupV0_lo_lo_hi_lo_36 = {regroupV0_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_2};
  wire [127:0]       regroupV0_lo_lo_hi_hi_36 = {regroupV0_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_2};
  wire [255:0]       regroupV0_lo_lo_hi_68 = {regroupV0_lo_lo_hi_hi_36, regroupV0_lo_lo_hi_lo_36};
  wire [511:0]       regroupV0_lo_lo_68 = {regroupV0_lo_lo_hi_68, regroupV0_lo_lo_lo_68};
  wire [127:0]       regroupV0_lo_hi_lo_lo_36 = {regroupV0_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_2};
  wire [127:0]       regroupV0_lo_hi_lo_hi_36 = {regroupV0_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_2};
  wire [255:0]       regroupV0_lo_hi_lo_68 = {regroupV0_lo_hi_lo_hi_36, regroupV0_lo_hi_lo_lo_36};
  wire [127:0]       regroupV0_lo_hi_hi_lo_36 = {regroupV0_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_2};
  wire [127:0]       regroupV0_lo_hi_hi_hi_36 = {regroupV0_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_2};
  wire [255:0]       regroupV0_lo_hi_hi_68 = {regroupV0_lo_hi_hi_hi_36, regroupV0_lo_hi_hi_lo_36};
  wire [511:0]       regroupV0_lo_hi_68 = {regroupV0_lo_hi_hi_68, regroupV0_lo_hi_lo_68};
  wire [1023:0]      regroupV0_lo_68 = {regroupV0_lo_hi_68, regroupV0_lo_lo_68};
  wire [127:0]       regroupV0_hi_lo_lo_lo_36 = {regroupV0_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_2};
  wire [127:0]       regroupV0_hi_lo_lo_hi_36 = {regroupV0_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_2};
  wire [255:0]       regroupV0_hi_lo_lo_68 = {regroupV0_hi_lo_lo_hi_36, regroupV0_hi_lo_lo_lo_36};
  wire [127:0]       regroupV0_hi_lo_hi_lo_36 = {regroupV0_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_2};
  wire [127:0]       regroupV0_hi_lo_hi_hi_36 = {regroupV0_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_2};
  wire [255:0]       regroupV0_hi_lo_hi_68 = {regroupV0_hi_lo_hi_hi_36, regroupV0_hi_lo_hi_lo_36};
  wire [511:0]       regroupV0_hi_lo_68 = {regroupV0_hi_lo_hi_68, regroupV0_hi_lo_lo_68};
  wire [127:0]       regroupV0_hi_hi_lo_lo_36 = {regroupV0_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_2};
  wire [127:0]       regroupV0_hi_hi_lo_hi_36 = {regroupV0_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_2};
  wire [255:0]       regroupV0_hi_hi_lo_68 = {regroupV0_hi_hi_lo_hi_36, regroupV0_hi_hi_lo_lo_36};
  wire [127:0]       regroupV0_hi_hi_hi_lo_36 = {regroupV0_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_2};
  wire [127:0]       regroupV0_hi_hi_hi_hi_36 = {regroupV0_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_2};
  wire [255:0]       regroupV0_hi_hi_hi_68 = {regroupV0_hi_hi_hi_hi_36, regroupV0_hi_hi_hi_lo_36};
  wire [511:0]       regroupV0_hi_hi_68 = {regroupV0_hi_hi_hi_68, regroupV0_hi_hi_lo_68};
  wire [1023:0]      regroupV0_hi_68 = {regroupV0_hi_hi_68, regroupV0_hi_lo_68};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_3 = {regroupV0_lo_68[32], regroupV0_lo_68[0]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_3 = {regroupV0_lo_68[96], regroupV0_lo_68[64]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_37 = {regroupV0_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_3 = {regroupV0_lo_68[160], regroupV0_lo_68[128]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_3 = {regroupV0_lo_68[224], regroupV0_lo_68[192]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_37 = {regroupV0_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_69 = {regroupV0_lo_lo_lo_hi_37, regroupV0_lo_lo_lo_lo_37};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_3 = {regroupV0_lo_68[288], regroupV0_lo_68[256]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_3 = {regroupV0_lo_68[352], regroupV0_lo_68[320]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_37 = {regroupV0_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_3 = {regroupV0_lo_68[416], regroupV0_lo_68[384]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_3 = {regroupV0_lo_68[480], regroupV0_lo_68[448]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_37 = {regroupV0_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_69 = {regroupV0_lo_lo_hi_hi_37, regroupV0_lo_lo_hi_lo_37};
  wire [15:0]        regroupV0_lo_lo_69 = {regroupV0_lo_lo_hi_69, regroupV0_lo_lo_lo_69};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_3 = {regroupV0_lo_68[544], regroupV0_lo_68[512]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_3 = {regroupV0_lo_68[608], regroupV0_lo_68[576]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_37 = {regroupV0_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_3 = {regroupV0_lo_68[672], regroupV0_lo_68[640]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_3 = {regroupV0_lo_68[736], regroupV0_lo_68[704]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_37 = {regroupV0_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_69 = {regroupV0_lo_hi_lo_hi_37, regroupV0_lo_hi_lo_lo_37};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_3 = {regroupV0_lo_68[800], regroupV0_lo_68[768]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_3 = {regroupV0_lo_68[864], regroupV0_lo_68[832]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_37 = {regroupV0_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_3 = {regroupV0_lo_68[928], regroupV0_lo_68[896]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_3 = {regroupV0_lo_68[992], regroupV0_lo_68[960]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_37 = {regroupV0_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_69 = {regroupV0_lo_hi_hi_hi_37, regroupV0_lo_hi_hi_lo_37};
  wire [15:0]        regroupV0_lo_hi_69 = {regroupV0_lo_hi_hi_69, regroupV0_lo_hi_lo_69};
  wire [31:0]        regroupV0_lo_69 = {regroupV0_lo_hi_69, regroupV0_lo_lo_69};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_3 = {regroupV0_hi_68[32], regroupV0_hi_68[0]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_3 = {regroupV0_hi_68[96], regroupV0_hi_68[64]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_37 = {regroupV0_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_3 = {regroupV0_hi_68[160], regroupV0_hi_68[128]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_3 = {regroupV0_hi_68[224], regroupV0_hi_68[192]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_37 = {regroupV0_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_69 = {regroupV0_hi_lo_lo_hi_37, regroupV0_hi_lo_lo_lo_37};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_3 = {regroupV0_hi_68[288], regroupV0_hi_68[256]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_3 = {regroupV0_hi_68[352], regroupV0_hi_68[320]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_37 = {regroupV0_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_3 = {regroupV0_hi_68[416], regroupV0_hi_68[384]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_3 = {regroupV0_hi_68[480], regroupV0_hi_68[448]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_37 = {regroupV0_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_69 = {regroupV0_hi_lo_hi_hi_37, regroupV0_hi_lo_hi_lo_37};
  wire [15:0]        regroupV0_hi_lo_69 = {regroupV0_hi_lo_hi_69, regroupV0_hi_lo_lo_69};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_3 = {regroupV0_hi_68[544], regroupV0_hi_68[512]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_3 = {regroupV0_hi_68[608], regroupV0_hi_68[576]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_37 = {regroupV0_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_3 = {regroupV0_hi_68[672], regroupV0_hi_68[640]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_3 = {regroupV0_hi_68[736], regroupV0_hi_68[704]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_37 = {regroupV0_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_69 = {regroupV0_hi_hi_lo_hi_37, regroupV0_hi_hi_lo_lo_37};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_3 = {regroupV0_hi_68[800], regroupV0_hi_68[768]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_3 = {regroupV0_hi_68[864], regroupV0_hi_68[832]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_37 = {regroupV0_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_3 = {regroupV0_hi_68[928], regroupV0_hi_68[896]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_3 = {regroupV0_hi_68[992], regroupV0_hi_68[960]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_37 = {regroupV0_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_69 = {regroupV0_hi_hi_hi_hi_37, regroupV0_hi_hi_hi_lo_37};
  wire [15:0]        regroupV0_hi_hi_69 = {regroupV0_hi_hi_hi_69, regroupV0_hi_hi_lo_69};
  wire [31:0]        regroupV0_hi_69 = {regroupV0_hi_hi_69, regroupV0_hi_lo_69};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_4 = {regroupV0_lo_68[33], regroupV0_lo_68[1]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_4 = {regroupV0_lo_68[97], regroupV0_lo_68[65]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_38 = {regroupV0_lo_lo_lo_lo_hi_4, regroupV0_lo_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_4 = {regroupV0_lo_68[161], regroupV0_lo_68[129]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_4 = {regroupV0_lo_68[225], regroupV0_lo_68[193]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_38 = {regroupV0_lo_lo_lo_hi_hi_4, regroupV0_lo_lo_lo_hi_lo_4};
  wire [7:0]         regroupV0_lo_lo_lo_70 = {regroupV0_lo_lo_lo_hi_38, regroupV0_lo_lo_lo_lo_38};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_4 = {regroupV0_lo_68[289], regroupV0_lo_68[257]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_4 = {regroupV0_lo_68[353], regroupV0_lo_68[321]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_38 = {regroupV0_lo_lo_hi_lo_hi_4, regroupV0_lo_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_4 = {regroupV0_lo_68[417], regroupV0_lo_68[385]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_4 = {regroupV0_lo_68[481], regroupV0_lo_68[449]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_38 = {regroupV0_lo_lo_hi_hi_hi_4, regroupV0_lo_lo_hi_hi_lo_4};
  wire [7:0]         regroupV0_lo_lo_hi_70 = {regroupV0_lo_lo_hi_hi_38, regroupV0_lo_lo_hi_lo_38};
  wire [15:0]        regroupV0_lo_lo_70 = {regroupV0_lo_lo_hi_70, regroupV0_lo_lo_lo_70};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_4 = {regroupV0_lo_68[545], regroupV0_lo_68[513]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_4 = {regroupV0_lo_68[609], regroupV0_lo_68[577]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_38 = {regroupV0_lo_hi_lo_lo_hi_4, regroupV0_lo_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_4 = {regroupV0_lo_68[673], regroupV0_lo_68[641]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_4 = {regroupV0_lo_68[737], regroupV0_lo_68[705]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_38 = {regroupV0_lo_hi_lo_hi_hi_4, regroupV0_lo_hi_lo_hi_lo_4};
  wire [7:0]         regroupV0_lo_hi_lo_70 = {regroupV0_lo_hi_lo_hi_38, regroupV0_lo_hi_lo_lo_38};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_4 = {regroupV0_lo_68[801], regroupV0_lo_68[769]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_4 = {regroupV0_lo_68[865], regroupV0_lo_68[833]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_38 = {regroupV0_lo_hi_hi_lo_hi_4, regroupV0_lo_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_4 = {regroupV0_lo_68[929], regroupV0_lo_68[897]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_4 = {regroupV0_lo_68[993], regroupV0_lo_68[961]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_38 = {regroupV0_lo_hi_hi_hi_hi_4, regroupV0_lo_hi_hi_hi_lo_4};
  wire [7:0]         regroupV0_lo_hi_hi_70 = {regroupV0_lo_hi_hi_hi_38, regroupV0_lo_hi_hi_lo_38};
  wire [15:0]        regroupV0_lo_hi_70 = {regroupV0_lo_hi_hi_70, regroupV0_lo_hi_lo_70};
  wire [31:0]        regroupV0_lo_70 = {regroupV0_lo_hi_70, regroupV0_lo_lo_70};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_4 = {regroupV0_hi_68[33], regroupV0_hi_68[1]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_4 = {regroupV0_hi_68[97], regroupV0_hi_68[65]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_38 = {regroupV0_hi_lo_lo_lo_hi_4, regroupV0_hi_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_4 = {regroupV0_hi_68[161], regroupV0_hi_68[129]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_4 = {regroupV0_hi_68[225], regroupV0_hi_68[193]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_38 = {regroupV0_hi_lo_lo_hi_hi_4, regroupV0_hi_lo_lo_hi_lo_4};
  wire [7:0]         regroupV0_hi_lo_lo_70 = {regroupV0_hi_lo_lo_hi_38, regroupV0_hi_lo_lo_lo_38};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_4 = {regroupV0_hi_68[289], regroupV0_hi_68[257]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_4 = {regroupV0_hi_68[353], regroupV0_hi_68[321]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_38 = {regroupV0_hi_lo_hi_lo_hi_4, regroupV0_hi_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_4 = {regroupV0_hi_68[417], regroupV0_hi_68[385]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_4 = {regroupV0_hi_68[481], regroupV0_hi_68[449]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_38 = {regroupV0_hi_lo_hi_hi_hi_4, regroupV0_hi_lo_hi_hi_lo_4};
  wire [7:0]         regroupV0_hi_lo_hi_70 = {regroupV0_hi_lo_hi_hi_38, regroupV0_hi_lo_hi_lo_38};
  wire [15:0]        regroupV0_hi_lo_70 = {regroupV0_hi_lo_hi_70, regroupV0_hi_lo_lo_70};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_4 = {regroupV0_hi_68[545], regroupV0_hi_68[513]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_4 = {regroupV0_hi_68[609], regroupV0_hi_68[577]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_38 = {regroupV0_hi_hi_lo_lo_hi_4, regroupV0_hi_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_4 = {regroupV0_hi_68[673], regroupV0_hi_68[641]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_4 = {regroupV0_hi_68[737], regroupV0_hi_68[705]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_38 = {regroupV0_hi_hi_lo_hi_hi_4, regroupV0_hi_hi_lo_hi_lo_4};
  wire [7:0]         regroupV0_hi_hi_lo_70 = {regroupV0_hi_hi_lo_hi_38, regroupV0_hi_hi_lo_lo_38};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_4 = {regroupV0_hi_68[801], regroupV0_hi_68[769]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_4 = {regroupV0_hi_68[865], regroupV0_hi_68[833]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_38 = {regroupV0_hi_hi_hi_lo_hi_4, regroupV0_hi_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_4 = {regroupV0_hi_68[929], regroupV0_hi_68[897]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_4 = {regroupV0_hi_68[993], regroupV0_hi_68[961]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_38 = {regroupV0_hi_hi_hi_hi_hi_4, regroupV0_hi_hi_hi_hi_lo_4};
  wire [7:0]         regroupV0_hi_hi_hi_70 = {regroupV0_hi_hi_hi_hi_38, regroupV0_hi_hi_hi_lo_38};
  wire [15:0]        regroupV0_hi_hi_70 = {regroupV0_hi_hi_hi_70, regroupV0_hi_hi_lo_70};
  wire [31:0]        regroupV0_hi_70 = {regroupV0_hi_hi_70, regroupV0_hi_lo_70};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_5 = {regroupV0_lo_68[34], regroupV0_lo_68[2]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_5 = {regroupV0_lo_68[98], regroupV0_lo_68[66]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_39 = {regroupV0_lo_lo_lo_lo_hi_5, regroupV0_lo_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_5 = {regroupV0_lo_68[162], regroupV0_lo_68[130]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_5 = {regroupV0_lo_68[226], regroupV0_lo_68[194]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_39 = {regroupV0_lo_lo_lo_hi_hi_5, regroupV0_lo_lo_lo_hi_lo_5};
  wire [7:0]         regroupV0_lo_lo_lo_71 = {regroupV0_lo_lo_lo_hi_39, regroupV0_lo_lo_lo_lo_39};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_5 = {regroupV0_lo_68[290], regroupV0_lo_68[258]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_5 = {regroupV0_lo_68[354], regroupV0_lo_68[322]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_39 = {regroupV0_lo_lo_hi_lo_hi_5, regroupV0_lo_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_5 = {regroupV0_lo_68[418], regroupV0_lo_68[386]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_5 = {regroupV0_lo_68[482], regroupV0_lo_68[450]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_39 = {regroupV0_lo_lo_hi_hi_hi_5, regroupV0_lo_lo_hi_hi_lo_5};
  wire [7:0]         regroupV0_lo_lo_hi_71 = {regroupV0_lo_lo_hi_hi_39, regroupV0_lo_lo_hi_lo_39};
  wire [15:0]        regroupV0_lo_lo_71 = {regroupV0_lo_lo_hi_71, regroupV0_lo_lo_lo_71};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_5 = {regroupV0_lo_68[546], regroupV0_lo_68[514]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_5 = {regroupV0_lo_68[610], regroupV0_lo_68[578]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_39 = {regroupV0_lo_hi_lo_lo_hi_5, regroupV0_lo_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_5 = {regroupV0_lo_68[674], regroupV0_lo_68[642]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_5 = {regroupV0_lo_68[738], regroupV0_lo_68[706]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_39 = {regroupV0_lo_hi_lo_hi_hi_5, regroupV0_lo_hi_lo_hi_lo_5};
  wire [7:0]         regroupV0_lo_hi_lo_71 = {regroupV0_lo_hi_lo_hi_39, regroupV0_lo_hi_lo_lo_39};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_5 = {regroupV0_lo_68[802], regroupV0_lo_68[770]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_5 = {regroupV0_lo_68[866], regroupV0_lo_68[834]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_39 = {regroupV0_lo_hi_hi_lo_hi_5, regroupV0_lo_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_5 = {regroupV0_lo_68[930], regroupV0_lo_68[898]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_5 = {regroupV0_lo_68[994], regroupV0_lo_68[962]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_39 = {regroupV0_lo_hi_hi_hi_hi_5, regroupV0_lo_hi_hi_hi_lo_5};
  wire [7:0]         regroupV0_lo_hi_hi_71 = {regroupV0_lo_hi_hi_hi_39, regroupV0_lo_hi_hi_lo_39};
  wire [15:0]        regroupV0_lo_hi_71 = {regroupV0_lo_hi_hi_71, regroupV0_lo_hi_lo_71};
  wire [31:0]        regroupV0_lo_71 = {regroupV0_lo_hi_71, regroupV0_lo_lo_71};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_5 = {regroupV0_hi_68[34], regroupV0_hi_68[2]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_5 = {regroupV0_hi_68[98], regroupV0_hi_68[66]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_39 = {regroupV0_hi_lo_lo_lo_hi_5, regroupV0_hi_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_5 = {regroupV0_hi_68[162], regroupV0_hi_68[130]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_5 = {regroupV0_hi_68[226], regroupV0_hi_68[194]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_39 = {regroupV0_hi_lo_lo_hi_hi_5, regroupV0_hi_lo_lo_hi_lo_5};
  wire [7:0]         regroupV0_hi_lo_lo_71 = {regroupV0_hi_lo_lo_hi_39, regroupV0_hi_lo_lo_lo_39};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_5 = {regroupV0_hi_68[290], regroupV0_hi_68[258]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_5 = {regroupV0_hi_68[354], regroupV0_hi_68[322]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_39 = {regroupV0_hi_lo_hi_lo_hi_5, regroupV0_hi_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_5 = {regroupV0_hi_68[418], regroupV0_hi_68[386]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_5 = {regroupV0_hi_68[482], regroupV0_hi_68[450]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_39 = {regroupV0_hi_lo_hi_hi_hi_5, regroupV0_hi_lo_hi_hi_lo_5};
  wire [7:0]         regroupV0_hi_lo_hi_71 = {regroupV0_hi_lo_hi_hi_39, regroupV0_hi_lo_hi_lo_39};
  wire [15:0]        regroupV0_hi_lo_71 = {regroupV0_hi_lo_hi_71, regroupV0_hi_lo_lo_71};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_5 = {regroupV0_hi_68[546], regroupV0_hi_68[514]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_5 = {regroupV0_hi_68[610], regroupV0_hi_68[578]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_39 = {regroupV0_hi_hi_lo_lo_hi_5, regroupV0_hi_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_5 = {regroupV0_hi_68[674], regroupV0_hi_68[642]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_5 = {regroupV0_hi_68[738], regroupV0_hi_68[706]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_39 = {regroupV0_hi_hi_lo_hi_hi_5, regroupV0_hi_hi_lo_hi_lo_5};
  wire [7:0]         regroupV0_hi_hi_lo_71 = {regroupV0_hi_hi_lo_hi_39, regroupV0_hi_hi_lo_lo_39};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_5 = {regroupV0_hi_68[802], regroupV0_hi_68[770]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_5 = {regroupV0_hi_68[866], regroupV0_hi_68[834]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_39 = {regroupV0_hi_hi_hi_lo_hi_5, regroupV0_hi_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_5 = {regroupV0_hi_68[930], regroupV0_hi_68[898]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_5 = {regroupV0_hi_68[994], regroupV0_hi_68[962]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_39 = {regroupV0_hi_hi_hi_hi_hi_5, regroupV0_hi_hi_hi_hi_lo_5};
  wire [7:0]         regroupV0_hi_hi_hi_71 = {regroupV0_hi_hi_hi_hi_39, regroupV0_hi_hi_hi_lo_39};
  wire [15:0]        regroupV0_hi_hi_71 = {regroupV0_hi_hi_hi_71, regroupV0_hi_hi_lo_71};
  wire [31:0]        regroupV0_hi_71 = {regroupV0_hi_hi_71, regroupV0_hi_lo_71};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_6 = {regroupV0_lo_68[35], regroupV0_lo_68[3]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_6 = {regroupV0_lo_68[99], regroupV0_lo_68[67]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_40 = {regroupV0_lo_lo_lo_lo_hi_6, regroupV0_lo_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_6 = {regroupV0_lo_68[163], regroupV0_lo_68[131]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_6 = {regroupV0_lo_68[227], regroupV0_lo_68[195]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_40 = {regroupV0_lo_lo_lo_hi_hi_6, regroupV0_lo_lo_lo_hi_lo_6};
  wire [7:0]         regroupV0_lo_lo_lo_72 = {regroupV0_lo_lo_lo_hi_40, regroupV0_lo_lo_lo_lo_40};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_6 = {regroupV0_lo_68[291], regroupV0_lo_68[259]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_6 = {regroupV0_lo_68[355], regroupV0_lo_68[323]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_40 = {regroupV0_lo_lo_hi_lo_hi_6, regroupV0_lo_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_6 = {regroupV0_lo_68[419], regroupV0_lo_68[387]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_6 = {regroupV0_lo_68[483], regroupV0_lo_68[451]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_40 = {regroupV0_lo_lo_hi_hi_hi_6, regroupV0_lo_lo_hi_hi_lo_6};
  wire [7:0]         regroupV0_lo_lo_hi_72 = {regroupV0_lo_lo_hi_hi_40, regroupV0_lo_lo_hi_lo_40};
  wire [15:0]        regroupV0_lo_lo_72 = {regroupV0_lo_lo_hi_72, regroupV0_lo_lo_lo_72};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_6 = {regroupV0_lo_68[547], regroupV0_lo_68[515]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_6 = {regroupV0_lo_68[611], regroupV0_lo_68[579]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_40 = {regroupV0_lo_hi_lo_lo_hi_6, regroupV0_lo_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_6 = {regroupV0_lo_68[675], regroupV0_lo_68[643]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_6 = {regroupV0_lo_68[739], regroupV0_lo_68[707]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_40 = {regroupV0_lo_hi_lo_hi_hi_6, regroupV0_lo_hi_lo_hi_lo_6};
  wire [7:0]         regroupV0_lo_hi_lo_72 = {regroupV0_lo_hi_lo_hi_40, regroupV0_lo_hi_lo_lo_40};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_6 = {regroupV0_lo_68[803], regroupV0_lo_68[771]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_6 = {regroupV0_lo_68[867], regroupV0_lo_68[835]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_40 = {regroupV0_lo_hi_hi_lo_hi_6, regroupV0_lo_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_6 = {regroupV0_lo_68[931], regroupV0_lo_68[899]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_6 = {regroupV0_lo_68[995], regroupV0_lo_68[963]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_40 = {regroupV0_lo_hi_hi_hi_hi_6, regroupV0_lo_hi_hi_hi_lo_6};
  wire [7:0]         regroupV0_lo_hi_hi_72 = {regroupV0_lo_hi_hi_hi_40, regroupV0_lo_hi_hi_lo_40};
  wire [15:0]        regroupV0_lo_hi_72 = {regroupV0_lo_hi_hi_72, regroupV0_lo_hi_lo_72};
  wire [31:0]        regroupV0_lo_72 = {regroupV0_lo_hi_72, regroupV0_lo_lo_72};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_6 = {regroupV0_hi_68[35], regroupV0_hi_68[3]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_6 = {regroupV0_hi_68[99], regroupV0_hi_68[67]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_40 = {regroupV0_hi_lo_lo_lo_hi_6, regroupV0_hi_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_6 = {regroupV0_hi_68[163], regroupV0_hi_68[131]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_6 = {regroupV0_hi_68[227], regroupV0_hi_68[195]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_40 = {regroupV0_hi_lo_lo_hi_hi_6, regroupV0_hi_lo_lo_hi_lo_6};
  wire [7:0]         regroupV0_hi_lo_lo_72 = {regroupV0_hi_lo_lo_hi_40, regroupV0_hi_lo_lo_lo_40};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_6 = {regroupV0_hi_68[291], regroupV0_hi_68[259]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_6 = {regroupV0_hi_68[355], regroupV0_hi_68[323]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_40 = {regroupV0_hi_lo_hi_lo_hi_6, regroupV0_hi_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_6 = {regroupV0_hi_68[419], regroupV0_hi_68[387]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_6 = {regroupV0_hi_68[483], regroupV0_hi_68[451]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_40 = {regroupV0_hi_lo_hi_hi_hi_6, regroupV0_hi_lo_hi_hi_lo_6};
  wire [7:0]         regroupV0_hi_lo_hi_72 = {regroupV0_hi_lo_hi_hi_40, regroupV0_hi_lo_hi_lo_40};
  wire [15:0]        regroupV0_hi_lo_72 = {regroupV0_hi_lo_hi_72, regroupV0_hi_lo_lo_72};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_6 = {regroupV0_hi_68[547], regroupV0_hi_68[515]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_6 = {regroupV0_hi_68[611], regroupV0_hi_68[579]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_40 = {regroupV0_hi_hi_lo_lo_hi_6, regroupV0_hi_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_6 = {regroupV0_hi_68[675], regroupV0_hi_68[643]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_6 = {regroupV0_hi_68[739], regroupV0_hi_68[707]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_40 = {regroupV0_hi_hi_lo_hi_hi_6, regroupV0_hi_hi_lo_hi_lo_6};
  wire [7:0]         regroupV0_hi_hi_lo_72 = {regroupV0_hi_hi_lo_hi_40, regroupV0_hi_hi_lo_lo_40};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_6 = {regroupV0_hi_68[803], regroupV0_hi_68[771]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_6 = {regroupV0_hi_68[867], regroupV0_hi_68[835]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_40 = {regroupV0_hi_hi_hi_lo_hi_6, regroupV0_hi_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_6 = {regroupV0_hi_68[931], regroupV0_hi_68[899]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_6 = {regroupV0_hi_68[995], regroupV0_hi_68[963]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_40 = {regroupV0_hi_hi_hi_hi_hi_6, regroupV0_hi_hi_hi_hi_lo_6};
  wire [7:0]         regroupV0_hi_hi_hi_72 = {regroupV0_hi_hi_hi_hi_40, regroupV0_hi_hi_hi_lo_40};
  wire [15:0]        regroupV0_hi_hi_72 = {regroupV0_hi_hi_hi_72, regroupV0_hi_hi_lo_72};
  wire [31:0]        regroupV0_hi_72 = {regroupV0_hi_hi_72, regroupV0_hi_lo_72};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_7 = {regroupV0_lo_68[36], regroupV0_lo_68[4]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_7 = {regroupV0_lo_68[100], regroupV0_lo_68[68]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_41 = {regroupV0_lo_lo_lo_lo_hi_7, regroupV0_lo_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_7 = {regroupV0_lo_68[164], regroupV0_lo_68[132]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_7 = {regroupV0_lo_68[228], regroupV0_lo_68[196]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_41 = {regroupV0_lo_lo_lo_hi_hi_7, regroupV0_lo_lo_lo_hi_lo_7};
  wire [7:0]         regroupV0_lo_lo_lo_73 = {regroupV0_lo_lo_lo_hi_41, regroupV0_lo_lo_lo_lo_41};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_7 = {regroupV0_lo_68[292], regroupV0_lo_68[260]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_7 = {regroupV0_lo_68[356], regroupV0_lo_68[324]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_41 = {regroupV0_lo_lo_hi_lo_hi_7, regroupV0_lo_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_7 = {regroupV0_lo_68[420], regroupV0_lo_68[388]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_7 = {regroupV0_lo_68[484], regroupV0_lo_68[452]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_41 = {regroupV0_lo_lo_hi_hi_hi_7, regroupV0_lo_lo_hi_hi_lo_7};
  wire [7:0]         regroupV0_lo_lo_hi_73 = {regroupV0_lo_lo_hi_hi_41, regroupV0_lo_lo_hi_lo_41};
  wire [15:0]        regroupV0_lo_lo_73 = {regroupV0_lo_lo_hi_73, regroupV0_lo_lo_lo_73};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_7 = {regroupV0_lo_68[548], regroupV0_lo_68[516]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_7 = {regroupV0_lo_68[612], regroupV0_lo_68[580]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_41 = {regroupV0_lo_hi_lo_lo_hi_7, regroupV0_lo_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_7 = {regroupV0_lo_68[676], regroupV0_lo_68[644]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_7 = {regroupV0_lo_68[740], regroupV0_lo_68[708]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_41 = {regroupV0_lo_hi_lo_hi_hi_7, regroupV0_lo_hi_lo_hi_lo_7};
  wire [7:0]         regroupV0_lo_hi_lo_73 = {regroupV0_lo_hi_lo_hi_41, regroupV0_lo_hi_lo_lo_41};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_7 = {regroupV0_lo_68[804], regroupV0_lo_68[772]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_7 = {regroupV0_lo_68[868], regroupV0_lo_68[836]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_41 = {regroupV0_lo_hi_hi_lo_hi_7, regroupV0_lo_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_7 = {regroupV0_lo_68[932], regroupV0_lo_68[900]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_7 = {regroupV0_lo_68[996], regroupV0_lo_68[964]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_41 = {regroupV0_lo_hi_hi_hi_hi_7, regroupV0_lo_hi_hi_hi_lo_7};
  wire [7:0]         regroupV0_lo_hi_hi_73 = {regroupV0_lo_hi_hi_hi_41, regroupV0_lo_hi_hi_lo_41};
  wire [15:0]        regroupV0_lo_hi_73 = {regroupV0_lo_hi_hi_73, regroupV0_lo_hi_lo_73};
  wire [31:0]        regroupV0_lo_73 = {regroupV0_lo_hi_73, regroupV0_lo_lo_73};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_7 = {regroupV0_hi_68[36], regroupV0_hi_68[4]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_7 = {regroupV0_hi_68[100], regroupV0_hi_68[68]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_41 = {regroupV0_hi_lo_lo_lo_hi_7, regroupV0_hi_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_7 = {regroupV0_hi_68[164], regroupV0_hi_68[132]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_7 = {regroupV0_hi_68[228], regroupV0_hi_68[196]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_41 = {regroupV0_hi_lo_lo_hi_hi_7, regroupV0_hi_lo_lo_hi_lo_7};
  wire [7:0]         regroupV0_hi_lo_lo_73 = {regroupV0_hi_lo_lo_hi_41, regroupV0_hi_lo_lo_lo_41};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_7 = {regroupV0_hi_68[292], regroupV0_hi_68[260]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_7 = {regroupV0_hi_68[356], regroupV0_hi_68[324]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_41 = {regroupV0_hi_lo_hi_lo_hi_7, regroupV0_hi_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_7 = {regroupV0_hi_68[420], regroupV0_hi_68[388]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_7 = {regroupV0_hi_68[484], regroupV0_hi_68[452]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_41 = {regroupV0_hi_lo_hi_hi_hi_7, regroupV0_hi_lo_hi_hi_lo_7};
  wire [7:0]         regroupV0_hi_lo_hi_73 = {regroupV0_hi_lo_hi_hi_41, regroupV0_hi_lo_hi_lo_41};
  wire [15:0]        regroupV0_hi_lo_73 = {regroupV0_hi_lo_hi_73, regroupV0_hi_lo_lo_73};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_7 = {regroupV0_hi_68[548], regroupV0_hi_68[516]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_7 = {regroupV0_hi_68[612], regroupV0_hi_68[580]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_41 = {regroupV0_hi_hi_lo_lo_hi_7, regroupV0_hi_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_7 = {regroupV0_hi_68[676], regroupV0_hi_68[644]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_7 = {regroupV0_hi_68[740], regroupV0_hi_68[708]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_41 = {regroupV0_hi_hi_lo_hi_hi_7, regroupV0_hi_hi_lo_hi_lo_7};
  wire [7:0]         regroupV0_hi_hi_lo_73 = {regroupV0_hi_hi_lo_hi_41, regroupV0_hi_hi_lo_lo_41};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_7 = {regroupV0_hi_68[804], regroupV0_hi_68[772]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_7 = {regroupV0_hi_68[868], regroupV0_hi_68[836]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_41 = {regroupV0_hi_hi_hi_lo_hi_7, regroupV0_hi_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_7 = {regroupV0_hi_68[932], regroupV0_hi_68[900]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_7 = {regroupV0_hi_68[996], regroupV0_hi_68[964]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_41 = {regroupV0_hi_hi_hi_hi_hi_7, regroupV0_hi_hi_hi_hi_lo_7};
  wire [7:0]         regroupV0_hi_hi_hi_73 = {regroupV0_hi_hi_hi_hi_41, regroupV0_hi_hi_hi_lo_41};
  wire [15:0]        regroupV0_hi_hi_73 = {regroupV0_hi_hi_hi_73, regroupV0_hi_hi_lo_73};
  wire [31:0]        regroupV0_hi_73 = {regroupV0_hi_hi_73, regroupV0_hi_lo_73};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_8 = {regroupV0_lo_68[37], regroupV0_lo_68[5]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_8 = {regroupV0_lo_68[101], regroupV0_lo_68[69]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_42 = {regroupV0_lo_lo_lo_lo_hi_8, regroupV0_lo_lo_lo_lo_lo_8};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_8 = {regroupV0_lo_68[165], regroupV0_lo_68[133]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_8 = {regroupV0_lo_68[229], regroupV0_lo_68[197]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_42 = {regroupV0_lo_lo_lo_hi_hi_8, regroupV0_lo_lo_lo_hi_lo_8};
  wire [7:0]         regroupV0_lo_lo_lo_74 = {regroupV0_lo_lo_lo_hi_42, regroupV0_lo_lo_lo_lo_42};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_8 = {regroupV0_lo_68[293], regroupV0_lo_68[261]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_8 = {regroupV0_lo_68[357], regroupV0_lo_68[325]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_42 = {regroupV0_lo_lo_hi_lo_hi_8, regroupV0_lo_lo_hi_lo_lo_8};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_8 = {regroupV0_lo_68[421], regroupV0_lo_68[389]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_8 = {regroupV0_lo_68[485], regroupV0_lo_68[453]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_42 = {regroupV0_lo_lo_hi_hi_hi_8, regroupV0_lo_lo_hi_hi_lo_8};
  wire [7:0]         regroupV0_lo_lo_hi_74 = {regroupV0_lo_lo_hi_hi_42, regroupV0_lo_lo_hi_lo_42};
  wire [15:0]        regroupV0_lo_lo_74 = {regroupV0_lo_lo_hi_74, regroupV0_lo_lo_lo_74};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_8 = {regroupV0_lo_68[549], regroupV0_lo_68[517]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_8 = {regroupV0_lo_68[613], regroupV0_lo_68[581]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_42 = {regroupV0_lo_hi_lo_lo_hi_8, regroupV0_lo_hi_lo_lo_lo_8};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_8 = {regroupV0_lo_68[677], regroupV0_lo_68[645]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_8 = {regroupV0_lo_68[741], regroupV0_lo_68[709]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_42 = {regroupV0_lo_hi_lo_hi_hi_8, regroupV0_lo_hi_lo_hi_lo_8};
  wire [7:0]         regroupV0_lo_hi_lo_74 = {regroupV0_lo_hi_lo_hi_42, regroupV0_lo_hi_lo_lo_42};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_8 = {regroupV0_lo_68[805], regroupV0_lo_68[773]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_8 = {regroupV0_lo_68[869], regroupV0_lo_68[837]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_42 = {regroupV0_lo_hi_hi_lo_hi_8, regroupV0_lo_hi_hi_lo_lo_8};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_8 = {regroupV0_lo_68[933], regroupV0_lo_68[901]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_8 = {regroupV0_lo_68[997], regroupV0_lo_68[965]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_42 = {regroupV0_lo_hi_hi_hi_hi_8, regroupV0_lo_hi_hi_hi_lo_8};
  wire [7:0]         regroupV0_lo_hi_hi_74 = {regroupV0_lo_hi_hi_hi_42, regroupV0_lo_hi_hi_lo_42};
  wire [15:0]        regroupV0_lo_hi_74 = {regroupV0_lo_hi_hi_74, regroupV0_lo_hi_lo_74};
  wire [31:0]        regroupV0_lo_74 = {regroupV0_lo_hi_74, regroupV0_lo_lo_74};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_8 = {regroupV0_hi_68[37], regroupV0_hi_68[5]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_8 = {regroupV0_hi_68[101], regroupV0_hi_68[69]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_42 = {regroupV0_hi_lo_lo_lo_hi_8, regroupV0_hi_lo_lo_lo_lo_8};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_8 = {regroupV0_hi_68[165], regroupV0_hi_68[133]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_8 = {regroupV0_hi_68[229], regroupV0_hi_68[197]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_42 = {regroupV0_hi_lo_lo_hi_hi_8, regroupV0_hi_lo_lo_hi_lo_8};
  wire [7:0]         regroupV0_hi_lo_lo_74 = {regroupV0_hi_lo_lo_hi_42, regroupV0_hi_lo_lo_lo_42};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_8 = {regroupV0_hi_68[293], regroupV0_hi_68[261]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_8 = {regroupV0_hi_68[357], regroupV0_hi_68[325]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_42 = {regroupV0_hi_lo_hi_lo_hi_8, regroupV0_hi_lo_hi_lo_lo_8};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_8 = {regroupV0_hi_68[421], regroupV0_hi_68[389]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_8 = {regroupV0_hi_68[485], regroupV0_hi_68[453]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_42 = {regroupV0_hi_lo_hi_hi_hi_8, regroupV0_hi_lo_hi_hi_lo_8};
  wire [7:0]         regroupV0_hi_lo_hi_74 = {regroupV0_hi_lo_hi_hi_42, regroupV0_hi_lo_hi_lo_42};
  wire [15:0]        regroupV0_hi_lo_74 = {regroupV0_hi_lo_hi_74, regroupV0_hi_lo_lo_74};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_8 = {regroupV0_hi_68[549], regroupV0_hi_68[517]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_8 = {regroupV0_hi_68[613], regroupV0_hi_68[581]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_42 = {regroupV0_hi_hi_lo_lo_hi_8, regroupV0_hi_hi_lo_lo_lo_8};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_8 = {regroupV0_hi_68[677], regroupV0_hi_68[645]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_8 = {regroupV0_hi_68[741], regroupV0_hi_68[709]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_42 = {regroupV0_hi_hi_lo_hi_hi_8, regroupV0_hi_hi_lo_hi_lo_8};
  wire [7:0]         regroupV0_hi_hi_lo_74 = {regroupV0_hi_hi_lo_hi_42, regroupV0_hi_hi_lo_lo_42};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_8 = {regroupV0_hi_68[805], regroupV0_hi_68[773]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_8 = {regroupV0_hi_68[869], regroupV0_hi_68[837]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_42 = {regroupV0_hi_hi_hi_lo_hi_8, regroupV0_hi_hi_hi_lo_lo_8};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_8 = {regroupV0_hi_68[933], regroupV0_hi_68[901]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_8 = {regroupV0_hi_68[997], regroupV0_hi_68[965]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_42 = {regroupV0_hi_hi_hi_hi_hi_8, regroupV0_hi_hi_hi_hi_lo_8};
  wire [7:0]         regroupV0_hi_hi_hi_74 = {regroupV0_hi_hi_hi_hi_42, regroupV0_hi_hi_hi_lo_42};
  wire [15:0]        regroupV0_hi_hi_74 = {regroupV0_hi_hi_hi_74, regroupV0_hi_hi_lo_74};
  wire [31:0]        regroupV0_hi_74 = {regroupV0_hi_hi_74, regroupV0_hi_lo_74};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_9 = {regroupV0_lo_68[38], regroupV0_lo_68[6]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_9 = {regroupV0_lo_68[102], regroupV0_lo_68[70]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_43 = {regroupV0_lo_lo_lo_lo_hi_9, regroupV0_lo_lo_lo_lo_lo_9};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_9 = {regroupV0_lo_68[166], regroupV0_lo_68[134]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_9 = {regroupV0_lo_68[230], regroupV0_lo_68[198]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_43 = {regroupV0_lo_lo_lo_hi_hi_9, regroupV0_lo_lo_lo_hi_lo_9};
  wire [7:0]         regroupV0_lo_lo_lo_75 = {regroupV0_lo_lo_lo_hi_43, regroupV0_lo_lo_lo_lo_43};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_9 = {regroupV0_lo_68[294], regroupV0_lo_68[262]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_9 = {regroupV0_lo_68[358], regroupV0_lo_68[326]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_43 = {regroupV0_lo_lo_hi_lo_hi_9, regroupV0_lo_lo_hi_lo_lo_9};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_9 = {regroupV0_lo_68[422], regroupV0_lo_68[390]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_9 = {regroupV0_lo_68[486], regroupV0_lo_68[454]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_43 = {regroupV0_lo_lo_hi_hi_hi_9, regroupV0_lo_lo_hi_hi_lo_9};
  wire [7:0]         regroupV0_lo_lo_hi_75 = {regroupV0_lo_lo_hi_hi_43, regroupV0_lo_lo_hi_lo_43};
  wire [15:0]        regroupV0_lo_lo_75 = {regroupV0_lo_lo_hi_75, regroupV0_lo_lo_lo_75};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_9 = {regroupV0_lo_68[550], regroupV0_lo_68[518]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_9 = {regroupV0_lo_68[614], regroupV0_lo_68[582]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_43 = {regroupV0_lo_hi_lo_lo_hi_9, regroupV0_lo_hi_lo_lo_lo_9};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_9 = {regroupV0_lo_68[678], regroupV0_lo_68[646]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_9 = {regroupV0_lo_68[742], regroupV0_lo_68[710]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_43 = {regroupV0_lo_hi_lo_hi_hi_9, regroupV0_lo_hi_lo_hi_lo_9};
  wire [7:0]         regroupV0_lo_hi_lo_75 = {regroupV0_lo_hi_lo_hi_43, regroupV0_lo_hi_lo_lo_43};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_9 = {regroupV0_lo_68[806], regroupV0_lo_68[774]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_9 = {regroupV0_lo_68[870], regroupV0_lo_68[838]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_43 = {regroupV0_lo_hi_hi_lo_hi_9, regroupV0_lo_hi_hi_lo_lo_9};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_9 = {regroupV0_lo_68[934], regroupV0_lo_68[902]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_9 = {regroupV0_lo_68[998], regroupV0_lo_68[966]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_43 = {regroupV0_lo_hi_hi_hi_hi_9, regroupV0_lo_hi_hi_hi_lo_9};
  wire [7:0]         regroupV0_lo_hi_hi_75 = {regroupV0_lo_hi_hi_hi_43, regroupV0_lo_hi_hi_lo_43};
  wire [15:0]        regroupV0_lo_hi_75 = {regroupV0_lo_hi_hi_75, regroupV0_lo_hi_lo_75};
  wire [31:0]        regroupV0_lo_75 = {regroupV0_lo_hi_75, regroupV0_lo_lo_75};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_9 = {regroupV0_hi_68[38], regroupV0_hi_68[6]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_9 = {regroupV0_hi_68[102], regroupV0_hi_68[70]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_43 = {regroupV0_hi_lo_lo_lo_hi_9, regroupV0_hi_lo_lo_lo_lo_9};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_9 = {regroupV0_hi_68[166], regroupV0_hi_68[134]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_9 = {regroupV0_hi_68[230], regroupV0_hi_68[198]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_43 = {regroupV0_hi_lo_lo_hi_hi_9, regroupV0_hi_lo_lo_hi_lo_9};
  wire [7:0]         regroupV0_hi_lo_lo_75 = {regroupV0_hi_lo_lo_hi_43, regroupV0_hi_lo_lo_lo_43};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_9 = {regroupV0_hi_68[294], regroupV0_hi_68[262]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_9 = {regroupV0_hi_68[358], regroupV0_hi_68[326]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_43 = {regroupV0_hi_lo_hi_lo_hi_9, regroupV0_hi_lo_hi_lo_lo_9};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_9 = {regroupV0_hi_68[422], regroupV0_hi_68[390]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_9 = {regroupV0_hi_68[486], regroupV0_hi_68[454]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_43 = {regroupV0_hi_lo_hi_hi_hi_9, regroupV0_hi_lo_hi_hi_lo_9};
  wire [7:0]         regroupV0_hi_lo_hi_75 = {regroupV0_hi_lo_hi_hi_43, regroupV0_hi_lo_hi_lo_43};
  wire [15:0]        regroupV0_hi_lo_75 = {regroupV0_hi_lo_hi_75, regroupV0_hi_lo_lo_75};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_9 = {regroupV0_hi_68[550], regroupV0_hi_68[518]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_9 = {regroupV0_hi_68[614], regroupV0_hi_68[582]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_43 = {regroupV0_hi_hi_lo_lo_hi_9, regroupV0_hi_hi_lo_lo_lo_9};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_9 = {regroupV0_hi_68[678], regroupV0_hi_68[646]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_9 = {regroupV0_hi_68[742], regroupV0_hi_68[710]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_43 = {regroupV0_hi_hi_lo_hi_hi_9, regroupV0_hi_hi_lo_hi_lo_9};
  wire [7:0]         regroupV0_hi_hi_lo_75 = {regroupV0_hi_hi_lo_hi_43, regroupV0_hi_hi_lo_lo_43};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_9 = {regroupV0_hi_68[806], regroupV0_hi_68[774]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_9 = {regroupV0_hi_68[870], regroupV0_hi_68[838]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_43 = {regroupV0_hi_hi_hi_lo_hi_9, regroupV0_hi_hi_hi_lo_lo_9};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_9 = {regroupV0_hi_68[934], regroupV0_hi_68[902]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_9 = {regroupV0_hi_68[998], regroupV0_hi_68[966]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_43 = {regroupV0_hi_hi_hi_hi_hi_9, regroupV0_hi_hi_hi_hi_lo_9};
  wire [7:0]         regroupV0_hi_hi_hi_75 = {regroupV0_hi_hi_hi_hi_43, regroupV0_hi_hi_hi_lo_43};
  wire [15:0]        regroupV0_hi_hi_75 = {regroupV0_hi_hi_hi_75, regroupV0_hi_hi_lo_75};
  wire [31:0]        regroupV0_hi_75 = {regroupV0_hi_hi_75, regroupV0_hi_lo_75};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_10 = {regroupV0_lo_68[39], regroupV0_lo_68[7]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_10 = {regroupV0_lo_68[103], regroupV0_lo_68[71]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_44 = {regroupV0_lo_lo_lo_lo_hi_10, regroupV0_lo_lo_lo_lo_lo_10};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_10 = {regroupV0_lo_68[167], regroupV0_lo_68[135]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_10 = {regroupV0_lo_68[231], regroupV0_lo_68[199]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_44 = {regroupV0_lo_lo_lo_hi_hi_10, regroupV0_lo_lo_lo_hi_lo_10};
  wire [7:0]         regroupV0_lo_lo_lo_76 = {regroupV0_lo_lo_lo_hi_44, regroupV0_lo_lo_lo_lo_44};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_10 = {regroupV0_lo_68[295], regroupV0_lo_68[263]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_10 = {regroupV0_lo_68[359], regroupV0_lo_68[327]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_44 = {regroupV0_lo_lo_hi_lo_hi_10, regroupV0_lo_lo_hi_lo_lo_10};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_10 = {regroupV0_lo_68[423], regroupV0_lo_68[391]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_10 = {regroupV0_lo_68[487], regroupV0_lo_68[455]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_44 = {regroupV0_lo_lo_hi_hi_hi_10, regroupV0_lo_lo_hi_hi_lo_10};
  wire [7:0]         regroupV0_lo_lo_hi_76 = {regroupV0_lo_lo_hi_hi_44, regroupV0_lo_lo_hi_lo_44};
  wire [15:0]        regroupV0_lo_lo_76 = {regroupV0_lo_lo_hi_76, regroupV0_lo_lo_lo_76};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_10 = {regroupV0_lo_68[551], regroupV0_lo_68[519]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_10 = {regroupV0_lo_68[615], regroupV0_lo_68[583]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_44 = {regroupV0_lo_hi_lo_lo_hi_10, regroupV0_lo_hi_lo_lo_lo_10};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_10 = {regroupV0_lo_68[679], regroupV0_lo_68[647]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_10 = {regroupV0_lo_68[743], regroupV0_lo_68[711]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_44 = {regroupV0_lo_hi_lo_hi_hi_10, regroupV0_lo_hi_lo_hi_lo_10};
  wire [7:0]         regroupV0_lo_hi_lo_76 = {regroupV0_lo_hi_lo_hi_44, regroupV0_lo_hi_lo_lo_44};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_10 = {regroupV0_lo_68[807], regroupV0_lo_68[775]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_10 = {regroupV0_lo_68[871], regroupV0_lo_68[839]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_44 = {regroupV0_lo_hi_hi_lo_hi_10, regroupV0_lo_hi_hi_lo_lo_10};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_10 = {regroupV0_lo_68[935], regroupV0_lo_68[903]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_10 = {regroupV0_lo_68[999], regroupV0_lo_68[967]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_44 = {regroupV0_lo_hi_hi_hi_hi_10, regroupV0_lo_hi_hi_hi_lo_10};
  wire [7:0]         regroupV0_lo_hi_hi_76 = {regroupV0_lo_hi_hi_hi_44, regroupV0_lo_hi_hi_lo_44};
  wire [15:0]        regroupV0_lo_hi_76 = {regroupV0_lo_hi_hi_76, regroupV0_lo_hi_lo_76};
  wire [31:0]        regroupV0_lo_76 = {regroupV0_lo_hi_76, regroupV0_lo_lo_76};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_10 = {regroupV0_hi_68[39], regroupV0_hi_68[7]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_10 = {regroupV0_hi_68[103], regroupV0_hi_68[71]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_44 = {regroupV0_hi_lo_lo_lo_hi_10, regroupV0_hi_lo_lo_lo_lo_10};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_10 = {regroupV0_hi_68[167], regroupV0_hi_68[135]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_10 = {regroupV0_hi_68[231], regroupV0_hi_68[199]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_44 = {regroupV0_hi_lo_lo_hi_hi_10, regroupV0_hi_lo_lo_hi_lo_10};
  wire [7:0]         regroupV0_hi_lo_lo_76 = {regroupV0_hi_lo_lo_hi_44, regroupV0_hi_lo_lo_lo_44};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_10 = {regroupV0_hi_68[295], regroupV0_hi_68[263]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_10 = {regroupV0_hi_68[359], regroupV0_hi_68[327]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_44 = {regroupV0_hi_lo_hi_lo_hi_10, regroupV0_hi_lo_hi_lo_lo_10};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_10 = {regroupV0_hi_68[423], regroupV0_hi_68[391]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_10 = {regroupV0_hi_68[487], regroupV0_hi_68[455]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_44 = {regroupV0_hi_lo_hi_hi_hi_10, regroupV0_hi_lo_hi_hi_lo_10};
  wire [7:0]         regroupV0_hi_lo_hi_76 = {regroupV0_hi_lo_hi_hi_44, regroupV0_hi_lo_hi_lo_44};
  wire [15:0]        regroupV0_hi_lo_76 = {regroupV0_hi_lo_hi_76, regroupV0_hi_lo_lo_76};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_10 = {regroupV0_hi_68[551], regroupV0_hi_68[519]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_10 = {regroupV0_hi_68[615], regroupV0_hi_68[583]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_44 = {regroupV0_hi_hi_lo_lo_hi_10, regroupV0_hi_hi_lo_lo_lo_10};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_10 = {regroupV0_hi_68[679], regroupV0_hi_68[647]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_10 = {regroupV0_hi_68[743], regroupV0_hi_68[711]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_44 = {regroupV0_hi_hi_lo_hi_hi_10, regroupV0_hi_hi_lo_hi_lo_10};
  wire [7:0]         regroupV0_hi_hi_lo_76 = {regroupV0_hi_hi_lo_hi_44, regroupV0_hi_hi_lo_lo_44};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_10 = {regroupV0_hi_68[807], regroupV0_hi_68[775]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_10 = {regroupV0_hi_68[871], regroupV0_hi_68[839]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_44 = {regroupV0_hi_hi_hi_lo_hi_10, regroupV0_hi_hi_hi_lo_lo_10};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_10 = {regroupV0_hi_68[935], regroupV0_hi_68[903]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_10 = {regroupV0_hi_68[999], regroupV0_hi_68[967]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_44 = {regroupV0_hi_hi_hi_hi_hi_10, regroupV0_hi_hi_hi_hi_lo_10};
  wire [7:0]         regroupV0_hi_hi_hi_76 = {regroupV0_hi_hi_hi_hi_44, regroupV0_hi_hi_hi_lo_44};
  wire [15:0]        regroupV0_hi_hi_76 = {regroupV0_hi_hi_hi_76, regroupV0_hi_hi_lo_76};
  wire [31:0]        regroupV0_hi_76 = {regroupV0_hi_hi_76, regroupV0_hi_lo_76};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_11 = {regroupV0_lo_68[40], regroupV0_lo_68[8]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_11 = {regroupV0_lo_68[104], regroupV0_lo_68[72]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_45 = {regroupV0_lo_lo_lo_lo_hi_11, regroupV0_lo_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_11 = {regroupV0_lo_68[168], regroupV0_lo_68[136]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_11 = {regroupV0_lo_68[232], regroupV0_lo_68[200]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_45 = {regroupV0_lo_lo_lo_hi_hi_11, regroupV0_lo_lo_lo_hi_lo_11};
  wire [7:0]         regroupV0_lo_lo_lo_77 = {regroupV0_lo_lo_lo_hi_45, regroupV0_lo_lo_lo_lo_45};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_11 = {regroupV0_lo_68[296], regroupV0_lo_68[264]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_11 = {regroupV0_lo_68[360], regroupV0_lo_68[328]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_45 = {regroupV0_lo_lo_hi_lo_hi_11, regroupV0_lo_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_11 = {regroupV0_lo_68[424], regroupV0_lo_68[392]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_11 = {regroupV0_lo_68[488], regroupV0_lo_68[456]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_45 = {regroupV0_lo_lo_hi_hi_hi_11, regroupV0_lo_lo_hi_hi_lo_11};
  wire [7:0]         regroupV0_lo_lo_hi_77 = {regroupV0_lo_lo_hi_hi_45, regroupV0_lo_lo_hi_lo_45};
  wire [15:0]        regroupV0_lo_lo_77 = {regroupV0_lo_lo_hi_77, regroupV0_lo_lo_lo_77};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_11 = {regroupV0_lo_68[552], regroupV0_lo_68[520]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_11 = {regroupV0_lo_68[616], regroupV0_lo_68[584]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_45 = {regroupV0_lo_hi_lo_lo_hi_11, regroupV0_lo_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_11 = {regroupV0_lo_68[680], regroupV0_lo_68[648]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_11 = {regroupV0_lo_68[744], regroupV0_lo_68[712]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_45 = {regroupV0_lo_hi_lo_hi_hi_11, regroupV0_lo_hi_lo_hi_lo_11};
  wire [7:0]         regroupV0_lo_hi_lo_77 = {regroupV0_lo_hi_lo_hi_45, regroupV0_lo_hi_lo_lo_45};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_11 = {regroupV0_lo_68[808], regroupV0_lo_68[776]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_11 = {regroupV0_lo_68[872], regroupV0_lo_68[840]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_45 = {regroupV0_lo_hi_hi_lo_hi_11, regroupV0_lo_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_11 = {regroupV0_lo_68[936], regroupV0_lo_68[904]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_11 = {regroupV0_lo_68[1000], regroupV0_lo_68[968]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_45 = {regroupV0_lo_hi_hi_hi_hi_11, regroupV0_lo_hi_hi_hi_lo_11};
  wire [7:0]         regroupV0_lo_hi_hi_77 = {regroupV0_lo_hi_hi_hi_45, regroupV0_lo_hi_hi_lo_45};
  wire [15:0]        regroupV0_lo_hi_77 = {regroupV0_lo_hi_hi_77, regroupV0_lo_hi_lo_77};
  wire [31:0]        regroupV0_lo_77 = {regroupV0_lo_hi_77, regroupV0_lo_lo_77};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_11 = {regroupV0_hi_68[40], regroupV0_hi_68[8]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_11 = {regroupV0_hi_68[104], regroupV0_hi_68[72]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_45 = {regroupV0_hi_lo_lo_lo_hi_11, regroupV0_hi_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_11 = {regroupV0_hi_68[168], regroupV0_hi_68[136]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_11 = {regroupV0_hi_68[232], regroupV0_hi_68[200]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_45 = {regroupV0_hi_lo_lo_hi_hi_11, regroupV0_hi_lo_lo_hi_lo_11};
  wire [7:0]         regroupV0_hi_lo_lo_77 = {regroupV0_hi_lo_lo_hi_45, regroupV0_hi_lo_lo_lo_45};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_11 = {regroupV0_hi_68[296], regroupV0_hi_68[264]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_11 = {regroupV0_hi_68[360], regroupV0_hi_68[328]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_45 = {regroupV0_hi_lo_hi_lo_hi_11, regroupV0_hi_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_11 = {regroupV0_hi_68[424], regroupV0_hi_68[392]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_11 = {regroupV0_hi_68[488], regroupV0_hi_68[456]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_45 = {regroupV0_hi_lo_hi_hi_hi_11, regroupV0_hi_lo_hi_hi_lo_11};
  wire [7:0]         regroupV0_hi_lo_hi_77 = {regroupV0_hi_lo_hi_hi_45, regroupV0_hi_lo_hi_lo_45};
  wire [15:0]        regroupV0_hi_lo_77 = {regroupV0_hi_lo_hi_77, regroupV0_hi_lo_lo_77};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_11 = {regroupV0_hi_68[552], regroupV0_hi_68[520]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_11 = {regroupV0_hi_68[616], regroupV0_hi_68[584]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_45 = {regroupV0_hi_hi_lo_lo_hi_11, regroupV0_hi_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_11 = {regroupV0_hi_68[680], regroupV0_hi_68[648]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_11 = {regroupV0_hi_68[744], regroupV0_hi_68[712]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_45 = {regroupV0_hi_hi_lo_hi_hi_11, regroupV0_hi_hi_lo_hi_lo_11};
  wire [7:0]         regroupV0_hi_hi_lo_77 = {regroupV0_hi_hi_lo_hi_45, regroupV0_hi_hi_lo_lo_45};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_11 = {regroupV0_hi_68[808], regroupV0_hi_68[776]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_11 = {regroupV0_hi_68[872], regroupV0_hi_68[840]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_45 = {regroupV0_hi_hi_hi_lo_hi_11, regroupV0_hi_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_11 = {regroupV0_hi_68[936], regroupV0_hi_68[904]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_11 = {regroupV0_hi_68[1000], regroupV0_hi_68[968]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_45 = {regroupV0_hi_hi_hi_hi_hi_11, regroupV0_hi_hi_hi_hi_lo_11};
  wire [7:0]         regroupV0_hi_hi_hi_77 = {regroupV0_hi_hi_hi_hi_45, regroupV0_hi_hi_hi_lo_45};
  wire [15:0]        regroupV0_hi_hi_77 = {regroupV0_hi_hi_hi_77, regroupV0_hi_hi_lo_77};
  wire [31:0]        regroupV0_hi_77 = {regroupV0_hi_hi_77, regroupV0_hi_lo_77};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_12 = {regroupV0_lo_68[41], regroupV0_lo_68[9]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_12 = {regroupV0_lo_68[105], regroupV0_lo_68[73]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_46 = {regroupV0_lo_lo_lo_lo_hi_12, regroupV0_lo_lo_lo_lo_lo_12};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_12 = {regroupV0_lo_68[169], regroupV0_lo_68[137]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_12 = {regroupV0_lo_68[233], regroupV0_lo_68[201]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_46 = {regroupV0_lo_lo_lo_hi_hi_12, regroupV0_lo_lo_lo_hi_lo_12};
  wire [7:0]         regroupV0_lo_lo_lo_78 = {regroupV0_lo_lo_lo_hi_46, regroupV0_lo_lo_lo_lo_46};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_12 = {regroupV0_lo_68[297], regroupV0_lo_68[265]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_12 = {regroupV0_lo_68[361], regroupV0_lo_68[329]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_46 = {regroupV0_lo_lo_hi_lo_hi_12, regroupV0_lo_lo_hi_lo_lo_12};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_12 = {regroupV0_lo_68[425], regroupV0_lo_68[393]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_12 = {regroupV0_lo_68[489], regroupV0_lo_68[457]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_46 = {regroupV0_lo_lo_hi_hi_hi_12, regroupV0_lo_lo_hi_hi_lo_12};
  wire [7:0]         regroupV0_lo_lo_hi_78 = {regroupV0_lo_lo_hi_hi_46, regroupV0_lo_lo_hi_lo_46};
  wire [15:0]        regroupV0_lo_lo_78 = {regroupV0_lo_lo_hi_78, regroupV0_lo_lo_lo_78};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_12 = {regroupV0_lo_68[553], regroupV0_lo_68[521]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_12 = {regroupV0_lo_68[617], regroupV0_lo_68[585]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_46 = {regroupV0_lo_hi_lo_lo_hi_12, regroupV0_lo_hi_lo_lo_lo_12};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_12 = {regroupV0_lo_68[681], regroupV0_lo_68[649]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_12 = {regroupV0_lo_68[745], regroupV0_lo_68[713]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_46 = {regroupV0_lo_hi_lo_hi_hi_12, regroupV0_lo_hi_lo_hi_lo_12};
  wire [7:0]         regroupV0_lo_hi_lo_78 = {regroupV0_lo_hi_lo_hi_46, regroupV0_lo_hi_lo_lo_46};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_12 = {regroupV0_lo_68[809], regroupV0_lo_68[777]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_12 = {regroupV0_lo_68[873], regroupV0_lo_68[841]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_46 = {regroupV0_lo_hi_hi_lo_hi_12, regroupV0_lo_hi_hi_lo_lo_12};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_12 = {regroupV0_lo_68[937], regroupV0_lo_68[905]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_12 = {regroupV0_lo_68[1001], regroupV0_lo_68[969]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_46 = {regroupV0_lo_hi_hi_hi_hi_12, regroupV0_lo_hi_hi_hi_lo_12};
  wire [7:0]         regroupV0_lo_hi_hi_78 = {regroupV0_lo_hi_hi_hi_46, regroupV0_lo_hi_hi_lo_46};
  wire [15:0]        regroupV0_lo_hi_78 = {regroupV0_lo_hi_hi_78, regroupV0_lo_hi_lo_78};
  wire [31:0]        regroupV0_lo_78 = {regroupV0_lo_hi_78, regroupV0_lo_lo_78};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_12 = {regroupV0_hi_68[41], regroupV0_hi_68[9]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_12 = {regroupV0_hi_68[105], regroupV0_hi_68[73]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_46 = {regroupV0_hi_lo_lo_lo_hi_12, regroupV0_hi_lo_lo_lo_lo_12};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_12 = {regroupV0_hi_68[169], regroupV0_hi_68[137]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_12 = {regroupV0_hi_68[233], regroupV0_hi_68[201]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_46 = {regroupV0_hi_lo_lo_hi_hi_12, regroupV0_hi_lo_lo_hi_lo_12};
  wire [7:0]         regroupV0_hi_lo_lo_78 = {regroupV0_hi_lo_lo_hi_46, regroupV0_hi_lo_lo_lo_46};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_12 = {regroupV0_hi_68[297], regroupV0_hi_68[265]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_12 = {regroupV0_hi_68[361], regroupV0_hi_68[329]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_46 = {regroupV0_hi_lo_hi_lo_hi_12, regroupV0_hi_lo_hi_lo_lo_12};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_12 = {regroupV0_hi_68[425], regroupV0_hi_68[393]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_12 = {regroupV0_hi_68[489], regroupV0_hi_68[457]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_46 = {regroupV0_hi_lo_hi_hi_hi_12, regroupV0_hi_lo_hi_hi_lo_12};
  wire [7:0]         regroupV0_hi_lo_hi_78 = {regroupV0_hi_lo_hi_hi_46, regroupV0_hi_lo_hi_lo_46};
  wire [15:0]        regroupV0_hi_lo_78 = {regroupV0_hi_lo_hi_78, regroupV0_hi_lo_lo_78};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_12 = {regroupV0_hi_68[553], regroupV0_hi_68[521]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_12 = {regroupV0_hi_68[617], regroupV0_hi_68[585]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_46 = {regroupV0_hi_hi_lo_lo_hi_12, regroupV0_hi_hi_lo_lo_lo_12};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_12 = {regroupV0_hi_68[681], regroupV0_hi_68[649]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_12 = {regroupV0_hi_68[745], regroupV0_hi_68[713]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_46 = {regroupV0_hi_hi_lo_hi_hi_12, regroupV0_hi_hi_lo_hi_lo_12};
  wire [7:0]         regroupV0_hi_hi_lo_78 = {regroupV0_hi_hi_lo_hi_46, regroupV0_hi_hi_lo_lo_46};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_12 = {regroupV0_hi_68[809], regroupV0_hi_68[777]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_12 = {regroupV0_hi_68[873], regroupV0_hi_68[841]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_46 = {regroupV0_hi_hi_hi_lo_hi_12, regroupV0_hi_hi_hi_lo_lo_12};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_12 = {regroupV0_hi_68[937], regroupV0_hi_68[905]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_12 = {regroupV0_hi_68[1001], regroupV0_hi_68[969]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_46 = {regroupV0_hi_hi_hi_hi_hi_12, regroupV0_hi_hi_hi_hi_lo_12};
  wire [7:0]         regroupV0_hi_hi_hi_78 = {regroupV0_hi_hi_hi_hi_46, regroupV0_hi_hi_hi_lo_46};
  wire [15:0]        regroupV0_hi_hi_78 = {regroupV0_hi_hi_hi_78, regroupV0_hi_hi_lo_78};
  wire [31:0]        regroupV0_hi_78 = {regroupV0_hi_hi_78, regroupV0_hi_lo_78};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_13 = {regroupV0_lo_68[42], regroupV0_lo_68[10]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_13 = {regroupV0_lo_68[106], regroupV0_lo_68[74]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_47 = {regroupV0_lo_lo_lo_lo_hi_13, regroupV0_lo_lo_lo_lo_lo_13};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_13 = {regroupV0_lo_68[170], regroupV0_lo_68[138]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_13 = {regroupV0_lo_68[234], regroupV0_lo_68[202]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_47 = {regroupV0_lo_lo_lo_hi_hi_13, regroupV0_lo_lo_lo_hi_lo_13};
  wire [7:0]         regroupV0_lo_lo_lo_79 = {regroupV0_lo_lo_lo_hi_47, regroupV0_lo_lo_lo_lo_47};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_13 = {regroupV0_lo_68[298], regroupV0_lo_68[266]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_13 = {regroupV0_lo_68[362], regroupV0_lo_68[330]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_47 = {regroupV0_lo_lo_hi_lo_hi_13, regroupV0_lo_lo_hi_lo_lo_13};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_13 = {regroupV0_lo_68[426], regroupV0_lo_68[394]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_13 = {regroupV0_lo_68[490], regroupV0_lo_68[458]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_47 = {regroupV0_lo_lo_hi_hi_hi_13, regroupV0_lo_lo_hi_hi_lo_13};
  wire [7:0]         regroupV0_lo_lo_hi_79 = {regroupV0_lo_lo_hi_hi_47, regroupV0_lo_lo_hi_lo_47};
  wire [15:0]        regroupV0_lo_lo_79 = {regroupV0_lo_lo_hi_79, regroupV0_lo_lo_lo_79};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_13 = {regroupV0_lo_68[554], regroupV0_lo_68[522]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_13 = {regroupV0_lo_68[618], regroupV0_lo_68[586]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_47 = {regroupV0_lo_hi_lo_lo_hi_13, regroupV0_lo_hi_lo_lo_lo_13};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_13 = {regroupV0_lo_68[682], regroupV0_lo_68[650]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_13 = {regroupV0_lo_68[746], regroupV0_lo_68[714]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_47 = {regroupV0_lo_hi_lo_hi_hi_13, regroupV0_lo_hi_lo_hi_lo_13};
  wire [7:0]         regroupV0_lo_hi_lo_79 = {regroupV0_lo_hi_lo_hi_47, regroupV0_lo_hi_lo_lo_47};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_13 = {regroupV0_lo_68[810], regroupV0_lo_68[778]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_13 = {regroupV0_lo_68[874], regroupV0_lo_68[842]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_47 = {regroupV0_lo_hi_hi_lo_hi_13, regroupV0_lo_hi_hi_lo_lo_13};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_13 = {regroupV0_lo_68[938], regroupV0_lo_68[906]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_13 = {regroupV0_lo_68[1002], regroupV0_lo_68[970]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_47 = {regroupV0_lo_hi_hi_hi_hi_13, regroupV0_lo_hi_hi_hi_lo_13};
  wire [7:0]         regroupV0_lo_hi_hi_79 = {regroupV0_lo_hi_hi_hi_47, regroupV0_lo_hi_hi_lo_47};
  wire [15:0]        regroupV0_lo_hi_79 = {regroupV0_lo_hi_hi_79, regroupV0_lo_hi_lo_79};
  wire [31:0]        regroupV0_lo_79 = {regroupV0_lo_hi_79, regroupV0_lo_lo_79};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_13 = {regroupV0_hi_68[42], regroupV0_hi_68[10]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_13 = {regroupV0_hi_68[106], regroupV0_hi_68[74]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_47 = {regroupV0_hi_lo_lo_lo_hi_13, regroupV0_hi_lo_lo_lo_lo_13};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_13 = {regroupV0_hi_68[170], regroupV0_hi_68[138]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_13 = {regroupV0_hi_68[234], regroupV0_hi_68[202]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_47 = {regroupV0_hi_lo_lo_hi_hi_13, regroupV0_hi_lo_lo_hi_lo_13};
  wire [7:0]         regroupV0_hi_lo_lo_79 = {regroupV0_hi_lo_lo_hi_47, regroupV0_hi_lo_lo_lo_47};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_13 = {regroupV0_hi_68[298], regroupV0_hi_68[266]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_13 = {regroupV0_hi_68[362], regroupV0_hi_68[330]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_47 = {regroupV0_hi_lo_hi_lo_hi_13, regroupV0_hi_lo_hi_lo_lo_13};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_13 = {regroupV0_hi_68[426], regroupV0_hi_68[394]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_13 = {regroupV0_hi_68[490], regroupV0_hi_68[458]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_47 = {regroupV0_hi_lo_hi_hi_hi_13, regroupV0_hi_lo_hi_hi_lo_13};
  wire [7:0]         regroupV0_hi_lo_hi_79 = {regroupV0_hi_lo_hi_hi_47, regroupV0_hi_lo_hi_lo_47};
  wire [15:0]        regroupV0_hi_lo_79 = {regroupV0_hi_lo_hi_79, regroupV0_hi_lo_lo_79};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_13 = {regroupV0_hi_68[554], regroupV0_hi_68[522]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_13 = {regroupV0_hi_68[618], regroupV0_hi_68[586]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_47 = {regroupV0_hi_hi_lo_lo_hi_13, regroupV0_hi_hi_lo_lo_lo_13};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_13 = {regroupV0_hi_68[682], regroupV0_hi_68[650]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_13 = {regroupV0_hi_68[746], regroupV0_hi_68[714]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_47 = {regroupV0_hi_hi_lo_hi_hi_13, regroupV0_hi_hi_lo_hi_lo_13};
  wire [7:0]         regroupV0_hi_hi_lo_79 = {regroupV0_hi_hi_lo_hi_47, regroupV0_hi_hi_lo_lo_47};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_13 = {regroupV0_hi_68[810], regroupV0_hi_68[778]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_13 = {regroupV0_hi_68[874], regroupV0_hi_68[842]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_47 = {regroupV0_hi_hi_hi_lo_hi_13, regroupV0_hi_hi_hi_lo_lo_13};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_13 = {regroupV0_hi_68[938], regroupV0_hi_68[906]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_13 = {regroupV0_hi_68[1002], regroupV0_hi_68[970]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_47 = {regroupV0_hi_hi_hi_hi_hi_13, regroupV0_hi_hi_hi_hi_lo_13};
  wire [7:0]         regroupV0_hi_hi_hi_79 = {regroupV0_hi_hi_hi_hi_47, regroupV0_hi_hi_hi_lo_47};
  wire [15:0]        regroupV0_hi_hi_79 = {regroupV0_hi_hi_hi_79, regroupV0_hi_hi_lo_79};
  wire [31:0]        regroupV0_hi_79 = {regroupV0_hi_hi_79, regroupV0_hi_lo_79};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_14 = {regroupV0_lo_68[43], regroupV0_lo_68[11]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_14 = {regroupV0_lo_68[107], regroupV0_lo_68[75]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_48 = {regroupV0_lo_lo_lo_lo_hi_14, regroupV0_lo_lo_lo_lo_lo_14};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_14 = {regroupV0_lo_68[171], regroupV0_lo_68[139]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_14 = {regroupV0_lo_68[235], regroupV0_lo_68[203]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_48 = {regroupV0_lo_lo_lo_hi_hi_14, regroupV0_lo_lo_lo_hi_lo_14};
  wire [7:0]         regroupV0_lo_lo_lo_80 = {regroupV0_lo_lo_lo_hi_48, regroupV0_lo_lo_lo_lo_48};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_14 = {regroupV0_lo_68[299], regroupV0_lo_68[267]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_14 = {regroupV0_lo_68[363], regroupV0_lo_68[331]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_48 = {regroupV0_lo_lo_hi_lo_hi_14, regroupV0_lo_lo_hi_lo_lo_14};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_14 = {regroupV0_lo_68[427], regroupV0_lo_68[395]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_14 = {regroupV0_lo_68[491], regroupV0_lo_68[459]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_48 = {regroupV0_lo_lo_hi_hi_hi_14, regroupV0_lo_lo_hi_hi_lo_14};
  wire [7:0]         regroupV0_lo_lo_hi_80 = {regroupV0_lo_lo_hi_hi_48, regroupV0_lo_lo_hi_lo_48};
  wire [15:0]        regroupV0_lo_lo_80 = {regroupV0_lo_lo_hi_80, regroupV0_lo_lo_lo_80};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_14 = {regroupV0_lo_68[555], regroupV0_lo_68[523]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_14 = {regroupV0_lo_68[619], regroupV0_lo_68[587]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_48 = {regroupV0_lo_hi_lo_lo_hi_14, regroupV0_lo_hi_lo_lo_lo_14};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_14 = {regroupV0_lo_68[683], regroupV0_lo_68[651]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_14 = {regroupV0_lo_68[747], regroupV0_lo_68[715]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_48 = {regroupV0_lo_hi_lo_hi_hi_14, regroupV0_lo_hi_lo_hi_lo_14};
  wire [7:0]         regroupV0_lo_hi_lo_80 = {regroupV0_lo_hi_lo_hi_48, regroupV0_lo_hi_lo_lo_48};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_14 = {regroupV0_lo_68[811], regroupV0_lo_68[779]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_14 = {regroupV0_lo_68[875], regroupV0_lo_68[843]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_48 = {regroupV0_lo_hi_hi_lo_hi_14, regroupV0_lo_hi_hi_lo_lo_14};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_14 = {regroupV0_lo_68[939], regroupV0_lo_68[907]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_14 = {regroupV0_lo_68[1003], regroupV0_lo_68[971]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_48 = {regroupV0_lo_hi_hi_hi_hi_14, regroupV0_lo_hi_hi_hi_lo_14};
  wire [7:0]         regroupV0_lo_hi_hi_80 = {regroupV0_lo_hi_hi_hi_48, regroupV0_lo_hi_hi_lo_48};
  wire [15:0]        regroupV0_lo_hi_80 = {regroupV0_lo_hi_hi_80, regroupV0_lo_hi_lo_80};
  wire [31:0]        regroupV0_lo_80 = {regroupV0_lo_hi_80, regroupV0_lo_lo_80};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_14 = {regroupV0_hi_68[43], regroupV0_hi_68[11]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_14 = {regroupV0_hi_68[107], regroupV0_hi_68[75]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_48 = {regroupV0_hi_lo_lo_lo_hi_14, regroupV0_hi_lo_lo_lo_lo_14};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_14 = {regroupV0_hi_68[171], regroupV0_hi_68[139]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_14 = {regroupV0_hi_68[235], regroupV0_hi_68[203]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_48 = {regroupV0_hi_lo_lo_hi_hi_14, regroupV0_hi_lo_lo_hi_lo_14};
  wire [7:0]         regroupV0_hi_lo_lo_80 = {regroupV0_hi_lo_lo_hi_48, regroupV0_hi_lo_lo_lo_48};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_14 = {regroupV0_hi_68[299], regroupV0_hi_68[267]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_14 = {regroupV0_hi_68[363], regroupV0_hi_68[331]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_48 = {regroupV0_hi_lo_hi_lo_hi_14, regroupV0_hi_lo_hi_lo_lo_14};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_14 = {regroupV0_hi_68[427], regroupV0_hi_68[395]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_14 = {regroupV0_hi_68[491], regroupV0_hi_68[459]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_48 = {regroupV0_hi_lo_hi_hi_hi_14, regroupV0_hi_lo_hi_hi_lo_14};
  wire [7:0]         regroupV0_hi_lo_hi_80 = {regroupV0_hi_lo_hi_hi_48, regroupV0_hi_lo_hi_lo_48};
  wire [15:0]        regroupV0_hi_lo_80 = {regroupV0_hi_lo_hi_80, regroupV0_hi_lo_lo_80};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_14 = {regroupV0_hi_68[555], regroupV0_hi_68[523]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_14 = {regroupV0_hi_68[619], regroupV0_hi_68[587]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_48 = {regroupV0_hi_hi_lo_lo_hi_14, regroupV0_hi_hi_lo_lo_lo_14};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_14 = {regroupV0_hi_68[683], regroupV0_hi_68[651]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_14 = {regroupV0_hi_68[747], regroupV0_hi_68[715]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_48 = {regroupV0_hi_hi_lo_hi_hi_14, regroupV0_hi_hi_lo_hi_lo_14};
  wire [7:0]         regroupV0_hi_hi_lo_80 = {regroupV0_hi_hi_lo_hi_48, regroupV0_hi_hi_lo_lo_48};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_14 = {regroupV0_hi_68[811], regroupV0_hi_68[779]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_14 = {regroupV0_hi_68[875], regroupV0_hi_68[843]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_48 = {regroupV0_hi_hi_hi_lo_hi_14, regroupV0_hi_hi_hi_lo_lo_14};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_14 = {regroupV0_hi_68[939], regroupV0_hi_68[907]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_14 = {regroupV0_hi_68[1003], regroupV0_hi_68[971]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_48 = {regroupV0_hi_hi_hi_hi_hi_14, regroupV0_hi_hi_hi_hi_lo_14};
  wire [7:0]         regroupV0_hi_hi_hi_80 = {regroupV0_hi_hi_hi_hi_48, regroupV0_hi_hi_hi_lo_48};
  wire [15:0]        regroupV0_hi_hi_80 = {regroupV0_hi_hi_hi_80, regroupV0_hi_hi_lo_80};
  wire [31:0]        regroupV0_hi_80 = {regroupV0_hi_hi_80, regroupV0_hi_lo_80};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_15 = {regroupV0_lo_68[44], regroupV0_lo_68[12]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_15 = {regroupV0_lo_68[108], regroupV0_lo_68[76]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_49 = {regroupV0_lo_lo_lo_lo_hi_15, regroupV0_lo_lo_lo_lo_lo_15};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_15 = {regroupV0_lo_68[172], regroupV0_lo_68[140]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_15 = {regroupV0_lo_68[236], regroupV0_lo_68[204]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_49 = {regroupV0_lo_lo_lo_hi_hi_15, regroupV0_lo_lo_lo_hi_lo_15};
  wire [7:0]         regroupV0_lo_lo_lo_81 = {regroupV0_lo_lo_lo_hi_49, regroupV0_lo_lo_lo_lo_49};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_15 = {regroupV0_lo_68[300], regroupV0_lo_68[268]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_15 = {regroupV0_lo_68[364], regroupV0_lo_68[332]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_49 = {regroupV0_lo_lo_hi_lo_hi_15, regroupV0_lo_lo_hi_lo_lo_15};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_15 = {regroupV0_lo_68[428], regroupV0_lo_68[396]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_15 = {regroupV0_lo_68[492], regroupV0_lo_68[460]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_49 = {regroupV0_lo_lo_hi_hi_hi_15, regroupV0_lo_lo_hi_hi_lo_15};
  wire [7:0]         regroupV0_lo_lo_hi_81 = {regroupV0_lo_lo_hi_hi_49, regroupV0_lo_lo_hi_lo_49};
  wire [15:0]        regroupV0_lo_lo_81 = {regroupV0_lo_lo_hi_81, regroupV0_lo_lo_lo_81};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_15 = {regroupV0_lo_68[556], regroupV0_lo_68[524]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_15 = {regroupV0_lo_68[620], regroupV0_lo_68[588]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_49 = {regroupV0_lo_hi_lo_lo_hi_15, regroupV0_lo_hi_lo_lo_lo_15};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_15 = {regroupV0_lo_68[684], regroupV0_lo_68[652]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_15 = {regroupV0_lo_68[748], regroupV0_lo_68[716]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_49 = {regroupV0_lo_hi_lo_hi_hi_15, regroupV0_lo_hi_lo_hi_lo_15};
  wire [7:0]         regroupV0_lo_hi_lo_81 = {regroupV0_lo_hi_lo_hi_49, regroupV0_lo_hi_lo_lo_49};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_15 = {regroupV0_lo_68[812], regroupV0_lo_68[780]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_15 = {regroupV0_lo_68[876], regroupV0_lo_68[844]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_49 = {regroupV0_lo_hi_hi_lo_hi_15, regroupV0_lo_hi_hi_lo_lo_15};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_15 = {regroupV0_lo_68[940], regroupV0_lo_68[908]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_15 = {regroupV0_lo_68[1004], regroupV0_lo_68[972]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_49 = {regroupV0_lo_hi_hi_hi_hi_15, regroupV0_lo_hi_hi_hi_lo_15};
  wire [7:0]         regroupV0_lo_hi_hi_81 = {regroupV0_lo_hi_hi_hi_49, regroupV0_lo_hi_hi_lo_49};
  wire [15:0]        regroupV0_lo_hi_81 = {regroupV0_lo_hi_hi_81, regroupV0_lo_hi_lo_81};
  wire [31:0]        regroupV0_lo_81 = {regroupV0_lo_hi_81, regroupV0_lo_lo_81};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_15 = {regroupV0_hi_68[44], regroupV0_hi_68[12]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_15 = {regroupV0_hi_68[108], regroupV0_hi_68[76]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_49 = {regroupV0_hi_lo_lo_lo_hi_15, regroupV0_hi_lo_lo_lo_lo_15};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_15 = {regroupV0_hi_68[172], regroupV0_hi_68[140]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_15 = {regroupV0_hi_68[236], regroupV0_hi_68[204]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_49 = {regroupV0_hi_lo_lo_hi_hi_15, regroupV0_hi_lo_lo_hi_lo_15};
  wire [7:0]         regroupV0_hi_lo_lo_81 = {regroupV0_hi_lo_lo_hi_49, regroupV0_hi_lo_lo_lo_49};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_15 = {regroupV0_hi_68[300], regroupV0_hi_68[268]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_15 = {regroupV0_hi_68[364], regroupV0_hi_68[332]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_49 = {regroupV0_hi_lo_hi_lo_hi_15, regroupV0_hi_lo_hi_lo_lo_15};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_15 = {regroupV0_hi_68[428], regroupV0_hi_68[396]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_15 = {regroupV0_hi_68[492], regroupV0_hi_68[460]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_49 = {regroupV0_hi_lo_hi_hi_hi_15, regroupV0_hi_lo_hi_hi_lo_15};
  wire [7:0]         regroupV0_hi_lo_hi_81 = {regroupV0_hi_lo_hi_hi_49, regroupV0_hi_lo_hi_lo_49};
  wire [15:0]        regroupV0_hi_lo_81 = {regroupV0_hi_lo_hi_81, regroupV0_hi_lo_lo_81};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_15 = {regroupV0_hi_68[556], regroupV0_hi_68[524]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_15 = {regroupV0_hi_68[620], regroupV0_hi_68[588]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_49 = {regroupV0_hi_hi_lo_lo_hi_15, regroupV0_hi_hi_lo_lo_lo_15};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_15 = {regroupV0_hi_68[684], regroupV0_hi_68[652]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_15 = {regroupV0_hi_68[748], regroupV0_hi_68[716]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_49 = {regroupV0_hi_hi_lo_hi_hi_15, regroupV0_hi_hi_lo_hi_lo_15};
  wire [7:0]         regroupV0_hi_hi_lo_81 = {regroupV0_hi_hi_lo_hi_49, regroupV0_hi_hi_lo_lo_49};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_15 = {regroupV0_hi_68[812], regroupV0_hi_68[780]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_15 = {regroupV0_hi_68[876], regroupV0_hi_68[844]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_49 = {regroupV0_hi_hi_hi_lo_hi_15, regroupV0_hi_hi_hi_lo_lo_15};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_15 = {regroupV0_hi_68[940], regroupV0_hi_68[908]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_15 = {regroupV0_hi_68[1004], regroupV0_hi_68[972]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_49 = {regroupV0_hi_hi_hi_hi_hi_15, regroupV0_hi_hi_hi_hi_lo_15};
  wire [7:0]         regroupV0_hi_hi_hi_81 = {regroupV0_hi_hi_hi_hi_49, regroupV0_hi_hi_hi_lo_49};
  wire [15:0]        regroupV0_hi_hi_81 = {regroupV0_hi_hi_hi_81, regroupV0_hi_hi_lo_81};
  wire [31:0]        regroupV0_hi_81 = {regroupV0_hi_hi_81, regroupV0_hi_lo_81};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_16 = {regroupV0_lo_68[45], regroupV0_lo_68[13]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_16 = {regroupV0_lo_68[109], regroupV0_lo_68[77]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_50 = {regroupV0_lo_lo_lo_lo_hi_16, regroupV0_lo_lo_lo_lo_lo_16};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_16 = {regroupV0_lo_68[173], regroupV0_lo_68[141]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_16 = {regroupV0_lo_68[237], regroupV0_lo_68[205]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_50 = {regroupV0_lo_lo_lo_hi_hi_16, regroupV0_lo_lo_lo_hi_lo_16};
  wire [7:0]         regroupV0_lo_lo_lo_82 = {regroupV0_lo_lo_lo_hi_50, regroupV0_lo_lo_lo_lo_50};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_16 = {regroupV0_lo_68[301], regroupV0_lo_68[269]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_16 = {regroupV0_lo_68[365], regroupV0_lo_68[333]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_50 = {regroupV0_lo_lo_hi_lo_hi_16, regroupV0_lo_lo_hi_lo_lo_16};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_16 = {regroupV0_lo_68[429], regroupV0_lo_68[397]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_16 = {regroupV0_lo_68[493], regroupV0_lo_68[461]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_50 = {regroupV0_lo_lo_hi_hi_hi_16, regroupV0_lo_lo_hi_hi_lo_16};
  wire [7:0]         regroupV0_lo_lo_hi_82 = {regroupV0_lo_lo_hi_hi_50, regroupV0_lo_lo_hi_lo_50};
  wire [15:0]        regroupV0_lo_lo_82 = {regroupV0_lo_lo_hi_82, regroupV0_lo_lo_lo_82};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_16 = {regroupV0_lo_68[557], regroupV0_lo_68[525]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_16 = {regroupV0_lo_68[621], regroupV0_lo_68[589]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_50 = {regroupV0_lo_hi_lo_lo_hi_16, regroupV0_lo_hi_lo_lo_lo_16};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_16 = {regroupV0_lo_68[685], regroupV0_lo_68[653]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_16 = {regroupV0_lo_68[749], regroupV0_lo_68[717]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_50 = {regroupV0_lo_hi_lo_hi_hi_16, regroupV0_lo_hi_lo_hi_lo_16};
  wire [7:0]         regroupV0_lo_hi_lo_82 = {regroupV0_lo_hi_lo_hi_50, regroupV0_lo_hi_lo_lo_50};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_16 = {regroupV0_lo_68[813], regroupV0_lo_68[781]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_16 = {regroupV0_lo_68[877], regroupV0_lo_68[845]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_50 = {regroupV0_lo_hi_hi_lo_hi_16, regroupV0_lo_hi_hi_lo_lo_16};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_16 = {regroupV0_lo_68[941], regroupV0_lo_68[909]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_16 = {regroupV0_lo_68[1005], regroupV0_lo_68[973]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_50 = {regroupV0_lo_hi_hi_hi_hi_16, regroupV0_lo_hi_hi_hi_lo_16};
  wire [7:0]         regroupV0_lo_hi_hi_82 = {regroupV0_lo_hi_hi_hi_50, regroupV0_lo_hi_hi_lo_50};
  wire [15:0]        regroupV0_lo_hi_82 = {regroupV0_lo_hi_hi_82, regroupV0_lo_hi_lo_82};
  wire [31:0]        regroupV0_lo_82 = {regroupV0_lo_hi_82, regroupV0_lo_lo_82};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_16 = {regroupV0_hi_68[45], regroupV0_hi_68[13]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_16 = {regroupV0_hi_68[109], regroupV0_hi_68[77]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_50 = {regroupV0_hi_lo_lo_lo_hi_16, regroupV0_hi_lo_lo_lo_lo_16};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_16 = {regroupV0_hi_68[173], regroupV0_hi_68[141]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_16 = {regroupV0_hi_68[237], regroupV0_hi_68[205]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_50 = {regroupV0_hi_lo_lo_hi_hi_16, regroupV0_hi_lo_lo_hi_lo_16};
  wire [7:0]         regroupV0_hi_lo_lo_82 = {regroupV0_hi_lo_lo_hi_50, regroupV0_hi_lo_lo_lo_50};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_16 = {regroupV0_hi_68[301], regroupV0_hi_68[269]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_16 = {regroupV0_hi_68[365], regroupV0_hi_68[333]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_50 = {regroupV0_hi_lo_hi_lo_hi_16, regroupV0_hi_lo_hi_lo_lo_16};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_16 = {regroupV0_hi_68[429], regroupV0_hi_68[397]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_16 = {regroupV0_hi_68[493], regroupV0_hi_68[461]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_50 = {regroupV0_hi_lo_hi_hi_hi_16, regroupV0_hi_lo_hi_hi_lo_16};
  wire [7:0]         regroupV0_hi_lo_hi_82 = {regroupV0_hi_lo_hi_hi_50, regroupV0_hi_lo_hi_lo_50};
  wire [15:0]        regroupV0_hi_lo_82 = {regroupV0_hi_lo_hi_82, regroupV0_hi_lo_lo_82};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_16 = {regroupV0_hi_68[557], regroupV0_hi_68[525]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_16 = {regroupV0_hi_68[621], regroupV0_hi_68[589]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_50 = {regroupV0_hi_hi_lo_lo_hi_16, regroupV0_hi_hi_lo_lo_lo_16};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_16 = {regroupV0_hi_68[685], regroupV0_hi_68[653]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_16 = {regroupV0_hi_68[749], regroupV0_hi_68[717]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_50 = {regroupV0_hi_hi_lo_hi_hi_16, regroupV0_hi_hi_lo_hi_lo_16};
  wire [7:0]         regroupV0_hi_hi_lo_82 = {regroupV0_hi_hi_lo_hi_50, regroupV0_hi_hi_lo_lo_50};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_16 = {regroupV0_hi_68[813], regroupV0_hi_68[781]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_16 = {regroupV0_hi_68[877], regroupV0_hi_68[845]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_50 = {regroupV0_hi_hi_hi_lo_hi_16, regroupV0_hi_hi_hi_lo_lo_16};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_16 = {regroupV0_hi_68[941], regroupV0_hi_68[909]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_16 = {regroupV0_hi_68[1005], regroupV0_hi_68[973]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_50 = {regroupV0_hi_hi_hi_hi_hi_16, regroupV0_hi_hi_hi_hi_lo_16};
  wire [7:0]         regroupV0_hi_hi_hi_82 = {regroupV0_hi_hi_hi_hi_50, regroupV0_hi_hi_hi_lo_50};
  wire [15:0]        regroupV0_hi_hi_82 = {regroupV0_hi_hi_hi_82, regroupV0_hi_hi_lo_82};
  wire [31:0]        regroupV0_hi_82 = {regroupV0_hi_hi_82, regroupV0_hi_lo_82};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_17 = {regroupV0_lo_68[46], regroupV0_lo_68[14]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_17 = {regroupV0_lo_68[110], regroupV0_lo_68[78]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_51 = {regroupV0_lo_lo_lo_lo_hi_17, regroupV0_lo_lo_lo_lo_lo_17};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_17 = {regroupV0_lo_68[174], regroupV0_lo_68[142]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_17 = {regroupV0_lo_68[238], regroupV0_lo_68[206]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_51 = {regroupV0_lo_lo_lo_hi_hi_17, regroupV0_lo_lo_lo_hi_lo_17};
  wire [7:0]         regroupV0_lo_lo_lo_83 = {regroupV0_lo_lo_lo_hi_51, regroupV0_lo_lo_lo_lo_51};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_17 = {regroupV0_lo_68[302], regroupV0_lo_68[270]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_17 = {regroupV0_lo_68[366], regroupV0_lo_68[334]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_51 = {regroupV0_lo_lo_hi_lo_hi_17, regroupV0_lo_lo_hi_lo_lo_17};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_17 = {regroupV0_lo_68[430], regroupV0_lo_68[398]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_17 = {regroupV0_lo_68[494], regroupV0_lo_68[462]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_51 = {regroupV0_lo_lo_hi_hi_hi_17, regroupV0_lo_lo_hi_hi_lo_17};
  wire [7:0]         regroupV0_lo_lo_hi_83 = {regroupV0_lo_lo_hi_hi_51, regroupV0_lo_lo_hi_lo_51};
  wire [15:0]        regroupV0_lo_lo_83 = {regroupV0_lo_lo_hi_83, regroupV0_lo_lo_lo_83};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_17 = {regroupV0_lo_68[558], regroupV0_lo_68[526]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_17 = {regroupV0_lo_68[622], regroupV0_lo_68[590]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_51 = {regroupV0_lo_hi_lo_lo_hi_17, regroupV0_lo_hi_lo_lo_lo_17};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_17 = {regroupV0_lo_68[686], regroupV0_lo_68[654]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_17 = {regroupV0_lo_68[750], regroupV0_lo_68[718]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_51 = {regroupV0_lo_hi_lo_hi_hi_17, regroupV0_lo_hi_lo_hi_lo_17};
  wire [7:0]         regroupV0_lo_hi_lo_83 = {regroupV0_lo_hi_lo_hi_51, regroupV0_lo_hi_lo_lo_51};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_17 = {regroupV0_lo_68[814], regroupV0_lo_68[782]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_17 = {regroupV0_lo_68[878], regroupV0_lo_68[846]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_51 = {regroupV0_lo_hi_hi_lo_hi_17, regroupV0_lo_hi_hi_lo_lo_17};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_17 = {regroupV0_lo_68[942], regroupV0_lo_68[910]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_17 = {regroupV0_lo_68[1006], regroupV0_lo_68[974]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_51 = {regroupV0_lo_hi_hi_hi_hi_17, regroupV0_lo_hi_hi_hi_lo_17};
  wire [7:0]         regroupV0_lo_hi_hi_83 = {regroupV0_lo_hi_hi_hi_51, regroupV0_lo_hi_hi_lo_51};
  wire [15:0]        regroupV0_lo_hi_83 = {regroupV0_lo_hi_hi_83, regroupV0_lo_hi_lo_83};
  wire [31:0]        regroupV0_lo_83 = {regroupV0_lo_hi_83, regroupV0_lo_lo_83};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_17 = {regroupV0_hi_68[46], regroupV0_hi_68[14]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_17 = {regroupV0_hi_68[110], regroupV0_hi_68[78]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_51 = {regroupV0_hi_lo_lo_lo_hi_17, regroupV0_hi_lo_lo_lo_lo_17};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_17 = {regroupV0_hi_68[174], regroupV0_hi_68[142]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_17 = {regroupV0_hi_68[238], regroupV0_hi_68[206]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_51 = {regroupV0_hi_lo_lo_hi_hi_17, regroupV0_hi_lo_lo_hi_lo_17};
  wire [7:0]         regroupV0_hi_lo_lo_83 = {regroupV0_hi_lo_lo_hi_51, regroupV0_hi_lo_lo_lo_51};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_17 = {regroupV0_hi_68[302], regroupV0_hi_68[270]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_17 = {regroupV0_hi_68[366], regroupV0_hi_68[334]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_51 = {regroupV0_hi_lo_hi_lo_hi_17, regroupV0_hi_lo_hi_lo_lo_17};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_17 = {regroupV0_hi_68[430], regroupV0_hi_68[398]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_17 = {regroupV0_hi_68[494], regroupV0_hi_68[462]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_51 = {regroupV0_hi_lo_hi_hi_hi_17, regroupV0_hi_lo_hi_hi_lo_17};
  wire [7:0]         regroupV0_hi_lo_hi_83 = {regroupV0_hi_lo_hi_hi_51, regroupV0_hi_lo_hi_lo_51};
  wire [15:0]        regroupV0_hi_lo_83 = {regroupV0_hi_lo_hi_83, regroupV0_hi_lo_lo_83};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_17 = {regroupV0_hi_68[558], regroupV0_hi_68[526]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_17 = {regroupV0_hi_68[622], regroupV0_hi_68[590]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_51 = {regroupV0_hi_hi_lo_lo_hi_17, regroupV0_hi_hi_lo_lo_lo_17};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_17 = {regroupV0_hi_68[686], regroupV0_hi_68[654]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_17 = {regroupV0_hi_68[750], regroupV0_hi_68[718]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_51 = {regroupV0_hi_hi_lo_hi_hi_17, regroupV0_hi_hi_lo_hi_lo_17};
  wire [7:0]         regroupV0_hi_hi_lo_83 = {regroupV0_hi_hi_lo_hi_51, regroupV0_hi_hi_lo_lo_51};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_17 = {regroupV0_hi_68[814], regroupV0_hi_68[782]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_17 = {regroupV0_hi_68[878], regroupV0_hi_68[846]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_51 = {regroupV0_hi_hi_hi_lo_hi_17, regroupV0_hi_hi_hi_lo_lo_17};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_17 = {regroupV0_hi_68[942], regroupV0_hi_68[910]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_17 = {regroupV0_hi_68[1006], regroupV0_hi_68[974]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_51 = {regroupV0_hi_hi_hi_hi_hi_17, regroupV0_hi_hi_hi_hi_lo_17};
  wire [7:0]         regroupV0_hi_hi_hi_83 = {regroupV0_hi_hi_hi_hi_51, regroupV0_hi_hi_hi_lo_51};
  wire [15:0]        regroupV0_hi_hi_83 = {regroupV0_hi_hi_hi_83, regroupV0_hi_hi_lo_83};
  wire [31:0]        regroupV0_hi_83 = {regroupV0_hi_hi_83, regroupV0_hi_lo_83};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_18 = {regroupV0_lo_68[47], regroupV0_lo_68[15]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_18 = {regroupV0_lo_68[111], regroupV0_lo_68[79]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_52 = {regroupV0_lo_lo_lo_lo_hi_18, regroupV0_lo_lo_lo_lo_lo_18};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_18 = {regroupV0_lo_68[175], regroupV0_lo_68[143]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_18 = {regroupV0_lo_68[239], regroupV0_lo_68[207]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_52 = {regroupV0_lo_lo_lo_hi_hi_18, regroupV0_lo_lo_lo_hi_lo_18};
  wire [7:0]         regroupV0_lo_lo_lo_84 = {regroupV0_lo_lo_lo_hi_52, regroupV0_lo_lo_lo_lo_52};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_18 = {regroupV0_lo_68[303], regroupV0_lo_68[271]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_18 = {regroupV0_lo_68[367], regroupV0_lo_68[335]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_52 = {regroupV0_lo_lo_hi_lo_hi_18, regroupV0_lo_lo_hi_lo_lo_18};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_18 = {regroupV0_lo_68[431], regroupV0_lo_68[399]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_18 = {regroupV0_lo_68[495], regroupV0_lo_68[463]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_52 = {regroupV0_lo_lo_hi_hi_hi_18, regroupV0_lo_lo_hi_hi_lo_18};
  wire [7:0]         regroupV0_lo_lo_hi_84 = {regroupV0_lo_lo_hi_hi_52, regroupV0_lo_lo_hi_lo_52};
  wire [15:0]        regroupV0_lo_lo_84 = {regroupV0_lo_lo_hi_84, regroupV0_lo_lo_lo_84};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_18 = {regroupV0_lo_68[559], regroupV0_lo_68[527]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_18 = {regroupV0_lo_68[623], regroupV0_lo_68[591]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_52 = {regroupV0_lo_hi_lo_lo_hi_18, regroupV0_lo_hi_lo_lo_lo_18};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_18 = {regroupV0_lo_68[687], regroupV0_lo_68[655]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_18 = {regroupV0_lo_68[751], regroupV0_lo_68[719]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_52 = {regroupV0_lo_hi_lo_hi_hi_18, regroupV0_lo_hi_lo_hi_lo_18};
  wire [7:0]         regroupV0_lo_hi_lo_84 = {regroupV0_lo_hi_lo_hi_52, regroupV0_lo_hi_lo_lo_52};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_18 = {regroupV0_lo_68[815], regroupV0_lo_68[783]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_18 = {regroupV0_lo_68[879], regroupV0_lo_68[847]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_52 = {regroupV0_lo_hi_hi_lo_hi_18, regroupV0_lo_hi_hi_lo_lo_18};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_18 = {regroupV0_lo_68[943], regroupV0_lo_68[911]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_18 = {regroupV0_lo_68[1007], regroupV0_lo_68[975]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_52 = {regroupV0_lo_hi_hi_hi_hi_18, regroupV0_lo_hi_hi_hi_lo_18};
  wire [7:0]         regroupV0_lo_hi_hi_84 = {regroupV0_lo_hi_hi_hi_52, regroupV0_lo_hi_hi_lo_52};
  wire [15:0]        regroupV0_lo_hi_84 = {regroupV0_lo_hi_hi_84, regroupV0_lo_hi_lo_84};
  wire [31:0]        regroupV0_lo_84 = {regroupV0_lo_hi_84, regroupV0_lo_lo_84};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_18 = {regroupV0_hi_68[47], regroupV0_hi_68[15]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_18 = {regroupV0_hi_68[111], regroupV0_hi_68[79]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_52 = {regroupV0_hi_lo_lo_lo_hi_18, regroupV0_hi_lo_lo_lo_lo_18};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_18 = {regroupV0_hi_68[175], regroupV0_hi_68[143]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_18 = {regroupV0_hi_68[239], regroupV0_hi_68[207]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_52 = {regroupV0_hi_lo_lo_hi_hi_18, regroupV0_hi_lo_lo_hi_lo_18};
  wire [7:0]         regroupV0_hi_lo_lo_84 = {regroupV0_hi_lo_lo_hi_52, regroupV0_hi_lo_lo_lo_52};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_18 = {regroupV0_hi_68[303], regroupV0_hi_68[271]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_18 = {regroupV0_hi_68[367], regroupV0_hi_68[335]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_52 = {regroupV0_hi_lo_hi_lo_hi_18, regroupV0_hi_lo_hi_lo_lo_18};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_18 = {regroupV0_hi_68[431], regroupV0_hi_68[399]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_18 = {regroupV0_hi_68[495], regroupV0_hi_68[463]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_52 = {regroupV0_hi_lo_hi_hi_hi_18, regroupV0_hi_lo_hi_hi_lo_18};
  wire [7:0]         regroupV0_hi_lo_hi_84 = {regroupV0_hi_lo_hi_hi_52, regroupV0_hi_lo_hi_lo_52};
  wire [15:0]        regroupV0_hi_lo_84 = {regroupV0_hi_lo_hi_84, regroupV0_hi_lo_lo_84};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_18 = {regroupV0_hi_68[559], regroupV0_hi_68[527]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_18 = {regroupV0_hi_68[623], regroupV0_hi_68[591]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_52 = {regroupV0_hi_hi_lo_lo_hi_18, regroupV0_hi_hi_lo_lo_lo_18};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_18 = {regroupV0_hi_68[687], regroupV0_hi_68[655]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_18 = {regroupV0_hi_68[751], regroupV0_hi_68[719]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_52 = {regroupV0_hi_hi_lo_hi_hi_18, regroupV0_hi_hi_lo_hi_lo_18};
  wire [7:0]         regroupV0_hi_hi_lo_84 = {regroupV0_hi_hi_lo_hi_52, regroupV0_hi_hi_lo_lo_52};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_18 = {regroupV0_hi_68[815], regroupV0_hi_68[783]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_18 = {regroupV0_hi_68[879], regroupV0_hi_68[847]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_52 = {regroupV0_hi_hi_hi_lo_hi_18, regroupV0_hi_hi_hi_lo_lo_18};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_18 = {regroupV0_hi_68[943], regroupV0_hi_68[911]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_18 = {regroupV0_hi_68[1007], regroupV0_hi_68[975]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_52 = {regroupV0_hi_hi_hi_hi_hi_18, regroupV0_hi_hi_hi_hi_lo_18};
  wire [7:0]         regroupV0_hi_hi_hi_84 = {regroupV0_hi_hi_hi_hi_52, regroupV0_hi_hi_hi_lo_52};
  wire [15:0]        regroupV0_hi_hi_84 = {regroupV0_hi_hi_hi_84, regroupV0_hi_hi_lo_84};
  wire [31:0]        regroupV0_hi_84 = {regroupV0_hi_hi_84, regroupV0_hi_lo_84};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_19 = {regroupV0_lo_68[48], regroupV0_lo_68[16]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_19 = {regroupV0_lo_68[112], regroupV0_lo_68[80]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_53 = {regroupV0_lo_lo_lo_lo_hi_19, regroupV0_lo_lo_lo_lo_lo_19};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_19 = {regroupV0_lo_68[176], regroupV0_lo_68[144]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_19 = {regroupV0_lo_68[240], regroupV0_lo_68[208]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_53 = {regroupV0_lo_lo_lo_hi_hi_19, regroupV0_lo_lo_lo_hi_lo_19};
  wire [7:0]         regroupV0_lo_lo_lo_85 = {regroupV0_lo_lo_lo_hi_53, regroupV0_lo_lo_lo_lo_53};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_19 = {regroupV0_lo_68[304], regroupV0_lo_68[272]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_19 = {regroupV0_lo_68[368], regroupV0_lo_68[336]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_53 = {regroupV0_lo_lo_hi_lo_hi_19, regroupV0_lo_lo_hi_lo_lo_19};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_19 = {regroupV0_lo_68[432], regroupV0_lo_68[400]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_19 = {regroupV0_lo_68[496], regroupV0_lo_68[464]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_53 = {regroupV0_lo_lo_hi_hi_hi_19, regroupV0_lo_lo_hi_hi_lo_19};
  wire [7:0]         regroupV0_lo_lo_hi_85 = {regroupV0_lo_lo_hi_hi_53, regroupV0_lo_lo_hi_lo_53};
  wire [15:0]        regroupV0_lo_lo_85 = {regroupV0_lo_lo_hi_85, regroupV0_lo_lo_lo_85};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_19 = {regroupV0_lo_68[560], regroupV0_lo_68[528]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_19 = {regroupV0_lo_68[624], regroupV0_lo_68[592]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_53 = {regroupV0_lo_hi_lo_lo_hi_19, regroupV0_lo_hi_lo_lo_lo_19};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_19 = {regroupV0_lo_68[688], regroupV0_lo_68[656]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_19 = {regroupV0_lo_68[752], regroupV0_lo_68[720]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_53 = {regroupV0_lo_hi_lo_hi_hi_19, regroupV0_lo_hi_lo_hi_lo_19};
  wire [7:0]         regroupV0_lo_hi_lo_85 = {regroupV0_lo_hi_lo_hi_53, regroupV0_lo_hi_lo_lo_53};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_19 = {regroupV0_lo_68[816], regroupV0_lo_68[784]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_19 = {regroupV0_lo_68[880], regroupV0_lo_68[848]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_53 = {regroupV0_lo_hi_hi_lo_hi_19, regroupV0_lo_hi_hi_lo_lo_19};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_19 = {regroupV0_lo_68[944], regroupV0_lo_68[912]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_19 = {regroupV0_lo_68[1008], regroupV0_lo_68[976]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_53 = {regroupV0_lo_hi_hi_hi_hi_19, regroupV0_lo_hi_hi_hi_lo_19};
  wire [7:0]         regroupV0_lo_hi_hi_85 = {regroupV0_lo_hi_hi_hi_53, regroupV0_lo_hi_hi_lo_53};
  wire [15:0]        regroupV0_lo_hi_85 = {regroupV0_lo_hi_hi_85, regroupV0_lo_hi_lo_85};
  wire [31:0]        regroupV0_lo_85 = {regroupV0_lo_hi_85, regroupV0_lo_lo_85};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_19 = {regroupV0_hi_68[48], regroupV0_hi_68[16]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_19 = {regroupV0_hi_68[112], regroupV0_hi_68[80]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_53 = {regroupV0_hi_lo_lo_lo_hi_19, regroupV0_hi_lo_lo_lo_lo_19};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_19 = {regroupV0_hi_68[176], regroupV0_hi_68[144]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_19 = {regroupV0_hi_68[240], regroupV0_hi_68[208]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_53 = {regroupV0_hi_lo_lo_hi_hi_19, regroupV0_hi_lo_lo_hi_lo_19};
  wire [7:0]         regroupV0_hi_lo_lo_85 = {regroupV0_hi_lo_lo_hi_53, regroupV0_hi_lo_lo_lo_53};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_19 = {regroupV0_hi_68[304], regroupV0_hi_68[272]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_19 = {regroupV0_hi_68[368], regroupV0_hi_68[336]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_53 = {regroupV0_hi_lo_hi_lo_hi_19, regroupV0_hi_lo_hi_lo_lo_19};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_19 = {regroupV0_hi_68[432], regroupV0_hi_68[400]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_19 = {regroupV0_hi_68[496], regroupV0_hi_68[464]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_53 = {regroupV0_hi_lo_hi_hi_hi_19, regroupV0_hi_lo_hi_hi_lo_19};
  wire [7:0]         regroupV0_hi_lo_hi_85 = {regroupV0_hi_lo_hi_hi_53, regroupV0_hi_lo_hi_lo_53};
  wire [15:0]        regroupV0_hi_lo_85 = {regroupV0_hi_lo_hi_85, regroupV0_hi_lo_lo_85};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_19 = {regroupV0_hi_68[560], regroupV0_hi_68[528]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_19 = {regroupV0_hi_68[624], regroupV0_hi_68[592]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_53 = {regroupV0_hi_hi_lo_lo_hi_19, regroupV0_hi_hi_lo_lo_lo_19};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_19 = {regroupV0_hi_68[688], regroupV0_hi_68[656]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_19 = {regroupV0_hi_68[752], regroupV0_hi_68[720]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_53 = {regroupV0_hi_hi_lo_hi_hi_19, regroupV0_hi_hi_lo_hi_lo_19};
  wire [7:0]         regroupV0_hi_hi_lo_85 = {regroupV0_hi_hi_lo_hi_53, regroupV0_hi_hi_lo_lo_53};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_19 = {regroupV0_hi_68[816], regroupV0_hi_68[784]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_19 = {regroupV0_hi_68[880], regroupV0_hi_68[848]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_53 = {regroupV0_hi_hi_hi_lo_hi_19, regroupV0_hi_hi_hi_lo_lo_19};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_19 = {regroupV0_hi_68[944], regroupV0_hi_68[912]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_19 = {regroupV0_hi_68[1008], regroupV0_hi_68[976]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_53 = {regroupV0_hi_hi_hi_hi_hi_19, regroupV0_hi_hi_hi_hi_lo_19};
  wire [7:0]         regroupV0_hi_hi_hi_85 = {regroupV0_hi_hi_hi_hi_53, regroupV0_hi_hi_hi_lo_53};
  wire [15:0]        regroupV0_hi_hi_85 = {regroupV0_hi_hi_hi_85, regroupV0_hi_hi_lo_85};
  wire [31:0]        regroupV0_hi_85 = {regroupV0_hi_hi_85, regroupV0_hi_lo_85};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_20 = {regroupV0_lo_68[49], regroupV0_lo_68[17]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_20 = {regroupV0_lo_68[113], regroupV0_lo_68[81]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_54 = {regroupV0_lo_lo_lo_lo_hi_20, regroupV0_lo_lo_lo_lo_lo_20};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_20 = {regroupV0_lo_68[177], regroupV0_lo_68[145]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_20 = {regroupV0_lo_68[241], regroupV0_lo_68[209]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_54 = {regroupV0_lo_lo_lo_hi_hi_20, regroupV0_lo_lo_lo_hi_lo_20};
  wire [7:0]         regroupV0_lo_lo_lo_86 = {regroupV0_lo_lo_lo_hi_54, regroupV0_lo_lo_lo_lo_54};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_20 = {regroupV0_lo_68[305], regroupV0_lo_68[273]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_20 = {regroupV0_lo_68[369], regroupV0_lo_68[337]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_54 = {regroupV0_lo_lo_hi_lo_hi_20, regroupV0_lo_lo_hi_lo_lo_20};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_20 = {regroupV0_lo_68[433], regroupV0_lo_68[401]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_20 = {regroupV0_lo_68[497], regroupV0_lo_68[465]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_54 = {regroupV0_lo_lo_hi_hi_hi_20, regroupV0_lo_lo_hi_hi_lo_20};
  wire [7:0]         regroupV0_lo_lo_hi_86 = {regroupV0_lo_lo_hi_hi_54, regroupV0_lo_lo_hi_lo_54};
  wire [15:0]        regroupV0_lo_lo_86 = {regroupV0_lo_lo_hi_86, regroupV0_lo_lo_lo_86};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_20 = {regroupV0_lo_68[561], regroupV0_lo_68[529]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_20 = {regroupV0_lo_68[625], regroupV0_lo_68[593]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_54 = {regroupV0_lo_hi_lo_lo_hi_20, regroupV0_lo_hi_lo_lo_lo_20};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_20 = {regroupV0_lo_68[689], regroupV0_lo_68[657]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_20 = {regroupV0_lo_68[753], regroupV0_lo_68[721]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_54 = {regroupV0_lo_hi_lo_hi_hi_20, regroupV0_lo_hi_lo_hi_lo_20};
  wire [7:0]         regroupV0_lo_hi_lo_86 = {regroupV0_lo_hi_lo_hi_54, regroupV0_lo_hi_lo_lo_54};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_20 = {regroupV0_lo_68[817], regroupV0_lo_68[785]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_20 = {regroupV0_lo_68[881], regroupV0_lo_68[849]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_54 = {regroupV0_lo_hi_hi_lo_hi_20, regroupV0_lo_hi_hi_lo_lo_20};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_20 = {regroupV0_lo_68[945], regroupV0_lo_68[913]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_20 = {regroupV0_lo_68[1009], regroupV0_lo_68[977]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_54 = {regroupV0_lo_hi_hi_hi_hi_20, regroupV0_lo_hi_hi_hi_lo_20};
  wire [7:0]         regroupV0_lo_hi_hi_86 = {regroupV0_lo_hi_hi_hi_54, regroupV0_lo_hi_hi_lo_54};
  wire [15:0]        regroupV0_lo_hi_86 = {regroupV0_lo_hi_hi_86, regroupV0_lo_hi_lo_86};
  wire [31:0]        regroupV0_lo_86 = {regroupV0_lo_hi_86, regroupV0_lo_lo_86};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_20 = {regroupV0_hi_68[49], regroupV0_hi_68[17]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_20 = {regroupV0_hi_68[113], regroupV0_hi_68[81]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_54 = {regroupV0_hi_lo_lo_lo_hi_20, regroupV0_hi_lo_lo_lo_lo_20};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_20 = {regroupV0_hi_68[177], regroupV0_hi_68[145]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_20 = {regroupV0_hi_68[241], regroupV0_hi_68[209]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_54 = {regroupV0_hi_lo_lo_hi_hi_20, regroupV0_hi_lo_lo_hi_lo_20};
  wire [7:0]         regroupV0_hi_lo_lo_86 = {regroupV0_hi_lo_lo_hi_54, regroupV0_hi_lo_lo_lo_54};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_20 = {regroupV0_hi_68[305], regroupV0_hi_68[273]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_20 = {regroupV0_hi_68[369], regroupV0_hi_68[337]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_54 = {regroupV0_hi_lo_hi_lo_hi_20, regroupV0_hi_lo_hi_lo_lo_20};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_20 = {regroupV0_hi_68[433], regroupV0_hi_68[401]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_20 = {regroupV0_hi_68[497], regroupV0_hi_68[465]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_54 = {regroupV0_hi_lo_hi_hi_hi_20, regroupV0_hi_lo_hi_hi_lo_20};
  wire [7:0]         regroupV0_hi_lo_hi_86 = {regroupV0_hi_lo_hi_hi_54, regroupV0_hi_lo_hi_lo_54};
  wire [15:0]        regroupV0_hi_lo_86 = {regroupV0_hi_lo_hi_86, regroupV0_hi_lo_lo_86};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_20 = {regroupV0_hi_68[561], regroupV0_hi_68[529]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_20 = {regroupV0_hi_68[625], regroupV0_hi_68[593]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_54 = {regroupV0_hi_hi_lo_lo_hi_20, regroupV0_hi_hi_lo_lo_lo_20};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_20 = {regroupV0_hi_68[689], regroupV0_hi_68[657]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_20 = {regroupV0_hi_68[753], regroupV0_hi_68[721]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_54 = {regroupV0_hi_hi_lo_hi_hi_20, regroupV0_hi_hi_lo_hi_lo_20};
  wire [7:0]         regroupV0_hi_hi_lo_86 = {regroupV0_hi_hi_lo_hi_54, regroupV0_hi_hi_lo_lo_54};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_20 = {regroupV0_hi_68[817], regroupV0_hi_68[785]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_20 = {regroupV0_hi_68[881], regroupV0_hi_68[849]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_54 = {regroupV0_hi_hi_hi_lo_hi_20, regroupV0_hi_hi_hi_lo_lo_20};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_20 = {regroupV0_hi_68[945], regroupV0_hi_68[913]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_20 = {regroupV0_hi_68[1009], regroupV0_hi_68[977]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_54 = {regroupV0_hi_hi_hi_hi_hi_20, regroupV0_hi_hi_hi_hi_lo_20};
  wire [7:0]         regroupV0_hi_hi_hi_86 = {regroupV0_hi_hi_hi_hi_54, regroupV0_hi_hi_hi_lo_54};
  wire [15:0]        regroupV0_hi_hi_86 = {regroupV0_hi_hi_hi_86, regroupV0_hi_hi_lo_86};
  wire [31:0]        regroupV0_hi_86 = {regroupV0_hi_hi_86, regroupV0_hi_lo_86};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_21 = {regroupV0_lo_68[50], regroupV0_lo_68[18]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_21 = {regroupV0_lo_68[114], regroupV0_lo_68[82]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_55 = {regroupV0_lo_lo_lo_lo_hi_21, regroupV0_lo_lo_lo_lo_lo_21};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_21 = {regroupV0_lo_68[178], regroupV0_lo_68[146]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_21 = {regroupV0_lo_68[242], regroupV0_lo_68[210]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_55 = {regroupV0_lo_lo_lo_hi_hi_21, regroupV0_lo_lo_lo_hi_lo_21};
  wire [7:0]         regroupV0_lo_lo_lo_87 = {regroupV0_lo_lo_lo_hi_55, regroupV0_lo_lo_lo_lo_55};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_21 = {regroupV0_lo_68[306], regroupV0_lo_68[274]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_21 = {regroupV0_lo_68[370], regroupV0_lo_68[338]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_55 = {regroupV0_lo_lo_hi_lo_hi_21, regroupV0_lo_lo_hi_lo_lo_21};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_21 = {regroupV0_lo_68[434], regroupV0_lo_68[402]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_21 = {regroupV0_lo_68[498], regroupV0_lo_68[466]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_55 = {regroupV0_lo_lo_hi_hi_hi_21, regroupV0_lo_lo_hi_hi_lo_21};
  wire [7:0]         regroupV0_lo_lo_hi_87 = {regroupV0_lo_lo_hi_hi_55, regroupV0_lo_lo_hi_lo_55};
  wire [15:0]        regroupV0_lo_lo_87 = {regroupV0_lo_lo_hi_87, regroupV0_lo_lo_lo_87};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_21 = {regroupV0_lo_68[562], regroupV0_lo_68[530]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_21 = {regroupV0_lo_68[626], regroupV0_lo_68[594]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_55 = {regroupV0_lo_hi_lo_lo_hi_21, regroupV0_lo_hi_lo_lo_lo_21};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_21 = {regroupV0_lo_68[690], regroupV0_lo_68[658]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_21 = {regroupV0_lo_68[754], regroupV0_lo_68[722]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_55 = {regroupV0_lo_hi_lo_hi_hi_21, regroupV0_lo_hi_lo_hi_lo_21};
  wire [7:0]         regroupV0_lo_hi_lo_87 = {regroupV0_lo_hi_lo_hi_55, regroupV0_lo_hi_lo_lo_55};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_21 = {regroupV0_lo_68[818], regroupV0_lo_68[786]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_21 = {regroupV0_lo_68[882], regroupV0_lo_68[850]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_55 = {regroupV0_lo_hi_hi_lo_hi_21, regroupV0_lo_hi_hi_lo_lo_21};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_21 = {regroupV0_lo_68[946], regroupV0_lo_68[914]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_21 = {regroupV0_lo_68[1010], regroupV0_lo_68[978]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_55 = {regroupV0_lo_hi_hi_hi_hi_21, regroupV0_lo_hi_hi_hi_lo_21};
  wire [7:0]         regroupV0_lo_hi_hi_87 = {regroupV0_lo_hi_hi_hi_55, regroupV0_lo_hi_hi_lo_55};
  wire [15:0]        regroupV0_lo_hi_87 = {regroupV0_lo_hi_hi_87, regroupV0_lo_hi_lo_87};
  wire [31:0]        regroupV0_lo_87 = {regroupV0_lo_hi_87, regroupV0_lo_lo_87};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_21 = {regroupV0_hi_68[50], regroupV0_hi_68[18]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_21 = {regroupV0_hi_68[114], regroupV0_hi_68[82]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_55 = {regroupV0_hi_lo_lo_lo_hi_21, regroupV0_hi_lo_lo_lo_lo_21};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_21 = {regroupV0_hi_68[178], regroupV0_hi_68[146]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_21 = {regroupV0_hi_68[242], regroupV0_hi_68[210]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_55 = {regroupV0_hi_lo_lo_hi_hi_21, regroupV0_hi_lo_lo_hi_lo_21};
  wire [7:0]         regroupV0_hi_lo_lo_87 = {regroupV0_hi_lo_lo_hi_55, regroupV0_hi_lo_lo_lo_55};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_21 = {regroupV0_hi_68[306], regroupV0_hi_68[274]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_21 = {regroupV0_hi_68[370], regroupV0_hi_68[338]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_55 = {regroupV0_hi_lo_hi_lo_hi_21, regroupV0_hi_lo_hi_lo_lo_21};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_21 = {regroupV0_hi_68[434], regroupV0_hi_68[402]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_21 = {regroupV0_hi_68[498], regroupV0_hi_68[466]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_55 = {regroupV0_hi_lo_hi_hi_hi_21, regroupV0_hi_lo_hi_hi_lo_21};
  wire [7:0]         regroupV0_hi_lo_hi_87 = {regroupV0_hi_lo_hi_hi_55, regroupV0_hi_lo_hi_lo_55};
  wire [15:0]        regroupV0_hi_lo_87 = {regroupV0_hi_lo_hi_87, regroupV0_hi_lo_lo_87};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_21 = {regroupV0_hi_68[562], regroupV0_hi_68[530]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_21 = {regroupV0_hi_68[626], regroupV0_hi_68[594]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_55 = {regroupV0_hi_hi_lo_lo_hi_21, regroupV0_hi_hi_lo_lo_lo_21};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_21 = {regroupV0_hi_68[690], regroupV0_hi_68[658]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_21 = {regroupV0_hi_68[754], regroupV0_hi_68[722]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_55 = {regroupV0_hi_hi_lo_hi_hi_21, regroupV0_hi_hi_lo_hi_lo_21};
  wire [7:0]         regroupV0_hi_hi_lo_87 = {regroupV0_hi_hi_lo_hi_55, regroupV0_hi_hi_lo_lo_55};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_21 = {regroupV0_hi_68[818], regroupV0_hi_68[786]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_21 = {regroupV0_hi_68[882], regroupV0_hi_68[850]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_55 = {regroupV0_hi_hi_hi_lo_hi_21, regroupV0_hi_hi_hi_lo_lo_21};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_21 = {regroupV0_hi_68[946], regroupV0_hi_68[914]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_21 = {regroupV0_hi_68[1010], regroupV0_hi_68[978]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_55 = {regroupV0_hi_hi_hi_hi_hi_21, regroupV0_hi_hi_hi_hi_lo_21};
  wire [7:0]         regroupV0_hi_hi_hi_87 = {regroupV0_hi_hi_hi_hi_55, regroupV0_hi_hi_hi_lo_55};
  wire [15:0]        regroupV0_hi_hi_87 = {regroupV0_hi_hi_hi_87, regroupV0_hi_hi_lo_87};
  wire [31:0]        regroupV0_hi_87 = {regroupV0_hi_hi_87, regroupV0_hi_lo_87};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_22 = {regroupV0_lo_68[51], regroupV0_lo_68[19]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_22 = {regroupV0_lo_68[115], regroupV0_lo_68[83]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_56 = {regroupV0_lo_lo_lo_lo_hi_22, regroupV0_lo_lo_lo_lo_lo_22};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_22 = {regroupV0_lo_68[179], regroupV0_lo_68[147]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_22 = {regroupV0_lo_68[243], regroupV0_lo_68[211]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_56 = {regroupV0_lo_lo_lo_hi_hi_22, regroupV0_lo_lo_lo_hi_lo_22};
  wire [7:0]         regroupV0_lo_lo_lo_88 = {regroupV0_lo_lo_lo_hi_56, regroupV0_lo_lo_lo_lo_56};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_22 = {regroupV0_lo_68[307], regroupV0_lo_68[275]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_22 = {regroupV0_lo_68[371], regroupV0_lo_68[339]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_56 = {regroupV0_lo_lo_hi_lo_hi_22, regroupV0_lo_lo_hi_lo_lo_22};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_22 = {regroupV0_lo_68[435], regroupV0_lo_68[403]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_22 = {regroupV0_lo_68[499], regroupV0_lo_68[467]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_56 = {regroupV0_lo_lo_hi_hi_hi_22, regroupV0_lo_lo_hi_hi_lo_22};
  wire [7:0]         regroupV0_lo_lo_hi_88 = {regroupV0_lo_lo_hi_hi_56, regroupV0_lo_lo_hi_lo_56};
  wire [15:0]        regroupV0_lo_lo_88 = {regroupV0_lo_lo_hi_88, regroupV0_lo_lo_lo_88};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_22 = {regroupV0_lo_68[563], regroupV0_lo_68[531]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_22 = {regroupV0_lo_68[627], regroupV0_lo_68[595]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_56 = {regroupV0_lo_hi_lo_lo_hi_22, regroupV0_lo_hi_lo_lo_lo_22};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_22 = {regroupV0_lo_68[691], regroupV0_lo_68[659]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_22 = {regroupV0_lo_68[755], regroupV0_lo_68[723]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_56 = {regroupV0_lo_hi_lo_hi_hi_22, regroupV0_lo_hi_lo_hi_lo_22};
  wire [7:0]         regroupV0_lo_hi_lo_88 = {regroupV0_lo_hi_lo_hi_56, regroupV0_lo_hi_lo_lo_56};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_22 = {regroupV0_lo_68[819], regroupV0_lo_68[787]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_22 = {regroupV0_lo_68[883], regroupV0_lo_68[851]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_56 = {regroupV0_lo_hi_hi_lo_hi_22, regroupV0_lo_hi_hi_lo_lo_22};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_22 = {regroupV0_lo_68[947], regroupV0_lo_68[915]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_22 = {regroupV0_lo_68[1011], regroupV0_lo_68[979]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_56 = {regroupV0_lo_hi_hi_hi_hi_22, regroupV0_lo_hi_hi_hi_lo_22};
  wire [7:0]         regroupV0_lo_hi_hi_88 = {regroupV0_lo_hi_hi_hi_56, regroupV0_lo_hi_hi_lo_56};
  wire [15:0]        regroupV0_lo_hi_88 = {regroupV0_lo_hi_hi_88, regroupV0_lo_hi_lo_88};
  wire [31:0]        regroupV0_lo_88 = {regroupV0_lo_hi_88, regroupV0_lo_lo_88};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_22 = {regroupV0_hi_68[51], regroupV0_hi_68[19]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_22 = {regroupV0_hi_68[115], regroupV0_hi_68[83]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_56 = {regroupV0_hi_lo_lo_lo_hi_22, regroupV0_hi_lo_lo_lo_lo_22};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_22 = {regroupV0_hi_68[179], regroupV0_hi_68[147]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_22 = {regroupV0_hi_68[243], regroupV0_hi_68[211]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_56 = {regroupV0_hi_lo_lo_hi_hi_22, regroupV0_hi_lo_lo_hi_lo_22};
  wire [7:0]         regroupV0_hi_lo_lo_88 = {regroupV0_hi_lo_lo_hi_56, regroupV0_hi_lo_lo_lo_56};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_22 = {regroupV0_hi_68[307], regroupV0_hi_68[275]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_22 = {regroupV0_hi_68[371], regroupV0_hi_68[339]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_56 = {regroupV0_hi_lo_hi_lo_hi_22, regroupV0_hi_lo_hi_lo_lo_22};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_22 = {regroupV0_hi_68[435], regroupV0_hi_68[403]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_22 = {regroupV0_hi_68[499], regroupV0_hi_68[467]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_56 = {regroupV0_hi_lo_hi_hi_hi_22, regroupV0_hi_lo_hi_hi_lo_22};
  wire [7:0]         regroupV0_hi_lo_hi_88 = {regroupV0_hi_lo_hi_hi_56, regroupV0_hi_lo_hi_lo_56};
  wire [15:0]        regroupV0_hi_lo_88 = {regroupV0_hi_lo_hi_88, regroupV0_hi_lo_lo_88};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_22 = {regroupV0_hi_68[563], regroupV0_hi_68[531]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_22 = {regroupV0_hi_68[627], regroupV0_hi_68[595]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_56 = {regroupV0_hi_hi_lo_lo_hi_22, regroupV0_hi_hi_lo_lo_lo_22};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_22 = {regroupV0_hi_68[691], regroupV0_hi_68[659]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_22 = {regroupV0_hi_68[755], regroupV0_hi_68[723]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_56 = {regroupV0_hi_hi_lo_hi_hi_22, regroupV0_hi_hi_lo_hi_lo_22};
  wire [7:0]         regroupV0_hi_hi_lo_88 = {regroupV0_hi_hi_lo_hi_56, regroupV0_hi_hi_lo_lo_56};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_22 = {regroupV0_hi_68[819], regroupV0_hi_68[787]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_22 = {regroupV0_hi_68[883], regroupV0_hi_68[851]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_56 = {regroupV0_hi_hi_hi_lo_hi_22, regroupV0_hi_hi_hi_lo_lo_22};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_22 = {regroupV0_hi_68[947], regroupV0_hi_68[915]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_22 = {regroupV0_hi_68[1011], regroupV0_hi_68[979]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_56 = {regroupV0_hi_hi_hi_hi_hi_22, regroupV0_hi_hi_hi_hi_lo_22};
  wire [7:0]         regroupV0_hi_hi_hi_88 = {regroupV0_hi_hi_hi_hi_56, regroupV0_hi_hi_hi_lo_56};
  wire [15:0]        regroupV0_hi_hi_88 = {regroupV0_hi_hi_hi_88, regroupV0_hi_hi_lo_88};
  wire [31:0]        regroupV0_hi_88 = {regroupV0_hi_hi_88, regroupV0_hi_lo_88};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_23 = {regroupV0_lo_68[52], regroupV0_lo_68[20]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_23 = {regroupV0_lo_68[116], regroupV0_lo_68[84]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_57 = {regroupV0_lo_lo_lo_lo_hi_23, regroupV0_lo_lo_lo_lo_lo_23};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_23 = {regroupV0_lo_68[180], regroupV0_lo_68[148]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_23 = {regroupV0_lo_68[244], regroupV0_lo_68[212]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_57 = {regroupV0_lo_lo_lo_hi_hi_23, regroupV0_lo_lo_lo_hi_lo_23};
  wire [7:0]         regroupV0_lo_lo_lo_89 = {regroupV0_lo_lo_lo_hi_57, regroupV0_lo_lo_lo_lo_57};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_23 = {regroupV0_lo_68[308], regroupV0_lo_68[276]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_23 = {regroupV0_lo_68[372], regroupV0_lo_68[340]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_57 = {regroupV0_lo_lo_hi_lo_hi_23, regroupV0_lo_lo_hi_lo_lo_23};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_23 = {regroupV0_lo_68[436], regroupV0_lo_68[404]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_23 = {regroupV0_lo_68[500], regroupV0_lo_68[468]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_57 = {regroupV0_lo_lo_hi_hi_hi_23, regroupV0_lo_lo_hi_hi_lo_23};
  wire [7:0]         regroupV0_lo_lo_hi_89 = {regroupV0_lo_lo_hi_hi_57, regroupV0_lo_lo_hi_lo_57};
  wire [15:0]        regroupV0_lo_lo_89 = {regroupV0_lo_lo_hi_89, regroupV0_lo_lo_lo_89};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_23 = {regroupV0_lo_68[564], regroupV0_lo_68[532]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_23 = {regroupV0_lo_68[628], regroupV0_lo_68[596]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_57 = {regroupV0_lo_hi_lo_lo_hi_23, regroupV0_lo_hi_lo_lo_lo_23};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_23 = {regroupV0_lo_68[692], regroupV0_lo_68[660]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_23 = {regroupV0_lo_68[756], regroupV0_lo_68[724]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_57 = {regroupV0_lo_hi_lo_hi_hi_23, regroupV0_lo_hi_lo_hi_lo_23};
  wire [7:0]         regroupV0_lo_hi_lo_89 = {regroupV0_lo_hi_lo_hi_57, regroupV0_lo_hi_lo_lo_57};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_23 = {regroupV0_lo_68[820], regroupV0_lo_68[788]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_23 = {regroupV0_lo_68[884], regroupV0_lo_68[852]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_57 = {regroupV0_lo_hi_hi_lo_hi_23, regroupV0_lo_hi_hi_lo_lo_23};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_23 = {regroupV0_lo_68[948], regroupV0_lo_68[916]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_23 = {regroupV0_lo_68[1012], regroupV0_lo_68[980]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_57 = {regroupV0_lo_hi_hi_hi_hi_23, regroupV0_lo_hi_hi_hi_lo_23};
  wire [7:0]         regroupV0_lo_hi_hi_89 = {regroupV0_lo_hi_hi_hi_57, regroupV0_lo_hi_hi_lo_57};
  wire [15:0]        regroupV0_lo_hi_89 = {regroupV0_lo_hi_hi_89, regroupV0_lo_hi_lo_89};
  wire [31:0]        regroupV0_lo_89 = {regroupV0_lo_hi_89, regroupV0_lo_lo_89};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_23 = {regroupV0_hi_68[52], regroupV0_hi_68[20]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_23 = {regroupV0_hi_68[116], regroupV0_hi_68[84]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_57 = {regroupV0_hi_lo_lo_lo_hi_23, regroupV0_hi_lo_lo_lo_lo_23};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_23 = {regroupV0_hi_68[180], regroupV0_hi_68[148]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_23 = {regroupV0_hi_68[244], regroupV0_hi_68[212]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_57 = {regroupV0_hi_lo_lo_hi_hi_23, regroupV0_hi_lo_lo_hi_lo_23};
  wire [7:0]         regroupV0_hi_lo_lo_89 = {regroupV0_hi_lo_lo_hi_57, regroupV0_hi_lo_lo_lo_57};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_23 = {regroupV0_hi_68[308], regroupV0_hi_68[276]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_23 = {regroupV0_hi_68[372], regroupV0_hi_68[340]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_57 = {regroupV0_hi_lo_hi_lo_hi_23, regroupV0_hi_lo_hi_lo_lo_23};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_23 = {regroupV0_hi_68[436], regroupV0_hi_68[404]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_23 = {regroupV0_hi_68[500], regroupV0_hi_68[468]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_57 = {regroupV0_hi_lo_hi_hi_hi_23, regroupV0_hi_lo_hi_hi_lo_23};
  wire [7:0]         regroupV0_hi_lo_hi_89 = {regroupV0_hi_lo_hi_hi_57, regroupV0_hi_lo_hi_lo_57};
  wire [15:0]        regroupV0_hi_lo_89 = {regroupV0_hi_lo_hi_89, regroupV0_hi_lo_lo_89};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_23 = {regroupV0_hi_68[564], regroupV0_hi_68[532]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_23 = {regroupV0_hi_68[628], regroupV0_hi_68[596]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_57 = {regroupV0_hi_hi_lo_lo_hi_23, regroupV0_hi_hi_lo_lo_lo_23};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_23 = {regroupV0_hi_68[692], regroupV0_hi_68[660]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_23 = {regroupV0_hi_68[756], regroupV0_hi_68[724]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_57 = {regroupV0_hi_hi_lo_hi_hi_23, regroupV0_hi_hi_lo_hi_lo_23};
  wire [7:0]         regroupV0_hi_hi_lo_89 = {regroupV0_hi_hi_lo_hi_57, regroupV0_hi_hi_lo_lo_57};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_23 = {regroupV0_hi_68[820], regroupV0_hi_68[788]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_23 = {regroupV0_hi_68[884], regroupV0_hi_68[852]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_57 = {regroupV0_hi_hi_hi_lo_hi_23, regroupV0_hi_hi_hi_lo_lo_23};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_23 = {regroupV0_hi_68[948], regroupV0_hi_68[916]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_23 = {regroupV0_hi_68[1012], regroupV0_hi_68[980]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_57 = {regroupV0_hi_hi_hi_hi_hi_23, regroupV0_hi_hi_hi_hi_lo_23};
  wire [7:0]         regroupV0_hi_hi_hi_89 = {regroupV0_hi_hi_hi_hi_57, regroupV0_hi_hi_hi_lo_57};
  wire [15:0]        regroupV0_hi_hi_89 = {regroupV0_hi_hi_hi_89, regroupV0_hi_hi_lo_89};
  wire [31:0]        regroupV0_hi_89 = {regroupV0_hi_hi_89, regroupV0_hi_lo_89};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_24 = {regroupV0_lo_68[53], regroupV0_lo_68[21]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_24 = {regroupV0_lo_68[117], regroupV0_lo_68[85]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_58 = {regroupV0_lo_lo_lo_lo_hi_24, regroupV0_lo_lo_lo_lo_lo_24};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_24 = {regroupV0_lo_68[181], regroupV0_lo_68[149]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_24 = {regroupV0_lo_68[245], regroupV0_lo_68[213]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_58 = {regroupV0_lo_lo_lo_hi_hi_24, regroupV0_lo_lo_lo_hi_lo_24};
  wire [7:0]         regroupV0_lo_lo_lo_90 = {regroupV0_lo_lo_lo_hi_58, regroupV0_lo_lo_lo_lo_58};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_24 = {regroupV0_lo_68[309], regroupV0_lo_68[277]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_24 = {regroupV0_lo_68[373], regroupV0_lo_68[341]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_58 = {regroupV0_lo_lo_hi_lo_hi_24, regroupV0_lo_lo_hi_lo_lo_24};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_24 = {regroupV0_lo_68[437], regroupV0_lo_68[405]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_24 = {regroupV0_lo_68[501], regroupV0_lo_68[469]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_58 = {regroupV0_lo_lo_hi_hi_hi_24, regroupV0_lo_lo_hi_hi_lo_24};
  wire [7:0]         regroupV0_lo_lo_hi_90 = {regroupV0_lo_lo_hi_hi_58, regroupV0_lo_lo_hi_lo_58};
  wire [15:0]        regroupV0_lo_lo_90 = {regroupV0_lo_lo_hi_90, regroupV0_lo_lo_lo_90};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_24 = {regroupV0_lo_68[565], regroupV0_lo_68[533]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_24 = {regroupV0_lo_68[629], regroupV0_lo_68[597]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_58 = {regroupV0_lo_hi_lo_lo_hi_24, regroupV0_lo_hi_lo_lo_lo_24};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_24 = {regroupV0_lo_68[693], regroupV0_lo_68[661]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_24 = {regroupV0_lo_68[757], regroupV0_lo_68[725]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_58 = {regroupV0_lo_hi_lo_hi_hi_24, regroupV0_lo_hi_lo_hi_lo_24};
  wire [7:0]         regroupV0_lo_hi_lo_90 = {regroupV0_lo_hi_lo_hi_58, regroupV0_lo_hi_lo_lo_58};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_24 = {regroupV0_lo_68[821], regroupV0_lo_68[789]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_24 = {regroupV0_lo_68[885], regroupV0_lo_68[853]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_58 = {regroupV0_lo_hi_hi_lo_hi_24, regroupV0_lo_hi_hi_lo_lo_24};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_24 = {regroupV0_lo_68[949], regroupV0_lo_68[917]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_24 = {regroupV0_lo_68[1013], regroupV0_lo_68[981]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_58 = {regroupV0_lo_hi_hi_hi_hi_24, regroupV0_lo_hi_hi_hi_lo_24};
  wire [7:0]         regroupV0_lo_hi_hi_90 = {regroupV0_lo_hi_hi_hi_58, regroupV0_lo_hi_hi_lo_58};
  wire [15:0]        regroupV0_lo_hi_90 = {regroupV0_lo_hi_hi_90, regroupV0_lo_hi_lo_90};
  wire [31:0]        regroupV0_lo_90 = {regroupV0_lo_hi_90, regroupV0_lo_lo_90};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_24 = {regroupV0_hi_68[53], regroupV0_hi_68[21]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_24 = {regroupV0_hi_68[117], regroupV0_hi_68[85]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_58 = {regroupV0_hi_lo_lo_lo_hi_24, regroupV0_hi_lo_lo_lo_lo_24};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_24 = {regroupV0_hi_68[181], regroupV0_hi_68[149]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_24 = {regroupV0_hi_68[245], regroupV0_hi_68[213]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_58 = {regroupV0_hi_lo_lo_hi_hi_24, regroupV0_hi_lo_lo_hi_lo_24};
  wire [7:0]         regroupV0_hi_lo_lo_90 = {regroupV0_hi_lo_lo_hi_58, regroupV0_hi_lo_lo_lo_58};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_24 = {regroupV0_hi_68[309], regroupV0_hi_68[277]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_24 = {regroupV0_hi_68[373], regroupV0_hi_68[341]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_58 = {regroupV0_hi_lo_hi_lo_hi_24, regroupV0_hi_lo_hi_lo_lo_24};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_24 = {regroupV0_hi_68[437], regroupV0_hi_68[405]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_24 = {regroupV0_hi_68[501], regroupV0_hi_68[469]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_58 = {regroupV0_hi_lo_hi_hi_hi_24, regroupV0_hi_lo_hi_hi_lo_24};
  wire [7:0]         regroupV0_hi_lo_hi_90 = {regroupV0_hi_lo_hi_hi_58, regroupV0_hi_lo_hi_lo_58};
  wire [15:0]        regroupV0_hi_lo_90 = {regroupV0_hi_lo_hi_90, regroupV0_hi_lo_lo_90};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_24 = {regroupV0_hi_68[565], regroupV0_hi_68[533]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_24 = {regroupV0_hi_68[629], regroupV0_hi_68[597]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_58 = {regroupV0_hi_hi_lo_lo_hi_24, regroupV0_hi_hi_lo_lo_lo_24};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_24 = {regroupV0_hi_68[693], regroupV0_hi_68[661]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_24 = {regroupV0_hi_68[757], regroupV0_hi_68[725]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_58 = {regroupV0_hi_hi_lo_hi_hi_24, regroupV0_hi_hi_lo_hi_lo_24};
  wire [7:0]         regroupV0_hi_hi_lo_90 = {regroupV0_hi_hi_lo_hi_58, regroupV0_hi_hi_lo_lo_58};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_24 = {regroupV0_hi_68[821], regroupV0_hi_68[789]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_24 = {regroupV0_hi_68[885], regroupV0_hi_68[853]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_58 = {regroupV0_hi_hi_hi_lo_hi_24, regroupV0_hi_hi_hi_lo_lo_24};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_24 = {regroupV0_hi_68[949], regroupV0_hi_68[917]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_24 = {regroupV0_hi_68[1013], regroupV0_hi_68[981]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_58 = {regroupV0_hi_hi_hi_hi_hi_24, regroupV0_hi_hi_hi_hi_lo_24};
  wire [7:0]         regroupV0_hi_hi_hi_90 = {regroupV0_hi_hi_hi_hi_58, regroupV0_hi_hi_hi_lo_58};
  wire [15:0]        regroupV0_hi_hi_90 = {regroupV0_hi_hi_hi_90, regroupV0_hi_hi_lo_90};
  wire [31:0]        regroupV0_hi_90 = {regroupV0_hi_hi_90, regroupV0_hi_lo_90};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_25 = {regroupV0_lo_68[54], regroupV0_lo_68[22]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_25 = {regroupV0_lo_68[118], regroupV0_lo_68[86]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_59 = {regroupV0_lo_lo_lo_lo_hi_25, regroupV0_lo_lo_lo_lo_lo_25};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_25 = {regroupV0_lo_68[182], regroupV0_lo_68[150]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_25 = {regroupV0_lo_68[246], regroupV0_lo_68[214]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_59 = {regroupV0_lo_lo_lo_hi_hi_25, regroupV0_lo_lo_lo_hi_lo_25};
  wire [7:0]         regroupV0_lo_lo_lo_91 = {regroupV0_lo_lo_lo_hi_59, regroupV0_lo_lo_lo_lo_59};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_25 = {regroupV0_lo_68[310], regroupV0_lo_68[278]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_25 = {regroupV0_lo_68[374], regroupV0_lo_68[342]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_59 = {regroupV0_lo_lo_hi_lo_hi_25, regroupV0_lo_lo_hi_lo_lo_25};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_25 = {regroupV0_lo_68[438], regroupV0_lo_68[406]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_25 = {regroupV0_lo_68[502], regroupV0_lo_68[470]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_59 = {regroupV0_lo_lo_hi_hi_hi_25, regroupV0_lo_lo_hi_hi_lo_25};
  wire [7:0]         regroupV0_lo_lo_hi_91 = {regroupV0_lo_lo_hi_hi_59, regroupV0_lo_lo_hi_lo_59};
  wire [15:0]        regroupV0_lo_lo_91 = {regroupV0_lo_lo_hi_91, regroupV0_lo_lo_lo_91};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_25 = {regroupV0_lo_68[566], regroupV0_lo_68[534]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_25 = {regroupV0_lo_68[630], regroupV0_lo_68[598]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_59 = {regroupV0_lo_hi_lo_lo_hi_25, regroupV0_lo_hi_lo_lo_lo_25};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_25 = {regroupV0_lo_68[694], regroupV0_lo_68[662]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_25 = {regroupV0_lo_68[758], regroupV0_lo_68[726]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_59 = {regroupV0_lo_hi_lo_hi_hi_25, regroupV0_lo_hi_lo_hi_lo_25};
  wire [7:0]         regroupV0_lo_hi_lo_91 = {regroupV0_lo_hi_lo_hi_59, regroupV0_lo_hi_lo_lo_59};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_25 = {regroupV0_lo_68[822], regroupV0_lo_68[790]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_25 = {regroupV0_lo_68[886], regroupV0_lo_68[854]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_59 = {regroupV0_lo_hi_hi_lo_hi_25, regroupV0_lo_hi_hi_lo_lo_25};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_25 = {regroupV0_lo_68[950], regroupV0_lo_68[918]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_25 = {regroupV0_lo_68[1014], regroupV0_lo_68[982]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_59 = {regroupV0_lo_hi_hi_hi_hi_25, regroupV0_lo_hi_hi_hi_lo_25};
  wire [7:0]         regroupV0_lo_hi_hi_91 = {regroupV0_lo_hi_hi_hi_59, regroupV0_lo_hi_hi_lo_59};
  wire [15:0]        regroupV0_lo_hi_91 = {regroupV0_lo_hi_hi_91, regroupV0_lo_hi_lo_91};
  wire [31:0]        regroupV0_lo_91 = {regroupV0_lo_hi_91, regroupV0_lo_lo_91};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_25 = {regroupV0_hi_68[54], regroupV0_hi_68[22]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_25 = {regroupV0_hi_68[118], regroupV0_hi_68[86]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_59 = {regroupV0_hi_lo_lo_lo_hi_25, regroupV0_hi_lo_lo_lo_lo_25};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_25 = {regroupV0_hi_68[182], regroupV0_hi_68[150]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_25 = {regroupV0_hi_68[246], regroupV0_hi_68[214]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_59 = {regroupV0_hi_lo_lo_hi_hi_25, regroupV0_hi_lo_lo_hi_lo_25};
  wire [7:0]         regroupV0_hi_lo_lo_91 = {regroupV0_hi_lo_lo_hi_59, regroupV0_hi_lo_lo_lo_59};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_25 = {regroupV0_hi_68[310], regroupV0_hi_68[278]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_25 = {regroupV0_hi_68[374], regroupV0_hi_68[342]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_59 = {regroupV0_hi_lo_hi_lo_hi_25, regroupV0_hi_lo_hi_lo_lo_25};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_25 = {regroupV0_hi_68[438], regroupV0_hi_68[406]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_25 = {regroupV0_hi_68[502], regroupV0_hi_68[470]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_59 = {regroupV0_hi_lo_hi_hi_hi_25, regroupV0_hi_lo_hi_hi_lo_25};
  wire [7:0]         regroupV0_hi_lo_hi_91 = {regroupV0_hi_lo_hi_hi_59, regroupV0_hi_lo_hi_lo_59};
  wire [15:0]        regroupV0_hi_lo_91 = {regroupV0_hi_lo_hi_91, regroupV0_hi_lo_lo_91};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_25 = {regroupV0_hi_68[566], regroupV0_hi_68[534]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_25 = {regroupV0_hi_68[630], regroupV0_hi_68[598]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_59 = {regroupV0_hi_hi_lo_lo_hi_25, regroupV0_hi_hi_lo_lo_lo_25};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_25 = {regroupV0_hi_68[694], regroupV0_hi_68[662]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_25 = {regroupV0_hi_68[758], regroupV0_hi_68[726]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_59 = {regroupV0_hi_hi_lo_hi_hi_25, regroupV0_hi_hi_lo_hi_lo_25};
  wire [7:0]         regroupV0_hi_hi_lo_91 = {regroupV0_hi_hi_lo_hi_59, regroupV0_hi_hi_lo_lo_59};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_25 = {regroupV0_hi_68[822], regroupV0_hi_68[790]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_25 = {regroupV0_hi_68[886], regroupV0_hi_68[854]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_59 = {regroupV0_hi_hi_hi_lo_hi_25, regroupV0_hi_hi_hi_lo_lo_25};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_25 = {regroupV0_hi_68[950], regroupV0_hi_68[918]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_25 = {regroupV0_hi_68[1014], regroupV0_hi_68[982]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_59 = {regroupV0_hi_hi_hi_hi_hi_25, regroupV0_hi_hi_hi_hi_lo_25};
  wire [7:0]         regroupV0_hi_hi_hi_91 = {regroupV0_hi_hi_hi_hi_59, regroupV0_hi_hi_hi_lo_59};
  wire [15:0]        regroupV0_hi_hi_91 = {regroupV0_hi_hi_hi_91, regroupV0_hi_hi_lo_91};
  wire [31:0]        regroupV0_hi_91 = {regroupV0_hi_hi_91, regroupV0_hi_lo_91};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_26 = {regroupV0_lo_68[55], regroupV0_lo_68[23]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_26 = {regroupV0_lo_68[119], regroupV0_lo_68[87]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_60 = {regroupV0_lo_lo_lo_lo_hi_26, regroupV0_lo_lo_lo_lo_lo_26};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_26 = {regroupV0_lo_68[183], regroupV0_lo_68[151]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_26 = {regroupV0_lo_68[247], regroupV0_lo_68[215]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_60 = {regroupV0_lo_lo_lo_hi_hi_26, regroupV0_lo_lo_lo_hi_lo_26};
  wire [7:0]         regroupV0_lo_lo_lo_92 = {regroupV0_lo_lo_lo_hi_60, regroupV0_lo_lo_lo_lo_60};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_26 = {regroupV0_lo_68[311], regroupV0_lo_68[279]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_26 = {regroupV0_lo_68[375], regroupV0_lo_68[343]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_60 = {regroupV0_lo_lo_hi_lo_hi_26, regroupV0_lo_lo_hi_lo_lo_26};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_26 = {regroupV0_lo_68[439], regroupV0_lo_68[407]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_26 = {regroupV0_lo_68[503], regroupV0_lo_68[471]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_60 = {regroupV0_lo_lo_hi_hi_hi_26, regroupV0_lo_lo_hi_hi_lo_26};
  wire [7:0]         regroupV0_lo_lo_hi_92 = {regroupV0_lo_lo_hi_hi_60, regroupV0_lo_lo_hi_lo_60};
  wire [15:0]        regroupV0_lo_lo_92 = {regroupV0_lo_lo_hi_92, regroupV0_lo_lo_lo_92};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_26 = {regroupV0_lo_68[567], regroupV0_lo_68[535]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_26 = {regroupV0_lo_68[631], regroupV0_lo_68[599]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_60 = {regroupV0_lo_hi_lo_lo_hi_26, regroupV0_lo_hi_lo_lo_lo_26};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_26 = {regroupV0_lo_68[695], regroupV0_lo_68[663]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_26 = {regroupV0_lo_68[759], regroupV0_lo_68[727]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_60 = {regroupV0_lo_hi_lo_hi_hi_26, regroupV0_lo_hi_lo_hi_lo_26};
  wire [7:0]         regroupV0_lo_hi_lo_92 = {regroupV0_lo_hi_lo_hi_60, regroupV0_lo_hi_lo_lo_60};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_26 = {regroupV0_lo_68[823], regroupV0_lo_68[791]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_26 = {regroupV0_lo_68[887], regroupV0_lo_68[855]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_60 = {regroupV0_lo_hi_hi_lo_hi_26, regroupV0_lo_hi_hi_lo_lo_26};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_26 = {regroupV0_lo_68[951], regroupV0_lo_68[919]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_26 = {regroupV0_lo_68[1015], regroupV0_lo_68[983]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_60 = {regroupV0_lo_hi_hi_hi_hi_26, regroupV0_lo_hi_hi_hi_lo_26};
  wire [7:0]         regroupV0_lo_hi_hi_92 = {regroupV0_lo_hi_hi_hi_60, regroupV0_lo_hi_hi_lo_60};
  wire [15:0]        regroupV0_lo_hi_92 = {regroupV0_lo_hi_hi_92, regroupV0_lo_hi_lo_92};
  wire [31:0]        regroupV0_lo_92 = {regroupV0_lo_hi_92, regroupV0_lo_lo_92};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_26 = {regroupV0_hi_68[55], regroupV0_hi_68[23]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_26 = {regroupV0_hi_68[119], regroupV0_hi_68[87]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_60 = {regroupV0_hi_lo_lo_lo_hi_26, regroupV0_hi_lo_lo_lo_lo_26};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_26 = {regroupV0_hi_68[183], regroupV0_hi_68[151]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_26 = {regroupV0_hi_68[247], regroupV0_hi_68[215]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_60 = {regroupV0_hi_lo_lo_hi_hi_26, regroupV0_hi_lo_lo_hi_lo_26};
  wire [7:0]         regroupV0_hi_lo_lo_92 = {regroupV0_hi_lo_lo_hi_60, regroupV0_hi_lo_lo_lo_60};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_26 = {regroupV0_hi_68[311], regroupV0_hi_68[279]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_26 = {regroupV0_hi_68[375], regroupV0_hi_68[343]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_60 = {regroupV0_hi_lo_hi_lo_hi_26, regroupV0_hi_lo_hi_lo_lo_26};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_26 = {regroupV0_hi_68[439], regroupV0_hi_68[407]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_26 = {regroupV0_hi_68[503], regroupV0_hi_68[471]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_60 = {regroupV0_hi_lo_hi_hi_hi_26, regroupV0_hi_lo_hi_hi_lo_26};
  wire [7:0]         regroupV0_hi_lo_hi_92 = {regroupV0_hi_lo_hi_hi_60, regroupV0_hi_lo_hi_lo_60};
  wire [15:0]        regroupV0_hi_lo_92 = {regroupV0_hi_lo_hi_92, regroupV0_hi_lo_lo_92};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_26 = {regroupV0_hi_68[567], regroupV0_hi_68[535]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_26 = {regroupV0_hi_68[631], regroupV0_hi_68[599]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_60 = {regroupV0_hi_hi_lo_lo_hi_26, regroupV0_hi_hi_lo_lo_lo_26};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_26 = {regroupV0_hi_68[695], regroupV0_hi_68[663]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_26 = {regroupV0_hi_68[759], regroupV0_hi_68[727]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_60 = {regroupV0_hi_hi_lo_hi_hi_26, regroupV0_hi_hi_lo_hi_lo_26};
  wire [7:0]         regroupV0_hi_hi_lo_92 = {regroupV0_hi_hi_lo_hi_60, regroupV0_hi_hi_lo_lo_60};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_26 = {regroupV0_hi_68[823], regroupV0_hi_68[791]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_26 = {regroupV0_hi_68[887], regroupV0_hi_68[855]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_60 = {regroupV0_hi_hi_hi_lo_hi_26, regroupV0_hi_hi_hi_lo_lo_26};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_26 = {regroupV0_hi_68[951], regroupV0_hi_68[919]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_26 = {regroupV0_hi_68[1015], regroupV0_hi_68[983]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_60 = {regroupV0_hi_hi_hi_hi_hi_26, regroupV0_hi_hi_hi_hi_lo_26};
  wire [7:0]         regroupV0_hi_hi_hi_92 = {regroupV0_hi_hi_hi_hi_60, regroupV0_hi_hi_hi_lo_60};
  wire [15:0]        regroupV0_hi_hi_92 = {regroupV0_hi_hi_hi_92, regroupV0_hi_hi_lo_92};
  wire [31:0]        regroupV0_hi_92 = {regroupV0_hi_hi_92, regroupV0_hi_lo_92};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_27 = {regroupV0_lo_68[56], regroupV0_lo_68[24]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_27 = {regroupV0_lo_68[120], regroupV0_lo_68[88]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_61 = {regroupV0_lo_lo_lo_lo_hi_27, regroupV0_lo_lo_lo_lo_lo_27};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_27 = {regroupV0_lo_68[184], regroupV0_lo_68[152]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_27 = {regroupV0_lo_68[248], regroupV0_lo_68[216]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_61 = {regroupV0_lo_lo_lo_hi_hi_27, regroupV0_lo_lo_lo_hi_lo_27};
  wire [7:0]         regroupV0_lo_lo_lo_93 = {regroupV0_lo_lo_lo_hi_61, regroupV0_lo_lo_lo_lo_61};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_27 = {regroupV0_lo_68[312], regroupV0_lo_68[280]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_27 = {regroupV0_lo_68[376], regroupV0_lo_68[344]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_61 = {regroupV0_lo_lo_hi_lo_hi_27, regroupV0_lo_lo_hi_lo_lo_27};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_27 = {regroupV0_lo_68[440], regroupV0_lo_68[408]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_27 = {regroupV0_lo_68[504], regroupV0_lo_68[472]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_61 = {regroupV0_lo_lo_hi_hi_hi_27, regroupV0_lo_lo_hi_hi_lo_27};
  wire [7:0]         regroupV0_lo_lo_hi_93 = {regroupV0_lo_lo_hi_hi_61, regroupV0_lo_lo_hi_lo_61};
  wire [15:0]        regroupV0_lo_lo_93 = {regroupV0_lo_lo_hi_93, regroupV0_lo_lo_lo_93};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_27 = {regroupV0_lo_68[568], regroupV0_lo_68[536]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_27 = {regroupV0_lo_68[632], regroupV0_lo_68[600]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_61 = {regroupV0_lo_hi_lo_lo_hi_27, regroupV0_lo_hi_lo_lo_lo_27};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_27 = {regroupV0_lo_68[696], regroupV0_lo_68[664]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_27 = {regroupV0_lo_68[760], regroupV0_lo_68[728]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_61 = {regroupV0_lo_hi_lo_hi_hi_27, regroupV0_lo_hi_lo_hi_lo_27};
  wire [7:0]         regroupV0_lo_hi_lo_93 = {regroupV0_lo_hi_lo_hi_61, regroupV0_lo_hi_lo_lo_61};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_27 = {regroupV0_lo_68[824], regroupV0_lo_68[792]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_27 = {regroupV0_lo_68[888], regroupV0_lo_68[856]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_61 = {regroupV0_lo_hi_hi_lo_hi_27, regroupV0_lo_hi_hi_lo_lo_27};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_27 = {regroupV0_lo_68[952], regroupV0_lo_68[920]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_27 = {regroupV0_lo_68[1016], regroupV0_lo_68[984]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_61 = {regroupV0_lo_hi_hi_hi_hi_27, regroupV0_lo_hi_hi_hi_lo_27};
  wire [7:0]         regroupV0_lo_hi_hi_93 = {regroupV0_lo_hi_hi_hi_61, regroupV0_lo_hi_hi_lo_61};
  wire [15:0]        regroupV0_lo_hi_93 = {regroupV0_lo_hi_hi_93, regroupV0_lo_hi_lo_93};
  wire [31:0]        regroupV0_lo_93 = {regroupV0_lo_hi_93, regroupV0_lo_lo_93};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_27 = {regroupV0_hi_68[56], regroupV0_hi_68[24]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_27 = {regroupV0_hi_68[120], regroupV0_hi_68[88]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_61 = {regroupV0_hi_lo_lo_lo_hi_27, regroupV0_hi_lo_lo_lo_lo_27};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_27 = {regroupV0_hi_68[184], regroupV0_hi_68[152]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_27 = {regroupV0_hi_68[248], regroupV0_hi_68[216]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_61 = {regroupV0_hi_lo_lo_hi_hi_27, regroupV0_hi_lo_lo_hi_lo_27};
  wire [7:0]         regroupV0_hi_lo_lo_93 = {regroupV0_hi_lo_lo_hi_61, regroupV0_hi_lo_lo_lo_61};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_27 = {regroupV0_hi_68[312], regroupV0_hi_68[280]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_27 = {regroupV0_hi_68[376], regroupV0_hi_68[344]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_61 = {regroupV0_hi_lo_hi_lo_hi_27, regroupV0_hi_lo_hi_lo_lo_27};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_27 = {regroupV0_hi_68[440], regroupV0_hi_68[408]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_27 = {regroupV0_hi_68[504], regroupV0_hi_68[472]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_61 = {regroupV0_hi_lo_hi_hi_hi_27, regroupV0_hi_lo_hi_hi_lo_27};
  wire [7:0]         regroupV0_hi_lo_hi_93 = {regroupV0_hi_lo_hi_hi_61, regroupV0_hi_lo_hi_lo_61};
  wire [15:0]        regroupV0_hi_lo_93 = {regroupV0_hi_lo_hi_93, regroupV0_hi_lo_lo_93};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_27 = {regroupV0_hi_68[568], regroupV0_hi_68[536]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_27 = {regroupV0_hi_68[632], regroupV0_hi_68[600]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_61 = {regroupV0_hi_hi_lo_lo_hi_27, regroupV0_hi_hi_lo_lo_lo_27};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_27 = {regroupV0_hi_68[696], regroupV0_hi_68[664]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_27 = {regroupV0_hi_68[760], regroupV0_hi_68[728]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_61 = {regroupV0_hi_hi_lo_hi_hi_27, regroupV0_hi_hi_lo_hi_lo_27};
  wire [7:0]         regroupV0_hi_hi_lo_93 = {regroupV0_hi_hi_lo_hi_61, regroupV0_hi_hi_lo_lo_61};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_27 = {regroupV0_hi_68[824], regroupV0_hi_68[792]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_27 = {regroupV0_hi_68[888], regroupV0_hi_68[856]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_61 = {regroupV0_hi_hi_hi_lo_hi_27, regroupV0_hi_hi_hi_lo_lo_27};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_27 = {regroupV0_hi_68[952], regroupV0_hi_68[920]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_27 = {regroupV0_hi_68[1016], regroupV0_hi_68[984]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_61 = {regroupV0_hi_hi_hi_hi_hi_27, regroupV0_hi_hi_hi_hi_lo_27};
  wire [7:0]         regroupV0_hi_hi_hi_93 = {regroupV0_hi_hi_hi_hi_61, regroupV0_hi_hi_hi_lo_61};
  wire [15:0]        regroupV0_hi_hi_93 = {regroupV0_hi_hi_hi_93, regroupV0_hi_hi_lo_93};
  wire [31:0]        regroupV0_hi_93 = {regroupV0_hi_hi_93, regroupV0_hi_lo_93};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_28 = {regroupV0_lo_68[57], regroupV0_lo_68[25]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_28 = {regroupV0_lo_68[121], regroupV0_lo_68[89]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_62 = {regroupV0_lo_lo_lo_lo_hi_28, regroupV0_lo_lo_lo_lo_lo_28};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_28 = {regroupV0_lo_68[185], regroupV0_lo_68[153]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_28 = {regroupV0_lo_68[249], regroupV0_lo_68[217]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_62 = {regroupV0_lo_lo_lo_hi_hi_28, regroupV0_lo_lo_lo_hi_lo_28};
  wire [7:0]         regroupV0_lo_lo_lo_94 = {regroupV0_lo_lo_lo_hi_62, regroupV0_lo_lo_lo_lo_62};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_28 = {regroupV0_lo_68[313], regroupV0_lo_68[281]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_28 = {regroupV0_lo_68[377], regroupV0_lo_68[345]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_62 = {regroupV0_lo_lo_hi_lo_hi_28, regroupV0_lo_lo_hi_lo_lo_28};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_28 = {regroupV0_lo_68[441], regroupV0_lo_68[409]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_28 = {regroupV0_lo_68[505], regroupV0_lo_68[473]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_62 = {regroupV0_lo_lo_hi_hi_hi_28, regroupV0_lo_lo_hi_hi_lo_28};
  wire [7:0]         regroupV0_lo_lo_hi_94 = {regroupV0_lo_lo_hi_hi_62, regroupV0_lo_lo_hi_lo_62};
  wire [15:0]        regroupV0_lo_lo_94 = {regroupV0_lo_lo_hi_94, regroupV0_lo_lo_lo_94};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_28 = {regroupV0_lo_68[569], regroupV0_lo_68[537]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_28 = {regroupV0_lo_68[633], regroupV0_lo_68[601]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_62 = {regroupV0_lo_hi_lo_lo_hi_28, regroupV0_lo_hi_lo_lo_lo_28};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_28 = {regroupV0_lo_68[697], regroupV0_lo_68[665]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_28 = {regroupV0_lo_68[761], regroupV0_lo_68[729]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_62 = {regroupV0_lo_hi_lo_hi_hi_28, regroupV0_lo_hi_lo_hi_lo_28};
  wire [7:0]         regroupV0_lo_hi_lo_94 = {regroupV0_lo_hi_lo_hi_62, regroupV0_lo_hi_lo_lo_62};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_28 = {regroupV0_lo_68[825], regroupV0_lo_68[793]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_28 = {regroupV0_lo_68[889], regroupV0_lo_68[857]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_62 = {regroupV0_lo_hi_hi_lo_hi_28, regroupV0_lo_hi_hi_lo_lo_28};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_28 = {regroupV0_lo_68[953], regroupV0_lo_68[921]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_28 = {regroupV0_lo_68[1017], regroupV0_lo_68[985]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_62 = {regroupV0_lo_hi_hi_hi_hi_28, regroupV0_lo_hi_hi_hi_lo_28};
  wire [7:0]         regroupV0_lo_hi_hi_94 = {regroupV0_lo_hi_hi_hi_62, regroupV0_lo_hi_hi_lo_62};
  wire [15:0]        regroupV0_lo_hi_94 = {regroupV0_lo_hi_hi_94, regroupV0_lo_hi_lo_94};
  wire [31:0]        regroupV0_lo_94 = {regroupV0_lo_hi_94, regroupV0_lo_lo_94};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_28 = {regroupV0_hi_68[57], regroupV0_hi_68[25]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_28 = {regroupV0_hi_68[121], regroupV0_hi_68[89]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_62 = {regroupV0_hi_lo_lo_lo_hi_28, regroupV0_hi_lo_lo_lo_lo_28};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_28 = {regroupV0_hi_68[185], regroupV0_hi_68[153]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_28 = {regroupV0_hi_68[249], regroupV0_hi_68[217]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_62 = {regroupV0_hi_lo_lo_hi_hi_28, regroupV0_hi_lo_lo_hi_lo_28};
  wire [7:0]         regroupV0_hi_lo_lo_94 = {regroupV0_hi_lo_lo_hi_62, regroupV0_hi_lo_lo_lo_62};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_28 = {regroupV0_hi_68[313], regroupV0_hi_68[281]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_28 = {regroupV0_hi_68[377], regroupV0_hi_68[345]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_62 = {regroupV0_hi_lo_hi_lo_hi_28, regroupV0_hi_lo_hi_lo_lo_28};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_28 = {regroupV0_hi_68[441], regroupV0_hi_68[409]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_28 = {regroupV0_hi_68[505], regroupV0_hi_68[473]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_62 = {regroupV0_hi_lo_hi_hi_hi_28, regroupV0_hi_lo_hi_hi_lo_28};
  wire [7:0]         regroupV0_hi_lo_hi_94 = {regroupV0_hi_lo_hi_hi_62, regroupV0_hi_lo_hi_lo_62};
  wire [15:0]        regroupV0_hi_lo_94 = {regroupV0_hi_lo_hi_94, regroupV0_hi_lo_lo_94};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_28 = {regroupV0_hi_68[569], regroupV0_hi_68[537]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_28 = {regroupV0_hi_68[633], regroupV0_hi_68[601]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_62 = {regroupV0_hi_hi_lo_lo_hi_28, regroupV0_hi_hi_lo_lo_lo_28};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_28 = {regroupV0_hi_68[697], regroupV0_hi_68[665]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_28 = {regroupV0_hi_68[761], regroupV0_hi_68[729]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_62 = {regroupV0_hi_hi_lo_hi_hi_28, regroupV0_hi_hi_lo_hi_lo_28};
  wire [7:0]         regroupV0_hi_hi_lo_94 = {regroupV0_hi_hi_lo_hi_62, regroupV0_hi_hi_lo_lo_62};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_28 = {regroupV0_hi_68[825], regroupV0_hi_68[793]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_28 = {regroupV0_hi_68[889], regroupV0_hi_68[857]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_62 = {regroupV0_hi_hi_hi_lo_hi_28, regroupV0_hi_hi_hi_lo_lo_28};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_28 = {regroupV0_hi_68[953], regroupV0_hi_68[921]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_28 = {regroupV0_hi_68[1017], regroupV0_hi_68[985]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_62 = {regroupV0_hi_hi_hi_hi_hi_28, regroupV0_hi_hi_hi_hi_lo_28};
  wire [7:0]         regroupV0_hi_hi_hi_94 = {regroupV0_hi_hi_hi_hi_62, regroupV0_hi_hi_hi_lo_62};
  wire [15:0]        regroupV0_hi_hi_94 = {regroupV0_hi_hi_hi_94, regroupV0_hi_hi_lo_94};
  wire [31:0]        regroupV0_hi_94 = {regroupV0_hi_hi_94, regroupV0_hi_lo_94};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_29 = {regroupV0_lo_68[58], regroupV0_lo_68[26]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_29 = {regroupV0_lo_68[122], regroupV0_lo_68[90]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_63 = {regroupV0_lo_lo_lo_lo_hi_29, regroupV0_lo_lo_lo_lo_lo_29};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_29 = {regroupV0_lo_68[186], regroupV0_lo_68[154]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_29 = {regroupV0_lo_68[250], regroupV0_lo_68[218]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_63 = {regroupV0_lo_lo_lo_hi_hi_29, regroupV0_lo_lo_lo_hi_lo_29};
  wire [7:0]         regroupV0_lo_lo_lo_95 = {regroupV0_lo_lo_lo_hi_63, regroupV0_lo_lo_lo_lo_63};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_29 = {regroupV0_lo_68[314], regroupV0_lo_68[282]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_29 = {regroupV0_lo_68[378], regroupV0_lo_68[346]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_63 = {regroupV0_lo_lo_hi_lo_hi_29, regroupV0_lo_lo_hi_lo_lo_29};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_29 = {regroupV0_lo_68[442], regroupV0_lo_68[410]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_29 = {regroupV0_lo_68[506], regroupV0_lo_68[474]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_63 = {regroupV0_lo_lo_hi_hi_hi_29, regroupV0_lo_lo_hi_hi_lo_29};
  wire [7:0]         regroupV0_lo_lo_hi_95 = {regroupV0_lo_lo_hi_hi_63, regroupV0_lo_lo_hi_lo_63};
  wire [15:0]        regroupV0_lo_lo_95 = {regroupV0_lo_lo_hi_95, regroupV0_lo_lo_lo_95};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_29 = {regroupV0_lo_68[570], regroupV0_lo_68[538]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_29 = {regroupV0_lo_68[634], regroupV0_lo_68[602]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_63 = {regroupV0_lo_hi_lo_lo_hi_29, regroupV0_lo_hi_lo_lo_lo_29};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_29 = {regroupV0_lo_68[698], regroupV0_lo_68[666]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_29 = {regroupV0_lo_68[762], regroupV0_lo_68[730]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_63 = {regroupV0_lo_hi_lo_hi_hi_29, regroupV0_lo_hi_lo_hi_lo_29};
  wire [7:0]         regroupV0_lo_hi_lo_95 = {regroupV0_lo_hi_lo_hi_63, regroupV0_lo_hi_lo_lo_63};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_29 = {regroupV0_lo_68[826], regroupV0_lo_68[794]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_29 = {regroupV0_lo_68[890], regroupV0_lo_68[858]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_63 = {regroupV0_lo_hi_hi_lo_hi_29, regroupV0_lo_hi_hi_lo_lo_29};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_29 = {regroupV0_lo_68[954], regroupV0_lo_68[922]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_29 = {regroupV0_lo_68[1018], regroupV0_lo_68[986]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_63 = {regroupV0_lo_hi_hi_hi_hi_29, regroupV0_lo_hi_hi_hi_lo_29};
  wire [7:0]         regroupV0_lo_hi_hi_95 = {regroupV0_lo_hi_hi_hi_63, regroupV0_lo_hi_hi_lo_63};
  wire [15:0]        regroupV0_lo_hi_95 = {regroupV0_lo_hi_hi_95, regroupV0_lo_hi_lo_95};
  wire [31:0]        regroupV0_lo_95 = {regroupV0_lo_hi_95, regroupV0_lo_lo_95};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_29 = {regroupV0_hi_68[58], regroupV0_hi_68[26]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_29 = {regroupV0_hi_68[122], regroupV0_hi_68[90]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_63 = {regroupV0_hi_lo_lo_lo_hi_29, regroupV0_hi_lo_lo_lo_lo_29};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_29 = {regroupV0_hi_68[186], regroupV0_hi_68[154]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_29 = {regroupV0_hi_68[250], regroupV0_hi_68[218]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_63 = {regroupV0_hi_lo_lo_hi_hi_29, regroupV0_hi_lo_lo_hi_lo_29};
  wire [7:0]         regroupV0_hi_lo_lo_95 = {regroupV0_hi_lo_lo_hi_63, regroupV0_hi_lo_lo_lo_63};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_29 = {regroupV0_hi_68[314], regroupV0_hi_68[282]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_29 = {regroupV0_hi_68[378], regroupV0_hi_68[346]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_63 = {regroupV0_hi_lo_hi_lo_hi_29, regroupV0_hi_lo_hi_lo_lo_29};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_29 = {regroupV0_hi_68[442], regroupV0_hi_68[410]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_29 = {regroupV0_hi_68[506], regroupV0_hi_68[474]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_63 = {regroupV0_hi_lo_hi_hi_hi_29, regroupV0_hi_lo_hi_hi_lo_29};
  wire [7:0]         regroupV0_hi_lo_hi_95 = {regroupV0_hi_lo_hi_hi_63, regroupV0_hi_lo_hi_lo_63};
  wire [15:0]        regroupV0_hi_lo_95 = {regroupV0_hi_lo_hi_95, regroupV0_hi_lo_lo_95};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_29 = {regroupV0_hi_68[570], regroupV0_hi_68[538]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_29 = {regroupV0_hi_68[634], regroupV0_hi_68[602]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_63 = {regroupV0_hi_hi_lo_lo_hi_29, regroupV0_hi_hi_lo_lo_lo_29};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_29 = {regroupV0_hi_68[698], regroupV0_hi_68[666]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_29 = {regroupV0_hi_68[762], regroupV0_hi_68[730]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_63 = {regroupV0_hi_hi_lo_hi_hi_29, regroupV0_hi_hi_lo_hi_lo_29};
  wire [7:0]         regroupV0_hi_hi_lo_95 = {regroupV0_hi_hi_lo_hi_63, regroupV0_hi_hi_lo_lo_63};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_29 = {regroupV0_hi_68[826], regroupV0_hi_68[794]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_29 = {regroupV0_hi_68[890], regroupV0_hi_68[858]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_63 = {regroupV0_hi_hi_hi_lo_hi_29, regroupV0_hi_hi_hi_lo_lo_29};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_29 = {regroupV0_hi_68[954], regroupV0_hi_68[922]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_29 = {regroupV0_hi_68[1018], regroupV0_hi_68[986]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_63 = {regroupV0_hi_hi_hi_hi_hi_29, regroupV0_hi_hi_hi_hi_lo_29};
  wire [7:0]         regroupV0_hi_hi_hi_95 = {regroupV0_hi_hi_hi_hi_63, regroupV0_hi_hi_hi_lo_63};
  wire [15:0]        regroupV0_hi_hi_95 = {regroupV0_hi_hi_hi_95, regroupV0_hi_hi_lo_95};
  wire [31:0]        regroupV0_hi_95 = {regroupV0_hi_hi_95, regroupV0_hi_lo_95};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_30 = {regroupV0_lo_68[59], regroupV0_lo_68[27]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_30 = {regroupV0_lo_68[123], regroupV0_lo_68[91]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_64 = {regroupV0_lo_lo_lo_lo_hi_30, regroupV0_lo_lo_lo_lo_lo_30};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_30 = {regroupV0_lo_68[187], regroupV0_lo_68[155]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_30 = {regroupV0_lo_68[251], regroupV0_lo_68[219]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_64 = {regroupV0_lo_lo_lo_hi_hi_30, regroupV0_lo_lo_lo_hi_lo_30};
  wire [7:0]         regroupV0_lo_lo_lo_96 = {regroupV0_lo_lo_lo_hi_64, regroupV0_lo_lo_lo_lo_64};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_30 = {regroupV0_lo_68[315], regroupV0_lo_68[283]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_30 = {regroupV0_lo_68[379], regroupV0_lo_68[347]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_64 = {regroupV0_lo_lo_hi_lo_hi_30, regroupV0_lo_lo_hi_lo_lo_30};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_30 = {regroupV0_lo_68[443], regroupV0_lo_68[411]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_30 = {regroupV0_lo_68[507], regroupV0_lo_68[475]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_64 = {regroupV0_lo_lo_hi_hi_hi_30, regroupV0_lo_lo_hi_hi_lo_30};
  wire [7:0]         regroupV0_lo_lo_hi_96 = {regroupV0_lo_lo_hi_hi_64, regroupV0_lo_lo_hi_lo_64};
  wire [15:0]        regroupV0_lo_lo_96 = {regroupV0_lo_lo_hi_96, regroupV0_lo_lo_lo_96};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_30 = {regroupV0_lo_68[571], regroupV0_lo_68[539]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_30 = {regroupV0_lo_68[635], regroupV0_lo_68[603]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_64 = {regroupV0_lo_hi_lo_lo_hi_30, regroupV0_lo_hi_lo_lo_lo_30};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_30 = {regroupV0_lo_68[699], regroupV0_lo_68[667]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_30 = {regroupV0_lo_68[763], regroupV0_lo_68[731]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_64 = {regroupV0_lo_hi_lo_hi_hi_30, regroupV0_lo_hi_lo_hi_lo_30};
  wire [7:0]         regroupV0_lo_hi_lo_96 = {regroupV0_lo_hi_lo_hi_64, regroupV0_lo_hi_lo_lo_64};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_30 = {regroupV0_lo_68[827], regroupV0_lo_68[795]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_30 = {regroupV0_lo_68[891], regroupV0_lo_68[859]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_64 = {regroupV0_lo_hi_hi_lo_hi_30, regroupV0_lo_hi_hi_lo_lo_30};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_30 = {regroupV0_lo_68[955], regroupV0_lo_68[923]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_30 = {regroupV0_lo_68[1019], regroupV0_lo_68[987]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_64 = {regroupV0_lo_hi_hi_hi_hi_30, regroupV0_lo_hi_hi_hi_lo_30};
  wire [7:0]         regroupV0_lo_hi_hi_96 = {regroupV0_lo_hi_hi_hi_64, regroupV0_lo_hi_hi_lo_64};
  wire [15:0]        regroupV0_lo_hi_96 = {regroupV0_lo_hi_hi_96, regroupV0_lo_hi_lo_96};
  wire [31:0]        regroupV0_lo_96 = {regroupV0_lo_hi_96, regroupV0_lo_lo_96};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_30 = {regroupV0_hi_68[59], regroupV0_hi_68[27]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_30 = {regroupV0_hi_68[123], regroupV0_hi_68[91]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_64 = {regroupV0_hi_lo_lo_lo_hi_30, regroupV0_hi_lo_lo_lo_lo_30};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_30 = {regroupV0_hi_68[187], regroupV0_hi_68[155]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_30 = {regroupV0_hi_68[251], regroupV0_hi_68[219]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_64 = {regroupV0_hi_lo_lo_hi_hi_30, regroupV0_hi_lo_lo_hi_lo_30};
  wire [7:0]         regroupV0_hi_lo_lo_96 = {regroupV0_hi_lo_lo_hi_64, regroupV0_hi_lo_lo_lo_64};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_30 = {regroupV0_hi_68[315], regroupV0_hi_68[283]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_30 = {regroupV0_hi_68[379], regroupV0_hi_68[347]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_64 = {regroupV0_hi_lo_hi_lo_hi_30, regroupV0_hi_lo_hi_lo_lo_30};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_30 = {regroupV0_hi_68[443], regroupV0_hi_68[411]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_30 = {regroupV0_hi_68[507], regroupV0_hi_68[475]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_64 = {regroupV0_hi_lo_hi_hi_hi_30, regroupV0_hi_lo_hi_hi_lo_30};
  wire [7:0]         regroupV0_hi_lo_hi_96 = {regroupV0_hi_lo_hi_hi_64, regroupV0_hi_lo_hi_lo_64};
  wire [15:0]        regroupV0_hi_lo_96 = {regroupV0_hi_lo_hi_96, regroupV0_hi_lo_lo_96};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_30 = {regroupV0_hi_68[571], regroupV0_hi_68[539]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_30 = {regroupV0_hi_68[635], regroupV0_hi_68[603]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_64 = {regroupV0_hi_hi_lo_lo_hi_30, regroupV0_hi_hi_lo_lo_lo_30};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_30 = {regroupV0_hi_68[699], regroupV0_hi_68[667]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_30 = {regroupV0_hi_68[763], regroupV0_hi_68[731]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_64 = {regroupV0_hi_hi_lo_hi_hi_30, regroupV0_hi_hi_lo_hi_lo_30};
  wire [7:0]         regroupV0_hi_hi_lo_96 = {regroupV0_hi_hi_lo_hi_64, regroupV0_hi_hi_lo_lo_64};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_30 = {regroupV0_hi_68[827], regroupV0_hi_68[795]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_30 = {regroupV0_hi_68[891], regroupV0_hi_68[859]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_64 = {regroupV0_hi_hi_hi_lo_hi_30, regroupV0_hi_hi_hi_lo_lo_30};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_30 = {regroupV0_hi_68[955], regroupV0_hi_68[923]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_30 = {regroupV0_hi_68[1019], regroupV0_hi_68[987]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_64 = {regroupV0_hi_hi_hi_hi_hi_30, regroupV0_hi_hi_hi_hi_lo_30};
  wire [7:0]         regroupV0_hi_hi_hi_96 = {regroupV0_hi_hi_hi_hi_64, regroupV0_hi_hi_hi_lo_64};
  wire [15:0]        regroupV0_hi_hi_96 = {regroupV0_hi_hi_hi_96, regroupV0_hi_hi_lo_96};
  wire [31:0]        regroupV0_hi_96 = {regroupV0_hi_hi_96, regroupV0_hi_lo_96};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_31 = {regroupV0_lo_68[60], regroupV0_lo_68[28]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_31 = {regroupV0_lo_68[124], regroupV0_lo_68[92]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_65 = {regroupV0_lo_lo_lo_lo_hi_31, regroupV0_lo_lo_lo_lo_lo_31};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_31 = {regroupV0_lo_68[188], regroupV0_lo_68[156]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_31 = {regroupV0_lo_68[252], regroupV0_lo_68[220]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_65 = {regroupV0_lo_lo_lo_hi_hi_31, regroupV0_lo_lo_lo_hi_lo_31};
  wire [7:0]         regroupV0_lo_lo_lo_97 = {regroupV0_lo_lo_lo_hi_65, regroupV0_lo_lo_lo_lo_65};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_31 = {regroupV0_lo_68[316], regroupV0_lo_68[284]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_31 = {regroupV0_lo_68[380], regroupV0_lo_68[348]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_65 = {regroupV0_lo_lo_hi_lo_hi_31, regroupV0_lo_lo_hi_lo_lo_31};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_31 = {regroupV0_lo_68[444], regroupV0_lo_68[412]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_31 = {regroupV0_lo_68[508], regroupV0_lo_68[476]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_65 = {regroupV0_lo_lo_hi_hi_hi_31, regroupV0_lo_lo_hi_hi_lo_31};
  wire [7:0]         regroupV0_lo_lo_hi_97 = {regroupV0_lo_lo_hi_hi_65, regroupV0_lo_lo_hi_lo_65};
  wire [15:0]        regroupV0_lo_lo_97 = {regroupV0_lo_lo_hi_97, regroupV0_lo_lo_lo_97};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_31 = {regroupV0_lo_68[572], regroupV0_lo_68[540]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_31 = {regroupV0_lo_68[636], regroupV0_lo_68[604]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_65 = {regroupV0_lo_hi_lo_lo_hi_31, regroupV0_lo_hi_lo_lo_lo_31};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_31 = {regroupV0_lo_68[700], regroupV0_lo_68[668]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_31 = {regroupV0_lo_68[764], regroupV0_lo_68[732]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_65 = {regroupV0_lo_hi_lo_hi_hi_31, regroupV0_lo_hi_lo_hi_lo_31};
  wire [7:0]         regroupV0_lo_hi_lo_97 = {regroupV0_lo_hi_lo_hi_65, regroupV0_lo_hi_lo_lo_65};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_31 = {regroupV0_lo_68[828], regroupV0_lo_68[796]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_31 = {regroupV0_lo_68[892], regroupV0_lo_68[860]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_65 = {regroupV0_lo_hi_hi_lo_hi_31, regroupV0_lo_hi_hi_lo_lo_31};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_31 = {regroupV0_lo_68[956], regroupV0_lo_68[924]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_31 = {regroupV0_lo_68[1020], regroupV0_lo_68[988]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_65 = {regroupV0_lo_hi_hi_hi_hi_31, regroupV0_lo_hi_hi_hi_lo_31};
  wire [7:0]         regroupV0_lo_hi_hi_97 = {regroupV0_lo_hi_hi_hi_65, regroupV0_lo_hi_hi_lo_65};
  wire [15:0]        regroupV0_lo_hi_97 = {regroupV0_lo_hi_hi_97, regroupV0_lo_hi_lo_97};
  wire [31:0]        regroupV0_lo_97 = {regroupV0_lo_hi_97, regroupV0_lo_lo_97};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_31 = {regroupV0_hi_68[60], regroupV0_hi_68[28]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_31 = {regroupV0_hi_68[124], regroupV0_hi_68[92]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_65 = {regroupV0_hi_lo_lo_lo_hi_31, regroupV0_hi_lo_lo_lo_lo_31};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_31 = {regroupV0_hi_68[188], regroupV0_hi_68[156]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_31 = {regroupV0_hi_68[252], regroupV0_hi_68[220]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_65 = {regroupV0_hi_lo_lo_hi_hi_31, regroupV0_hi_lo_lo_hi_lo_31};
  wire [7:0]         regroupV0_hi_lo_lo_97 = {regroupV0_hi_lo_lo_hi_65, regroupV0_hi_lo_lo_lo_65};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_31 = {regroupV0_hi_68[316], regroupV0_hi_68[284]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_31 = {regroupV0_hi_68[380], regroupV0_hi_68[348]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_65 = {regroupV0_hi_lo_hi_lo_hi_31, regroupV0_hi_lo_hi_lo_lo_31};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_31 = {regroupV0_hi_68[444], regroupV0_hi_68[412]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_31 = {regroupV0_hi_68[508], regroupV0_hi_68[476]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_65 = {regroupV0_hi_lo_hi_hi_hi_31, regroupV0_hi_lo_hi_hi_lo_31};
  wire [7:0]         regroupV0_hi_lo_hi_97 = {regroupV0_hi_lo_hi_hi_65, regroupV0_hi_lo_hi_lo_65};
  wire [15:0]        regroupV0_hi_lo_97 = {regroupV0_hi_lo_hi_97, regroupV0_hi_lo_lo_97};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_31 = {regroupV0_hi_68[572], regroupV0_hi_68[540]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_31 = {regroupV0_hi_68[636], regroupV0_hi_68[604]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_65 = {regroupV0_hi_hi_lo_lo_hi_31, regroupV0_hi_hi_lo_lo_lo_31};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_31 = {regroupV0_hi_68[700], regroupV0_hi_68[668]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_31 = {regroupV0_hi_68[764], regroupV0_hi_68[732]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_65 = {regroupV0_hi_hi_lo_hi_hi_31, regroupV0_hi_hi_lo_hi_lo_31};
  wire [7:0]         regroupV0_hi_hi_lo_97 = {regroupV0_hi_hi_lo_hi_65, regroupV0_hi_hi_lo_lo_65};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_31 = {regroupV0_hi_68[828], regroupV0_hi_68[796]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_31 = {regroupV0_hi_68[892], regroupV0_hi_68[860]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_65 = {regroupV0_hi_hi_hi_lo_hi_31, regroupV0_hi_hi_hi_lo_lo_31};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_31 = {regroupV0_hi_68[956], regroupV0_hi_68[924]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_31 = {regroupV0_hi_68[1020], regroupV0_hi_68[988]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_65 = {regroupV0_hi_hi_hi_hi_hi_31, regroupV0_hi_hi_hi_hi_lo_31};
  wire [7:0]         regroupV0_hi_hi_hi_97 = {regroupV0_hi_hi_hi_hi_65, regroupV0_hi_hi_hi_lo_65};
  wire [15:0]        regroupV0_hi_hi_97 = {regroupV0_hi_hi_hi_97, regroupV0_hi_hi_lo_97};
  wire [31:0]        regroupV0_hi_97 = {regroupV0_hi_hi_97, regroupV0_hi_lo_97};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_32 = {regroupV0_lo_68[61], regroupV0_lo_68[29]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_32 = {regroupV0_lo_68[125], regroupV0_lo_68[93]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_66 = {regroupV0_lo_lo_lo_lo_hi_32, regroupV0_lo_lo_lo_lo_lo_32};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_32 = {regroupV0_lo_68[189], regroupV0_lo_68[157]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_32 = {regroupV0_lo_68[253], regroupV0_lo_68[221]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_66 = {regroupV0_lo_lo_lo_hi_hi_32, regroupV0_lo_lo_lo_hi_lo_32};
  wire [7:0]         regroupV0_lo_lo_lo_98 = {regroupV0_lo_lo_lo_hi_66, regroupV0_lo_lo_lo_lo_66};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_32 = {regroupV0_lo_68[317], regroupV0_lo_68[285]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_32 = {regroupV0_lo_68[381], regroupV0_lo_68[349]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_66 = {regroupV0_lo_lo_hi_lo_hi_32, regroupV0_lo_lo_hi_lo_lo_32};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_32 = {regroupV0_lo_68[445], regroupV0_lo_68[413]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_32 = {regroupV0_lo_68[509], regroupV0_lo_68[477]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_66 = {regroupV0_lo_lo_hi_hi_hi_32, regroupV0_lo_lo_hi_hi_lo_32};
  wire [7:0]         regroupV0_lo_lo_hi_98 = {regroupV0_lo_lo_hi_hi_66, regroupV0_lo_lo_hi_lo_66};
  wire [15:0]        regroupV0_lo_lo_98 = {regroupV0_lo_lo_hi_98, regroupV0_lo_lo_lo_98};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_32 = {regroupV0_lo_68[573], regroupV0_lo_68[541]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_32 = {regroupV0_lo_68[637], regroupV0_lo_68[605]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_66 = {regroupV0_lo_hi_lo_lo_hi_32, regroupV0_lo_hi_lo_lo_lo_32};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_32 = {regroupV0_lo_68[701], regroupV0_lo_68[669]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_32 = {regroupV0_lo_68[765], regroupV0_lo_68[733]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_66 = {regroupV0_lo_hi_lo_hi_hi_32, regroupV0_lo_hi_lo_hi_lo_32};
  wire [7:0]         regroupV0_lo_hi_lo_98 = {regroupV0_lo_hi_lo_hi_66, regroupV0_lo_hi_lo_lo_66};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_32 = {regroupV0_lo_68[829], regroupV0_lo_68[797]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_32 = {regroupV0_lo_68[893], regroupV0_lo_68[861]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_66 = {regroupV0_lo_hi_hi_lo_hi_32, regroupV0_lo_hi_hi_lo_lo_32};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_32 = {regroupV0_lo_68[957], regroupV0_lo_68[925]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_32 = {regroupV0_lo_68[1021], regroupV0_lo_68[989]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_66 = {regroupV0_lo_hi_hi_hi_hi_32, regroupV0_lo_hi_hi_hi_lo_32};
  wire [7:0]         regroupV0_lo_hi_hi_98 = {regroupV0_lo_hi_hi_hi_66, regroupV0_lo_hi_hi_lo_66};
  wire [15:0]        regroupV0_lo_hi_98 = {regroupV0_lo_hi_hi_98, regroupV0_lo_hi_lo_98};
  wire [31:0]        regroupV0_lo_98 = {regroupV0_lo_hi_98, regroupV0_lo_lo_98};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_32 = {regroupV0_hi_68[61], regroupV0_hi_68[29]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_32 = {regroupV0_hi_68[125], regroupV0_hi_68[93]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_66 = {regroupV0_hi_lo_lo_lo_hi_32, regroupV0_hi_lo_lo_lo_lo_32};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_32 = {regroupV0_hi_68[189], regroupV0_hi_68[157]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_32 = {regroupV0_hi_68[253], regroupV0_hi_68[221]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_66 = {regroupV0_hi_lo_lo_hi_hi_32, regroupV0_hi_lo_lo_hi_lo_32};
  wire [7:0]         regroupV0_hi_lo_lo_98 = {regroupV0_hi_lo_lo_hi_66, regroupV0_hi_lo_lo_lo_66};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_32 = {regroupV0_hi_68[317], regroupV0_hi_68[285]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_32 = {regroupV0_hi_68[381], regroupV0_hi_68[349]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_66 = {regroupV0_hi_lo_hi_lo_hi_32, regroupV0_hi_lo_hi_lo_lo_32};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_32 = {regroupV0_hi_68[445], regroupV0_hi_68[413]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_32 = {regroupV0_hi_68[509], regroupV0_hi_68[477]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_66 = {regroupV0_hi_lo_hi_hi_hi_32, regroupV0_hi_lo_hi_hi_lo_32};
  wire [7:0]         regroupV0_hi_lo_hi_98 = {regroupV0_hi_lo_hi_hi_66, regroupV0_hi_lo_hi_lo_66};
  wire [15:0]        regroupV0_hi_lo_98 = {regroupV0_hi_lo_hi_98, regroupV0_hi_lo_lo_98};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_32 = {regroupV0_hi_68[573], regroupV0_hi_68[541]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_32 = {regroupV0_hi_68[637], regroupV0_hi_68[605]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_66 = {regroupV0_hi_hi_lo_lo_hi_32, regroupV0_hi_hi_lo_lo_lo_32};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_32 = {regroupV0_hi_68[701], regroupV0_hi_68[669]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_32 = {regroupV0_hi_68[765], regroupV0_hi_68[733]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_66 = {regroupV0_hi_hi_lo_hi_hi_32, regroupV0_hi_hi_lo_hi_lo_32};
  wire [7:0]         regroupV0_hi_hi_lo_98 = {regroupV0_hi_hi_lo_hi_66, regroupV0_hi_hi_lo_lo_66};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_32 = {regroupV0_hi_68[829], regroupV0_hi_68[797]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_32 = {regroupV0_hi_68[893], regroupV0_hi_68[861]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_66 = {regroupV0_hi_hi_hi_lo_hi_32, regroupV0_hi_hi_hi_lo_lo_32};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_32 = {regroupV0_hi_68[957], regroupV0_hi_68[925]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_32 = {regroupV0_hi_68[1021], regroupV0_hi_68[989]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_66 = {regroupV0_hi_hi_hi_hi_hi_32, regroupV0_hi_hi_hi_hi_lo_32};
  wire [7:0]         regroupV0_hi_hi_hi_98 = {regroupV0_hi_hi_hi_hi_66, regroupV0_hi_hi_hi_lo_66};
  wire [15:0]        regroupV0_hi_hi_98 = {regroupV0_hi_hi_hi_98, regroupV0_hi_hi_lo_98};
  wire [31:0]        regroupV0_hi_98 = {regroupV0_hi_hi_98, regroupV0_hi_lo_98};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_33 = {regroupV0_lo_68[62], regroupV0_lo_68[30]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_33 = {regroupV0_lo_68[126], regroupV0_lo_68[94]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_67 = {regroupV0_lo_lo_lo_lo_hi_33, regroupV0_lo_lo_lo_lo_lo_33};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_33 = {regroupV0_lo_68[190], regroupV0_lo_68[158]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_33 = {regroupV0_lo_68[254], regroupV0_lo_68[222]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_67 = {regroupV0_lo_lo_lo_hi_hi_33, regroupV0_lo_lo_lo_hi_lo_33};
  wire [7:0]         regroupV0_lo_lo_lo_99 = {regroupV0_lo_lo_lo_hi_67, regroupV0_lo_lo_lo_lo_67};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_33 = {regroupV0_lo_68[318], regroupV0_lo_68[286]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_33 = {regroupV0_lo_68[382], regroupV0_lo_68[350]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_67 = {regroupV0_lo_lo_hi_lo_hi_33, regroupV0_lo_lo_hi_lo_lo_33};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_33 = {regroupV0_lo_68[446], regroupV0_lo_68[414]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_33 = {regroupV0_lo_68[510], regroupV0_lo_68[478]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_67 = {regroupV0_lo_lo_hi_hi_hi_33, regroupV0_lo_lo_hi_hi_lo_33};
  wire [7:0]         regroupV0_lo_lo_hi_99 = {regroupV0_lo_lo_hi_hi_67, regroupV0_lo_lo_hi_lo_67};
  wire [15:0]        regroupV0_lo_lo_99 = {regroupV0_lo_lo_hi_99, regroupV0_lo_lo_lo_99};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_33 = {regroupV0_lo_68[574], regroupV0_lo_68[542]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_33 = {regroupV0_lo_68[638], regroupV0_lo_68[606]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_67 = {regroupV0_lo_hi_lo_lo_hi_33, regroupV0_lo_hi_lo_lo_lo_33};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_33 = {regroupV0_lo_68[702], regroupV0_lo_68[670]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_33 = {regroupV0_lo_68[766], regroupV0_lo_68[734]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_67 = {regroupV0_lo_hi_lo_hi_hi_33, regroupV0_lo_hi_lo_hi_lo_33};
  wire [7:0]         regroupV0_lo_hi_lo_99 = {regroupV0_lo_hi_lo_hi_67, regroupV0_lo_hi_lo_lo_67};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_33 = {regroupV0_lo_68[830], regroupV0_lo_68[798]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_33 = {regroupV0_lo_68[894], regroupV0_lo_68[862]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_67 = {regroupV0_lo_hi_hi_lo_hi_33, regroupV0_lo_hi_hi_lo_lo_33};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_33 = {regroupV0_lo_68[958], regroupV0_lo_68[926]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_33 = {regroupV0_lo_68[1022], regroupV0_lo_68[990]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_67 = {regroupV0_lo_hi_hi_hi_hi_33, regroupV0_lo_hi_hi_hi_lo_33};
  wire [7:0]         regroupV0_lo_hi_hi_99 = {regroupV0_lo_hi_hi_hi_67, regroupV0_lo_hi_hi_lo_67};
  wire [15:0]        regroupV0_lo_hi_99 = {regroupV0_lo_hi_hi_99, regroupV0_lo_hi_lo_99};
  wire [31:0]        regroupV0_lo_99 = {regroupV0_lo_hi_99, regroupV0_lo_lo_99};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_33 = {regroupV0_hi_68[62], regroupV0_hi_68[30]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_33 = {regroupV0_hi_68[126], regroupV0_hi_68[94]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_67 = {regroupV0_hi_lo_lo_lo_hi_33, regroupV0_hi_lo_lo_lo_lo_33};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_33 = {regroupV0_hi_68[190], regroupV0_hi_68[158]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_33 = {regroupV0_hi_68[254], regroupV0_hi_68[222]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_67 = {regroupV0_hi_lo_lo_hi_hi_33, regroupV0_hi_lo_lo_hi_lo_33};
  wire [7:0]         regroupV0_hi_lo_lo_99 = {regroupV0_hi_lo_lo_hi_67, regroupV0_hi_lo_lo_lo_67};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_33 = {regroupV0_hi_68[318], regroupV0_hi_68[286]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_33 = {regroupV0_hi_68[382], regroupV0_hi_68[350]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_67 = {regroupV0_hi_lo_hi_lo_hi_33, regroupV0_hi_lo_hi_lo_lo_33};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_33 = {regroupV0_hi_68[446], regroupV0_hi_68[414]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_33 = {regroupV0_hi_68[510], regroupV0_hi_68[478]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_67 = {regroupV0_hi_lo_hi_hi_hi_33, regroupV0_hi_lo_hi_hi_lo_33};
  wire [7:0]         regroupV0_hi_lo_hi_99 = {regroupV0_hi_lo_hi_hi_67, regroupV0_hi_lo_hi_lo_67};
  wire [15:0]        regroupV0_hi_lo_99 = {regroupV0_hi_lo_hi_99, regroupV0_hi_lo_lo_99};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_33 = {regroupV0_hi_68[574], regroupV0_hi_68[542]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_33 = {regroupV0_hi_68[638], regroupV0_hi_68[606]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_67 = {regroupV0_hi_hi_lo_lo_hi_33, regroupV0_hi_hi_lo_lo_lo_33};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_33 = {regroupV0_hi_68[702], regroupV0_hi_68[670]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_33 = {regroupV0_hi_68[766], regroupV0_hi_68[734]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_67 = {regroupV0_hi_hi_lo_hi_hi_33, regroupV0_hi_hi_lo_hi_lo_33};
  wire [7:0]         regroupV0_hi_hi_lo_99 = {regroupV0_hi_hi_lo_hi_67, regroupV0_hi_hi_lo_lo_67};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_33 = {regroupV0_hi_68[830], regroupV0_hi_68[798]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_33 = {regroupV0_hi_68[894], regroupV0_hi_68[862]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_67 = {regroupV0_hi_hi_hi_lo_hi_33, regroupV0_hi_hi_hi_lo_lo_33};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_33 = {regroupV0_hi_68[958], regroupV0_hi_68[926]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_33 = {regroupV0_hi_68[1022], regroupV0_hi_68[990]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_67 = {regroupV0_hi_hi_hi_hi_hi_33, regroupV0_hi_hi_hi_hi_lo_33};
  wire [7:0]         regroupV0_hi_hi_hi_99 = {regroupV0_hi_hi_hi_hi_67, regroupV0_hi_hi_hi_lo_67};
  wire [15:0]        regroupV0_hi_hi_99 = {regroupV0_hi_hi_hi_99, regroupV0_hi_hi_lo_99};
  wire [31:0]        regroupV0_hi_99 = {regroupV0_hi_hi_99, regroupV0_hi_lo_99};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_34 = {regroupV0_lo_68[63], regroupV0_lo_68[31]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_34 = {regroupV0_lo_68[127], regroupV0_lo_68[95]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_68 = {regroupV0_lo_lo_lo_lo_hi_34, regroupV0_lo_lo_lo_lo_lo_34};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_34 = {regroupV0_lo_68[191], regroupV0_lo_68[159]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_34 = {regroupV0_lo_68[255], regroupV0_lo_68[223]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_68 = {regroupV0_lo_lo_lo_hi_hi_34, regroupV0_lo_lo_lo_hi_lo_34};
  wire [7:0]         regroupV0_lo_lo_lo_100 = {regroupV0_lo_lo_lo_hi_68, regroupV0_lo_lo_lo_lo_68};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_34 = {regroupV0_lo_68[319], regroupV0_lo_68[287]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_34 = {regroupV0_lo_68[383], regroupV0_lo_68[351]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_68 = {regroupV0_lo_lo_hi_lo_hi_34, regroupV0_lo_lo_hi_lo_lo_34};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_34 = {regroupV0_lo_68[447], regroupV0_lo_68[415]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_34 = {regroupV0_lo_68[511], regroupV0_lo_68[479]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_68 = {regroupV0_lo_lo_hi_hi_hi_34, regroupV0_lo_lo_hi_hi_lo_34};
  wire [7:0]         regroupV0_lo_lo_hi_100 = {regroupV0_lo_lo_hi_hi_68, regroupV0_lo_lo_hi_lo_68};
  wire [15:0]        regroupV0_lo_lo_100 = {regroupV0_lo_lo_hi_100, regroupV0_lo_lo_lo_100};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_34 = {regroupV0_lo_68[575], regroupV0_lo_68[543]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_34 = {regroupV0_lo_68[639], regroupV0_lo_68[607]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_68 = {regroupV0_lo_hi_lo_lo_hi_34, regroupV0_lo_hi_lo_lo_lo_34};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_34 = {regroupV0_lo_68[703], regroupV0_lo_68[671]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_34 = {regroupV0_lo_68[767], regroupV0_lo_68[735]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_68 = {regroupV0_lo_hi_lo_hi_hi_34, regroupV0_lo_hi_lo_hi_lo_34};
  wire [7:0]         regroupV0_lo_hi_lo_100 = {regroupV0_lo_hi_lo_hi_68, regroupV0_lo_hi_lo_lo_68};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_34 = {regroupV0_lo_68[831], regroupV0_lo_68[799]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_34 = {regroupV0_lo_68[895], regroupV0_lo_68[863]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_68 = {regroupV0_lo_hi_hi_lo_hi_34, regroupV0_lo_hi_hi_lo_lo_34};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_34 = {regroupV0_lo_68[959], regroupV0_lo_68[927]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_34 = {regroupV0_lo_68[1023], regroupV0_lo_68[991]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_68 = {regroupV0_lo_hi_hi_hi_hi_34, regroupV0_lo_hi_hi_hi_lo_34};
  wire [7:0]         regroupV0_lo_hi_hi_100 = {regroupV0_lo_hi_hi_hi_68, regroupV0_lo_hi_hi_lo_68};
  wire [15:0]        regroupV0_lo_hi_100 = {regroupV0_lo_hi_hi_100, regroupV0_lo_hi_lo_100};
  wire [31:0]        regroupV0_lo_100 = {regroupV0_lo_hi_100, regroupV0_lo_lo_100};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_34 = {regroupV0_hi_68[63], regroupV0_hi_68[31]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_34 = {regroupV0_hi_68[127], regroupV0_hi_68[95]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_68 = {regroupV0_hi_lo_lo_lo_hi_34, regroupV0_hi_lo_lo_lo_lo_34};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_34 = {regroupV0_hi_68[191], regroupV0_hi_68[159]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_34 = {regroupV0_hi_68[255], regroupV0_hi_68[223]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_68 = {regroupV0_hi_lo_lo_hi_hi_34, regroupV0_hi_lo_lo_hi_lo_34};
  wire [7:0]         regroupV0_hi_lo_lo_100 = {regroupV0_hi_lo_lo_hi_68, regroupV0_hi_lo_lo_lo_68};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_34 = {regroupV0_hi_68[319], regroupV0_hi_68[287]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_34 = {regroupV0_hi_68[383], regroupV0_hi_68[351]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_68 = {regroupV0_hi_lo_hi_lo_hi_34, regroupV0_hi_lo_hi_lo_lo_34};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_34 = {regroupV0_hi_68[447], regroupV0_hi_68[415]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_34 = {regroupV0_hi_68[511], regroupV0_hi_68[479]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_68 = {regroupV0_hi_lo_hi_hi_hi_34, regroupV0_hi_lo_hi_hi_lo_34};
  wire [7:0]         regroupV0_hi_lo_hi_100 = {regroupV0_hi_lo_hi_hi_68, regroupV0_hi_lo_hi_lo_68};
  wire [15:0]        regroupV0_hi_lo_100 = {regroupV0_hi_lo_hi_100, regroupV0_hi_lo_lo_100};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_34 = {regroupV0_hi_68[575], regroupV0_hi_68[543]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_34 = {regroupV0_hi_68[639], regroupV0_hi_68[607]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_68 = {regroupV0_hi_hi_lo_lo_hi_34, regroupV0_hi_hi_lo_lo_lo_34};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_34 = {regroupV0_hi_68[703], regroupV0_hi_68[671]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_34 = {regroupV0_hi_68[767], regroupV0_hi_68[735]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_68 = {regroupV0_hi_hi_lo_hi_hi_34, regroupV0_hi_hi_lo_hi_lo_34};
  wire [7:0]         regroupV0_hi_hi_lo_100 = {regroupV0_hi_hi_lo_hi_68, regroupV0_hi_hi_lo_lo_68};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_34 = {regroupV0_hi_68[831], regroupV0_hi_68[799]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_34 = {regroupV0_hi_68[895], regroupV0_hi_68[863]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_68 = {regroupV0_hi_hi_hi_lo_hi_34, regroupV0_hi_hi_hi_lo_lo_34};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_34 = {regroupV0_hi_68[959], regroupV0_hi_68[927]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_34 = {regroupV0_hi_68[1023], regroupV0_hi_68[991]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_68 = {regroupV0_hi_hi_hi_hi_hi_34, regroupV0_hi_hi_hi_hi_lo_34};
  wire [7:0]         regroupV0_hi_hi_hi_100 = {regroupV0_hi_hi_hi_hi_68, regroupV0_hi_hi_hi_lo_68};
  wire [15:0]        regroupV0_hi_hi_100 = {regroupV0_hi_hi_hi_100, regroupV0_hi_hi_lo_100};
  wire [31:0]        regroupV0_hi_100 = {regroupV0_hi_hi_100, regroupV0_hi_lo_100};
  wire [127:0]       regroupV0_lo_lo_lo_lo_69 = {regroupV0_hi_70, regroupV0_lo_70, regroupV0_hi_69, regroupV0_lo_69};
  wire [127:0]       regroupV0_lo_lo_lo_hi_69 = {regroupV0_hi_72, regroupV0_lo_72, regroupV0_hi_71, regroupV0_lo_71};
  wire [255:0]       regroupV0_lo_lo_lo_101 = {regroupV0_lo_lo_lo_hi_69, regroupV0_lo_lo_lo_lo_69};
  wire [127:0]       regroupV0_lo_lo_hi_lo_69 = {regroupV0_hi_74, regroupV0_lo_74, regroupV0_hi_73, regroupV0_lo_73};
  wire [127:0]       regroupV0_lo_lo_hi_hi_69 = {regroupV0_hi_76, regroupV0_lo_76, regroupV0_hi_75, regroupV0_lo_75};
  wire [255:0]       regroupV0_lo_lo_hi_101 = {regroupV0_lo_lo_hi_hi_69, regroupV0_lo_lo_hi_lo_69};
  wire [511:0]       regroupV0_lo_lo_101 = {regroupV0_lo_lo_hi_101, regroupV0_lo_lo_lo_101};
  wire [127:0]       regroupV0_lo_hi_lo_lo_69 = {regroupV0_hi_78, regroupV0_lo_78, regroupV0_hi_77, regroupV0_lo_77};
  wire [127:0]       regroupV0_lo_hi_lo_hi_69 = {regroupV0_hi_80, regroupV0_lo_80, regroupV0_hi_79, regroupV0_lo_79};
  wire [255:0]       regroupV0_lo_hi_lo_101 = {regroupV0_lo_hi_lo_hi_69, regroupV0_lo_hi_lo_lo_69};
  wire [127:0]       regroupV0_lo_hi_hi_lo_69 = {regroupV0_hi_82, regroupV0_lo_82, regroupV0_hi_81, regroupV0_lo_81};
  wire [127:0]       regroupV0_lo_hi_hi_hi_69 = {regroupV0_hi_84, regroupV0_lo_84, regroupV0_hi_83, regroupV0_lo_83};
  wire [255:0]       regroupV0_lo_hi_hi_101 = {regroupV0_lo_hi_hi_hi_69, regroupV0_lo_hi_hi_lo_69};
  wire [511:0]       regroupV0_lo_hi_101 = {regroupV0_lo_hi_hi_101, regroupV0_lo_hi_lo_101};
  wire [1023:0]      regroupV0_lo_101 = {regroupV0_lo_hi_101, regroupV0_lo_lo_101};
  wire [127:0]       regroupV0_hi_lo_lo_lo_69 = {regroupV0_hi_86, regroupV0_lo_86, regroupV0_hi_85, regroupV0_lo_85};
  wire [127:0]       regroupV0_hi_lo_lo_hi_69 = {regroupV0_hi_88, regroupV0_lo_88, regroupV0_hi_87, regroupV0_lo_87};
  wire [255:0]       regroupV0_hi_lo_lo_101 = {regroupV0_hi_lo_lo_hi_69, regroupV0_hi_lo_lo_lo_69};
  wire [127:0]       regroupV0_hi_lo_hi_lo_69 = {regroupV0_hi_90, regroupV0_lo_90, regroupV0_hi_89, regroupV0_lo_89};
  wire [127:0]       regroupV0_hi_lo_hi_hi_69 = {regroupV0_hi_92, regroupV0_lo_92, regroupV0_hi_91, regroupV0_lo_91};
  wire [255:0]       regroupV0_hi_lo_hi_101 = {regroupV0_hi_lo_hi_hi_69, regroupV0_hi_lo_hi_lo_69};
  wire [511:0]       regroupV0_hi_lo_101 = {regroupV0_hi_lo_hi_101, regroupV0_hi_lo_lo_101};
  wire [127:0]       regroupV0_hi_hi_lo_lo_69 = {regroupV0_hi_94, regroupV0_lo_94, regroupV0_hi_93, regroupV0_lo_93};
  wire [127:0]       regroupV0_hi_hi_lo_hi_69 = {regroupV0_hi_96, regroupV0_lo_96, regroupV0_hi_95, regroupV0_lo_95};
  wire [255:0]       regroupV0_hi_hi_lo_101 = {regroupV0_hi_hi_lo_hi_69, regroupV0_hi_hi_lo_lo_69};
  wire [127:0]       regroupV0_hi_hi_hi_lo_69 = {regroupV0_hi_98, regroupV0_lo_98, regroupV0_hi_97, regroupV0_lo_97};
  wire [127:0]       regroupV0_hi_hi_hi_hi_69 = {regroupV0_hi_100, regroupV0_lo_100, regroupV0_hi_99, regroupV0_lo_99};
  wire [255:0]       regroupV0_hi_hi_hi_101 = {regroupV0_hi_hi_hi_hi_69, regroupV0_hi_hi_hi_lo_69};
  wire [511:0]       regroupV0_hi_hi_101 = {regroupV0_hi_hi_hi_101, regroupV0_hi_hi_lo_101};
  wire [1023:0]      regroupV0_hi_101 = {regroupV0_hi_hi_101, regroupV0_hi_lo_101};
  wire [2047:0]      regroupV0_2 = {regroupV0_hi_101, regroupV0_lo_101};
  wire [3:0]         _v0SelectBySew_T = 4'h1 << laneMaskSewSelect_0;
  wire [63:0]        v0SelectBySew = (_v0SelectBySew_T[0] ? regroupV0_0[63:0] : 64'h0) | (_v0SelectBySew_T[1] ? regroupV0_1[63:0] : 64'h0) | (_v0SelectBySew_T[2] ? regroupV0_2[63:0] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_9 = 4'h1 << laneMaskSewSelect_1;
  wire [63:0]        v0SelectBySew_1 = (_v0SelectBySew_T_9[0] ? regroupV0_0[127:64] : 64'h0) | (_v0SelectBySew_T_9[1] ? regroupV0_1[127:64] : 64'h0) | (_v0SelectBySew_T_9[2] ? regroupV0_2[127:64] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_18 = 4'h1 << laneMaskSewSelect_2;
  wire [63:0]        v0SelectBySew_2 = (_v0SelectBySew_T_18[0] ? regroupV0_0[191:128] : 64'h0) | (_v0SelectBySew_T_18[1] ? regroupV0_1[191:128] : 64'h0) | (_v0SelectBySew_T_18[2] ? regroupV0_2[191:128] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_27 = 4'h1 << laneMaskSewSelect_3;
  wire [63:0]        v0SelectBySew_3 = (_v0SelectBySew_T_27[0] ? regroupV0_0[255:192] : 64'h0) | (_v0SelectBySew_T_27[1] ? regroupV0_1[255:192] : 64'h0) | (_v0SelectBySew_T_27[2] ? regroupV0_2[255:192] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_36 = 4'h1 << laneMaskSewSelect_4;
  wire [63:0]        v0SelectBySew_4 = (_v0SelectBySew_T_36[0] ? regroupV0_0[319:256] : 64'h0) | (_v0SelectBySew_T_36[1] ? regroupV0_1[319:256] : 64'h0) | (_v0SelectBySew_T_36[2] ? regroupV0_2[319:256] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_45 = 4'h1 << laneMaskSewSelect_5;
  wire [63:0]        v0SelectBySew_5 = (_v0SelectBySew_T_45[0] ? regroupV0_0[383:320] : 64'h0) | (_v0SelectBySew_T_45[1] ? regroupV0_1[383:320] : 64'h0) | (_v0SelectBySew_T_45[2] ? regroupV0_2[383:320] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_54 = 4'h1 << laneMaskSewSelect_6;
  wire [63:0]        v0SelectBySew_6 = (_v0SelectBySew_T_54[0] ? regroupV0_0[447:384] : 64'h0) | (_v0SelectBySew_T_54[1] ? regroupV0_1[447:384] : 64'h0) | (_v0SelectBySew_T_54[2] ? regroupV0_2[447:384] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_63 = 4'h1 << laneMaskSewSelect_7;
  wire [63:0]        v0SelectBySew_7 = (_v0SelectBySew_T_63[0] ? regroupV0_0[511:448] : 64'h0) | (_v0SelectBySew_T_63[1] ? regroupV0_1[511:448] : 64'h0) | (_v0SelectBySew_T_63[2] ? regroupV0_2[511:448] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_72 = 4'h1 << laneMaskSewSelect_8;
  wire [63:0]        v0SelectBySew_8 = (_v0SelectBySew_T_72[0] ? regroupV0_0[575:512] : 64'h0) | (_v0SelectBySew_T_72[1] ? regroupV0_1[575:512] : 64'h0) | (_v0SelectBySew_T_72[2] ? regroupV0_2[575:512] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_81 = 4'h1 << laneMaskSewSelect_9;
  wire [63:0]        v0SelectBySew_9 = (_v0SelectBySew_T_81[0] ? regroupV0_0[639:576] : 64'h0) | (_v0SelectBySew_T_81[1] ? regroupV0_1[639:576] : 64'h0) | (_v0SelectBySew_T_81[2] ? regroupV0_2[639:576] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_90 = 4'h1 << laneMaskSewSelect_10;
  wire [63:0]        v0SelectBySew_10 = (_v0SelectBySew_T_90[0] ? regroupV0_0[703:640] : 64'h0) | (_v0SelectBySew_T_90[1] ? regroupV0_1[703:640] : 64'h0) | (_v0SelectBySew_T_90[2] ? regroupV0_2[703:640] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_99 = 4'h1 << laneMaskSewSelect_11;
  wire [63:0]        v0SelectBySew_11 = (_v0SelectBySew_T_99[0] ? regroupV0_0[767:704] : 64'h0) | (_v0SelectBySew_T_99[1] ? regroupV0_1[767:704] : 64'h0) | (_v0SelectBySew_T_99[2] ? regroupV0_2[767:704] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_108 = 4'h1 << laneMaskSewSelect_12;
  wire [63:0]        v0SelectBySew_12 = (_v0SelectBySew_T_108[0] ? regroupV0_0[831:768] : 64'h0) | (_v0SelectBySew_T_108[1] ? regroupV0_1[831:768] : 64'h0) | (_v0SelectBySew_T_108[2] ? regroupV0_2[831:768] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_117 = 4'h1 << laneMaskSewSelect_13;
  wire [63:0]        v0SelectBySew_13 = (_v0SelectBySew_T_117[0] ? regroupV0_0[895:832] : 64'h0) | (_v0SelectBySew_T_117[1] ? regroupV0_1[895:832] : 64'h0) | (_v0SelectBySew_T_117[2] ? regroupV0_2[895:832] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_126 = 4'h1 << laneMaskSewSelect_14;
  wire [63:0]        v0SelectBySew_14 = (_v0SelectBySew_T_126[0] ? regroupV0_0[959:896] : 64'h0) | (_v0SelectBySew_T_126[1] ? regroupV0_1[959:896] : 64'h0) | (_v0SelectBySew_T_126[2] ? regroupV0_2[959:896] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_135 = 4'h1 << laneMaskSewSelect_15;
  wire [63:0]        v0SelectBySew_15 = (_v0SelectBySew_T_135[0] ? regroupV0_0[1023:960] : 64'h0) | (_v0SelectBySew_T_135[1] ? regroupV0_1[1023:960] : 64'h0) | (_v0SelectBySew_T_135[2] ? regroupV0_2[1023:960] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_144 = 4'h1 << laneMaskSewSelect_16;
  wire [63:0]        v0SelectBySew_16 = (_v0SelectBySew_T_144[0] ? regroupV0_0[1087:1024] : 64'h0) | (_v0SelectBySew_T_144[1] ? regroupV0_1[1087:1024] : 64'h0) | (_v0SelectBySew_T_144[2] ? regroupV0_2[1087:1024] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_153 = 4'h1 << laneMaskSewSelect_17;
  wire [63:0]        v0SelectBySew_17 = (_v0SelectBySew_T_153[0] ? regroupV0_0[1151:1088] : 64'h0) | (_v0SelectBySew_T_153[1] ? regroupV0_1[1151:1088] : 64'h0) | (_v0SelectBySew_T_153[2] ? regroupV0_2[1151:1088] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_162 = 4'h1 << laneMaskSewSelect_18;
  wire [63:0]        v0SelectBySew_18 = (_v0SelectBySew_T_162[0] ? regroupV0_0[1215:1152] : 64'h0) | (_v0SelectBySew_T_162[1] ? regroupV0_1[1215:1152] : 64'h0) | (_v0SelectBySew_T_162[2] ? regroupV0_2[1215:1152] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_171 = 4'h1 << laneMaskSewSelect_19;
  wire [63:0]        v0SelectBySew_19 = (_v0SelectBySew_T_171[0] ? regroupV0_0[1279:1216] : 64'h0) | (_v0SelectBySew_T_171[1] ? regroupV0_1[1279:1216] : 64'h0) | (_v0SelectBySew_T_171[2] ? regroupV0_2[1279:1216] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_180 = 4'h1 << laneMaskSewSelect_20;
  wire [63:0]        v0SelectBySew_20 = (_v0SelectBySew_T_180[0] ? regroupV0_0[1343:1280] : 64'h0) | (_v0SelectBySew_T_180[1] ? regroupV0_1[1343:1280] : 64'h0) | (_v0SelectBySew_T_180[2] ? regroupV0_2[1343:1280] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_189 = 4'h1 << laneMaskSewSelect_21;
  wire [63:0]        v0SelectBySew_21 = (_v0SelectBySew_T_189[0] ? regroupV0_0[1407:1344] : 64'h0) | (_v0SelectBySew_T_189[1] ? regroupV0_1[1407:1344] : 64'h0) | (_v0SelectBySew_T_189[2] ? regroupV0_2[1407:1344] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_198 = 4'h1 << laneMaskSewSelect_22;
  wire [63:0]        v0SelectBySew_22 = (_v0SelectBySew_T_198[0] ? regroupV0_0[1471:1408] : 64'h0) | (_v0SelectBySew_T_198[1] ? regroupV0_1[1471:1408] : 64'h0) | (_v0SelectBySew_T_198[2] ? regroupV0_2[1471:1408] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_207 = 4'h1 << laneMaskSewSelect_23;
  wire [63:0]        v0SelectBySew_23 = (_v0SelectBySew_T_207[0] ? regroupV0_0[1535:1472] : 64'h0) | (_v0SelectBySew_T_207[1] ? regroupV0_1[1535:1472] : 64'h0) | (_v0SelectBySew_T_207[2] ? regroupV0_2[1535:1472] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_216 = 4'h1 << laneMaskSewSelect_24;
  wire [63:0]        v0SelectBySew_24 = (_v0SelectBySew_T_216[0] ? regroupV0_0[1599:1536] : 64'h0) | (_v0SelectBySew_T_216[1] ? regroupV0_1[1599:1536] : 64'h0) | (_v0SelectBySew_T_216[2] ? regroupV0_2[1599:1536] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_225 = 4'h1 << laneMaskSewSelect_25;
  wire [63:0]        v0SelectBySew_25 = (_v0SelectBySew_T_225[0] ? regroupV0_0[1663:1600] : 64'h0) | (_v0SelectBySew_T_225[1] ? regroupV0_1[1663:1600] : 64'h0) | (_v0SelectBySew_T_225[2] ? regroupV0_2[1663:1600] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_234 = 4'h1 << laneMaskSewSelect_26;
  wire [63:0]        v0SelectBySew_26 = (_v0SelectBySew_T_234[0] ? regroupV0_0[1727:1664] : 64'h0) | (_v0SelectBySew_T_234[1] ? regroupV0_1[1727:1664] : 64'h0) | (_v0SelectBySew_T_234[2] ? regroupV0_2[1727:1664] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_243 = 4'h1 << laneMaskSewSelect_27;
  wire [63:0]        v0SelectBySew_27 = (_v0SelectBySew_T_243[0] ? regroupV0_0[1791:1728] : 64'h0) | (_v0SelectBySew_T_243[1] ? regroupV0_1[1791:1728] : 64'h0) | (_v0SelectBySew_T_243[2] ? regroupV0_2[1791:1728] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_252 = 4'h1 << laneMaskSewSelect_28;
  wire [63:0]        v0SelectBySew_28 = (_v0SelectBySew_T_252[0] ? regroupV0_0[1855:1792] : 64'h0) | (_v0SelectBySew_T_252[1] ? regroupV0_1[1855:1792] : 64'h0) | (_v0SelectBySew_T_252[2] ? regroupV0_2[1855:1792] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_261 = 4'h1 << laneMaskSewSelect_29;
  wire [63:0]        v0SelectBySew_29 = (_v0SelectBySew_T_261[0] ? regroupV0_0[1919:1856] : 64'h0) | (_v0SelectBySew_T_261[1] ? regroupV0_1[1919:1856] : 64'h0) | (_v0SelectBySew_T_261[2] ? regroupV0_2[1919:1856] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_270 = 4'h1 << laneMaskSewSelect_30;
  wire [63:0]        v0SelectBySew_30 = (_v0SelectBySew_T_270[0] ? regroupV0_0[1983:1920] : 64'h0) | (_v0SelectBySew_T_270[1] ? regroupV0_1[1983:1920] : 64'h0) | (_v0SelectBySew_T_270[2] ? regroupV0_2[1983:1920] : 64'h0);
  wire [3:0]         _v0SelectBySew_T_279 = 4'h1 << laneMaskSewSelect_31;
  wire [63:0]        v0SelectBySew_31 = (_v0SelectBySew_T_279[0] ? regroupV0_0[2047:1984] : 64'h0) | (_v0SelectBySew_T_279[1] ? regroupV0_1[2047:1984] : 64'h0) | (_v0SelectBySew_T_279[2] ? regroupV0_2[2047:1984] : 64'h0);
  wire [3:0]         intLMULInput = 4'h1 << instReq_bits_vlmul[1:0];
  wire [13:0]        _dataPosition_T_1 = {3'h0, instReq_bits_readFromScala[10:0]} << instReq_bits_sew;
  wire [10:0]        dataPosition = _dataPosition_T_1[10:0];
  wire [3:0]         _sewOHInput_T = 4'h1 << instReq_bits_sew;
  wire [2:0]         sewOHInput = _sewOHInput_T[2:0];
  wire [1:0]         dataOffset = {dataPosition[1] & (|(sewOHInput[1:0])), dataPosition[0] & sewOHInput[0]};
  wire [4:0]         accessLane = dataPosition[6:2];
  wire [3:0]         dataGroup = dataPosition[10:7];
  wire               offset = dataGroup[0];
  wire [2:0]         accessRegGrowth = dataGroup[3:1];
  wire [2:0]         reallyGrowth = accessRegGrowth;
  wire [5:0]         decimalProportion = {offset, accessLane};
  wire [2:0]         decimal = decimalProportion[5:3];
  wire               notNeedRead = |{instReq_bits_vlmul[2] & decimal >= intLMULInput[3:1] | ~(instReq_bits_vlmul[2]) & {1'h0, accessRegGrowth} >= intLMULInput, instReq_bits_readFromScala[31:11]};
  reg  [1:0]         gatherReadState;
  wire               gatherSRead = gatherReadState == 2'h1;
  wire               gatherWaiteRead = gatherReadState == 2'h2;
  assign gatherResponse = &gatherReadState;
  wire               gatherData_valid_0 = gatherResponse;
  reg  [1:0]         gatherDatOffset;
  reg  [4:0]         gatherLane;
  reg                gatherOffset;
  reg  [2:0]         gatherGrowth;
  reg  [2:0]         instReg_instructionIndex;
  wire [2:0]         exeResp_0_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_1_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_2_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_3_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_4_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_5_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_6_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_7_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_8_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_9_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_10_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_11_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_12_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_13_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_14_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_15_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_16_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_17_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_18_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_19_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_20_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_21_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_22_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_23_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_24_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_25_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_26_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_27_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_28_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_29_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_30_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_31_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_0_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_1_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_2_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_3_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_4_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_5_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_6_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_7_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_8_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_9_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_10_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_11_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_12_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_13_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_14_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_15_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_16_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_17_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_18_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_19_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_20_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_21_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_22_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_23_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_24_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_25_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_26_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_27_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_28_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_29_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_30_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_31_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         writeRequest_0_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_1_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_2_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_3_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_4_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_5_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_6_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_7_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_8_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_9_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_10_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_11_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_12_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_13_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_14_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_15_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_16_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_17_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_18_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_19_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_20_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_21_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_22_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_23_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_24_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_25_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_26_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_27_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_28_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_29_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_30_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_31_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_0_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_1_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_2_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_3_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_4_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_5_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_6_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_7_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_8_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_9_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_10_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_11_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_12_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_13_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_14_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_15_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_16_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_17_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_18_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_19_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_20_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_21_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_22_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_23_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_24_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_25_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_26_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_27_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_28_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_29_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_30_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_31_enq_bits_index = instReg_instructionIndex;
  reg                instReg_decodeResult_specialSlot;
  reg  [4:0]         instReg_decodeResult_topUop;
  reg                instReg_decodeResult_popCount;
  reg                instReg_decodeResult_ffo;
  reg                instReg_decodeResult_average;
  reg                instReg_decodeResult_reverse;
  reg                instReg_decodeResult_dontNeedExecuteInLane;
  reg                instReg_decodeResult_scheduler;
  reg                instReg_decodeResult_sReadVD;
  reg                instReg_decodeResult_vtype;
  reg                instReg_decodeResult_sWrite;
  reg                instReg_decodeResult_crossRead;
  reg                instReg_decodeResult_crossWrite;
  reg                instReg_decodeResult_maskUnit;
  reg                instReg_decodeResult_special;
  reg                instReg_decodeResult_saturate;
  reg                instReg_decodeResult_vwmacc;
  reg                instReg_decodeResult_readOnly;
  reg                instReg_decodeResult_maskSource;
  reg                instReg_decodeResult_maskDestination;
  reg                instReg_decodeResult_maskLogic;
  reg  [3:0]         instReg_decodeResult_uop;
  reg                instReg_decodeResult_iota;
  reg                instReg_decodeResult_mv;
  reg                instReg_decodeResult_extend;
  reg                instReg_decodeResult_unOrderWrite;
  reg                instReg_decodeResult_compress;
  reg                instReg_decodeResult_gather16;
  reg                instReg_decodeResult_gather;
  reg                instReg_decodeResult_slid;
  reg                instReg_decodeResult_targetRd;
  reg                instReg_decodeResult_widenReduce;
  reg                instReg_decodeResult_red;
  reg                instReg_decodeResult_nr;
  reg                instReg_decodeResult_itype;
  reg                instReg_decodeResult_unsigned1;
  reg                instReg_decodeResult_unsigned0;
  reg                instReg_decodeResult_other;
  reg                instReg_decodeResult_multiCycle;
  reg                instReg_decodeResult_divider;
  reg                instReg_decodeResult_multiplier;
  reg                instReg_decodeResult_shift;
  reg                instReg_decodeResult_adder;
  reg                instReg_decodeResult_logic;
  reg  [31:0]        instReg_readFromScala;
  reg  [1:0]         instReg_sew;
  reg  [2:0]         instReg_vlmul;
  reg                instReg_maskType;
  reg  [2:0]         instReg_vxrm;
  reg  [4:0]         instReg_vs2;
  reg  [4:0]         instReg_vs1;
  reg  [4:0]         instReg_vd;
  wire [4:0]         writeRequest_0_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_1_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_2_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_3_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_4_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_5_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_6_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_7_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_8_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_9_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_10_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_11_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_12_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_13_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_14_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_15_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_16_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_17_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_18_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_19_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_20_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_21_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_22_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_23_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_24_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_25_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_26_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_27_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_28_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_29_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_30_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_31_writeData_vd = instReg_vd;
  reg  [11:0]        instReg_vl;
  wire [11:0]        reduceLastDataNeed_byteForVl = instReg_vl;
  wire               enqMvRD = instReq_bits_decodeResult_topUop == 5'hB;
  reg                instVlValid;
  wire               gatherRequestFire = gatherReadState == 2'h0 & gatherRead & ~instVlValid;
  wire               viotaReq = instReq_bits_decodeResult_topUop == 5'h8;
  reg                readVS1Reg_dataValid;
  reg                readVS1Reg_requestSend;
  reg                readVS1Reg_sendToExecution;
  reg  [31:0]        readVS1Reg_data;
  reg  [3:0]         readVS1Reg_readIndex;
  wire [3:0]         _sew1H_T = 4'h1 << instReg_sew;
  wire [2:0]         sew1H = _sew1H_T[2:0];
  wire [3:0]         unitType = 4'h1 << instReg_decodeResult_topUop[4:3];
  wire [3:0]         subType = 4'h1 << instReg_decodeResult_topUop[2:1];
  wire               readType = unitType[0];
  wire               gather16 = instReg_decodeResult_topUop == 5'h5;
  wire               maskDestinationType = instReg_decodeResult_topUop == 5'h18;
  wire               compress = instReg_decodeResult_topUop[4:1] == 4'h4;
  wire               viota = instReg_decodeResult_topUop == 5'h8;
  wire               mv = instReg_decodeResult_topUop[4:1] == 4'h5;
  wire               mvRd = instReg_decodeResult_topUop == 5'hB;
  wire               mvVd = instReg_decodeResult_topUop == 5'hA;
  wire               orderReduce = {instReg_decodeResult_topUop[4:2], instReg_decodeResult_topUop[0]} == 4'hB;
  wire               ffo = instReg_decodeResult_topUop[4:1] == 4'h7;
  wire               extendType = unitType[3] & (subType[2] | subType[1]);
  wire               readValid = readType & instVlValid;
  wire               noSource = mv | viota;
  wire               allGroupExecute = maskDestinationType | unitType[2] | compress | ffo;
  wire               useDefaultSew = readType & ~gather16;
  wire [1:0]         _dataSplitSew_T_11 = useDefaultSew ? instReg_sew : 2'h0;
  wire [1:0]         dataSplitSew = {_dataSplitSew_T_11[1], _dataSplitSew_T_11[0] | unitType[3] & subType[1] | gather16} | {allGroupExecute, 1'h0};
  wire               sourceDataUseDefaultSew = ~(unitType[3] | gather16);
  wire [1:0]         _sourceDataEEW_T_6 = (sourceDataUseDefaultSew ? instReg_sew : 2'h0) | (unitType[3] ? instReg_sew >> subType[2:1] : 2'h0);
  wire [1:0]         sourceDataEEW = {_sourceDataEEW_T_6[1], _sourceDataEEW_T_6[0] | gather16};
  wire [3:0]         executeIndexGrowth = 4'h1 << dataSplitSew;
  wire [1:0]         lastExecuteIndex = {2{executeIndexGrowth[0]}} | {executeIndexGrowth[1], 1'h0};
  wire [3:0]         _sourceDataEEW1H_T = 4'h1 << sourceDataEEW;
  wire [2:0]         sourceDataEEW1H = _sourceDataEEW1H_T[2:0];
  wire [10:0]        lastElementIndex = instReg_vl[10:0] - {10'h0, |instReg_vl};
  wire [10:0]        processingVl_lastByteIndex = lastElementIndex;
  wire               maskFormatSource = ffo | maskDestinationType;
  wire [6:0]         processingVl_lastGroupRemaining = processingVl_lastByteIndex[6:0];
  wire [3:0]         processingVl_0_1 = processingVl_lastByteIndex[10:7];
  wire [4:0]         processingVl_lastLaneIndex = processingVl_lastGroupRemaining[6:2];
  wire [31:0]        _processingVl_lastGroupDataNeed_T = 32'h1 << processingVl_lastLaneIndex;
  wire [30:0]        _GEN_31 = _processingVl_lastGroupDataNeed_T[30:0] | _processingVl_lastGroupDataNeed_T[31:1];
  wire [29:0]        _GEN_32 = _GEN_31[29:0] | {_processingVl_lastGroupDataNeed_T[31], _GEN_31[30:2]};
  wire [27:0]        _GEN_33 = _GEN_32[27:0] | {_processingVl_lastGroupDataNeed_T[31], _GEN_31[30], _GEN_32[29:4]};
  wire [23:0]        _GEN_34 = _GEN_33[23:0] | {_processingVl_lastGroupDataNeed_T[31], _GEN_31[30], _GEN_32[29:28], _GEN_33[27:8]};
  wire [31:0]        processingVl_0_2 =
    {_processingVl_lastGroupDataNeed_T[31], _GEN_31[30], _GEN_32[29:28], _GEN_33[27:24], _GEN_34[23:16], _GEN_34[15:0] | {_processingVl_lastGroupDataNeed_T[31], _GEN_31[30], _GEN_32[29:28], _GEN_33[27:24], _GEN_34[23:16]}};
  wire [11:0]        processingVl_lastByteIndex_1 = {lastElementIndex, 1'h0};
  wire [6:0]         processingVl_lastGroupRemaining_1 = processingVl_lastByteIndex_1[6:0];
  wire [4:0]         processingVl_1_1 = processingVl_lastByteIndex_1[11:7];
  wire [4:0]         processingVl_lastLaneIndex_1 = processingVl_lastGroupRemaining_1[6:2];
  wire [31:0]        _processingVl_lastGroupDataNeed_T_11 = 32'h1 << processingVl_lastLaneIndex_1;
  wire [30:0]        _GEN_35 = _processingVl_lastGroupDataNeed_T_11[30:0] | _processingVl_lastGroupDataNeed_T_11[31:1];
  wire [29:0]        _GEN_36 = _GEN_35[29:0] | {_processingVl_lastGroupDataNeed_T_11[31], _GEN_35[30:2]};
  wire [27:0]        _GEN_37 = _GEN_36[27:0] | {_processingVl_lastGroupDataNeed_T_11[31], _GEN_35[30], _GEN_36[29:4]};
  wire [23:0]        _GEN_38 = _GEN_37[23:0] | {_processingVl_lastGroupDataNeed_T_11[31], _GEN_35[30], _GEN_36[29:28], _GEN_37[27:8]};
  wire [31:0]        processingVl_1_2 =
    {_processingVl_lastGroupDataNeed_T_11[31], _GEN_35[30], _GEN_36[29:28], _GEN_37[27:24], _GEN_38[23:16], _GEN_38[15:0] | {_processingVl_lastGroupDataNeed_T_11[31], _GEN_35[30], _GEN_36[29:28], _GEN_37[27:24], _GEN_38[23:16]}};
  wire [12:0]        processingVl_lastByteIndex_2 = {lastElementIndex, 2'h0};
  wire [6:0]         processingVl_lastGroupRemaining_2 = processingVl_lastByteIndex_2[6:0];
  wire [5:0]         processingVl_2_1 = processingVl_lastByteIndex_2[12:7];
  wire [4:0]         processingVl_lastLaneIndex_2 = processingVl_lastGroupRemaining_2[6:2];
  wire [31:0]        _processingVl_lastGroupDataNeed_T_22 = 32'h1 << processingVl_lastLaneIndex_2;
  wire [30:0]        _GEN_39 = _processingVl_lastGroupDataNeed_T_22[30:0] | _processingVl_lastGroupDataNeed_T_22[31:1];
  wire [29:0]        _GEN_40 = _GEN_39[29:0] | {_processingVl_lastGroupDataNeed_T_22[31], _GEN_39[30:2]};
  wire [27:0]        _GEN_41 = _GEN_40[27:0] | {_processingVl_lastGroupDataNeed_T_22[31], _GEN_39[30], _GEN_40[29:4]};
  wire [23:0]        _GEN_42 = _GEN_41[23:0] | {_processingVl_lastGroupDataNeed_T_22[31], _GEN_39[30], _GEN_40[29:28], _GEN_41[27:8]};
  wire [31:0]        processingVl_2_2 =
    {_processingVl_lastGroupDataNeed_T_22[31], _GEN_39[30], _GEN_40[29:28], _GEN_41[27:24], _GEN_42[23:16], _GEN_42[15:0] | {_processingVl_lastGroupDataNeed_T_22[31], _GEN_39[30], _GEN_40[29:28], _GEN_41[27:24], _GEN_42[23:16]}};
  wire [9:0]         processingMaskVl_lastGroupRemaining = lastElementIndex[9:0];
  wire [9:0]         elementTailForMaskDestination = lastElementIndex[9:0];
  wire               processingMaskVl_lastGroupMisAlign = |processingMaskVl_lastGroupRemaining;
  wire               processingMaskVl_0_1 = lastElementIndex[10];
  wire [4:0]         processingMaskVl_lastLaneIndex = processingMaskVl_lastGroupRemaining[9:5] - {4'h0, processingMaskVl_lastGroupRemaining[4:0] == 5'h0};
  wire [31:0]        _processingMaskVl_dataNeedForPL_T = 32'h1 << processingMaskVl_lastLaneIndex;
  wire [30:0]        _GEN_43 = _processingMaskVl_dataNeedForPL_T[30:0] | _processingMaskVl_dataNeedForPL_T[31:1];
  wire [29:0]        _GEN_44 = _GEN_43[29:0] | {_processingMaskVl_dataNeedForPL_T[31], _GEN_43[30:2]};
  wire [27:0]        _GEN_45 = _GEN_44[27:0] | {_processingMaskVl_dataNeedForPL_T[31], _GEN_43[30], _GEN_44[29:4]};
  wire [23:0]        _GEN_46 = _GEN_45[23:0] | {_processingMaskVl_dataNeedForPL_T[31], _GEN_43[30], _GEN_44[29:28], _GEN_45[27:8]};
  wire [31:0]        processingMaskVl_dataNeedForPL =
    {_processingMaskVl_dataNeedForPL_T[31], _GEN_43[30], _GEN_44[29:28], _GEN_45[27:24], _GEN_46[23:16], _GEN_46[15:0] | {_processingMaskVl_dataNeedForPL_T[31], _GEN_43[30], _GEN_44[29:28], _GEN_45[27:24], _GEN_46[23:16]}};
  wire               processingMaskVl_dataNeedForNPL_misAlign = |(processingMaskVl_lastGroupRemaining[1:0]);
  wire [8:0]         processingMaskVl_dataNeedForNPL_datapathSize = {1'h0, processingMaskVl_lastGroupRemaining[9:2]} + {8'h0, processingMaskVl_dataNeedForNPL_misAlign};
  wire               processingMaskVl_dataNeedForNPL_allNeed = |(processingMaskVl_dataNeedForNPL_datapathSize[8:5]);
  wire [4:0]         processingMaskVl_dataNeedForNPL_lastLaneIndex = processingMaskVl_dataNeedForNPL_datapathSize[4:0];
  wire [31:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T = 32'h1 << processingMaskVl_dataNeedForNPL_lastLaneIndex;
  wire [31:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_3 = _processingMaskVl_dataNeedForNPL_dataNeed_T | {_processingMaskVl_dataNeedForNPL_dataNeed_T[30:0], 1'h0};
  wire [31:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_6 = _processingMaskVl_dataNeedForNPL_dataNeed_T_3 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_3[29:0], 2'h0};
  wire [31:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_9 = _processingMaskVl_dataNeedForNPL_dataNeed_T_6 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_6[27:0], 4'h0};
  wire [31:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_12 = _processingMaskVl_dataNeedForNPL_dataNeed_T_9 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_9[23:0], 8'h0};
  wire [31:0]        processingMaskVl_dataNeedForNPL_dataNeed = ~(_processingMaskVl_dataNeedForNPL_dataNeed_T_12 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_12[15:0], 16'h0}) | {32{processingMaskVl_dataNeedForNPL_allNeed}};
  wire               processingMaskVl_dataNeedForNPL_misAlign_1 = processingMaskVl_lastGroupRemaining[0];
  wire [9:0]         processingMaskVl_dataNeedForNPL_datapathSize_1 = {1'h0, processingMaskVl_lastGroupRemaining[9:1]} + {9'h0, processingMaskVl_dataNeedForNPL_misAlign_1};
  wire               processingMaskVl_dataNeedForNPL_allNeed_1 = |(processingMaskVl_dataNeedForNPL_datapathSize_1[9:5]);
  wire [4:0]         processingMaskVl_dataNeedForNPL_lastLaneIndex_1 = processingMaskVl_dataNeedForNPL_datapathSize_1[4:0];
  wire [31:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_19 = 32'h1 << processingMaskVl_dataNeedForNPL_lastLaneIndex_1;
  wire [31:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_22 = _processingMaskVl_dataNeedForNPL_dataNeed_T_19 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_19[30:0], 1'h0};
  wire [31:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_25 = _processingMaskVl_dataNeedForNPL_dataNeed_T_22 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_22[29:0], 2'h0};
  wire [31:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_28 = _processingMaskVl_dataNeedForNPL_dataNeed_T_25 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_25[27:0], 4'h0};
  wire [31:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_31 = _processingMaskVl_dataNeedForNPL_dataNeed_T_28 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_28[23:0], 8'h0};
  wire [31:0]        processingMaskVl_dataNeedForNPL_dataNeed_1 = ~(_processingMaskVl_dataNeedForNPL_dataNeed_T_31 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_31[15:0], 16'h0}) | {32{processingMaskVl_dataNeedForNPL_allNeed_1}};
  wire [10:0]        processingMaskVl_dataNeedForNPL_datapathSize_2 = {1'h0, processingMaskVl_lastGroupRemaining};
  wire               processingMaskVl_dataNeedForNPL_allNeed_2 = |(processingMaskVl_dataNeedForNPL_datapathSize_2[10:5]);
  wire [4:0]         processingMaskVl_dataNeedForNPL_lastLaneIndex_2 = processingMaskVl_dataNeedForNPL_datapathSize_2[4:0];
  wire [31:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_38 = 32'h1 << processingMaskVl_dataNeedForNPL_lastLaneIndex_2;
  wire [31:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_41 = _processingMaskVl_dataNeedForNPL_dataNeed_T_38 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_38[30:0], 1'h0};
  wire [31:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_44 = _processingMaskVl_dataNeedForNPL_dataNeed_T_41 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_41[29:0], 2'h0};
  wire [31:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_47 = _processingMaskVl_dataNeedForNPL_dataNeed_T_44 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_44[27:0], 4'h0};
  wire [31:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_50 = _processingMaskVl_dataNeedForNPL_dataNeed_T_47 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_47[23:0], 8'h0};
  wire [31:0]        processingMaskVl_dataNeedForNPL_dataNeed_2 = ~(_processingMaskVl_dataNeedForNPL_dataNeed_T_50 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_50[15:0], 16'h0}) | {32{processingMaskVl_dataNeedForNPL_allNeed_2}};
  wire [31:0]        processingMaskVl_dataNeedForNPL =
    (sew1H[0] ? processingMaskVl_dataNeedForNPL_dataNeed : 32'h0) | (sew1H[1] ? processingMaskVl_dataNeedForNPL_dataNeed_1 : 32'h0) | (sew1H[2] ? processingMaskVl_dataNeedForNPL_dataNeed_2 : 32'h0);
  wire [31:0]        processingMaskVl_0_2 = ffo ? processingMaskVl_dataNeedForPL : processingMaskVl_dataNeedForNPL;
  wire               reduceLastDataNeed_vlMSB = |(reduceLastDataNeed_byteForVl[11:7]);
  wire [6:0]         reduceLastDataNeed_vlLSB = instReg_vl[6:0];
  wire [6:0]         reduceLastDataNeed_vlLSB_1 = instReg_vl[6:0];
  wire [6:0]         reduceLastDataNeed_vlLSB_2 = instReg_vl[6:0];
  wire [4:0]         reduceLastDataNeed_lsbDSize = reduceLastDataNeed_vlLSB[6:2] - {4'h0, reduceLastDataNeed_vlLSB[1:0] == 2'h0};
  wire [31:0]        _reduceLastDataNeed_T = 32'h1 << reduceLastDataNeed_lsbDSize;
  wire [30:0]        _GEN_47 = _reduceLastDataNeed_T[30:0] | _reduceLastDataNeed_T[31:1];
  wire [29:0]        _GEN_48 = _GEN_47[29:0] | {_reduceLastDataNeed_T[31], _GEN_47[30:2]};
  wire [27:0]        _GEN_49 = _GEN_48[27:0] | {_reduceLastDataNeed_T[31], _GEN_47[30], _GEN_48[29:4]};
  wire [23:0]        _GEN_50 = _GEN_49[23:0] | {_reduceLastDataNeed_T[31], _GEN_47[30], _GEN_48[29:28], _GEN_49[27:8]};
  wire [12:0]        reduceLastDataNeed_byteForVl_1 = {instReg_vl, 1'h0};
  wire               reduceLastDataNeed_vlMSB_1 = |(reduceLastDataNeed_byteForVl_1[12:7]);
  wire [4:0]         reduceLastDataNeed_lsbDSize_1 = reduceLastDataNeed_vlLSB_1[6:2] - {4'h0, reduceLastDataNeed_vlLSB_1[1:0] == 2'h0};
  wire [31:0]        _reduceLastDataNeed_T_14 = 32'h1 << reduceLastDataNeed_lsbDSize_1;
  wire [30:0]        _GEN_51 = _reduceLastDataNeed_T_14[30:0] | _reduceLastDataNeed_T_14[31:1];
  wire [29:0]        _GEN_52 = _GEN_51[29:0] | {_reduceLastDataNeed_T_14[31], _GEN_51[30:2]};
  wire [27:0]        _GEN_53 = _GEN_52[27:0] | {_reduceLastDataNeed_T_14[31], _GEN_51[30], _GEN_52[29:4]};
  wire [23:0]        _GEN_54 = _GEN_53[23:0] | {_reduceLastDataNeed_T_14[31], _GEN_51[30], _GEN_52[29:28], _GEN_53[27:8]};
  wire [13:0]        reduceLastDataNeed_byteForVl_2 = {instReg_vl, 2'h0};
  wire               reduceLastDataNeed_vlMSB_2 = |(reduceLastDataNeed_byteForVl_2[13:7]);
  wire [4:0]         reduceLastDataNeed_lsbDSize_2 = reduceLastDataNeed_vlLSB_2[6:2] - {4'h0, reduceLastDataNeed_vlLSB_2[1:0] == 2'h0};
  wire [31:0]        _reduceLastDataNeed_T_28 = 32'h1 << reduceLastDataNeed_lsbDSize_2;
  wire [30:0]        _GEN_55 = _reduceLastDataNeed_T_28[30:0] | _reduceLastDataNeed_T_28[31:1];
  wire [29:0]        _GEN_56 = _GEN_55[29:0] | {_reduceLastDataNeed_T_28[31], _GEN_55[30:2]};
  wire [27:0]        _GEN_57 = _GEN_56[27:0] | {_reduceLastDataNeed_T_28[31], _GEN_55[30], _GEN_56[29:4]};
  wire [23:0]        _GEN_58 = _GEN_57[23:0] | {_reduceLastDataNeed_T_28[31], _GEN_55[30], _GEN_56[29:28], _GEN_57[27:8]};
  wire [31:0]        reduceLastDataNeed =
    (sew1H[0]
       ? {_reduceLastDataNeed_T[31], _GEN_47[30], _GEN_48[29:28], _GEN_49[27:24], _GEN_50[23:16], _GEN_50[15:0] | {_reduceLastDataNeed_T[31], _GEN_47[30], _GEN_48[29:28], _GEN_49[27:24], _GEN_50[23:16]}} | {32{reduceLastDataNeed_vlMSB}}
       : 32'h0)
    | (sew1H[1]
         ? {_reduceLastDataNeed_T_14[31], _GEN_51[30], _GEN_52[29:28], _GEN_53[27:24], _GEN_54[23:16], _GEN_54[15:0] | {_reduceLastDataNeed_T_14[31], _GEN_51[30], _GEN_52[29:28], _GEN_53[27:24], _GEN_54[23:16]}}
           | {32{reduceLastDataNeed_vlMSB_1}}
         : 32'h0)
    | (sew1H[2]
         ? {_reduceLastDataNeed_T_28[31], _GEN_55[30], _GEN_56[29:28], _GEN_57[27:24], _GEN_58[23:16], _GEN_58[15:0] | {_reduceLastDataNeed_T_28[31], _GEN_55[30], _GEN_56[29:28], _GEN_57[27:24], _GEN_58[23:16]}}
           | {32{reduceLastDataNeed_vlMSB_2}}
         : 32'h0);
  wire [1:0]         dataSourceSew = unitType[3] ? instReg_sew - instReg_decodeResult_topUop[2:1] : gather16 ? 2'h1 : instReg_sew;
  wire [3:0]         _dataSourceSew1H_T = 4'h1 << dataSourceSew;
  wire [2:0]         dataSourceSew1H = _dataSourceSew1H_T[2:0];
  wire               unorderReduce = ~orderReduce & unitType[2];
  wire               normalFormat = ~maskFormatSource & ~unorderReduce & ~mv;
  wire [5:0]         lastGroupForInstruction =
    {1'h0, {1'h0, {3'h0, maskFormatSource & processingMaskVl_0_1} | (normalFormat & dataSourceSew1H[0] ? processingVl_0_1 : 4'h0)} | (normalFormat & dataSourceSew1H[1] ? processingVl_1_1 : 5'h0)}
    | (normalFormat & dataSourceSew1H[2] ? processingVl_2_1 : 6'h0);
  wire [5:0]         popDataNeed_dataPathGroups = lastElementIndex[10:5];
  wire [4:0]         popDataNeed_lastLaneIndex = popDataNeed_dataPathGroups[4:0];
  wire               popDataNeed_lagerThanDLen = popDataNeed_dataPathGroups[5];
  wire [31:0]        _popDataNeed_T = 32'h1 << popDataNeed_lastLaneIndex;
  wire [30:0]        _GEN_59 = _popDataNeed_T[30:0] | _popDataNeed_T[31:1];
  wire [29:0]        _GEN_60 = _GEN_59[29:0] | {_popDataNeed_T[31], _GEN_59[30:2]};
  wire [27:0]        _GEN_61 = _GEN_60[27:0] | {_popDataNeed_T[31], _GEN_59[30], _GEN_60[29:4]};
  wire [23:0]        _GEN_62 = _GEN_61[23:0] | {_popDataNeed_T[31], _GEN_59[30], _GEN_60[29:28], _GEN_61[27:8]};
  wire [31:0]        popDataNeed =
    {_popDataNeed_T[31], _GEN_59[30], _GEN_60[29:28], _GEN_61[27:24], _GEN_62[23:16], _GEN_62[15:0] | {_popDataNeed_T[31], _GEN_59[30], _GEN_60[29:28], _GEN_61[27:24], _GEN_62[23:16]}} | {32{popDataNeed_lagerThanDLen}};
  wire [31:0]        lastGroupDataNeed =
    (unorderReduce & instReg_decodeResult_popCount ? popDataNeed : 32'h0) | (unorderReduce & ~instReg_decodeResult_popCount ? reduceLastDataNeed : 32'h0) | (maskFormatSource ? processingMaskVl_0_2 : 32'h0)
    | (normalFormat & dataSourceSew1H[0] ? processingVl_0_2 : 32'h0) | (normalFormat & dataSourceSew1H[1] ? processingVl_1_2 : 32'h0) | (normalFormat & dataSourceSew1H[2] ? processingVl_2_2 : 32'h0);
  wire [3:0]         exeRequestQueue_queue_dataIn_lo = {exeRequestQueue_0_enq_bits_index, exeRequestQueue_0_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi = {exeRequestQueue_0_enq_bits_source1, exeRequestQueue_0_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn = {exeRequestQueue_queue_dataIn_hi, exeRequestQueue_queue_dataIn_lo};
  wire               exeRequestQueue_queue_dataOut_ffo = _exeRequestQueue_queue_fifo_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_index = _exeRequestQueue_queue_fifo_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_source2 = _exeRequestQueue_queue_fifo_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_source1 = _exeRequestQueue_queue_fifo_data_out[67:36];
  wire               exeRequestQueue_0_enq_ready = ~_exeRequestQueue_queue_fifo_full;
  wire               exeRequestQueue_0_deq_ready;
  wire               exeRequestQueue_0_deq_valid = ~_exeRequestQueue_queue_fifo_empty | exeRequestQueue_0_enq_valid;
  wire [31:0]        exeRequestQueue_0_deq_bits_source1 = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_source1 : exeRequestQueue_queue_dataOut_source1;
  wire [31:0]        exeRequestQueue_0_deq_bits_source2 = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_source2 : exeRequestQueue_queue_dataOut_source2;
  wire [2:0]         exeRequestQueue_0_deq_bits_index = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_index : exeRequestQueue_queue_dataOut_index;
  wire               exeRequestQueue_0_deq_bits_ffo = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_ffo : exeRequestQueue_queue_dataOut_ffo;
  wire               tokenIO_0_maskRequestRelease_0 = exeRequestQueue_0_deq_ready & exeRequestQueue_0_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_1 = {exeRequestQueue_1_enq_bits_index, exeRequestQueue_1_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_1 = {exeRequestQueue_1_enq_bits_source1, exeRequestQueue_1_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_1 = {exeRequestQueue_queue_dataIn_hi_1, exeRequestQueue_queue_dataIn_lo_1};
  wire               exeRequestQueue_queue_dataOut_1_ffo = _exeRequestQueue_queue_fifo_1_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_1_index = _exeRequestQueue_queue_fifo_1_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_1_source2 = _exeRequestQueue_queue_fifo_1_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_1_source1 = _exeRequestQueue_queue_fifo_1_data_out[67:36];
  wire               exeRequestQueue_1_enq_ready = ~_exeRequestQueue_queue_fifo_1_full;
  wire               exeRequestQueue_1_deq_ready;
  wire               exeRequestQueue_1_deq_valid = ~_exeRequestQueue_queue_fifo_1_empty | exeRequestQueue_1_enq_valid;
  wire [31:0]        exeRequestQueue_1_deq_bits_source1 = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_source1 : exeRequestQueue_queue_dataOut_1_source1;
  wire [31:0]        exeRequestQueue_1_deq_bits_source2 = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_source2 : exeRequestQueue_queue_dataOut_1_source2;
  wire [2:0]         exeRequestQueue_1_deq_bits_index = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_index : exeRequestQueue_queue_dataOut_1_index;
  wire               exeRequestQueue_1_deq_bits_ffo = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_ffo : exeRequestQueue_queue_dataOut_1_ffo;
  wire               tokenIO_1_maskRequestRelease_0 = exeRequestQueue_1_deq_ready & exeRequestQueue_1_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_2 = {exeRequestQueue_2_enq_bits_index, exeRequestQueue_2_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_2 = {exeRequestQueue_2_enq_bits_source1, exeRequestQueue_2_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_2 = {exeRequestQueue_queue_dataIn_hi_2, exeRequestQueue_queue_dataIn_lo_2};
  wire               exeRequestQueue_queue_dataOut_2_ffo = _exeRequestQueue_queue_fifo_2_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_2_index = _exeRequestQueue_queue_fifo_2_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_2_source2 = _exeRequestQueue_queue_fifo_2_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_2_source1 = _exeRequestQueue_queue_fifo_2_data_out[67:36];
  wire               exeRequestQueue_2_enq_ready = ~_exeRequestQueue_queue_fifo_2_full;
  wire               exeRequestQueue_2_deq_ready;
  wire               exeRequestQueue_2_deq_valid = ~_exeRequestQueue_queue_fifo_2_empty | exeRequestQueue_2_enq_valid;
  wire [31:0]        exeRequestQueue_2_deq_bits_source1 = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_source1 : exeRequestQueue_queue_dataOut_2_source1;
  wire [31:0]        exeRequestQueue_2_deq_bits_source2 = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_source2 : exeRequestQueue_queue_dataOut_2_source2;
  wire [2:0]         exeRequestQueue_2_deq_bits_index = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_index : exeRequestQueue_queue_dataOut_2_index;
  wire               exeRequestQueue_2_deq_bits_ffo = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_ffo : exeRequestQueue_queue_dataOut_2_ffo;
  wire               tokenIO_2_maskRequestRelease_0 = exeRequestQueue_2_deq_ready & exeRequestQueue_2_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_3 = {exeRequestQueue_3_enq_bits_index, exeRequestQueue_3_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_3 = {exeRequestQueue_3_enq_bits_source1, exeRequestQueue_3_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_3 = {exeRequestQueue_queue_dataIn_hi_3, exeRequestQueue_queue_dataIn_lo_3};
  wire               exeRequestQueue_queue_dataOut_3_ffo = _exeRequestQueue_queue_fifo_3_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_3_index = _exeRequestQueue_queue_fifo_3_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_3_source2 = _exeRequestQueue_queue_fifo_3_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_3_source1 = _exeRequestQueue_queue_fifo_3_data_out[67:36];
  wire               exeRequestQueue_3_enq_ready = ~_exeRequestQueue_queue_fifo_3_full;
  wire               exeRequestQueue_3_deq_ready;
  wire               exeRequestQueue_3_deq_valid = ~_exeRequestQueue_queue_fifo_3_empty | exeRequestQueue_3_enq_valid;
  wire [31:0]        exeRequestQueue_3_deq_bits_source1 = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_source1 : exeRequestQueue_queue_dataOut_3_source1;
  wire [31:0]        exeRequestQueue_3_deq_bits_source2 = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_source2 : exeRequestQueue_queue_dataOut_3_source2;
  wire [2:0]         exeRequestQueue_3_deq_bits_index = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_index : exeRequestQueue_queue_dataOut_3_index;
  wire               exeRequestQueue_3_deq_bits_ffo = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_ffo : exeRequestQueue_queue_dataOut_3_ffo;
  wire               tokenIO_3_maskRequestRelease_0 = exeRequestQueue_3_deq_ready & exeRequestQueue_3_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_4 = {exeRequestQueue_4_enq_bits_index, exeRequestQueue_4_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_4 = {exeRequestQueue_4_enq_bits_source1, exeRequestQueue_4_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_4 = {exeRequestQueue_queue_dataIn_hi_4, exeRequestQueue_queue_dataIn_lo_4};
  wire               exeRequestQueue_queue_dataOut_4_ffo = _exeRequestQueue_queue_fifo_4_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_4_index = _exeRequestQueue_queue_fifo_4_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_4_source2 = _exeRequestQueue_queue_fifo_4_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_4_source1 = _exeRequestQueue_queue_fifo_4_data_out[67:36];
  wire               exeRequestQueue_4_enq_ready = ~_exeRequestQueue_queue_fifo_4_full;
  wire               exeRequestQueue_4_deq_ready;
  wire               exeRequestQueue_4_deq_valid = ~_exeRequestQueue_queue_fifo_4_empty | exeRequestQueue_4_enq_valid;
  wire [31:0]        exeRequestQueue_4_deq_bits_source1 = _exeRequestQueue_queue_fifo_4_empty ? exeRequestQueue_4_enq_bits_source1 : exeRequestQueue_queue_dataOut_4_source1;
  wire [31:0]        exeRequestQueue_4_deq_bits_source2 = _exeRequestQueue_queue_fifo_4_empty ? exeRequestQueue_4_enq_bits_source2 : exeRequestQueue_queue_dataOut_4_source2;
  wire [2:0]         exeRequestQueue_4_deq_bits_index = _exeRequestQueue_queue_fifo_4_empty ? exeRequestQueue_4_enq_bits_index : exeRequestQueue_queue_dataOut_4_index;
  wire               exeRequestQueue_4_deq_bits_ffo = _exeRequestQueue_queue_fifo_4_empty ? exeRequestQueue_4_enq_bits_ffo : exeRequestQueue_queue_dataOut_4_ffo;
  wire               tokenIO_4_maskRequestRelease_0 = exeRequestQueue_4_deq_ready & exeRequestQueue_4_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_5 = {exeRequestQueue_5_enq_bits_index, exeRequestQueue_5_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_5 = {exeRequestQueue_5_enq_bits_source1, exeRequestQueue_5_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_5 = {exeRequestQueue_queue_dataIn_hi_5, exeRequestQueue_queue_dataIn_lo_5};
  wire               exeRequestQueue_queue_dataOut_5_ffo = _exeRequestQueue_queue_fifo_5_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_5_index = _exeRequestQueue_queue_fifo_5_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_5_source2 = _exeRequestQueue_queue_fifo_5_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_5_source1 = _exeRequestQueue_queue_fifo_5_data_out[67:36];
  wire               exeRequestQueue_5_enq_ready = ~_exeRequestQueue_queue_fifo_5_full;
  wire               exeRequestQueue_5_deq_ready;
  wire               exeRequestQueue_5_deq_valid = ~_exeRequestQueue_queue_fifo_5_empty | exeRequestQueue_5_enq_valid;
  wire [31:0]        exeRequestQueue_5_deq_bits_source1 = _exeRequestQueue_queue_fifo_5_empty ? exeRequestQueue_5_enq_bits_source1 : exeRequestQueue_queue_dataOut_5_source1;
  wire [31:0]        exeRequestQueue_5_deq_bits_source2 = _exeRequestQueue_queue_fifo_5_empty ? exeRequestQueue_5_enq_bits_source2 : exeRequestQueue_queue_dataOut_5_source2;
  wire [2:0]         exeRequestQueue_5_deq_bits_index = _exeRequestQueue_queue_fifo_5_empty ? exeRequestQueue_5_enq_bits_index : exeRequestQueue_queue_dataOut_5_index;
  wire               exeRequestQueue_5_deq_bits_ffo = _exeRequestQueue_queue_fifo_5_empty ? exeRequestQueue_5_enq_bits_ffo : exeRequestQueue_queue_dataOut_5_ffo;
  wire               tokenIO_5_maskRequestRelease_0 = exeRequestQueue_5_deq_ready & exeRequestQueue_5_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_6 = {exeRequestQueue_6_enq_bits_index, exeRequestQueue_6_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_6 = {exeRequestQueue_6_enq_bits_source1, exeRequestQueue_6_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_6 = {exeRequestQueue_queue_dataIn_hi_6, exeRequestQueue_queue_dataIn_lo_6};
  wire               exeRequestQueue_queue_dataOut_6_ffo = _exeRequestQueue_queue_fifo_6_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_6_index = _exeRequestQueue_queue_fifo_6_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_6_source2 = _exeRequestQueue_queue_fifo_6_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_6_source1 = _exeRequestQueue_queue_fifo_6_data_out[67:36];
  wire               exeRequestQueue_6_enq_ready = ~_exeRequestQueue_queue_fifo_6_full;
  wire               exeRequestQueue_6_deq_ready;
  wire               exeRequestQueue_6_deq_valid = ~_exeRequestQueue_queue_fifo_6_empty | exeRequestQueue_6_enq_valid;
  wire [31:0]        exeRequestQueue_6_deq_bits_source1 = _exeRequestQueue_queue_fifo_6_empty ? exeRequestQueue_6_enq_bits_source1 : exeRequestQueue_queue_dataOut_6_source1;
  wire [31:0]        exeRequestQueue_6_deq_bits_source2 = _exeRequestQueue_queue_fifo_6_empty ? exeRequestQueue_6_enq_bits_source2 : exeRequestQueue_queue_dataOut_6_source2;
  wire [2:0]         exeRequestQueue_6_deq_bits_index = _exeRequestQueue_queue_fifo_6_empty ? exeRequestQueue_6_enq_bits_index : exeRequestQueue_queue_dataOut_6_index;
  wire               exeRequestQueue_6_deq_bits_ffo = _exeRequestQueue_queue_fifo_6_empty ? exeRequestQueue_6_enq_bits_ffo : exeRequestQueue_queue_dataOut_6_ffo;
  wire               tokenIO_6_maskRequestRelease_0 = exeRequestQueue_6_deq_ready & exeRequestQueue_6_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_7 = {exeRequestQueue_7_enq_bits_index, exeRequestQueue_7_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_7 = {exeRequestQueue_7_enq_bits_source1, exeRequestQueue_7_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_7 = {exeRequestQueue_queue_dataIn_hi_7, exeRequestQueue_queue_dataIn_lo_7};
  wire               exeRequestQueue_queue_dataOut_7_ffo = _exeRequestQueue_queue_fifo_7_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_7_index = _exeRequestQueue_queue_fifo_7_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_7_source2 = _exeRequestQueue_queue_fifo_7_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_7_source1 = _exeRequestQueue_queue_fifo_7_data_out[67:36];
  wire               exeRequestQueue_7_enq_ready = ~_exeRequestQueue_queue_fifo_7_full;
  wire               exeRequestQueue_7_deq_ready;
  wire               exeRequestQueue_7_deq_valid = ~_exeRequestQueue_queue_fifo_7_empty | exeRequestQueue_7_enq_valid;
  wire [31:0]        exeRequestQueue_7_deq_bits_source1 = _exeRequestQueue_queue_fifo_7_empty ? exeRequestQueue_7_enq_bits_source1 : exeRequestQueue_queue_dataOut_7_source1;
  wire [31:0]        exeRequestQueue_7_deq_bits_source2 = _exeRequestQueue_queue_fifo_7_empty ? exeRequestQueue_7_enq_bits_source2 : exeRequestQueue_queue_dataOut_7_source2;
  wire [2:0]         exeRequestQueue_7_deq_bits_index = _exeRequestQueue_queue_fifo_7_empty ? exeRequestQueue_7_enq_bits_index : exeRequestQueue_queue_dataOut_7_index;
  wire               exeRequestQueue_7_deq_bits_ffo = _exeRequestQueue_queue_fifo_7_empty ? exeRequestQueue_7_enq_bits_ffo : exeRequestQueue_queue_dataOut_7_ffo;
  wire               tokenIO_7_maskRequestRelease_0 = exeRequestQueue_7_deq_ready & exeRequestQueue_7_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_8 = {exeRequestQueue_8_enq_bits_index, exeRequestQueue_8_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_8 = {exeRequestQueue_8_enq_bits_source1, exeRequestQueue_8_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_8 = {exeRequestQueue_queue_dataIn_hi_8, exeRequestQueue_queue_dataIn_lo_8};
  wire               exeRequestQueue_queue_dataOut_8_ffo = _exeRequestQueue_queue_fifo_8_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_8_index = _exeRequestQueue_queue_fifo_8_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_8_source2 = _exeRequestQueue_queue_fifo_8_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_8_source1 = _exeRequestQueue_queue_fifo_8_data_out[67:36];
  wire               exeRequestQueue_8_enq_ready = ~_exeRequestQueue_queue_fifo_8_full;
  wire               exeRequestQueue_8_deq_ready;
  wire               exeRequestQueue_8_deq_valid = ~_exeRequestQueue_queue_fifo_8_empty | exeRequestQueue_8_enq_valid;
  wire [31:0]        exeRequestQueue_8_deq_bits_source1 = _exeRequestQueue_queue_fifo_8_empty ? exeRequestQueue_8_enq_bits_source1 : exeRequestQueue_queue_dataOut_8_source1;
  wire [31:0]        exeRequestQueue_8_deq_bits_source2 = _exeRequestQueue_queue_fifo_8_empty ? exeRequestQueue_8_enq_bits_source2 : exeRequestQueue_queue_dataOut_8_source2;
  wire [2:0]         exeRequestQueue_8_deq_bits_index = _exeRequestQueue_queue_fifo_8_empty ? exeRequestQueue_8_enq_bits_index : exeRequestQueue_queue_dataOut_8_index;
  wire               exeRequestQueue_8_deq_bits_ffo = _exeRequestQueue_queue_fifo_8_empty ? exeRequestQueue_8_enq_bits_ffo : exeRequestQueue_queue_dataOut_8_ffo;
  wire               tokenIO_8_maskRequestRelease_0 = exeRequestQueue_8_deq_ready & exeRequestQueue_8_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_9 = {exeRequestQueue_9_enq_bits_index, exeRequestQueue_9_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_9 = {exeRequestQueue_9_enq_bits_source1, exeRequestQueue_9_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_9 = {exeRequestQueue_queue_dataIn_hi_9, exeRequestQueue_queue_dataIn_lo_9};
  wire               exeRequestQueue_queue_dataOut_9_ffo = _exeRequestQueue_queue_fifo_9_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_9_index = _exeRequestQueue_queue_fifo_9_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_9_source2 = _exeRequestQueue_queue_fifo_9_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_9_source1 = _exeRequestQueue_queue_fifo_9_data_out[67:36];
  wire               exeRequestQueue_9_enq_ready = ~_exeRequestQueue_queue_fifo_9_full;
  wire               exeRequestQueue_9_deq_ready;
  wire               exeRequestQueue_9_deq_valid = ~_exeRequestQueue_queue_fifo_9_empty | exeRequestQueue_9_enq_valid;
  wire [31:0]        exeRequestQueue_9_deq_bits_source1 = _exeRequestQueue_queue_fifo_9_empty ? exeRequestQueue_9_enq_bits_source1 : exeRequestQueue_queue_dataOut_9_source1;
  wire [31:0]        exeRequestQueue_9_deq_bits_source2 = _exeRequestQueue_queue_fifo_9_empty ? exeRequestQueue_9_enq_bits_source2 : exeRequestQueue_queue_dataOut_9_source2;
  wire [2:0]         exeRequestQueue_9_deq_bits_index = _exeRequestQueue_queue_fifo_9_empty ? exeRequestQueue_9_enq_bits_index : exeRequestQueue_queue_dataOut_9_index;
  wire               exeRequestQueue_9_deq_bits_ffo = _exeRequestQueue_queue_fifo_9_empty ? exeRequestQueue_9_enq_bits_ffo : exeRequestQueue_queue_dataOut_9_ffo;
  wire               tokenIO_9_maskRequestRelease_0 = exeRequestQueue_9_deq_ready & exeRequestQueue_9_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_10 = {exeRequestQueue_10_enq_bits_index, exeRequestQueue_10_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_10 = {exeRequestQueue_10_enq_bits_source1, exeRequestQueue_10_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_10 = {exeRequestQueue_queue_dataIn_hi_10, exeRequestQueue_queue_dataIn_lo_10};
  wire               exeRequestQueue_queue_dataOut_10_ffo = _exeRequestQueue_queue_fifo_10_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_10_index = _exeRequestQueue_queue_fifo_10_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_10_source2 = _exeRequestQueue_queue_fifo_10_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_10_source1 = _exeRequestQueue_queue_fifo_10_data_out[67:36];
  wire               exeRequestQueue_10_enq_ready = ~_exeRequestQueue_queue_fifo_10_full;
  wire               exeRequestQueue_10_deq_ready;
  wire               exeRequestQueue_10_deq_valid = ~_exeRequestQueue_queue_fifo_10_empty | exeRequestQueue_10_enq_valid;
  wire [31:0]        exeRequestQueue_10_deq_bits_source1 = _exeRequestQueue_queue_fifo_10_empty ? exeRequestQueue_10_enq_bits_source1 : exeRequestQueue_queue_dataOut_10_source1;
  wire [31:0]        exeRequestQueue_10_deq_bits_source2 = _exeRequestQueue_queue_fifo_10_empty ? exeRequestQueue_10_enq_bits_source2 : exeRequestQueue_queue_dataOut_10_source2;
  wire [2:0]         exeRequestQueue_10_deq_bits_index = _exeRequestQueue_queue_fifo_10_empty ? exeRequestQueue_10_enq_bits_index : exeRequestQueue_queue_dataOut_10_index;
  wire               exeRequestQueue_10_deq_bits_ffo = _exeRequestQueue_queue_fifo_10_empty ? exeRequestQueue_10_enq_bits_ffo : exeRequestQueue_queue_dataOut_10_ffo;
  wire               tokenIO_10_maskRequestRelease_0 = exeRequestQueue_10_deq_ready & exeRequestQueue_10_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_11 = {exeRequestQueue_11_enq_bits_index, exeRequestQueue_11_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_11 = {exeRequestQueue_11_enq_bits_source1, exeRequestQueue_11_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_11 = {exeRequestQueue_queue_dataIn_hi_11, exeRequestQueue_queue_dataIn_lo_11};
  wire               exeRequestQueue_queue_dataOut_11_ffo = _exeRequestQueue_queue_fifo_11_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_11_index = _exeRequestQueue_queue_fifo_11_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_11_source2 = _exeRequestQueue_queue_fifo_11_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_11_source1 = _exeRequestQueue_queue_fifo_11_data_out[67:36];
  wire               exeRequestQueue_11_enq_ready = ~_exeRequestQueue_queue_fifo_11_full;
  wire               exeRequestQueue_11_deq_ready;
  wire               exeRequestQueue_11_deq_valid = ~_exeRequestQueue_queue_fifo_11_empty | exeRequestQueue_11_enq_valid;
  wire [31:0]        exeRequestQueue_11_deq_bits_source1 = _exeRequestQueue_queue_fifo_11_empty ? exeRequestQueue_11_enq_bits_source1 : exeRequestQueue_queue_dataOut_11_source1;
  wire [31:0]        exeRequestQueue_11_deq_bits_source2 = _exeRequestQueue_queue_fifo_11_empty ? exeRequestQueue_11_enq_bits_source2 : exeRequestQueue_queue_dataOut_11_source2;
  wire [2:0]         exeRequestQueue_11_deq_bits_index = _exeRequestQueue_queue_fifo_11_empty ? exeRequestQueue_11_enq_bits_index : exeRequestQueue_queue_dataOut_11_index;
  wire               exeRequestQueue_11_deq_bits_ffo = _exeRequestQueue_queue_fifo_11_empty ? exeRequestQueue_11_enq_bits_ffo : exeRequestQueue_queue_dataOut_11_ffo;
  wire               tokenIO_11_maskRequestRelease_0 = exeRequestQueue_11_deq_ready & exeRequestQueue_11_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_12 = {exeRequestQueue_12_enq_bits_index, exeRequestQueue_12_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_12 = {exeRequestQueue_12_enq_bits_source1, exeRequestQueue_12_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_12 = {exeRequestQueue_queue_dataIn_hi_12, exeRequestQueue_queue_dataIn_lo_12};
  wire               exeRequestQueue_queue_dataOut_12_ffo = _exeRequestQueue_queue_fifo_12_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_12_index = _exeRequestQueue_queue_fifo_12_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_12_source2 = _exeRequestQueue_queue_fifo_12_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_12_source1 = _exeRequestQueue_queue_fifo_12_data_out[67:36];
  wire               exeRequestQueue_12_enq_ready = ~_exeRequestQueue_queue_fifo_12_full;
  wire               exeRequestQueue_12_deq_ready;
  wire               exeRequestQueue_12_deq_valid = ~_exeRequestQueue_queue_fifo_12_empty | exeRequestQueue_12_enq_valid;
  wire [31:0]        exeRequestQueue_12_deq_bits_source1 = _exeRequestQueue_queue_fifo_12_empty ? exeRequestQueue_12_enq_bits_source1 : exeRequestQueue_queue_dataOut_12_source1;
  wire [31:0]        exeRequestQueue_12_deq_bits_source2 = _exeRequestQueue_queue_fifo_12_empty ? exeRequestQueue_12_enq_bits_source2 : exeRequestQueue_queue_dataOut_12_source2;
  wire [2:0]         exeRequestQueue_12_deq_bits_index = _exeRequestQueue_queue_fifo_12_empty ? exeRequestQueue_12_enq_bits_index : exeRequestQueue_queue_dataOut_12_index;
  wire               exeRequestQueue_12_deq_bits_ffo = _exeRequestQueue_queue_fifo_12_empty ? exeRequestQueue_12_enq_bits_ffo : exeRequestQueue_queue_dataOut_12_ffo;
  wire               tokenIO_12_maskRequestRelease_0 = exeRequestQueue_12_deq_ready & exeRequestQueue_12_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_13 = {exeRequestQueue_13_enq_bits_index, exeRequestQueue_13_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_13 = {exeRequestQueue_13_enq_bits_source1, exeRequestQueue_13_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_13 = {exeRequestQueue_queue_dataIn_hi_13, exeRequestQueue_queue_dataIn_lo_13};
  wire               exeRequestQueue_queue_dataOut_13_ffo = _exeRequestQueue_queue_fifo_13_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_13_index = _exeRequestQueue_queue_fifo_13_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_13_source2 = _exeRequestQueue_queue_fifo_13_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_13_source1 = _exeRequestQueue_queue_fifo_13_data_out[67:36];
  wire               exeRequestQueue_13_enq_ready = ~_exeRequestQueue_queue_fifo_13_full;
  wire               exeRequestQueue_13_deq_ready;
  wire               exeRequestQueue_13_deq_valid = ~_exeRequestQueue_queue_fifo_13_empty | exeRequestQueue_13_enq_valid;
  wire [31:0]        exeRequestQueue_13_deq_bits_source1 = _exeRequestQueue_queue_fifo_13_empty ? exeRequestQueue_13_enq_bits_source1 : exeRequestQueue_queue_dataOut_13_source1;
  wire [31:0]        exeRequestQueue_13_deq_bits_source2 = _exeRequestQueue_queue_fifo_13_empty ? exeRequestQueue_13_enq_bits_source2 : exeRequestQueue_queue_dataOut_13_source2;
  wire [2:0]         exeRequestQueue_13_deq_bits_index = _exeRequestQueue_queue_fifo_13_empty ? exeRequestQueue_13_enq_bits_index : exeRequestQueue_queue_dataOut_13_index;
  wire               exeRequestQueue_13_deq_bits_ffo = _exeRequestQueue_queue_fifo_13_empty ? exeRequestQueue_13_enq_bits_ffo : exeRequestQueue_queue_dataOut_13_ffo;
  wire               tokenIO_13_maskRequestRelease_0 = exeRequestQueue_13_deq_ready & exeRequestQueue_13_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_14 = {exeRequestQueue_14_enq_bits_index, exeRequestQueue_14_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_14 = {exeRequestQueue_14_enq_bits_source1, exeRequestQueue_14_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_14 = {exeRequestQueue_queue_dataIn_hi_14, exeRequestQueue_queue_dataIn_lo_14};
  wire               exeRequestQueue_queue_dataOut_14_ffo = _exeRequestQueue_queue_fifo_14_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_14_index = _exeRequestQueue_queue_fifo_14_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_14_source2 = _exeRequestQueue_queue_fifo_14_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_14_source1 = _exeRequestQueue_queue_fifo_14_data_out[67:36];
  wire               exeRequestQueue_14_enq_ready = ~_exeRequestQueue_queue_fifo_14_full;
  wire               exeRequestQueue_14_deq_ready;
  wire               exeRequestQueue_14_deq_valid = ~_exeRequestQueue_queue_fifo_14_empty | exeRequestQueue_14_enq_valid;
  wire [31:0]        exeRequestQueue_14_deq_bits_source1 = _exeRequestQueue_queue_fifo_14_empty ? exeRequestQueue_14_enq_bits_source1 : exeRequestQueue_queue_dataOut_14_source1;
  wire [31:0]        exeRequestQueue_14_deq_bits_source2 = _exeRequestQueue_queue_fifo_14_empty ? exeRequestQueue_14_enq_bits_source2 : exeRequestQueue_queue_dataOut_14_source2;
  wire [2:0]         exeRequestQueue_14_deq_bits_index = _exeRequestQueue_queue_fifo_14_empty ? exeRequestQueue_14_enq_bits_index : exeRequestQueue_queue_dataOut_14_index;
  wire               exeRequestQueue_14_deq_bits_ffo = _exeRequestQueue_queue_fifo_14_empty ? exeRequestQueue_14_enq_bits_ffo : exeRequestQueue_queue_dataOut_14_ffo;
  wire               tokenIO_14_maskRequestRelease_0 = exeRequestQueue_14_deq_ready & exeRequestQueue_14_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_15 = {exeRequestQueue_15_enq_bits_index, exeRequestQueue_15_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_15 = {exeRequestQueue_15_enq_bits_source1, exeRequestQueue_15_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_15 = {exeRequestQueue_queue_dataIn_hi_15, exeRequestQueue_queue_dataIn_lo_15};
  wire               exeRequestQueue_queue_dataOut_15_ffo = _exeRequestQueue_queue_fifo_15_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_15_index = _exeRequestQueue_queue_fifo_15_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_15_source2 = _exeRequestQueue_queue_fifo_15_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_15_source1 = _exeRequestQueue_queue_fifo_15_data_out[67:36];
  wire               exeRequestQueue_15_enq_ready = ~_exeRequestQueue_queue_fifo_15_full;
  wire               exeRequestQueue_15_deq_ready;
  wire               exeRequestQueue_15_deq_valid = ~_exeRequestQueue_queue_fifo_15_empty | exeRequestQueue_15_enq_valid;
  wire [31:0]        exeRequestQueue_15_deq_bits_source1 = _exeRequestQueue_queue_fifo_15_empty ? exeRequestQueue_15_enq_bits_source1 : exeRequestQueue_queue_dataOut_15_source1;
  wire [31:0]        exeRequestQueue_15_deq_bits_source2 = _exeRequestQueue_queue_fifo_15_empty ? exeRequestQueue_15_enq_bits_source2 : exeRequestQueue_queue_dataOut_15_source2;
  wire [2:0]         exeRequestQueue_15_deq_bits_index = _exeRequestQueue_queue_fifo_15_empty ? exeRequestQueue_15_enq_bits_index : exeRequestQueue_queue_dataOut_15_index;
  wire               exeRequestQueue_15_deq_bits_ffo = _exeRequestQueue_queue_fifo_15_empty ? exeRequestQueue_15_enq_bits_ffo : exeRequestQueue_queue_dataOut_15_ffo;
  wire               tokenIO_15_maskRequestRelease_0 = exeRequestQueue_15_deq_ready & exeRequestQueue_15_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_16 = {exeRequestQueue_16_enq_bits_index, exeRequestQueue_16_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_16 = {exeRequestQueue_16_enq_bits_source1, exeRequestQueue_16_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_16 = {exeRequestQueue_queue_dataIn_hi_16, exeRequestQueue_queue_dataIn_lo_16};
  wire               exeRequestQueue_queue_dataOut_16_ffo = _exeRequestQueue_queue_fifo_16_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_16_index = _exeRequestQueue_queue_fifo_16_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_16_source2 = _exeRequestQueue_queue_fifo_16_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_16_source1 = _exeRequestQueue_queue_fifo_16_data_out[67:36];
  wire               exeRequestQueue_16_enq_ready = ~_exeRequestQueue_queue_fifo_16_full;
  wire               exeRequestQueue_16_deq_ready;
  wire               exeRequestQueue_16_deq_valid = ~_exeRequestQueue_queue_fifo_16_empty | exeRequestQueue_16_enq_valid;
  wire [31:0]        exeRequestQueue_16_deq_bits_source1 = _exeRequestQueue_queue_fifo_16_empty ? exeRequestQueue_16_enq_bits_source1 : exeRequestQueue_queue_dataOut_16_source1;
  wire [31:0]        exeRequestQueue_16_deq_bits_source2 = _exeRequestQueue_queue_fifo_16_empty ? exeRequestQueue_16_enq_bits_source2 : exeRequestQueue_queue_dataOut_16_source2;
  wire [2:0]         exeRequestQueue_16_deq_bits_index = _exeRequestQueue_queue_fifo_16_empty ? exeRequestQueue_16_enq_bits_index : exeRequestQueue_queue_dataOut_16_index;
  wire               exeRequestQueue_16_deq_bits_ffo = _exeRequestQueue_queue_fifo_16_empty ? exeRequestQueue_16_enq_bits_ffo : exeRequestQueue_queue_dataOut_16_ffo;
  wire               tokenIO_16_maskRequestRelease_0 = exeRequestQueue_16_deq_ready & exeRequestQueue_16_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_17 = {exeRequestQueue_17_enq_bits_index, exeRequestQueue_17_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_17 = {exeRequestQueue_17_enq_bits_source1, exeRequestQueue_17_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_17 = {exeRequestQueue_queue_dataIn_hi_17, exeRequestQueue_queue_dataIn_lo_17};
  wire               exeRequestQueue_queue_dataOut_17_ffo = _exeRequestQueue_queue_fifo_17_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_17_index = _exeRequestQueue_queue_fifo_17_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_17_source2 = _exeRequestQueue_queue_fifo_17_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_17_source1 = _exeRequestQueue_queue_fifo_17_data_out[67:36];
  wire               exeRequestQueue_17_enq_ready = ~_exeRequestQueue_queue_fifo_17_full;
  wire               exeRequestQueue_17_deq_ready;
  wire               exeRequestQueue_17_deq_valid = ~_exeRequestQueue_queue_fifo_17_empty | exeRequestQueue_17_enq_valid;
  wire [31:0]        exeRequestQueue_17_deq_bits_source1 = _exeRequestQueue_queue_fifo_17_empty ? exeRequestQueue_17_enq_bits_source1 : exeRequestQueue_queue_dataOut_17_source1;
  wire [31:0]        exeRequestQueue_17_deq_bits_source2 = _exeRequestQueue_queue_fifo_17_empty ? exeRequestQueue_17_enq_bits_source2 : exeRequestQueue_queue_dataOut_17_source2;
  wire [2:0]         exeRequestQueue_17_deq_bits_index = _exeRequestQueue_queue_fifo_17_empty ? exeRequestQueue_17_enq_bits_index : exeRequestQueue_queue_dataOut_17_index;
  wire               exeRequestQueue_17_deq_bits_ffo = _exeRequestQueue_queue_fifo_17_empty ? exeRequestQueue_17_enq_bits_ffo : exeRequestQueue_queue_dataOut_17_ffo;
  wire               tokenIO_17_maskRequestRelease_0 = exeRequestQueue_17_deq_ready & exeRequestQueue_17_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_18 = {exeRequestQueue_18_enq_bits_index, exeRequestQueue_18_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_18 = {exeRequestQueue_18_enq_bits_source1, exeRequestQueue_18_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_18 = {exeRequestQueue_queue_dataIn_hi_18, exeRequestQueue_queue_dataIn_lo_18};
  wire               exeRequestQueue_queue_dataOut_18_ffo = _exeRequestQueue_queue_fifo_18_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_18_index = _exeRequestQueue_queue_fifo_18_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_18_source2 = _exeRequestQueue_queue_fifo_18_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_18_source1 = _exeRequestQueue_queue_fifo_18_data_out[67:36];
  wire               exeRequestQueue_18_enq_ready = ~_exeRequestQueue_queue_fifo_18_full;
  wire               exeRequestQueue_18_deq_ready;
  wire               exeRequestQueue_18_deq_valid = ~_exeRequestQueue_queue_fifo_18_empty | exeRequestQueue_18_enq_valid;
  wire [31:0]        exeRequestQueue_18_deq_bits_source1 = _exeRequestQueue_queue_fifo_18_empty ? exeRequestQueue_18_enq_bits_source1 : exeRequestQueue_queue_dataOut_18_source1;
  wire [31:0]        exeRequestQueue_18_deq_bits_source2 = _exeRequestQueue_queue_fifo_18_empty ? exeRequestQueue_18_enq_bits_source2 : exeRequestQueue_queue_dataOut_18_source2;
  wire [2:0]         exeRequestQueue_18_deq_bits_index = _exeRequestQueue_queue_fifo_18_empty ? exeRequestQueue_18_enq_bits_index : exeRequestQueue_queue_dataOut_18_index;
  wire               exeRequestQueue_18_deq_bits_ffo = _exeRequestQueue_queue_fifo_18_empty ? exeRequestQueue_18_enq_bits_ffo : exeRequestQueue_queue_dataOut_18_ffo;
  wire               tokenIO_18_maskRequestRelease_0 = exeRequestQueue_18_deq_ready & exeRequestQueue_18_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_19 = {exeRequestQueue_19_enq_bits_index, exeRequestQueue_19_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_19 = {exeRequestQueue_19_enq_bits_source1, exeRequestQueue_19_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_19 = {exeRequestQueue_queue_dataIn_hi_19, exeRequestQueue_queue_dataIn_lo_19};
  wire               exeRequestQueue_queue_dataOut_19_ffo = _exeRequestQueue_queue_fifo_19_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_19_index = _exeRequestQueue_queue_fifo_19_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_19_source2 = _exeRequestQueue_queue_fifo_19_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_19_source1 = _exeRequestQueue_queue_fifo_19_data_out[67:36];
  wire               exeRequestQueue_19_enq_ready = ~_exeRequestQueue_queue_fifo_19_full;
  wire               exeRequestQueue_19_deq_ready;
  wire               exeRequestQueue_19_deq_valid = ~_exeRequestQueue_queue_fifo_19_empty | exeRequestQueue_19_enq_valid;
  wire [31:0]        exeRequestQueue_19_deq_bits_source1 = _exeRequestQueue_queue_fifo_19_empty ? exeRequestQueue_19_enq_bits_source1 : exeRequestQueue_queue_dataOut_19_source1;
  wire [31:0]        exeRequestQueue_19_deq_bits_source2 = _exeRequestQueue_queue_fifo_19_empty ? exeRequestQueue_19_enq_bits_source2 : exeRequestQueue_queue_dataOut_19_source2;
  wire [2:0]         exeRequestQueue_19_deq_bits_index = _exeRequestQueue_queue_fifo_19_empty ? exeRequestQueue_19_enq_bits_index : exeRequestQueue_queue_dataOut_19_index;
  wire               exeRequestQueue_19_deq_bits_ffo = _exeRequestQueue_queue_fifo_19_empty ? exeRequestQueue_19_enq_bits_ffo : exeRequestQueue_queue_dataOut_19_ffo;
  wire               tokenIO_19_maskRequestRelease_0 = exeRequestQueue_19_deq_ready & exeRequestQueue_19_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_20 = {exeRequestQueue_20_enq_bits_index, exeRequestQueue_20_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_20 = {exeRequestQueue_20_enq_bits_source1, exeRequestQueue_20_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_20 = {exeRequestQueue_queue_dataIn_hi_20, exeRequestQueue_queue_dataIn_lo_20};
  wire               exeRequestQueue_queue_dataOut_20_ffo = _exeRequestQueue_queue_fifo_20_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_20_index = _exeRequestQueue_queue_fifo_20_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_20_source2 = _exeRequestQueue_queue_fifo_20_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_20_source1 = _exeRequestQueue_queue_fifo_20_data_out[67:36];
  wire               exeRequestQueue_20_enq_ready = ~_exeRequestQueue_queue_fifo_20_full;
  wire               exeRequestQueue_20_deq_ready;
  wire               exeRequestQueue_20_deq_valid = ~_exeRequestQueue_queue_fifo_20_empty | exeRequestQueue_20_enq_valid;
  wire [31:0]        exeRequestQueue_20_deq_bits_source1 = _exeRequestQueue_queue_fifo_20_empty ? exeRequestQueue_20_enq_bits_source1 : exeRequestQueue_queue_dataOut_20_source1;
  wire [31:0]        exeRequestQueue_20_deq_bits_source2 = _exeRequestQueue_queue_fifo_20_empty ? exeRequestQueue_20_enq_bits_source2 : exeRequestQueue_queue_dataOut_20_source2;
  wire [2:0]         exeRequestQueue_20_deq_bits_index = _exeRequestQueue_queue_fifo_20_empty ? exeRequestQueue_20_enq_bits_index : exeRequestQueue_queue_dataOut_20_index;
  wire               exeRequestQueue_20_deq_bits_ffo = _exeRequestQueue_queue_fifo_20_empty ? exeRequestQueue_20_enq_bits_ffo : exeRequestQueue_queue_dataOut_20_ffo;
  wire               tokenIO_20_maskRequestRelease_0 = exeRequestQueue_20_deq_ready & exeRequestQueue_20_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_21 = {exeRequestQueue_21_enq_bits_index, exeRequestQueue_21_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_21 = {exeRequestQueue_21_enq_bits_source1, exeRequestQueue_21_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_21 = {exeRequestQueue_queue_dataIn_hi_21, exeRequestQueue_queue_dataIn_lo_21};
  wire               exeRequestQueue_queue_dataOut_21_ffo = _exeRequestQueue_queue_fifo_21_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_21_index = _exeRequestQueue_queue_fifo_21_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_21_source2 = _exeRequestQueue_queue_fifo_21_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_21_source1 = _exeRequestQueue_queue_fifo_21_data_out[67:36];
  wire               exeRequestQueue_21_enq_ready = ~_exeRequestQueue_queue_fifo_21_full;
  wire               exeRequestQueue_21_deq_ready;
  wire               exeRequestQueue_21_deq_valid = ~_exeRequestQueue_queue_fifo_21_empty | exeRequestQueue_21_enq_valid;
  wire [31:0]        exeRequestQueue_21_deq_bits_source1 = _exeRequestQueue_queue_fifo_21_empty ? exeRequestQueue_21_enq_bits_source1 : exeRequestQueue_queue_dataOut_21_source1;
  wire [31:0]        exeRequestQueue_21_deq_bits_source2 = _exeRequestQueue_queue_fifo_21_empty ? exeRequestQueue_21_enq_bits_source2 : exeRequestQueue_queue_dataOut_21_source2;
  wire [2:0]         exeRequestQueue_21_deq_bits_index = _exeRequestQueue_queue_fifo_21_empty ? exeRequestQueue_21_enq_bits_index : exeRequestQueue_queue_dataOut_21_index;
  wire               exeRequestQueue_21_deq_bits_ffo = _exeRequestQueue_queue_fifo_21_empty ? exeRequestQueue_21_enq_bits_ffo : exeRequestQueue_queue_dataOut_21_ffo;
  wire               tokenIO_21_maskRequestRelease_0 = exeRequestQueue_21_deq_ready & exeRequestQueue_21_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_22 = {exeRequestQueue_22_enq_bits_index, exeRequestQueue_22_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_22 = {exeRequestQueue_22_enq_bits_source1, exeRequestQueue_22_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_22 = {exeRequestQueue_queue_dataIn_hi_22, exeRequestQueue_queue_dataIn_lo_22};
  wire               exeRequestQueue_queue_dataOut_22_ffo = _exeRequestQueue_queue_fifo_22_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_22_index = _exeRequestQueue_queue_fifo_22_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_22_source2 = _exeRequestQueue_queue_fifo_22_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_22_source1 = _exeRequestQueue_queue_fifo_22_data_out[67:36];
  wire               exeRequestQueue_22_enq_ready = ~_exeRequestQueue_queue_fifo_22_full;
  wire               exeRequestQueue_22_deq_ready;
  wire               exeRequestQueue_22_deq_valid = ~_exeRequestQueue_queue_fifo_22_empty | exeRequestQueue_22_enq_valid;
  wire [31:0]        exeRequestQueue_22_deq_bits_source1 = _exeRequestQueue_queue_fifo_22_empty ? exeRequestQueue_22_enq_bits_source1 : exeRequestQueue_queue_dataOut_22_source1;
  wire [31:0]        exeRequestQueue_22_deq_bits_source2 = _exeRequestQueue_queue_fifo_22_empty ? exeRequestQueue_22_enq_bits_source2 : exeRequestQueue_queue_dataOut_22_source2;
  wire [2:0]         exeRequestQueue_22_deq_bits_index = _exeRequestQueue_queue_fifo_22_empty ? exeRequestQueue_22_enq_bits_index : exeRequestQueue_queue_dataOut_22_index;
  wire               exeRequestQueue_22_deq_bits_ffo = _exeRequestQueue_queue_fifo_22_empty ? exeRequestQueue_22_enq_bits_ffo : exeRequestQueue_queue_dataOut_22_ffo;
  wire               tokenIO_22_maskRequestRelease_0 = exeRequestQueue_22_deq_ready & exeRequestQueue_22_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_23 = {exeRequestQueue_23_enq_bits_index, exeRequestQueue_23_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_23 = {exeRequestQueue_23_enq_bits_source1, exeRequestQueue_23_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_23 = {exeRequestQueue_queue_dataIn_hi_23, exeRequestQueue_queue_dataIn_lo_23};
  wire               exeRequestQueue_queue_dataOut_23_ffo = _exeRequestQueue_queue_fifo_23_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_23_index = _exeRequestQueue_queue_fifo_23_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_23_source2 = _exeRequestQueue_queue_fifo_23_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_23_source1 = _exeRequestQueue_queue_fifo_23_data_out[67:36];
  wire               exeRequestQueue_23_enq_ready = ~_exeRequestQueue_queue_fifo_23_full;
  wire               exeRequestQueue_23_deq_ready;
  wire               exeRequestQueue_23_deq_valid = ~_exeRequestQueue_queue_fifo_23_empty | exeRequestQueue_23_enq_valid;
  wire [31:0]        exeRequestQueue_23_deq_bits_source1 = _exeRequestQueue_queue_fifo_23_empty ? exeRequestQueue_23_enq_bits_source1 : exeRequestQueue_queue_dataOut_23_source1;
  wire [31:0]        exeRequestQueue_23_deq_bits_source2 = _exeRequestQueue_queue_fifo_23_empty ? exeRequestQueue_23_enq_bits_source2 : exeRequestQueue_queue_dataOut_23_source2;
  wire [2:0]         exeRequestQueue_23_deq_bits_index = _exeRequestQueue_queue_fifo_23_empty ? exeRequestQueue_23_enq_bits_index : exeRequestQueue_queue_dataOut_23_index;
  wire               exeRequestQueue_23_deq_bits_ffo = _exeRequestQueue_queue_fifo_23_empty ? exeRequestQueue_23_enq_bits_ffo : exeRequestQueue_queue_dataOut_23_ffo;
  wire               tokenIO_23_maskRequestRelease_0 = exeRequestQueue_23_deq_ready & exeRequestQueue_23_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_24 = {exeRequestQueue_24_enq_bits_index, exeRequestQueue_24_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_24 = {exeRequestQueue_24_enq_bits_source1, exeRequestQueue_24_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_24 = {exeRequestQueue_queue_dataIn_hi_24, exeRequestQueue_queue_dataIn_lo_24};
  wire               exeRequestQueue_queue_dataOut_24_ffo = _exeRequestQueue_queue_fifo_24_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_24_index = _exeRequestQueue_queue_fifo_24_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_24_source2 = _exeRequestQueue_queue_fifo_24_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_24_source1 = _exeRequestQueue_queue_fifo_24_data_out[67:36];
  wire               exeRequestQueue_24_enq_ready = ~_exeRequestQueue_queue_fifo_24_full;
  wire               exeRequestQueue_24_deq_ready;
  wire               exeRequestQueue_24_deq_valid = ~_exeRequestQueue_queue_fifo_24_empty | exeRequestQueue_24_enq_valid;
  wire [31:0]        exeRequestQueue_24_deq_bits_source1 = _exeRequestQueue_queue_fifo_24_empty ? exeRequestQueue_24_enq_bits_source1 : exeRequestQueue_queue_dataOut_24_source1;
  wire [31:0]        exeRequestQueue_24_deq_bits_source2 = _exeRequestQueue_queue_fifo_24_empty ? exeRequestQueue_24_enq_bits_source2 : exeRequestQueue_queue_dataOut_24_source2;
  wire [2:0]         exeRequestQueue_24_deq_bits_index = _exeRequestQueue_queue_fifo_24_empty ? exeRequestQueue_24_enq_bits_index : exeRequestQueue_queue_dataOut_24_index;
  wire               exeRequestQueue_24_deq_bits_ffo = _exeRequestQueue_queue_fifo_24_empty ? exeRequestQueue_24_enq_bits_ffo : exeRequestQueue_queue_dataOut_24_ffo;
  wire               tokenIO_24_maskRequestRelease_0 = exeRequestQueue_24_deq_ready & exeRequestQueue_24_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_25 = {exeRequestQueue_25_enq_bits_index, exeRequestQueue_25_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_25 = {exeRequestQueue_25_enq_bits_source1, exeRequestQueue_25_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_25 = {exeRequestQueue_queue_dataIn_hi_25, exeRequestQueue_queue_dataIn_lo_25};
  wire               exeRequestQueue_queue_dataOut_25_ffo = _exeRequestQueue_queue_fifo_25_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_25_index = _exeRequestQueue_queue_fifo_25_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_25_source2 = _exeRequestQueue_queue_fifo_25_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_25_source1 = _exeRequestQueue_queue_fifo_25_data_out[67:36];
  wire               exeRequestQueue_25_enq_ready = ~_exeRequestQueue_queue_fifo_25_full;
  wire               exeRequestQueue_25_deq_ready;
  wire               exeRequestQueue_25_deq_valid = ~_exeRequestQueue_queue_fifo_25_empty | exeRequestQueue_25_enq_valid;
  wire [31:0]        exeRequestQueue_25_deq_bits_source1 = _exeRequestQueue_queue_fifo_25_empty ? exeRequestQueue_25_enq_bits_source1 : exeRequestQueue_queue_dataOut_25_source1;
  wire [31:0]        exeRequestQueue_25_deq_bits_source2 = _exeRequestQueue_queue_fifo_25_empty ? exeRequestQueue_25_enq_bits_source2 : exeRequestQueue_queue_dataOut_25_source2;
  wire [2:0]         exeRequestQueue_25_deq_bits_index = _exeRequestQueue_queue_fifo_25_empty ? exeRequestQueue_25_enq_bits_index : exeRequestQueue_queue_dataOut_25_index;
  wire               exeRequestQueue_25_deq_bits_ffo = _exeRequestQueue_queue_fifo_25_empty ? exeRequestQueue_25_enq_bits_ffo : exeRequestQueue_queue_dataOut_25_ffo;
  wire               tokenIO_25_maskRequestRelease_0 = exeRequestQueue_25_deq_ready & exeRequestQueue_25_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_26 = {exeRequestQueue_26_enq_bits_index, exeRequestQueue_26_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_26 = {exeRequestQueue_26_enq_bits_source1, exeRequestQueue_26_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_26 = {exeRequestQueue_queue_dataIn_hi_26, exeRequestQueue_queue_dataIn_lo_26};
  wire               exeRequestQueue_queue_dataOut_26_ffo = _exeRequestQueue_queue_fifo_26_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_26_index = _exeRequestQueue_queue_fifo_26_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_26_source2 = _exeRequestQueue_queue_fifo_26_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_26_source1 = _exeRequestQueue_queue_fifo_26_data_out[67:36];
  wire               exeRequestQueue_26_enq_ready = ~_exeRequestQueue_queue_fifo_26_full;
  wire               exeRequestQueue_26_deq_ready;
  wire               exeRequestQueue_26_deq_valid = ~_exeRequestQueue_queue_fifo_26_empty | exeRequestQueue_26_enq_valid;
  wire [31:0]        exeRequestQueue_26_deq_bits_source1 = _exeRequestQueue_queue_fifo_26_empty ? exeRequestQueue_26_enq_bits_source1 : exeRequestQueue_queue_dataOut_26_source1;
  wire [31:0]        exeRequestQueue_26_deq_bits_source2 = _exeRequestQueue_queue_fifo_26_empty ? exeRequestQueue_26_enq_bits_source2 : exeRequestQueue_queue_dataOut_26_source2;
  wire [2:0]         exeRequestQueue_26_deq_bits_index = _exeRequestQueue_queue_fifo_26_empty ? exeRequestQueue_26_enq_bits_index : exeRequestQueue_queue_dataOut_26_index;
  wire               exeRequestQueue_26_deq_bits_ffo = _exeRequestQueue_queue_fifo_26_empty ? exeRequestQueue_26_enq_bits_ffo : exeRequestQueue_queue_dataOut_26_ffo;
  wire               tokenIO_26_maskRequestRelease_0 = exeRequestQueue_26_deq_ready & exeRequestQueue_26_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_27 = {exeRequestQueue_27_enq_bits_index, exeRequestQueue_27_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_27 = {exeRequestQueue_27_enq_bits_source1, exeRequestQueue_27_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_27 = {exeRequestQueue_queue_dataIn_hi_27, exeRequestQueue_queue_dataIn_lo_27};
  wire               exeRequestQueue_queue_dataOut_27_ffo = _exeRequestQueue_queue_fifo_27_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_27_index = _exeRequestQueue_queue_fifo_27_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_27_source2 = _exeRequestQueue_queue_fifo_27_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_27_source1 = _exeRequestQueue_queue_fifo_27_data_out[67:36];
  wire               exeRequestQueue_27_enq_ready = ~_exeRequestQueue_queue_fifo_27_full;
  wire               exeRequestQueue_27_deq_ready;
  wire               exeRequestQueue_27_deq_valid = ~_exeRequestQueue_queue_fifo_27_empty | exeRequestQueue_27_enq_valid;
  wire [31:0]        exeRequestQueue_27_deq_bits_source1 = _exeRequestQueue_queue_fifo_27_empty ? exeRequestQueue_27_enq_bits_source1 : exeRequestQueue_queue_dataOut_27_source1;
  wire [31:0]        exeRequestQueue_27_deq_bits_source2 = _exeRequestQueue_queue_fifo_27_empty ? exeRequestQueue_27_enq_bits_source2 : exeRequestQueue_queue_dataOut_27_source2;
  wire [2:0]         exeRequestQueue_27_deq_bits_index = _exeRequestQueue_queue_fifo_27_empty ? exeRequestQueue_27_enq_bits_index : exeRequestQueue_queue_dataOut_27_index;
  wire               exeRequestQueue_27_deq_bits_ffo = _exeRequestQueue_queue_fifo_27_empty ? exeRequestQueue_27_enq_bits_ffo : exeRequestQueue_queue_dataOut_27_ffo;
  wire               tokenIO_27_maskRequestRelease_0 = exeRequestQueue_27_deq_ready & exeRequestQueue_27_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_28 = {exeRequestQueue_28_enq_bits_index, exeRequestQueue_28_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_28 = {exeRequestQueue_28_enq_bits_source1, exeRequestQueue_28_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_28 = {exeRequestQueue_queue_dataIn_hi_28, exeRequestQueue_queue_dataIn_lo_28};
  wire               exeRequestQueue_queue_dataOut_28_ffo = _exeRequestQueue_queue_fifo_28_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_28_index = _exeRequestQueue_queue_fifo_28_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_28_source2 = _exeRequestQueue_queue_fifo_28_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_28_source1 = _exeRequestQueue_queue_fifo_28_data_out[67:36];
  wire               exeRequestQueue_28_enq_ready = ~_exeRequestQueue_queue_fifo_28_full;
  wire               exeRequestQueue_28_deq_ready;
  wire               exeRequestQueue_28_deq_valid = ~_exeRequestQueue_queue_fifo_28_empty | exeRequestQueue_28_enq_valid;
  wire [31:0]        exeRequestQueue_28_deq_bits_source1 = _exeRequestQueue_queue_fifo_28_empty ? exeRequestQueue_28_enq_bits_source1 : exeRequestQueue_queue_dataOut_28_source1;
  wire [31:0]        exeRequestQueue_28_deq_bits_source2 = _exeRequestQueue_queue_fifo_28_empty ? exeRequestQueue_28_enq_bits_source2 : exeRequestQueue_queue_dataOut_28_source2;
  wire [2:0]         exeRequestQueue_28_deq_bits_index = _exeRequestQueue_queue_fifo_28_empty ? exeRequestQueue_28_enq_bits_index : exeRequestQueue_queue_dataOut_28_index;
  wire               exeRequestQueue_28_deq_bits_ffo = _exeRequestQueue_queue_fifo_28_empty ? exeRequestQueue_28_enq_bits_ffo : exeRequestQueue_queue_dataOut_28_ffo;
  wire               tokenIO_28_maskRequestRelease_0 = exeRequestQueue_28_deq_ready & exeRequestQueue_28_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_29 = {exeRequestQueue_29_enq_bits_index, exeRequestQueue_29_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_29 = {exeRequestQueue_29_enq_bits_source1, exeRequestQueue_29_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_29 = {exeRequestQueue_queue_dataIn_hi_29, exeRequestQueue_queue_dataIn_lo_29};
  wire               exeRequestQueue_queue_dataOut_29_ffo = _exeRequestQueue_queue_fifo_29_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_29_index = _exeRequestQueue_queue_fifo_29_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_29_source2 = _exeRequestQueue_queue_fifo_29_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_29_source1 = _exeRequestQueue_queue_fifo_29_data_out[67:36];
  wire               exeRequestQueue_29_enq_ready = ~_exeRequestQueue_queue_fifo_29_full;
  wire               exeRequestQueue_29_deq_ready;
  wire               exeRequestQueue_29_deq_valid = ~_exeRequestQueue_queue_fifo_29_empty | exeRequestQueue_29_enq_valid;
  wire [31:0]        exeRequestQueue_29_deq_bits_source1 = _exeRequestQueue_queue_fifo_29_empty ? exeRequestQueue_29_enq_bits_source1 : exeRequestQueue_queue_dataOut_29_source1;
  wire [31:0]        exeRequestQueue_29_deq_bits_source2 = _exeRequestQueue_queue_fifo_29_empty ? exeRequestQueue_29_enq_bits_source2 : exeRequestQueue_queue_dataOut_29_source2;
  wire [2:0]         exeRequestQueue_29_deq_bits_index = _exeRequestQueue_queue_fifo_29_empty ? exeRequestQueue_29_enq_bits_index : exeRequestQueue_queue_dataOut_29_index;
  wire               exeRequestQueue_29_deq_bits_ffo = _exeRequestQueue_queue_fifo_29_empty ? exeRequestQueue_29_enq_bits_ffo : exeRequestQueue_queue_dataOut_29_ffo;
  wire               tokenIO_29_maskRequestRelease_0 = exeRequestQueue_29_deq_ready & exeRequestQueue_29_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_30 = {exeRequestQueue_30_enq_bits_index, exeRequestQueue_30_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_30 = {exeRequestQueue_30_enq_bits_source1, exeRequestQueue_30_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_30 = {exeRequestQueue_queue_dataIn_hi_30, exeRequestQueue_queue_dataIn_lo_30};
  wire               exeRequestQueue_queue_dataOut_30_ffo = _exeRequestQueue_queue_fifo_30_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_30_index = _exeRequestQueue_queue_fifo_30_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_30_source2 = _exeRequestQueue_queue_fifo_30_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_30_source1 = _exeRequestQueue_queue_fifo_30_data_out[67:36];
  wire               exeRequestQueue_30_enq_ready = ~_exeRequestQueue_queue_fifo_30_full;
  wire               exeRequestQueue_30_deq_ready;
  wire               exeRequestQueue_30_deq_valid = ~_exeRequestQueue_queue_fifo_30_empty | exeRequestQueue_30_enq_valid;
  wire [31:0]        exeRequestQueue_30_deq_bits_source1 = _exeRequestQueue_queue_fifo_30_empty ? exeRequestQueue_30_enq_bits_source1 : exeRequestQueue_queue_dataOut_30_source1;
  wire [31:0]        exeRequestQueue_30_deq_bits_source2 = _exeRequestQueue_queue_fifo_30_empty ? exeRequestQueue_30_enq_bits_source2 : exeRequestQueue_queue_dataOut_30_source2;
  wire [2:0]         exeRequestQueue_30_deq_bits_index = _exeRequestQueue_queue_fifo_30_empty ? exeRequestQueue_30_enq_bits_index : exeRequestQueue_queue_dataOut_30_index;
  wire               exeRequestQueue_30_deq_bits_ffo = _exeRequestQueue_queue_fifo_30_empty ? exeRequestQueue_30_enq_bits_ffo : exeRequestQueue_queue_dataOut_30_ffo;
  wire               tokenIO_30_maskRequestRelease_0 = exeRequestQueue_30_deq_ready & exeRequestQueue_30_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_31 = {exeRequestQueue_31_enq_bits_index, exeRequestQueue_31_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_31 = {exeRequestQueue_31_enq_bits_source1, exeRequestQueue_31_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_31 = {exeRequestQueue_queue_dataIn_hi_31, exeRequestQueue_queue_dataIn_lo_31};
  wire               exeRequestQueue_queue_dataOut_31_ffo = _exeRequestQueue_queue_fifo_31_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_31_index = _exeRequestQueue_queue_fifo_31_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_31_source2 = _exeRequestQueue_queue_fifo_31_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_31_source1 = _exeRequestQueue_queue_fifo_31_data_out[67:36];
  wire               exeRequestQueue_31_enq_ready = ~_exeRequestQueue_queue_fifo_31_full;
  wire               exeRequestQueue_31_deq_ready;
  wire               exeRequestQueue_31_deq_valid = ~_exeRequestQueue_queue_fifo_31_empty | exeRequestQueue_31_enq_valid;
  wire [31:0]        exeRequestQueue_31_deq_bits_source1 = _exeRequestQueue_queue_fifo_31_empty ? exeRequestQueue_31_enq_bits_source1 : exeRequestQueue_queue_dataOut_31_source1;
  wire [31:0]        exeRequestQueue_31_deq_bits_source2 = _exeRequestQueue_queue_fifo_31_empty ? exeRequestQueue_31_enq_bits_source2 : exeRequestQueue_queue_dataOut_31_source2;
  wire [2:0]         exeRequestQueue_31_deq_bits_index = _exeRequestQueue_queue_fifo_31_empty ? exeRequestQueue_31_enq_bits_index : exeRequestQueue_queue_dataOut_31_index;
  wire               exeRequestQueue_31_deq_bits_ffo = _exeRequestQueue_queue_fifo_31_empty ? exeRequestQueue_31_enq_bits_ffo : exeRequestQueue_queue_dataOut_31_ffo;
  wire               tokenIO_31_maskRequestRelease_0 = exeRequestQueue_31_deq_ready & exeRequestQueue_31_deq_valid;
  reg                exeReqReg_0_valid;
  reg  [31:0]        exeReqReg_0_bits_source1;
  reg  [31:0]        exeReqReg_0_bits_source2;
  reg  [2:0]         exeReqReg_0_bits_index;
  reg                exeReqReg_0_bits_ffo;
  reg                exeReqReg_1_valid;
  reg  [31:0]        exeReqReg_1_bits_source1;
  reg  [31:0]        exeReqReg_1_bits_source2;
  reg  [2:0]         exeReqReg_1_bits_index;
  reg                exeReqReg_1_bits_ffo;
  reg                exeReqReg_2_valid;
  reg  [31:0]        exeReqReg_2_bits_source1;
  reg  [31:0]        exeReqReg_2_bits_source2;
  reg  [2:0]         exeReqReg_2_bits_index;
  reg                exeReqReg_2_bits_ffo;
  reg                exeReqReg_3_valid;
  reg  [31:0]        exeReqReg_3_bits_source1;
  reg  [31:0]        exeReqReg_3_bits_source2;
  reg  [2:0]         exeReqReg_3_bits_index;
  reg                exeReqReg_3_bits_ffo;
  reg                exeReqReg_4_valid;
  reg  [31:0]        exeReqReg_4_bits_source1;
  reg  [31:0]        exeReqReg_4_bits_source2;
  reg  [2:0]         exeReqReg_4_bits_index;
  reg                exeReqReg_4_bits_ffo;
  reg                exeReqReg_5_valid;
  reg  [31:0]        exeReqReg_5_bits_source1;
  reg  [31:0]        exeReqReg_5_bits_source2;
  reg  [2:0]         exeReqReg_5_bits_index;
  reg                exeReqReg_5_bits_ffo;
  reg                exeReqReg_6_valid;
  reg  [31:0]        exeReqReg_6_bits_source1;
  reg  [31:0]        exeReqReg_6_bits_source2;
  reg  [2:0]         exeReqReg_6_bits_index;
  reg                exeReqReg_6_bits_ffo;
  reg                exeReqReg_7_valid;
  reg  [31:0]        exeReqReg_7_bits_source1;
  reg  [31:0]        exeReqReg_7_bits_source2;
  reg  [2:0]         exeReqReg_7_bits_index;
  reg                exeReqReg_7_bits_ffo;
  reg                exeReqReg_8_valid;
  reg  [31:0]        exeReqReg_8_bits_source1;
  reg  [31:0]        exeReqReg_8_bits_source2;
  reg  [2:0]         exeReqReg_8_bits_index;
  reg                exeReqReg_8_bits_ffo;
  reg                exeReqReg_9_valid;
  reg  [31:0]        exeReqReg_9_bits_source1;
  reg  [31:0]        exeReqReg_9_bits_source2;
  reg  [2:0]         exeReqReg_9_bits_index;
  reg                exeReqReg_9_bits_ffo;
  reg                exeReqReg_10_valid;
  reg  [31:0]        exeReqReg_10_bits_source1;
  reg  [31:0]        exeReqReg_10_bits_source2;
  reg  [2:0]         exeReqReg_10_bits_index;
  reg                exeReqReg_10_bits_ffo;
  reg                exeReqReg_11_valid;
  reg  [31:0]        exeReqReg_11_bits_source1;
  reg  [31:0]        exeReqReg_11_bits_source2;
  reg  [2:0]         exeReqReg_11_bits_index;
  reg                exeReqReg_11_bits_ffo;
  reg                exeReqReg_12_valid;
  reg  [31:0]        exeReqReg_12_bits_source1;
  reg  [31:0]        exeReqReg_12_bits_source2;
  reg  [2:0]         exeReqReg_12_bits_index;
  reg                exeReqReg_12_bits_ffo;
  reg                exeReqReg_13_valid;
  reg  [31:0]        exeReqReg_13_bits_source1;
  reg  [31:0]        exeReqReg_13_bits_source2;
  reg  [2:0]         exeReqReg_13_bits_index;
  reg                exeReqReg_13_bits_ffo;
  reg                exeReqReg_14_valid;
  reg  [31:0]        exeReqReg_14_bits_source1;
  reg  [31:0]        exeReqReg_14_bits_source2;
  reg  [2:0]         exeReqReg_14_bits_index;
  reg                exeReqReg_14_bits_ffo;
  reg                exeReqReg_15_valid;
  reg  [31:0]        exeReqReg_15_bits_source1;
  reg  [31:0]        exeReqReg_15_bits_source2;
  reg  [2:0]         exeReqReg_15_bits_index;
  reg                exeReqReg_15_bits_ffo;
  reg                exeReqReg_16_valid;
  reg  [31:0]        exeReqReg_16_bits_source1;
  reg  [31:0]        exeReqReg_16_bits_source2;
  reg  [2:0]         exeReqReg_16_bits_index;
  reg                exeReqReg_16_bits_ffo;
  reg                exeReqReg_17_valid;
  reg  [31:0]        exeReqReg_17_bits_source1;
  reg  [31:0]        exeReqReg_17_bits_source2;
  reg  [2:0]         exeReqReg_17_bits_index;
  reg                exeReqReg_17_bits_ffo;
  reg                exeReqReg_18_valid;
  reg  [31:0]        exeReqReg_18_bits_source1;
  reg  [31:0]        exeReqReg_18_bits_source2;
  reg  [2:0]         exeReqReg_18_bits_index;
  reg                exeReqReg_18_bits_ffo;
  reg                exeReqReg_19_valid;
  reg  [31:0]        exeReqReg_19_bits_source1;
  reg  [31:0]        exeReqReg_19_bits_source2;
  reg  [2:0]         exeReqReg_19_bits_index;
  reg                exeReqReg_19_bits_ffo;
  reg                exeReqReg_20_valid;
  reg  [31:0]        exeReqReg_20_bits_source1;
  reg  [31:0]        exeReqReg_20_bits_source2;
  reg  [2:0]         exeReqReg_20_bits_index;
  reg                exeReqReg_20_bits_ffo;
  reg                exeReqReg_21_valid;
  reg  [31:0]        exeReqReg_21_bits_source1;
  reg  [31:0]        exeReqReg_21_bits_source2;
  reg  [2:0]         exeReqReg_21_bits_index;
  reg                exeReqReg_21_bits_ffo;
  reg                exeReqReg_22_valid;
  reg  [31:0]        exeReqReg_22_bits_source1;
  reg  [31:0]        exeReqReg_22_bits_source2;
  reg  [2:0]         exeReqReg_22_bits_index;
  reg                exeReqReg_22_bits_ffo;
  reg                exeReqReg_23_valid;
  reg  [31:0]        exeReqReg_23_bits_source1;
  reg  [31:0]        exeReqReg_23_bits_source2;
  reg  [2:0]         exeReqReg_23_bits_index;
  reg                exeReqReg_23_bits_ffo;
  reg                exeReqReg_24_valid;
  reg  [31:0]        exeReqReg_24_bits_source1;
  reg  [31:0]        exeReqReg_24_bits_source2;
  reg  [2:0]         exeReqReg_24_bits_index;
  reg                exeReqReg_24_bits_ffo;
  reg                exeReqReg_25_valid;
  reg  [31:0]        exeReqReg_25_bits_source1;
  reg  [31:0]        exeReqReg_25_bits_source2;
  reg  [2:0]         exeReqReg_25_bits_index;
  reg                exeReqReg_25_bits_ffo;
  reg                exeReqReg_26_valid;
  reg  [31:0]        exeReqReg_26_bits_source1;
  reg  [31:0]        exeReqReg_26_bits_source2;
  reg  [2:0]         exeReqReg_26_bits_index;
  reg                exeReqReg_26_bits_ffo;
  reg                exeReqReg_27_valid;
  reg  [31:0]        exeReqReg_27_bits_source1;
  reg  [31:0]        exeReqReg_27_bits_source2;
  reg  [2:0]         exeReqReg_27_bits_index;
  reg                exeReqReg_27_bits_ffo;
  reg                exeReqReg_28_valid;
  reg  [31:0]        exeReqReg_28_bits_source1;
  reg  [31:0]        exeReqReg_28_bits_source2;
  reg  [2:0]         exeReqReg_28_bits_index;
  reg                exeReqReg_28_bits_ffo;
  reg                exeReqReg_29_valid;
  reg  [31:0]        exeReqReg_29_bits_source1;
  reg  [31:0]        exeReqReg_29_bits_source2;
  reg  [2:0]         exeReqReg_29_bits_index;
  reg                exeReqReg_29_bits_ffo;
  reg                exeReqReg_30_valid;
  reg  [31:0]        exeReqReg_30_bits_source1;
  reg  [31:0]        exeReqReg_30_bits_source2;
  reg  [2:0]         exeReqReg_30_bits_index;
  reg                exeReqReg_30_bits_ffo;
  reg                exeReqReg_31_valid;
  reg  [31:0]        exeReqReg_31_bits_source1;
  reg  [31:0]        exeReqReg_31_bits_source2;
  reg  [2:0]         exeReqReg_31_bits_index;
  reg                exeReqReg_31_bits_ffo;
  reg  [4:0]         requestCounter;
  wire [5:0]         _GEN_63 = {1'h0, requestCounter};
  wire               counterValid = _GEN_63 <= lastGroupForInstruction;
  wire               lastGroup = _GEN_63 == lastGroupForInstruction | ~orderReduce & unitType[2] | mv;
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_lo_lo = {slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi, slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_lo_hi = {slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi, slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_lo_lo = {slideAddressGen_slideMaskInput_lo_lo_lo_hi, slideAddressGen_slideMaskInput_lo_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_hi_lo = {slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi, slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_hi_hi = {slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi, slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_lo_hi = {slideAddressGen_slideMaskInput_lo_lo_hi_hi, slideAddressGen_slideMaskInput_lo_lo_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_lo_lo = {slideAddressGen_slideMaskInput_lo_lo_hi, slideAddressGen_slideMaskInput_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_lo_lo = {slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi, slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_lo_hi = {slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi, slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_hi_lo = {slideAddressGen_slideMaskInput_lo_hi_lo_hi, slideAddressGen_slideMaskInput_lo_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_hi_lo = {slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi, slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_hi_hi = {slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi, slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_hi_hi = {slideAddressGen_slideMaskInput_lo_hi_hi_hi, slideAddressGen_slideMaskInput_lo_hi_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_lo_hi = {slideAddressGen_slideMaskInput_lo_hi_hi, slideAddressGen_slideMaskInput_lo_hi_lo};
  wire [1023:0]      slideAddressGen_slideMaskInput_lo = {slideAddressGen_slideMaskInput_lo_hi, slideAddressGen_slideMaskInput_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_lo_lo = {slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi, slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_lo_hi = {slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi, slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_lo_lo = {slideAddressGen_slideMaskInput_hi_lo_lo_hi, slideAddressGen_slideMaskInput_hi_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_hi_lo = {slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi, slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_hi_hi = {slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi, slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_lo_hi = {slideAddressGen_slideMaskInput_hi_lo_hi_hi, slideAddressGen_slideMaskInput_hi_lo_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_hi_lo = {slideAddressGen_slideMaskInput_hi_lo_hi, slideAddressGen_slideMaskInput_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_lo_lo = {slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi, slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_lo_hi = {slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi, slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_hi_lo = {slideAddressGen_slideMaskInput_hi_hi_lo_hi, slideAddressGen_slideMaskInput_hi_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_hi_lo = {slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi, slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_hi_hi = {slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi, slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_hi_hi = {slideAddressGen_slideMaskInput_hi_hi_hi_hi, slideAddressGen_slideMaskInput_hi_hi_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_hi_hi = {slideAddressGen_slideMaskInput_hi_hi_hi, slideAddressGen_slideMaskInput_hi_hi_lo};
  wire [1023:0]      slideAddressGen_slideMaskInput_hi = {slideAddressGen_slideMaskInput_hi_hi, slideAddressGen_slideMaskInput_hi_lo};
  wire [63:0][31:0]  _GEN_64 =
    {{slideAddressGen_slideMaskInput_hi[1023:992]},
     {slideAddressGen_slideMaskInput_hi[991:960]},
     {slideAddressGen_slideMaskInput_hi[959:928]},
     {slideAddressGen_slideMaskInput_hi[927:896]},
     {slideAddressGen_slideMaskInput_hi[895:864]},
     {slideAddressGen_slideMaskInput_hi[863:832]},
     {slideAddressGen_slideMaskInput_hi[831:800]},
     {slideAddressGen_slideMaskInput_hi[799:768]},
     {slideAddressGen_slideMaskInput_hi[767:736]},
     {slideAddressGen_slideMaskInput_hi[735:704]},
     {slideAddressGen_slideMaskInput_hi[703:672]},
     {slideAddressGen_slideMaskInput_hi[671:640]},
     {slideAddressGen_slideMaskInput_hi[639:608]},
     {slideAddressGen_slideMaskInput_hi[607:576]},
     {slideAddressGen_slideMaskInput_hi[575:544]},
     {slideAddressGen_slideMaskInput_hi[543:512]},
     {slideAddressGen_slideMaskInput_hi[511:480]},
     {slideAddressGen_slideMaskInput_hi[479:448]},
     {slideAddressGen_slideMaskInput_hi[447:416]},
     {slideAddressGen_slideMaskInput_hi[415:384]},
     {slideAddressGen_slideMaskInput_hi[383:352]},
     {slideAddressGen_slideMaskInput_hi[351:320]},
     {slideAddressGen_slideMaskInput_hi[319:288]},
     {slideAddressGen_slideMaskInput_hi[287:256]},
     {slideAddressGen_slideMaskInput_hi[255:224]},
     {slideAddressGen_slideMaskInput_hi[223:192]},
     {slideAddressGen_slideMaskInput_hi[191:160]},
     {slideAddressGen_slideMaskInput_hi[159:128]},
     {slideAddressGen_slideMaskInput_hi[127:96]},
     {slideAddressGen_slideMaskInput_hi[95:64]},
     {slideAddressGen_slideMaskInput_hi[63:32]},
     {slideAddressGen_slideMaskInput_hi[31:0]},
     {slideAddressGen_slideMaskInput_lo[1023:992]},
     {slideAddressGen_slideMaskInput_lo[991:960]},
     {slideAddressGen_slideMaskInput_lo[959:928]},
     {slideAddressGen_slideMaskInput_lo[927:896]},
     {slideAddressGen_slideMaskInput_lo[895:864]},
     {slideAddressGen_slideMaskInput_lo[863:832]},
     {slideAddressGen_slideMaskInput_lo[831:800]},
     {slideAddressGen_slideMaskInput_lo[799:768]},
     {slideAddressGen_slideMaskInput_lo[767:736]},
     {slideAddressGen_slideMaskInput_lo[735:704]},
     {slideAddressGen_slideMaskInput_lo[703:672]},
     {slideAddressGen_slideMaskInput_lo[671:640]},
     {slideAddressGen_slideMaskInput_lo[639:608]},
     {slideAddressGen_slideMaskInput_lo[607:576]},
     {slideAddressGen_slideMaskInput_lo[575:544]},
     {slideAddressGen_slideMaskInput_lo[543:512]},
     {slideAddressGen_slideMaskInput_lo[511:480]},
     {slideAddressGen_slideMaskInput_lo[479:448]},
     {slideAddressGen_slideMaskInput_lo[447:416]},
     {slideAddressGen_slideMaskInput_lo[415:384]},
     {slideAddressGen_slideMaskInput_lo[383:352]},
     {slideAddressGen_slideMaskInput_lo[351:320]},
     {slideAddressGen_slideMaskInput_lo[319:288]},
     {slideAddressGen_slideMaskInput_lo[287:256]},
     {slideAddressGen_slideMaskInput_lo[255:224]},
     {slideAddressGen_slideMaskInput_lo[223:192]},
     {slideAddressGen_slideMaskInput_lo[191:160]},
     {slideAddressGen_slideMaskInput_lo[159:128]},
     {slideAddressGen_slideMaskInput_lo[127:96]},
     {slideAddressGen_slideMaskInput_lo[95:64]},
     {slideAddressGen_slideMaskInput_lo[63:32]},
     {slideAddressGen_slideMaskInput_lo[31:0]}};
  wire               lastExecuteGroupDeq;
  wire               viotaCounterAdd;
  wire               groupCounterAdd = noSource ? viotaCounterAdd : lastExecuteGroupDeq;
  wire [31:0]        groupDataNeed = lastGroup ? lastGroupDataNeed : 32'hFFFFFFFF;
  reg  [1:0]         executeIndex;
  reg  [31:0]        readIssueStageState_groupReadState;
  reg  [31:0]        readIssueStageState_needRead;
  wire [31:0]        readWaitQueue_enq_bits_needRead = readIssueStageState_needRead;
  reg  [31:0]        readIssueStageState_elementValid;
  wire [31:0]        readWaitQueue_enq_bits_sourceValid = readIssueStageState_elementValid;
  reg  [31:0]        readIssueStageState_replaceVs1;
  wire [31:0]        readWaitQueue_enq_bits_replaceVs1 = readIssueStageState_replaceVs1;
  reg  [31:0]        readIssueStageState_readOffset;
  reg  [4:0]         readIssueStageState_accessLane_0;
  reg  [4:0]         readIssueStageState_accessLane_1;
  wire [4:0]         selectExecuteReq_1_bits_readLane = readIssueStageState_accessLane_1;
  reg  [4:0]         readIssueStageState_accessLane_2;
  wire [4:0]         selectExecuteReq_2_bits_readLane = readIssueStageState_accessLane_2;
  reg  [4:0]         readIssueStageState_accessLane_3;
  wire [4:0]         selectExecuteReq_3_bits_readLane = readIssueStageState_accessLane_3;
  reg  [4:0]         readIssueStageState_accessLane_4;
  wire [4:0]         selectExecuteReq_4_bits_readLane = readIssueStageState_accessLane_4;
  reg  [4:0]         readIssueStageState_accessLane_5;
  wire [4:0]         selectExecuteReq_5_bits_readLane = readIssueStageState_accessLane_5;
  reg  [4:0]         readIssueStageState_accessLane_6;
  wire [4:0]         selectExecuteReq_6_bits_readLane = readIssueStageState_accessLane_6;
  reg  [4:0]         readIssueStageState_accessLane_7;
  wire [4:0]         selectExecuteReq_7_bits_readLane = readIssueStageState_accessLane_7;
  reg  [4:0]         readIssueStageState_accessLane_8;
  wire [4:0]         selectExecuteReq_8_bits_readLane = readIssueStageState_accessLane_8;
  reg  [4:0]         readIssueStageState_accessLane_9;
  wire [4:0]         selectExecuteReq_9_bits_readLane = readIssueStageState_accessLane_9;
  reg  [4:0]         readIssueStageState_accessLane_10;
  wire [4:0]         selectExecuteReq_10_bits_readLane = readIssueStageState_accessLane_10;
  reg  [4:0]         readIssueStageState_accessLane_11;
  wire [4:0]         selectExecuteReq_11_bits_readLane = readIssueStageState_accessLane_11;
  reg  [4:0]         readIssueStageState_accessLane_12;
  wire [4:0]         selectExecuteReq_12_bits_readLane = readIssueStageState_accessLane_12;
  reg  [4:0]         readIssueStageState_accessLane_13;
  wire [4:0]         selectExecuteReq_13_bits_readLane = readIssueStageState_accessLane_13;
  reg  [4:0]         readIssueStageState_accessLane_14;
  wire [4:0]         selectExecuteReq_14_bits_readLane = readIssueStageState_accessLane_14;
  reg  [4:0]         readIssueStageState_accessLane_15;
  wire [4:0]         selectExecuteReq_15_bits_readLane = readIssueStageState_accessLane_15;
  reg  [4:0]         readIssueStageState_accessLane_16;
  wire [4:0]         selectExecuteReq_16_bits_readLane = readIssueStageState_accessLane_16;
  reg  [4:0]         readIssueStageState_accessLane_17;
  wire [4:0]         selectExecuteReq_17_bits_readLane = readIssueStageState_accessLane_17;
  reg  [4:0]         readIssueStageState_accessLane_18;
  wire [4:0]         selectExecuteReq_18_bits_readLane = readIssueStageState_accessLane_18;
  reg  [4:0]         readIssueStageState_accessLane_19;
  wire [4:0]         selectExecuteReq_19_bits_readLane = readIssueStageState_accessLane_19;
  reg  [4:0]         readIssueStageState_accessLane_20;
  wire [4:0]         selectExecuteReq_20_bits_readLane = readIssueStageState_accessLane_20;
  reg  [4:0]         readIssueStageState_accessLane_21;
  wire [4:0]         selectExecuteReq_21_bits_readLane = readIssueStageState_accessLane_21;
  reg  [4:0]         readIssueStageState_accessLane_22;
  wire [4:0]         selectExecuteReq_22_bits_readLane = readIssueStageState_accessLane_22;
  reg  [4:0]         readIssueStageState_accessLane_23;
  wire [4:0]         selectExecuteReq_23_bits_readLane = readIssueStageState_accessLane_23;
  reg  [4:0]         readIssueStageState_accessLane_24;
  wire [4:0]         selectExecuteReq_24_bits_readLane = readIssueStageState_accessLane_24;
  reg  [4:0]         readIssueStageState_accessLane_25;
  wire [4:0]         selectExecuteReq_25_bits_readLane = readIssueStageState_accessLane_25;
  reg  [4:0]         readIssueStageState_accessLane_26;
  wire [4:0]         selectExecuteReq_26_bits_readLane = readIssueStageState_accessLane_26;
  reg  [4:0]         readIssueStageState_accessLane_27;
  wire [4:0]         selectExecuteReq_27_bits_readLane = readIssueStageState_accessLane_27;
  reg  [4:0]         readIssueStageState_accessLane_28;
  wire [4:0]         selectExecuteReq_28_bits_readLane = readIssueStageState_accessLane_28;
  reg  [4:0]         readIssueStageState_accessLane_29;
  wire [4:0]         selectExecuteReq_29_bits_readLane = readIssueStageState_accessLane_29;
  reg  [4:0]         readIssueStageState_accessLane_30;
  wire [4:0]         selectExecuteReq_30_bits_readLane = readIssueStageState_accessLane_30;
  reg  [4:0]         readIssueStageState_accessLane_31;
  wire [4:0]         selectExecuteReq_31_bits_readLane = readIssueStageState_accessLane_31;
  reg  [2:0]         readIssueStageState_vsGrowth_0;
  reg  [2:0]         readIssueStageState_vsGrowth_1;
  reg  [2:0]         readIssueStageState_vsGrowth_2;
  reg  [2:0]         readIssueStageState_vsGrowth_3;
  reg  [2:0]         readIssueStageState_vsGrowth_4;
  reg  [2:0]         readIssueStageState_vsGrowth_5;
  reg  [2:0]         readIssueStageState_vsGrowth_6;
  reg  [2:0]         readIssueStageState_vsGrowth_7;
  reg  [2:0]         readIssueStageState_vsGrowth_8;
  reg  [2:0]         readIssueStageState_vsGrowth_9;
  reg  [2:0]         readIssueStageState_vsGrowth_10;
  reg  [2:0]         readIssueStageState_vsGrowth_11;
  reg  [2:0]         readIssueStageState_vsGrowth_12;
  reg  [2:0]         readIssueStageState_vsGrowth_13;
  reg  [2:0]         readIssueStageState_vsGrowth_14;
  reg  [2:0]         readIssueStageState_vsGrowth_15;
  reg  [2:0]         readIssueStageState_vsGrowth_16;
  reg  [2:0]         readIssueStageState_vsGrowth_17;
  reg  [2:0]         readIssueStageState_vsGrowth_18;
  reg  [2:0]         readIssueStageState_vsGrowth_19;
  reg  [2:0]         readIssueStageState_vsGrowth_20;
  reg  [2:0]         readIssueStageState_vsGrowth_21;
  reg  [2:0]         readIssueStageState_vsGrowth_22;
  reg  [2:0]         readIssueStageState_vsGrowth_23;
  reg  [2:0]         readIssueStageState_vsGrowth_24;
  reg  [2:0]         readIssueStageState_vsGrowth_25;
  reg  [2:0]         readIssueStageState_vsGrowth_26;
  reg  [2:0]         readIssueStageState_vsGrowth_27;
  reg  [2:0]         readIssueStageState_vsGrowth_28;
  reg  [2:0]         readIssueStageState_vsGrowth_29;
  reg  [2:0]         readIssueStageState_vsGrowth_30;
  reg  [2:0]         readIssueStageState_vsGrowth_31;
  reg  [6:0]         readIssueStageState_executeGroup;
  wire [6:0]         readWaitQueue_enq_bits_executeGroup = readIssueStageState_executeGroup;
  reg  [63:0]        readIssueStageState_readDataOffset;
  reg                readIssueStageState_last;
  wire               readWaitQueue_enq_bits_last = readIssueStageState_last;
  reg                readIssueStageValid;
  wire [5:0]         accessCountQueue_enq_bits_0 = accessCountEnq_0;
  wire [5:0]         accessCountQueue_enq_bits_1 = accessCountEnq_1;
  wire [5:0]         accessCountQueue_enq_bits_2 = accessCountEnq_2;
  wire [5:0]         accessCountQueue_enq_bits_3 = accessCountEnq_3;
  wire [5:0]         accessCountQueue_enq_bits_4 = accessCountEnq_4;
  wire [5:0]         accessCountQueue_enq_bits_5 = accessCountEnq_5;
  wire [5:0]         accessCountQueue_enq_bits_6 = accessCountEnq_6;
  wire [5:0]         accessCountQueue_enq_bits_7 = accessCountEnq_7;
  wire [5:0]         accessCountQueue_enq_bits_8 = accessCountEnq_8;
  wire [5:0]         accessCountQueue_enq_bits_9 = accessCountEnq_9;
  wire [5:0]         accessCountQueue_enq_bits_10 = accessCountEnq_10;
  wire [5:0]         accessCountQueue_enq_bits_11 = accessCountEnq_11;
  wire [5:0]         accessCountQueue_enq_bits_12 = accessCountEnq_12;
  wire [5:0]         accessCountQueue_enq_bits_13 = accessCountEnq_13;
  wire [5:0]         accessCountQueue_enq_bits_14 = accessCountEnq_14;
  wire [5:0]         accessCountQueue_enq_bits_15 = accessCountEnq_15;
  wire [5:0]         accessCountQueue_enq_bits_16 = accessCountEnq_16;
  wire [5:0]         accessCountQueue_enq_bits_17 = accessCountEnq_17;
  wire [5:0]         accessCountQueue_enq_bits_18 = accessCountEnq_18;
  wire [5:0]         accessCountQueue_enq_bits_19 = accessCountEnq_19;
  wire [5:0]         accessCountQueue_enq_bits_20 = accessCountEnq_20;
  wire [5:0]         accessCountQueue_enq_bits_21 = accessCountEnq_21;
  wire [5:0]         accessCountQueue_enq_bits_22 = accessCountEnq_22;
  wire [5:0]         accessCountQueue_enq_bits_23 = accessCountEnq_23;
  wire [5:0]         accessCountQueue_enq_bits_24 = accessCountEnq_24;
  wire [5:0]         accessCountQueue_enq_bits_25 = accessCountEnq_25;
  wire [5:0]         accessCountQueue_enq_bits_26 = accessCountEnq_26;
  wire [5:0]         accessCountQueue_enq_bits_27 = accessCountEnq_27;
  wire [5:0]         accessCountQueue_enq_bits_28 = accessCountEnq_28;
  wire [5:0]         accessCountQueue_enq_bits_29 = accessCountEnq_29;
  wire [5:0]         accessCountQueue_enq_bits_30 = accessCountEnq_30;
  wire [5:0]         accessCountQueue_enq_bits_31 = accessCountEnq_31;
  wire               readIssueStageEnq;
  wire               accessCountQueue_deq_valid;
  assign accessCountQueue_deq_valid = ~_accessCountQueue_fifo_empty;
  wire [5:0]         accessCountQueue_dataOut_0;
  wire [5:0]         accessCountQueue_dataOut_1;
  wire [5:0]         accessCountQueue_dataOut_2;
  wire [5:0]         accessCountQueue_dataOut_3;
  wire [5:0]         accessCountQueue_dataOut_4;
  wire [5:0]         accessCountQueue_dataOut_5;
  wire [5:0]         accessCountQueue_dataOut_6;
  wire [5:0]         accessCountQueue_dataOut_7;
  wire [5:0]         accessCountQueue_dataOut_8;
  wire [5:0]         accessCountQueue_dataOut_9;
  wire [5:0]         accessCountQueue_dataOut_10;
  wire [5:0]         accessCountQueue_dataOut_11;
  wire [5:0]         accessCountQueue_dataOut_12;
  wire [5:0]         accessCountQueue_dataOut_13;
  wire [5:0]         accessCountQueue_dataOut_14;
  wire [5:0]         accessCountQueue_dataOut_15;
  wire [5:0]         accessCountQueue_dataOut_16;
  wire [5:0]         accessCountQueue_dataOut_17;
  wire [5:0]         accessCountQueue_dataOut_18;
  wire [5:0]         accessCountQueue_dataOut_19;
  wire [5:0]         accessCountQueue_dataOut_20;
  wire [5:0]         accessCountQueue_dataOut_21;
  wire [5:0]         accessCountQueue_dataOut_22;
  wire [5:0]         accessCountQueue_dataOut_23;
  wire [5:0]         accessCountQueue_dataOut_24;
  wire [5:0]         accessCountQueue_dataOut_25;
  wire [5:0]         accessCountQueue_dataOut_26;
  wire [5:0]         accessCountQueue_dataOut_27;
  wire [5:0]         accessCountQueue_dataOut_28;
  wire [5:0]         accessCountQueue_dataOut_29;
  wire [5:0]         accessCountQueue_dataOut_30;
  wire [5:0]         accessCountQueue_dataOut_31;
  wire [11:0]        accessCountQueue_dataIn_lo_lo_lo_lo = {accessCountQueue_enq_bits_1, accessCountQueue_enq_bits_0};
  wire [11:0]        accessCountQueue_dataIn_lo_lo_lo_hi = {accessCountQueue_enq_bits_3, accessCountQueue_enq_bits_2};
  wire [23:0]        accessCountQueue_dataIn_lo_lo_lo = {accessCountQueue_dataIn_lo_lo_lo_hi, accessCountQueue_dataIn_lo_lo_lo_lo};
  wire [11:0]        accessCountQueue_dataIn_lo_lo_hi_lo = {accessCountQueue_enq_bits_5, accessCountQueue_enq_bits_4};
  wire [11:0]        accessCountQueue_dataIn_lo_lo_hi_hi = {accessCountQueue_enq_bits_7, accessCountQueue_enq_bits_6};
  wire [23:0]        accessCountQueue_dataIn_lo_lo_hi = {accessCountQueue_dataIn_lo_lo_hi_hi, accessCountQueue_dataIn_lo_lo_hi_lo};
  wire [47:0]        accessCountQueue_dataIn_lo_lo = {accessCountQueue_dataIn_lo_lo_hi, accessCountQueue_dataIn_lo_lo_lo};
  wire [11:0]        accessCountQueue_dataIn_lo_hi_lo_lo = {accessCountQueue_enq_bits_9, accessCountQueue_enq_bits_8};
  wire [11:0]        accessCountQueue_dataIn_lo_hi_lo_hi = {accessCountQueue_enq_bits_11, accessCountQueue_enq_bits_10};
  wire [23:0]        accessCountQueue_dataIn_lo_hi_lo = {accessCountQueue_dataIn_lo_hi_lo_hi, accessCountQueue_dataIn_lo_hi_lo_lo};
  wire [11:0]        accessCountQueue_dataIn_lo_hi_hi_lo = {accessCountQueue_enq_bits_13, accessCountQueue_enq_bits_12};
  wire [11:0]        accessCountQueue_dataIn_lo_hi_hi_hi = {accessCountQueue_enq_bits_15, accessCountQueue_enq_bits_14};
  wire [23:0]        accessCountQueue_dataIn_lo_hi_hi = {accessCountQueue_dataIn_lo_hi_hi_hi, accessCountQueue_dataIn_lo_hi_hi_lo};
  wire [47:0]        accessCountQueue_dataIn_lo_hi = {accessCountQueue_dataIn_lo_hi_hi, accessCountQueue_dataIn_lo_hi_lo};
  wire [95:0]        accessCountQueue_dataIn_lo = {accessCountQueue_dataIn_lo_hi, accessCountQueue_dataIn_lo_lo};
  wire [11:0]        accessCountQueue_dataIn_hi_lo_lo_lo = {accessCountQueue_enq_bits_17, accessCountQueue_enq_bits_16};
  wire [11:0]        accessCountQueue_dataIn_hi_lo_lo_hi = {accessCountQueue_enq_bits_19, accessCountQueue_enq_bits_18};
  wire [23:0]        accessCountQueue_dataIn_hi_lo_lo = {accessCountQueue_dataIn_hi_lo_lo_hi, accessCountQueue_dataIn_hi_lo_lo_lo};
  wire [11:0]        accessCountQueue_dataIn_hi_lo_hi_lo = {accessCountQueue_enq_bits_21, accessCountQueue_enq_bits_20};
  wire [11:0]        accessCountQueue_dataIn_hi_lo_hi_hi = {accessCountQueue_enq_bits_23, accessCountQueue_enq_bits_22};
  wire [23:0]        accessCountQueue_dataIn_hi_lo_hi = {accessCountQueue_dataIn_hi_lo_hi_hi, accessCountQueue_dataIn_hi_lo_hi_lo};
  wire [47:0]        accessCountQueue_dataIn_hi_lo = {accessCountQueue_dataIn_hi_lo_hi, accessCountQueue_dataIn_hi_lo_lo};
  wire [11:0]        accessCountQueue_dataIn_hi_hi_lo_lo = {accessCountQueue_enq_bits_25, accessCountQueue_enq_bits_24};
  wire [11:0]        accessCountQueue_dataIn_hi_hi_lo_hi = {accessCountQueue_enq_bits_27, accessCountQueue_enq_bits_26};
  wire [23:0]        accessCountQueue_dataIn_hi_hi_lo = {accessCountQueue_dataIn_hi_hi_lo_hi, accessCountQueue_dataIn_hi_hi_lo_lo};
  wire [11:0]        accessCountQueue_dataIn_hi_hi_hi_lo = {accessCountQueue_enq_bits_29, accessCountQueue_enq_bits_28};
  wire [11:0]        accessCountQueue_dataIn_hi_hi_hi_hi = {accessCountQueue_enq_bits_31, accessCountQueue_enq_bits_30};
  wire [23:0]        accessCountQueue_dataIn_hi_hi_hi = {accessCountQueue_dataIn_hi_hi_hi_hi, accessCountQueue_dataIn_hi_hi_hi_lo};
  wire [47:0]        accessCountQueue_dataIn_hi_hi = {accessCountQueue_dataIn_hi_hi_hi, accessCountQueue_dataIn_hi_hi_lo};
  wire [95:0]        accessCountQueue_dataIn_hi = {accessCountQueue_dataIn_hi_hi, accessCountQueue_dataIn_hi_lo};
  wire [191:0]       accessCountQueue_dataIn = {accessCountQueue_dataIn_hi, accessCountQueue_dataIn_lo};
  assign accessCountQueue_dataOut_0 = _accessCountQueue_fifo_data_out[5:0];
  assign accessCountQueue_dataOut_1 = _accessCountQueue_fifo_data_out[11:6];
  assign accessCountQueue_dataOut_2 = _accessCountQueue_fifo_data_out[17:12];
  assign accessCountQueue_dataOut_3 = _accessCountQueue_fifo_data_out[23:18];
  assign accessCountQueue_dataOut_4 = _accessCountQueue_fifo_data_out[29:24];
  assign accessCountQueue_dataOut_5 = _accessCountQueue_fifo_data_out[35:30];
  assign accessCountQueue_dataOut_6 = _accessCountQueue_fifo_data_out[41:36];
  assign accessCountQueue_dataOut_7 = _accessCountQueue_fifo_data_out[47:42];
  assign accessCountQueue_dataOut_8 = _accessCountQueue_fifo_data_out[53:48];
  assign accessCountQueue_dataOut_9 = _accessCountQueue_fifo_data_out[59:54];
  assign accessCountQueue_dataOut_10 = _accessCountQueue_fifo_data_out[65:60];
  assign accessCountQueue_dataOut_11 = _accessCountQueue_fifo_data_out[71:66];
  assign accessCountQueue_dataOut_12 = _accessCountQueue_fifo_data_out[77:72];
  assign accessCountQueue_dataOut_13 = _accessCountQueue_fifo_data_out[83:78];
  assign accessCountQueue_dataOut_14 = _accessCountQueue_fifo_data_out[89:84];
  assign accessCountQueue_dataOut_15 = _accessCountQueue_fifo_data_out[95:90];
  assign accessCountQueue_dataOut_16 = _accessCountQueue_fifo_data_out[101:96];
  assign accessCountQueue_dataOut_17 = _accessCountQueue_fifo_data_out[107:102];
  assign accessCountQueue_dataOut_18 = _accessCountQueue_fifo_data_out[113:108];
  assign accessCountQueue_dataOut_19 = _accessCountQueue_fifo_data_out[119:114];
  assign accessCountQueue_dataOut_20 = _accessCountQueue_fifo_data_out[125:120];
  assign accessCountQueue_dataOut_21 = _accessCountQueue_fifo_data_out[131:126];
  assign accessCountQueue_dataOut_22 = _accessCountQueue_fifo_data_out[137:132];
  assign accessCountQueue_dataOut_23 = _accessCountQueue_fifo_data_out[143:138];
  assign accessCountQueue_dataOut_24 = _accessCountQueue_fifo_data_out[149:144];
  assign accessCountQueue_dataOut_25 = _accessCountQueue_fifo_data_out[155:150];
  assign accessCountQueue_dataOut_26 = _accessCountQueue_fifo_data_out[161:156];
  assign accessCountQueue_dataOut_27 = _accessCountQueue_fifo_data_out[167:162];
  assign accessCountQueue_dataOut_28 = _accessCountQueue_fifo_data_out[173:168];
  assign accessCountQueue_dataOut_29 = _accessCountQueue_fifo_data_out[179:174];
  assign accessCountQueue_dataOut_30 = _accessCountQueue_fifo_data_out[185:180];
  assign accessCountQueue_dataOut_31 = _accessCountQueue_fifo_data_out[191:186];
  wire [5:0]         accessCountQueue_deq_bits_0 = accessCountQueue_dataOut_0;
  wire [5:0]         accessCountQueue_deq_bits_1 = accessCountQueue_dataOut_1;
  wire [5:0]         accessCountQueue_deq_bits_2 = accessCountQueue_dataOut_2;
  wire [5:0]         accessCountQueue_deq_bits_3 = accessCountQueue_dataOut_3;
  wire [5:0]         accessCountQueue_deq_bits_4 = accessCountQueue_dataOut_4;
  wire [5:0]         accessCountQueue_deq_bits_5 = accessCountQueue_dataOut_5;
  wire [5:0]         accessCountQueue_deq_bits_6 = accessCountQueue_dataOut_6;
  wire [5:0]         accessCountQueue_deq_bits_7 = accessCountQueue_dataOut_7;
  wire [5:0]         accessCountQueue_deq_bits_8 = accessCountQueue_dataOut_8;
  wire [5:0]         accessCountQueue_deq_bits_9 = accessCountQueue_dataOut_9;
  wire [5:0]         accessCountQueue_deq_bits_10 = accessCountQueue_dataOut_10;
  wire [5:0]         accessCountQueue_deq_bits_11 = accessCountQueue_dataOut_11;
  wire [5:0]         accessCountQueue_deq_bits_12 = accessCountQueue_dataOut_12;
  wire [5:0]         accessCountQueue_deq_bits_13 = accessCountQueue_dataOut_13;
  wire [5:0]         accessCountQueue_deq_bits_14 = accessCountQueue_dataOut_14;
  wire [5:0]         accessCountQueue_deq_bits_15 = accessCountQueue_dataOut_15;
  wire [5:0]         accessCountQueue_deq_bits_16 = accessCountQueue_dataOut_16;
  wire [5:0]         accessCountQueue_deq_bits_17 = accessCountQueue_dataOut_17;
  wire [5:0]         accessCountQueue_deq_bits_18 = accessCountQueue_dataOut_18;
  wire [5:0]         accessCountQueue_deq_bits_19 = accessCountQueue_dataOut_19;
  wire [5:0]         accessCountQueue_deq_bits_20 = accessCountQueue_dataOut_20;
  wire [5:0]         accessCountQueue_deq_bits_21 = accessCountQueue_dataOut_21;
  wire [5:0]         accessCountQueue_deq_bits_22 = accessCountQueue_dataOut_22;
  wire [5:0]         accessCountQueue_deq_bits_23 = accessCountQueue_dataOut_23;
  wire [5:0]         accessCountQueue_deq_bits_24 = accessCountQueue_dataOut_24;
  wire [5:0]         accessCountQueue_deq_bits_25 = accessCountQueue_dataOut_25;
  wire [5:0]         accessCountQueue_deq_bits_26 = accessCountQueue_dataOut_26;
  wire [5:0]         accessCountQueue_deq_bits_27 = accessCountQueue_dataOut_27;
  wire [5:0]         accessCountQueue_deq_bits_28 = accessCountQueue_dataOut_28;
  wire [5:0]         accessCountQueue_deq_bits_29 = accessCountQueue_dataOut_29;
  wire [5:0]         accessCountQueue_deq_bits_30 = accessCountQueue_dataOut_30;
  wire [5:0]         accessCountQueue_deq_bits_31 = accessCountQueue_dataOut_31;
  wire               accessCountQueue_enq_ready = ~_accessCountQueue_fifo_full;
  wire               accessCountQueue_enq_valid;
  wire               accessCountQueue_deq_ready;
  wire [6:0]         _extendGroupCount_T_1 = {requestCounter, executeIndex};
  wire [6:0]         _executeGroup_T_8 = executeIndexGrowth[0] ? _extendGroupCount_T_1 : 7'h0;
  wire [5:0]         _GEN_65 = _executeGroup_T_8[5:0] | (executeIndexGrowth[1] ? {requestCounter, executeIndex[1]} : 6'h0);
  wire [6:0]         executeGroup = {_executeGroup_T_8[6], _GEN_65[5], _GEN_65[4:0] | (executeIndexGrowth[2] ? requestCounter : 5'h0)};
  wire               vlMisAlign;
  assign vlMisAlign = |(instReg_vl[4:0]);
  wire [6:0]         lastexecuteGroup = instReg_vl[11:5] - {6'h0, ~vlMisAlign};
  wire               isVlBoundary = executeGroup == lastexecuteGroup;
  wire               validExecuteGroup = executeGroup <= lastexecuteGroup;
  wire [31:0]        _maskSplit_vlBoundaryCorrection_T_55 = 32'h1 << instReg_vl[4:0];
  wire [31:0]        _vlBoundaryCorrection_T_5 = _maskSplit_vlBoundaryCorrection_T_55 | {_maskSplit_vlBoundaryCorrection_T_55[30:0], 1'h0};
  wire [31:0]        _vlBoundaryCorrection_T_8 = _vlBoundaryCorrection_T_5 | {_vlBoundaryCorrection_T_5[29:0], 2'h0};
  wire [31:0]        _vlBoundaryCorrection_T_11 = _vlBoundaryCorrection_T_8 | {_vlBoundaryCorrection_T_8[27:0], 4'h0};
  wire [31:0]        _vlBoundaryCorrection_T_14 = _vlBoundaryCorrection_T_11 | {_vlBoundaryCorrection_T_11[23:0], 8'h0};
  wire [31:0]        vlBoundaryCorrection = ~({32{vlMisAlign & isVlBoundary}} & (_vlBoundaryCorrection_T_14 | {_vlBoundaryCorrection_T_14[15:0], 16'h0})) & {32{validExecuteGroup}};
  wire [127:0]       selectReadStageMask_lo_lo_lo_lo = {selectReadStageMask_lo_lo_lo_lo_hi, selectReadStageMask_lo_lo_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_lo_lo_hi = {selectReadStageMask_lo_lo_lo_hi_hi, selectReadStageMask_lo_lo_lo_hi_lo};
  wire [255:0]       selectReadStageMask_lo_lo_lo = {selectReadStageMask_lo_lo_lo_hi, selectReadStageMask_lo_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_lo_hi_lo = {selectReadStageMask_lo_lo_hi_lo_hi, selectReadStageMask_lo_lo_hi_lo_lo};
  wire [127:0]       selectReadStageMask_lo_lo_hi_hi = {selectReadStageMask_lo_lo_hi_hi_hi, selectReadStageMask_lo_lo_hi_hi_lo};
  wire [255:0]       selectReadStageMask_lo_lo_hi = {selectReadStageMask_lo_lo_hi_hi, selectReadStageMask_lo_lo_hi_lo};
  wire [511:0]       selectReadStageMask_lo_lo = {selectReadStageMask_lo_lo_hi, selectReadStageMask_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_lo_lo = {selectReadStageMask_lo_hi_lo_lo_hi, selectReadStageMask_lo_hi_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_lo_hi = {selectReadStageMask_lo_hi_lo_hi_hi, selectReadStageMask_lo_hi_lo_hi_lo};
  wire [255:0]       selectReadStageMask_lo_hi_lo = {selectReadStageMask_lo_hi_lo_hi, selectReadStageMask_lo_hi_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_hi_lo = {selectReadStageMask_lo_hi_hi_lo_hi, selectReadStageMask_lo_hi_hi_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_hi_hi = {selectReadStageMask_lo_hi_hi_hi_hi, selectReadStageMask_lo_hi_hi_hi_lo};
  wire [255:0]       selectReadStageMask_lo_hi_hi = {selectReadStageMask_lo_hi_hi_hi, selectReadStageMask_lo_hi_hi_lo};
  wire [511:0]       selectReadStageMask_lo_hi = {selectReadStageMask_lo_hi_hi, selectReadStageMask_lo_hi_lo};
  wire [1023:0]      selectReadStageMask_lo = {selectReadStageMask_lo_hi, selectReadStageMask_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_lo_lo = {selectReadStageMask_hi_lo_lo_lo_hi, selectReadStageMask_hi_lo_lo_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_lo_hi = {selectReadStageMask_hi_lo_lo_hi_hi, selectReadStageMask_hi_lo_lo_hi_lo};
  wire [255:0]       selectReadStageMask_hi_lo_lo = {selectReadStageMask_hi_lo_lo_hi, selectReadStageMask_hi_lo_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_hi_lo = {selectReadStageMask_hi_lo_hi_lo_hi, selectReadStageMask_hi_lo_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_hi_hi = {selectReadStageMask_hi_lo_hi_hi_hi, selectReadStageMask_hi_lo_hi_hi_lo};
  wire [255:0]       selectReadStageMask_hi_lo_hi = {selectReadStageMask_hi_lo_hi_hi, selectReadStageMask_hi_lo_hi_lo};
  wire [511:0]       selectReadStageMask_hi_lo = {selectReadStageMask_hi_lo_hi, selectReadStageMask_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_lo_lo = {selectReadStageMask_hi_hi_lo_lo_hi, selectReadStageMask_hi_hi_lo_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_lo_hi = {selectReadStageMask_hi_hi_lo_hi_hi, selectReadStageMask_hi_hi_lo_hi_lo};
  wire [255:0]       selectReadStageMask_hi_hi_lo = {selectReadStageMask_hi_hi_lo_hi, selectReadStageMask_hi_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_hi_lo = {selectReadStageMask_hi_hi_hi_lo_hi, selectReadStageMask_hi_hi_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_hi_hi = {selectReadStageMask_hi_hi_hi_hi_hi, selectReadStageMask_hi_hi_hi_hi_lo};
  wire [255:0]       selectReadStageMask_hi_hi_hi = {selectReadStageMask_hi_hi_hi_hi, selectReadStageMask_hi_hi_hi_lo};
  wire [511:0]       selectReadStageMask_hi_hi = {selectReadStageMask_hi_hi_hi, selectReadStageMask_hi_hi_lo};
  wire [1023:0]      selectReadStageMask_hi = {selectReadStageMask_hi_hi, selectReadStageMask_hi_lo};
  wire [63:0][31:0]  _GEN_66 =
    {{selectReadStageMask_hi[1023:992]},
     {selectReadStageMask_hi[991:960]},
     {selectReadStageMask_hi[959:928]},
     {selectReadStageMask_hi[927:896]},
     {selectReadStageMask_hi[895:864]},
     {selectReadStageMask_hi[863:832]},
     {selectReadStageMask_hi[831:800]},
     {selectReadStageMask_hi[799:768]},
     {selectReadStageMask_hi[767:736]},
     {selectReadStageMask_hi[735:704]},
     {selectReadStageMask_hi[703:672]},
     {selectReadStageMask_hi[671:640]},
     {selectReadStageMask_hi[639:608]},
     {selectReadStageMask_hi[607:576]},
     {selectReadStageMask_hi[575:544]},
     {selectReadStageMask_hi[543:512]},
     {selectReadStageMask_hi[511:480]},
     {selectReadStageMask_hi[479:448]},
     {selectReadStageMask_hi[447:416]},
     {selectReadStageMask_hi[415:384]},
     {selectReadStageMask_hi[383:352]},
     {selectReadStageMask_hi[351:320]},
     {selectReadStageMask_hi[319:288]},
     {selectReadStageMask_hi[287:256]},
     {selectReadStageMask_hi[255:224]},
     {selectReadStageMask_hi[223:192]},
     {selectReadStageMask_hi[191:160]},
     {selectReadStageMask_hi[159:128]},
     {selectReadStageMask_hi[127:96]},
     {selectReadStageMask_hi[95:64]},
     {selectReadStageMask_hi[63:32]},
     {selectReadStageMask_hi[31:0]},
     {selectReadStageMask_lo[1023:992]},
     {selectReadStageMask_lo[991:960]},
     {selectReadStageMask_lo[959:928]},
     {selectReadStageMask_lo[927:896]},
     {selectReadStageMask_lo[895:864]},
     {selectReadStageMask_lo[863:832]},
     {selectReadStageMask_lo[831:800]},
     {selectReadStageMask_lo[799:768]},
     {selectReadStageMask_lo[767:736]},
     {selectReadStageMask_lo[735:704]},
     {selectReadStageMask_lo[703:672]},
     {selectReadStageMask_lo[671:640]},
     {selectReadStageMask_lo[639:608]},
     {selectReadStageMask_lo[607:576]},
     {selectReadStageMask_lo[575:544]},
     {selectReadStageMask_lo[543:512]},
     {selectReadStageMask_lo[511:480]},
     {selectReadStageMask_lo[479:448]},
     {selectReadStageMask_lo[447:416]},
     {selectReadStageMask_lo[415:384]},
     {selectReadStageMask_lo[383:352]},
     {selectReadStageMask_lo[351:320]},
     {selectReadStageMask_lo[319:288]},
     {selectReadStageMask_lo[287:256]},
     {selectReadStageMask_lo[255:224]},
     {selectReadStageMask_lo[223:192]},
     {selectReadStageMask_lo[191:160]},
     {selectReadStageMask_lo[159:128]},
     {selectReadStageMask_lo[127:96]},
     {selectReadStageMask_lo[95:64]},
     {selectReadStageMask_lo[63:32]},
     {selectReadStageMask_lo[31:0]}};
  wire [31:0]        readMaskCorrection = (instReg_maskType ? _GEN_66[executeGroup[5:0]] : 32'hFFFFFFFF) & vlBoundaryCorrection;
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_lo = {maskSplit_maskSelect_lo_lo_lo_lo_hi, maskSplit_maskSelect_lo_lo_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_hi = {maskSplit_maskSelect_lo_lo_lo_hi_hi, maskSplit_maskSelect_lo_lo_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_lo_lo = {maskSplit_maskSelect_lo_lo_lo_hi, maskSplit_maskSelect_lo_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_lo = {maskSplit_maskSelect_lo_lo_hi_lo_hi, maskSplit_maskSelect_lo_lo_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_hi = {maskSplit_maskSelect_lo_lo_hi_hi_hi, maskSplit_maskSelect_lo_lo_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_lo_hi = {maskSplit_maskSelect_lo_lo_hi_hi, maskSplit_maskSelect_lo_lo_hi_lo};
  wire [511:0]       maskSplit_maskSelect_lo_lo = {maskSplit_maskSelect_lo_lo_hi, maskSplit_maskSelect_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_lo = {maskSplit_maskSelect_lo_hi_lo_lo_hi, maskSplit_maskSelect_lo_hi_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_hi = {maskSplit_maskSelect_lo_hi_lo_hi_hi, maskSplit_maskSelect_lo_hi_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_hi_lo = {maskSplit_maskSelect_lo_hi_lo_hi, maskSplit_maskSelect_lo_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_lo = {maskSplit_maskSelect_lo_hi_hi_lo_hi, maskSplit_maskSelect_lo_hi_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_hi = {maskSplit_maskSelect_lo_hi_hi_hi_hi, maskSplit_maskSelect_lo_hi_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_hi_hi = {maskSplit_maskSelect_lo_hi_hi_hi, maskSplit_maskSelect_lo_hi_hi_lo};
  wire [511:0]       maskSplit_maskSelect_lo_hi = {maskSplit_maskSelect_lo_hi_hi, maskSplit_maskSelect_lo_hi_lo};
  wire [1023:0]      maskSplit_maskSelect_lo = {maskSplit_maskSelect_lo_hi, maskSplit_maskSelect_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_lo = {maskSplit_maskSelect_hi_lo_lo_lo_hi, maskSplit_maskSelect_hi_lo_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_hi = {maskSplit_maskSelect_hi_lo_lo_hi_hi, maskSplit_maskSelect_hi_lo_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_lo_lo = {maskSplit_maskSelect_hi_lo_lo_hi, maskSplit_maskSelect_hi_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_lo = {maskSplit_maskSelect_hi_lo_hi_lo_hi, maskSplit_maskSelect_hi_lo_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_hi = {maskSplit_maskSelect_hi_lo_hi_hi_hi, maskSplit_maskSelect_hi_lo_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_lo_hi = {maskSplit_maskSelect_hi_lo_hi_hi, maskSplit_maskSelect_hi_lo_hi_lo};
  wire [511:0]       maskSplit_maskSelect_hi_lo = {maskSplit_maskSelect_hi_lo_hi, maskSplit_maskSelect_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_lo = {maskSplit_maskSelect_hi_hi_lo_lo_hi, maskSplit_maskSelect_hi_hi_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_hi = {maskSplit_maskSelect_hi_hi_lo_hi_hi, maskSplit_maskSelect_hi_hi_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_hi_lo = {maskSplit_maskSelect_hi_hi_lo_hi, maskSplit_maskSelect_hi_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_lo = {maskSplit_maskSelect_hi_hi_hi_lo_hi, maskSplit_maskSelect_hi_hi_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_hi = {maskSplit_maskSelect_hi_hi_hi_hi_hi, maskSplit_maskSelect_hi_hi_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_hi_hi = {maskSplit_maskSelect_hi_hi_hi_hi, maskSplit_maskSelect_hi_hi_hi_lo};
  wire [511:0]       maskSplit_maskSelect_hi_hi = {maskSplit_maskSelect_hi_hi_hi, maskSplit_maskSelect_hi_hi_lo};
  wire [1023:0]      maskSplit_maskSelect_hi = {maskSplit_maskSelect_hi_hi, maskSplit_maskSelect_hi_lo};
  wire [4:0]         executeGroupCounter;
  wire               maskSplit_vlMisAlign = |(instReg_vl[6:0]);
  wire [4:0]         maskSplit_lastexecuteGroup = instReg_vl[11:7] - {4'h0, ~maskSplit_vlMisAlign};
  wire               maskSplit_isVlBoundary = executeGroupCounter == maskSplit_lastexecuteGroup;
  wire               maskSplit_validExecuteGroup = executeGroupCounter <= maskSplit_lastexecuteGroup;
  wire [127:0]       _maskSplit_vlBoundaryCorrection_T_2 = 128'h1 << instReg_vl[6:0];
  wire [127:0]       _maskSplit_vlBoundaryCorrection_T_5 = _maskSplit_vlBoundaryCorrection_T_2 | {_maskSplit_vlBoundaryCorrection_T_2[126:0], 1'h0};
  wire [127:0]       _maskSplit_vlBoundaryCorrection_T_8 = _maskSplit_vlBoundaryCorrection_T_5 | {_maskSplit_vlBoundaryCorrection_T_5[125:0], 2'h0};
  wire [127:0]       _maskSplit_vlBoundaryCorrection_T_11 = _maskSplit_vlBoundaryCorrection_T_8 | {_maskSplit_vlBoundaryCorrection_T_8[123:0], 4'h0};
  wire [127:0]       _maskSplit_vlBoundaryCorrection_T_14 = _maskSplit_vlBoundaryCorrection_T_11 | {_maskSplit_vlBoundaryCorrection_T_11[119:0], 8'h0};
  wire [127:0]       _maskSplit_vlBoundaryCorrection_T_17 = _maskSplit_vlBoundaryCorrection_T_14 | {_maskSplit_vlBoundaryCorrection_T_14[111:0], 16'h0};
  wire [127:0]       _maskSplit_vlBoundaryCorrection_T_20 = _maskSplit_vlBoundaryCorrection_T_17 | {_maskSplit_vlBoundaryCorrection_T_17[95:0], 32'h0};
  wire [127:0]       maskSplit_vlBoundaryCorrection =
    ~({128{maskSplit_vlMisAlign & maskSplit_isVlBoundary}} & (_maskSplit_vlBoundaryCorrection_T_20 | {_maskSplit_vlBoundaryCorrection_T_20[63:0], 64'h0})) & {128{maskSplit_validExecuteGroup}};
  wire [15:0][127:0] _GEN_67 =
    {{maskSplit_maskSelect_hi[1023:896]},
     {maskSplit_maskSelect_hi[895:768]},
     {maskSplit_maskSelect_hi[767:640]},
     {maskSplit_maskSelect_hi[639:512]},
     {maskSplit_maskSelect_hi[511:384]},
     {maskSplit_maskSelect_hi[383:256]},
     {maskSplit_maskSelect_hi[255:128]},
     {maskSplit_maskSelect_hi[127:0]},
     {maskSplit_maskSelect_lo[1023:896]},
     {maskSplit_maskSelect_lo[895:768]},
     {maskSplit_maskSelect_lo[767:640]},
     {maskSplit_maskSelect_lo[639:512]},
     {maskSplit_maskSelect_lo[511:384]},
     {maskSplit_maskSelect_lo[383:256]},
     {maskSplit_maskSelect_lo[255:128]},
     {maskSplit_maskSelect_lo[127:0]}};
  wire [127:0]       maskSplit_0_2 = (instReg_maskType ? _GEN_67[executeGroupCounter[3:0]] : 128'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF) & maskSplit_vlBoundaryCorrection;
  wire [1:0]         maskSplit_byteMask_lo_lo_lo_lo_lo_lo = maskSplit_0_2[1:0];
  wire [1:0]         maskSplit_byteMask_lo_lo_lo_lo_lo_hi = maskSplit_0_2[3:2];
  wire [3:0]         maskSplit_byteMask_lo_lo_lo_lo_lo = {maskSplit_byteMask_lo_lo_lo_lo_lo_hi, maskSplit_byteMask_lo_lo_lo_lo_lo_lo};
  wire [1:0]         maskSplit_byteMask_lo_lo_lo_lo_hi_lo = maskSplit_0_2[5:4];
  wire [1:0]         maskSplit_byteMask_lo_lo_lo_lo_hi_hi = maskSplit_0_2[7:6];
  wire [3:0]         maskSplit_byteMask_lo_lo_lo_lo_hi = {maskSplit_byteMask_lo_lo_lo_lo_hi_hi, maskSplit_byteMask_lo_lo_lo_lo_hi_lo};
  wire [7:0]         maskSplit_byteMask_lo_lo_lo_lo = {maskSplit_byteMask_lo_lo_lo_lo_hi, maskSplit_byteMask_lo_lo_lo_lo_lo};
  wire [1:0]         maskSplit_byteMask_lo_lo_lo_hi_lo_lo = maskSplit_0_2[9:8];
  wire [1:0]         maskSplit_byteMask_lo_lo_lo_hi_lo_hi = maskSplit_0_2[11:10];
  wire [3:0]         maskSplit_byteMask_lo_lo_lo_hi_lo = {maskSplit_byteMask_lo_lo_lo_hi_lo_hi, maskSplit_byteMask_lo_lo_lo_hi_lo_lo};
  wire [1:0]         maskSplit_byteMask_lo_lo_lo_hi_hi_lo = maskSplit_0_2[13:12];
  wire [1:0]         maskSplit_byteMask_lo_lo_lo_hi_hi_hi = maskSplit_0_2[15:14];
  wire [3:0]         maskSplit_byteMask_lo_lo_lo_hi_hi = {maskSplit_byteMask_lo_lo_lo_hi_hi_hi, maskSplit_byteMask_lo_lo_lo_hi_hi_lo};
  wire [7:0]         maskSplit_byteMask_lo_lo_lo_hi = {maskSplit_byteMask_lo_lo_lo_hi_hi, maskSplit_byteMask_lo_lo_lo_hi_lo};
  wire [15:0]        maskSplit_byteMask_lo_lo_lo = {maskSplit_byteMask_lo_lo_lo_hi, maskSplit_byteMask_lo_lo_lo_lo};
  wire [1:0]         maskSplit_byteMask_lo_lo_hi_lo_lo_lo = maskSplit_0_2[17:16];
  wire [1:0]         maskSplit_byteMask_lo_lo_hi_lo_lo_hi = maskSplit_0_2[19:18];
  wire [3:0]         maskSplit_byteMask_lo_lo_hi_lo_lo = {maskSplit_byteMask_lo_lo_hi_lo_lo_hi, maskSplit_byteMask_lo_lo_hi_lo_lo_lo};
  wire [1:0]         maskSplit_byteMask_lo_lo_hi_lo_hi_lo = maskSplit_0_2[21:20];
  wire [1:0]         maskSplit_byteMask_lo_lo_hi_lo_hi_hi = maskSplit_0_2[23:22];
  wire [3:0]         maskSplit_byteMask_lo_lo_hi_lo_hi = {maskSplit_byteMask_lo_lo_hi_lo_hi_hi, maskSplit_byteMask_lo_lo_hi_lo_hi_lo};
  wire [7:0]         maskSplit_byteMask_lo_lo_hi_lo = {maskSplit_byteMask_lo_lo_hi_lo_hi, maskSplit_byteMask_lo_lo_hi_lo_lo};
  wire [1:0]         maskSplit_byteMask_lo_lo_hi_hi_lo_lo = maskSplit_0_2[25:24];
  wire [1:0]         maskSplit_byteMask_lo_lo_hi_hi_lo_hi = maskSplit_0_2[27:26];
  wire [3:0]         maskSplit_byteMask_lo_lo_hi_hi_lo = {maskSplit_byteMask_lo_lo_hi_hi_lo_hi, maskSplit_byteMask_lo_lo_hi_hi_lo_lo};
  wire [1:0]         maskSplit_byteMask_lo_lo_hi_hi_hi_lo = maskSplit_0_2[29:28];
  wire [1:0]         maskSplit_byteMask_lo_lo_hi_hi_hi_hi = maskSplit_0_2[31:30];
  wire [3:0]         maskSplit_byteMask_lo_lo_hi_hi_hi = {maskSplit_byteMask_lo_lo_hi_hi_hi_hi, maskSplit_byteMask_lo_lo_hi_hi_hi_lo};
  wire [7:0]         maskSplit_byteMask_lo_lo_hi_hi = {maskSplit_byteMask_lo_lo_hi_hi_hi, maskSplit_byteMask_lo_lo_hi_hi_lo};
  wire [15:0]        maskSplit_byteMask_lo_lo_hi = {maskSplit_byteMask_lo_lo_hi_hi, maskSplit_byteMask_lo_lo_hi_lo};
  wire [31:0]        maskSplit_byteMask_lo_lo = {maskSplit_byteMask_lo_lo_hi, maskSplit_byteMask_lo_lo_lo};
  wire [1:0]         maskSplit_byteMask_lo_hi_lo_lo_lo_lo = maskSplit_0_2[33:32];
  wire [1:0]         maskSplit_byteMask_lo_hi_lo_lo_lo_hi = maskSplit_0_2[35:34];
  wire [3:0]         maskSplit_byteMask_lo_hi_lo_lo_lo = {maskSplit_byteMask_lo_hi_lo_lo_lo_hi, maskSplit_byteMask_lo_hi_lo_lo_lo_lo};
  wire [1:0]         maskSplit_byteMask_lo_hi_lo_lo_hi_lo = maskSplit_0_2[37:36];
  wire [1:0]         maskSplit_byteMask_lo_hi_lo_lo_hi_hi = maskSplit_0_2[39:38];
  wire [3:0]         maskSplit_byteMask_lo_hi_lo_lo_hi = {maskSplit_byteMask_lo_hi_lo_lo_hi_hi, maskSplit_byteMask_lo_hi_lo_lo_hi_lo};
  wire [7:0]         maskSplit_byteMask_lo_hi_lo_lo = {maskSplit_byteMask_lo_hi_lo_lo_hi, maskSplit_byteMask_lo_hi_lo_lo_lo};
  wire [1:0]         maskSplit_byteMask_lo_hi_lo_hi_lo_lo = maskSplit_0_2[41:40];
  wire [1:0]         maskSplit_byteMask_lo_hi_lo_hi_lo_hi = maskSplit_0_2[43:42];
  wire [3:0]         maskSplit_byteMask_lo_hi_lo_hi_lo = {maskSplit_byteMask_lo_hi_lo_hi_lo_hi, maskSplit_byteMask_lo_hi_lo_hi_lo_lo};
  wire [1:0]         maskSplit_byteMask_lo_hi_lo_hi_hi_lo = maskSplit_0_2[45:44];
  wire [1:0]         maskSplit_byteMask_lo_hi_lo_hi_hi_hi = maskSplit_0_2[47:46];
  wire [3:0]         maskSplit_byteMask_lo_hi_lo_hi_hi = {maskSplit_byteMask_lo_hi_lo_hi_hi_hi, maskSplit_byteMask_lo_hi_lo_hi_hi_lo};
  wire [7:0]         maskSplit_byteMask_lo_hi_lo_hi = {maskSplit_byteMask_lo_hi_lo_hi_hi, maskSplit_byteMask_lo_hi_lo_hi_lo};
  wire [15:0]        maskSplit_byteMask_lo_hi_lo = {maskSplit_byteMask_lo_hi_lo_hi, maskSplit_byteMask_lo_hi_lo_lo};
  wire [1:0]         maskSplit_byteMask_lo_hi_hi_lo_lo_lo = maskSplit_0_2[49:48];
  wire [1:0]         maskSplit_byteMask_lo_hi_hi_lo_lo_hi = maskSplit_0_2[51:50];
  wire [3:0]         maskSplit_byteMask_lo_hi_hi_lo_lo = {maskSplit_byteMask_lo_hi_hi_lo_lo_hi, maskSplit_byteMask_lo_hi_hi_lo_lo_lo};
  wire [1:0]         maskSplit_byteMask_lo_hi_hi_lo_hi_lo = maskSplit_0_2[53:52];
  wire [1:0]         maskSplit_byteMask_lo_hi_hi_lo_hi_hi = maskSplit_0_2[55:54];
  wire [3:0]         maskSplit_byteMask_lo_hi_hi_lo_hi = {maskSplit_byteMask_lo_hi_hi_lo_hi_hi, maskSplit_byteMask_lo_hi_hi_lo_hi_lo};
  wire [7:0]         maskSplit_byteMask_lo_hi_hi_lo = {maskSplit_byteMask_lo_hi_hi_lo_hi, maskSplit_byteMask_lo_hi_hi_lo_lo};
  wire [1:0]         maskSplit_byteMask_lo_hi_hi_hi_lo_lo = maskSplit_0_2[57:56];
  wire [1:0]         maskSplit_byteMask_lo_hi_hi_hi_lo_hi = maskSplit_0_2[59:58];
  wire [3:0]         maskSplit_byteMask_lo_hi_hi_hi_lo = {maskSplit_byteMask_lo_hi_hi_hi_lo_hi, maskSplit_byteMask_lo_hi_hi_hi_lo_lo};
  wire [1:0]         maskSplit_byteMask_lo_hi_hi_hi_hi_lo = maskSplit_0_2[61:60];
  wire [1:0]         maskSplit_byteMask_lo_hi_hi_hi_hi_hi = maskSplit_0_2[63:62];
  wire [3:0]         maskSplit_byteMask_lo_hi_hi_hi_hi = {maskSplit_byteMask_lo_hi_hi_hi_hi_hi, maskSplit_byteMask_lo_hi_hi_hi_hi_lo};
  wire [7:0]         maskSplit_byteMask_lo_hi_hi_hi = {maskSplit_byteMask_lo_hi_hi_hi_hi, maskSplit_byteMask_lo_hi_hi_hi_lo};
  wire [15:0]        maskSplit_byteMask_lo_hi_hi = {maskSplit_byteMask_lo_hi_hi_hi, maskSplit_byteMask_lo_hi_hi_lo};
  wire [31:0]        maskSplit_byteMask_lo_hi = {maskSplit_byteMask_lo_hi_hi, maskSplit_byteMask_lo_hi_lo};
  wire [63:0]        maskSplit_byteMask_lo = {maskSplit_byteMask_lo_hi, maskSplit_byteMask_lo_lo};
  wire [1:0]         maskSplit_byteMask_hi_lo_lo_lo_lo_lo = maskSplit_0_2[65:64];
  wire [1:0]         maskSplit_byteMask_hi_lo_lo_lo_lo_hi = maskSplit_0_2[67:66];
  wire [3:0]         maskSplit_byteMask_hi_lo_lo_lo_lo = {maskSplit_byteMask_hi_lo_lo_lo_lo_hi, maskSplit_byteMask_hi_lo_lo_lo_lo_lo};
  wire [1:0]         maskSplit_byteMask_hi_lo_lo_lo_hi_lo = maskSplit_0_2[69:68];
  wire [1:0]         maskSplit_byteMask_hi_lo_lo_lo_hi_hi = maskSplit_0_2[71:70];
  wire [3:0]         maskSplit_byteMask_hi_lo_lo_lo_hi = {maskSplit_byteMask_hi_lo_lo_lo_hi_hi, maskSplit_byteMask_hi_lo_lo_lo_hi_lo};
  wire [7:0]         maskSplit_byteMask_hi_lo_lo_lo = {maskSplit_byteMask_hi_lo_lo_lo_hi, maskSplit_byteMask_hi_lo_lo_lo_lo};
  wire [1:0]         maskSplit_byteMask_hi_lo_lo_hi_lo_lo = maskSplit_0_2[73:72];
  wire [1:0]         maskSplit_byteMask_hi_lo_lo_hi_lo_hi = maskSplit_0_2[75:74];
  wire [3:0]         maskSplit_byteMask_hi_lo_lo_hi_lo = {maskSplit_byteMask_hi_lo_lo_hi_lo_hi, maskSplit_byteMask_hi_lo_lo_hi_lo_lo};
  wire [1:0]         maskSplit_byteMask_hi_lo_lo_hi_hi_lo = maskSplit_0_2[77:76];
  wire [1:0]         maskSplit_byteMask_hi_lo_lo_hi_hi_hi = maskSplit_0_2[79:78];
  wire [3:0]         maskSplit_byteMask_hi_lo_lo_hi_hi = {maskSplit_byteMask_hi_lo_lo_hi_hi_hi, maskSplit_byteMask_hi_lo_lo_hi_hi_lo};
  wire [7:0]         maskSplit_byteMask_hi_lo_lo_hi = {maskSplit_byteMask_hi_lo_lo_hi_hi, maskSplit_byteMask_hi_lo_lo_hi_lo};
  wire [15:0]        maskSplit_byteMask_hi_lo_lo = {maskSplit_byteMask_hi_lo_lo_hi, maskSplit_byteMask_hi_lo_lo_lo};
  wire [1:0]         maskSplit_byteMask_hi_lo_hi_lo_lo_lo = maskSplit_0_2[81:80];
  wire [1:0]         maskSplit_byteMask_hi_lo_hi_lo_lo_hi = maskSplit_0_2[83:82];
  wire [3:0]         maskSplit_byteMask_hi_lo_hi_lo_lo = {maskSplit_byteMask_hi_lo_hi_lo_lo_hi, maskSplit_byteMask_hi_lo_hi_lo_lo_lo};
  wire [1:0]         maskSplit_byteMask_hi_lo_hi_lo_hi_lo = maskSplit_0_2[85:84];
  wire [1:0]         maskSplit_byteMask_hi_lo_hi_lo_hi_hi = maskSplit_0_2[87:86];
  wire [3:0]         maskSplit_byteMask_hi_lo_hi_lo_hi = {maskSplit_byteMask_hi_lo_hi_lo_hi_hi, maskSplit_byteMask_hi_lo_hi_lo_hi_lo};
  wire [7:0]         maskSplit_byteMask_hi_lo_hi_lo = {maskSplit_byteMask_hi_lo_hi_lo_hi, maskSplit_byteMask_hi_lo_hi_lo_lo};
  wire [1:0]         maskSplit_byteMask_hi_lo_hi_hi_lo_lo = maskSplit_0_2[89:88];
  wire [1:0]         maskSplit_byteMask_hi_lo_hi_hi_lo_hi = maskSplit_0_2[91:90];
  wire [3:0]         maskSplit_byteMask_hi_lo_hi_hi_lo = {maskSplit_byteMask_hi_lo_hi_hi_lo_hi, maskSplit_byteMask_hi_lo_hi_hi_lo_lo};
  wire [1:0]         maskSplit_byteMask_hi_lo_hi_hi_hi_lo = maskSplit_0_2[93:92];
  wire [1:0]         maskSplit_byteMask_hi_lo_hi_hi_hi_hi = maskSplit_0_2[95:94];
  wire [3:0]         maskSplit_byteMask_hi_lo_hi_hi_hi = {maskSplit_byteMask_hi_lo_hi_hi_hi_hi, maskSplit_byteMask_hi_lo_hi_hi_hi_lo};
  wire [7:0]         maskSplit_byteMask_hi_lo_hi_hi = {maskSplit_byteMask_hi_lo_hi_hi_hi, maskSplit_byteMask_hi_lo_hi_hi_lo};
  wire [15:0]        maskSplit_byteMask_hi_lo_hi = {maskSplit_byteMask_hi_lo_hi_hi, maskSplit_byteMask_hi_lo_hi_lo};
  wire [31:0]        maskSplit_byteMask_hi_lo = {maskSplit_byteMask_hi_lo_hi, maskSplit_byteMask_hi_lo_lo};
  wire [1:0]         maskSplit_byteMask_hi_hi_lo_lo_lo_lo = maskSplit_0_2[97:96];
  wire [1:0]         maskSplit_byteMask_hi_hi_lo_lo_lo_hi = maskSplit_0_2[99:98];
  wire [3:0]         maskSplit_byteMask_hi_hi_lo_lo_lo = {maskSplit_byteMask_hi_hi_lo_lo_lo_hi, maskSplit_byteMask_hi_hi_lo_lo_lo_lo};
  wire [1:0]         maskSplit_byteMask_hi_hi_lo_lo_hi_lo = maskSplit_0_2[101:100];
  wire [1:0]         maskSplit_byteMask_hi_hi_lo_lo_hi_hi = maskSplit_0_2[103:102];
  wire [3:0]         maskSplit_byteMask_hi_hi_lo_lo_hi = {maskSplit_byteMask_hi_hi_lo_lo_hi_hi, maskSplit_byteMask_hi_hi_lo_lo_hi_lo};
  wire [7:0]         maskSplit_byteMask_hi_hi_lo_lo = {maskSplit_byteMask_hi_hi_lo_lo_hi, maskSplit_byteMask_hi_hi_lo_lo_lo};
  wire [1:0]         maskSplit_byteMask_hi_hi_lo_hi_lo_lo = maskSplit_0_2[105:104];
  wire [1:0]         maskSplit_byteMask_hi_hi_lo_hi_lo_hi = maskSplit_0_2[107:106];
  wire [3:0]         maskSplit_byteMask_hi_hi_lo_hi_lo = {maskSplit_byteMask_hi_hi_lo_hi_lo_hi, maskSplit_byteMask_hi_hi_lo_hi_lo_lo};
  wire [1:0]         maskSplit_byteMask_hi_hi_lo_hi_hi_lo = maskSplit_0_2[109:108];
  wire [1:0]         maskSplit_byteMask_hi_hi_lo_hi_hi_hi = maskSplit_0_2[111:110];
  wire [3:0]         maskSplit_byteMask_hi_hi_lo_hi_hi = {maskSplit_byteMask_hi_hi_lo_hi_hi_hi, maskSplit_byteMask_hi_hi_lo_hi_hi_lo};
  wire [7:0]         maskSplit_byteMask_hi_hi_lo_hi = {maskSplit_byteMask_hi_hi_lo_hi_hi, maskSplit_byteMask_hi_hi_lo_hi_lo};
  wire [15:0]        maskSplit_byteMask_hi_hi_lo = {maskSplit_byteMask_hi_hi_lo_hi, maskSplit_byteMask_hi_hi_lo_lo};
  wire [1:0]         maskSplit_byteMask_hi_hi_hi_lo_lo_lo = maskSplit_0_2[113:112];
  wire [1:0]         maskSplit_byteMask_hi_hi_hi_lo_lo_hi = maskSplit_0_2[115:114];
  wire [3:0]         maskSplit_byteMask_hi_hi_hi_lo_lo = {maskSplit_byteMask_hi_hi_hi_lo_lo_hi, maskSplit_byteMask_hi_hi_hi_lo_lo_lo};
  wire [1:0]         maskSplit_byteMask_hi_hi_hi_lo_hi_lo = maskSplit_0_2[117:116];
  wire [1:0]         maskSplit_byteMask_hi_hi_hi_lo_hi_hi = maskSplit_0_2[119:118];
  wire [3:0]         maskSplit_byteMask_hi_hi_hi_lo_hi = {maskSplit_byteMask_hi_hi_hi_lo_hi_hi, maskSplit_byteMask_hi_hi_hi_lo_hi_lo};
  wire [7:0]         maskSplit_byteMask_hi_hi_hi_lo = {maskSplit_byteMask_hi_hi_hi_lo_hi, maskSplit_byteMask_hi_hi_hi_lo_lo};
  wire [1:0]         maskSplit_byteMask_hi_hi_hi_hi_lo_lo = maskSplit_0_2[121:120];
  wire [1:0]         maskSplit_byteMask_hi_hi_hi_hi_lo_hi = maskSplit_0_2[123:122];
  wire [3:0]         maskSplit_byteMask_hi_hi_hi_hi_lo = {maskSplit_byteMask_hi_hi_hi_hi_lo_hi, maskSplit_byteMask_hi_hi_hi_hi_lo_lo};
  wire [1:0]         maskSplit_byteMask_hi_hi_hi_hi_hi_lo = maskSplit_0_2[125:124];
  wire [1:0]         maskSplit_byteMask_hi_hi_hi_hi_hi_hi = maskSplit_0_2[127:126];
  wire [3:0]         maskSplit_byteMask_hi_hi_hi_hi_hi = {maskSplit_byteMask_hi_hi_hi_hi_hi_hi, maskSplit_byteMask_hi_hi_hi_hi_hi_lo};
  wire [7:0]         maskSplit_byteMask_hi_hi_hi_hi = {maskSplit_byteMask_hi_hi_hi_hi_hi, maskSplit_byteMask_hi_hi_hi_hi_lo};
  wire [15:0]        maskSplit_byteMask_hi_hi_hi = {maskSplit_byteMask_hi_hi_hi_hi, maskSplit_byteMask_hi_hi_hi_lo};
  wire [31:0]        maskSplit_byteMask_hi_hi = {maskSplit_byteMask_hi_hi_hi, maskSplit_byteMask_hi_hi_lo};
  wire [63:0]        maskSplit_byteMask_hi = {maskSplit_byteMask_hi_hi, maskSplit_byteMask_hi_lo};
  wire [127:0]       maskSplit_0_1 = {maskSplit_byteMask_hi, maskSplit_byteMask_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_lo_1 = {maskSplit_maskSelect_lo_lo_lo_lo_hi_1, maskSplit_maskSelect_lo_lo_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_hi_1 = {maskSplit_maskSelect_lo_lo_lo_hi_hi_1, maskSplit_maskSelect_lo_lo_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_lo_lo_1 = {maskSplit_maskSelect_lo_lo_lo_hi_1, maskSplit_maskSelect_lo_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_lo_1 = {maskSplit_maskSelect_lo_lo_hi_lo_hi_1, maskSplit_maskSelect_lo_lo_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_hi_1 = {maskSplit_maskSelect_lo_lo_hi_hi_hi_1, maskSplit_maskSelect_lo_lo_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_lo_hi_1 = {maskSplit_maskSelect_lo_lo_hi_hi_1, maskSplit_maskSelect_lo_lo_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_lo_lo_1 = {maskSplit_maskSelect_lo_lo_hi_1, maskSplit_maskSelect_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_lo_1 = {maskSplit_maskSelect_lo_hi_lo_lo_hi_1, maskSplit_maskSelect_lo_hi_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_hi_1 = {maskSplit_maskSelect_lo_hi_lo_hi_hi_1, maskSplit_maskSelect_lo_hi_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_hi_lo_1 = {maskSplit_maskSelect_lo_hi_lo_hi_1, maskSplit_maskSelect_lo_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_lo_1 = {maskSplit_maskSelect_lo_hi_hi_lo_hi_1, maskSplit_maskSelect_lo_hi_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_hi_1 = {maskSplit_maskSelect_lo_hi_hi_hi_hi_1, maskSplit_maskSelect_lo_hi_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_hi_hi_1 = {maskSplit_maskSelect_lo_hi_hi_hi_1, maskSplit_maskSelect_lo_hi_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_lo_hi_1 = {maskSplit_maskSelect_lo_hi_hi_1, maskSplit_maskSelect_lo_hi_lo_1};
  wire [1023:0]      maskSplit_maskSelect_lo_1 = {maskSplit_maskSelect_lo_hi_1, maskSplit_maskSelect_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_lo_1 = {maskSplit_maskSelect_hi_lo_lo_lo_hi_1, maskSplit_maskSelect_hi_lo_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_hi_1 = {maskSplit_maskSelect_hi_lo_lo_hi_hi_1, maskSplit_maskSelect_hi_lo_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_lo_lo_1 = {maskSplit_maskSelect_hi_lo_lo_hi_1, maskSplit_maskSelect_hi_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_lo_1 = {maskSplit_maskSelect_hi_lo_hi_lo_hi_1, maskSplit_maskSelect_hi_lo_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_hi_1 = {maskSplit_maskSelect_hi_lo_hi_hi_hi_1, maskSplit_maskSelect_hi_lo_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_lo_hi_1 = {maskSplit_maskSelect_hi_lo_hi_hi_1, maskSplit_maskSelect_hi_lo_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_hi_lo_1 = {maskSplit_maskSelect_hi_lo_hi_1, maskSplit_maskSelect_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_lo_1 = {maskSplit_maskSelect_hi_hi_lo_lo_hi_1, maskSplit_maskSelect_hi_hi_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_hi_1 = {maskSplit_maskSelect_hi_hi_lo_hi_hi_1, maskSplit_maskSelect_hi_hi_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_hi_lo_1 = {maskSplit_maskSelect_hi_hi_lo_hi_1, maskSplit_maskSelect_hi_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_lo_1 = {maskSplit_maskSelect_hi_hi_hi_lo_hi_1, maskSplit_maskSelect_hi_hi_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_hi_1 = {maskSplit_maskSelect_hi_hi_hi_hi_hi_1, maskSplit_maskSelect_hi_hi_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_hi_hi_1 = {maskSplit_maskSelect_hi_hi_hi_hi_1, maskSplit_maskSelect_hi_hi_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_hi_hi_1 = {maskSplit_maskSelect_hi_hi_hi_1, maskSplit_maskSelect_hi_hi_lo_1};
  wire [1023:0]      maskSplit_maskSelect_hi_1 = {maskSplit_maskSelect_hi_hi_1, maskSplit_maskSelect_hi_lo_1};
  wire               maskSplit_vlMisAlign_1 = |(instReg_vl[5:0]);
  wire [5:0]         maskSplit_lastexecuteGroup_1 = instReg_vl[11:6] - {5'h0, ~maskSplit_vlMisAlign_1};
  wire [5:0]         _GEN_68 = {1'h0, executeGroupCounter};
  wire               maskSplit_isVlBoundary_1 = _GEN_68 == maskSplit_lastexecuteGroup_1;
  wire               maskSplit_validExecuteGroup_1 = _GEN_68 <= maskSplit_lastexecuteGroup_1;
  wire [63:0]        _maskSplit_vlBoundaryCorrection_T_30 = 64'h1 << instReg_vl[5:0];
  wire [63:0]        _maskSplit_vlBoundaryCorrection_T_33 = _maskSplit_vlBoundaryCorrection_T_30 | {_maskSplit_vlBoundaryCorrection_T_30[62:0], 1'h0};
  wire [63:0]        _maskSplit_vlBoundaryCorrection_T_36 = _maskSplit_vlBoundaryCorrection_T_33 | {_maskSplit_vlBoundaryCorrection_T_33[61:0], 2'h0};
  wire [63:0]        _maskSplit_vlBoundaryCorrection_T_39 = _maskSplit_vlBoundaryCorrection_T_36 | {_maskSplit_vlBoundaryCorrection_T_36[59:0], 4'h0};
  wire [63:0]        _maskSplit_vlBoundaryCorrection_T_42 = _maskSplit_vlBoundaryCorrection_T_39 | {_maskSplit_vlBoundaryCorrection_T_39[55:0], 8'h0};
  wire [63:0]        _maskSplit_vlBoundaryCorrection_T_45 = _maskSplit_vlBoundaryCorrection_T_42 | {_maskSplit_vlBoundaryCorrection_T_42[47:0], 16'h0};
  wire [63:0]        maskSplit_vlBoundaryCorrection_1 =
    ~({64{maskSplit_vlMisAlign_1 & maskSplit_isVlBoundary_1}} & (_maskSplit_vlBoundaryCorrection_T_45 | {_maskSplit_vlBoundaryCorrection_T_45[31:0], 32'h0})) & {64{maskSplit_validExecuteGroup_1}};
  wire [31:0][63:0]  _GEN_69 =
    {{maskSplit_maskSelect_hi_1[1023:960]},
     {maskSplit_maskSelect_hi_1[959:896]},
     {maskSplit_maskSelect_hi_1[895:832]},
     {maskSplit_maskSelect_hi_1[831:768]},
     {maskSplit_maskSelect_hi_1[767:704]},
     {maskSplit_maskSelect_hi_1[703:640]},
     {maskSplit_maskSelect_hi_1[639:576]},
     {maskSplit_maskSelect_hi_1[575:512]},
     {maskSplit_maskSelect_hi_1[511:448]},
     {maskSplit_maskSelect_hi_1[447:384]},
     {maskSplit_maskSelect_hi_1[383:320]},
     {maskSplit_maskSelect_hi_1[319:256]},
     {maskSplit_maskSelect_hi_1[255:192]},
     {maskSplit_maskSelect_hi_1[191:128]},
     {maskSplit_maskSelect_hi_1[127:64]},
     {maskSplit_maskSelect_hi_1[63:0]},
     {maskSplit_maskSelect_lo_1[1023:960]},
     {maskSplit_maskSelect_lo_1[959:896]},
     {maskSplit_maskSelect_lo_1[895:832]},
     {maskSplit_maskSelect_lo_1[831:768]},
     {maskSplit_maskSelect_lo_1[767:704]},
     {maskSplit_maskSelect_lo_1[703:640]},
     {maskSplit_maskSelect_lo_1[639:576]},
     {maskSplit_maskSelect_lo_1[575:512]},
     {maskSplit_maskSelect_lo_1[511:448]},
     {maskSplit_maskSelect_lo_1[447:384]},
     {maskSplit_maskSelect_lo_1[383:320]},
     {maskSplit_maskSelect_lo_1[319:256]},
     {maskSplit_maskSelect_lo_1[255:192]},
     {maskSplit_maskSelect_lo_1[191:128]},
     {maskSplit_maskSelect_lo_1[127:64]},
     {maskSplit_maskSelect_lo_1[63:0]}};
  wire [63:0]        maskSplit_1_2 = (instReg_maskType ? _GEN_69[executeGroupCounter] : 64'hFFFFFFFFFFFFFFFF) & maskSplit_vlBoundaryCorrection_1;
  wire [3:0]         maskSplit_byteMask_lo_lo_lo_lo_lo_1 = {{2{maskSplit_1_2[1]}}, {2{maskSplit_1_2[0]}}};
  wire [3:0]         maskSplit_byteMask_lo_lo_lo_lo_hi_1 = {{2{maskSplit_1_2[3]}}, {2{maskSplit_1_2[2]}}};
  wire [7:0]         maskSplit_byteMask_lo_lo_lo_lo_1 = {maskSplit_byteMask_lo_lo_lo_lo_hi_1, maskSplit_byteMask_lo_lo_lo_lo_lo_1};
  wire [3:0]         maskSplit_byteMask_lo_lo_lo_hi_lo_1 = {{2{maskSplit_1_2[5]}}, {2{maskSplit_1_2[4]}}};
  wire [3:0]         maskSplit_byteMask_lo_lo_lo_hi_hi_1 = {{2{maskSplit_1_2[7]}}, {2{maskSplit_1_2[6]}}};
  wire [7:0]         maskSplit_byteMask_lo_lo_lo_hi_1 = {maskSplit_byteMask_lo_lo_lo_hi_hi_1, maskSplit_byteMask_lo_lo_lo_hi_lo_1};
  wire [15:0]        maskSplit_byteMask_lo_lo_lo_1 = {maskSplit_byteMask_lo_lo_lo_hi_1, maskSplit_byteMask_lo_lo_lo_lo_1};
  wire [3:0]         maskSplit_byteMask_lo_lo_hi_lo_lo_1 = {{2{maskSplit_1_2[9]}}, {2{maskSplit_1_2[8]}}};
  wire [3:0]         maskSplit_byteMask_lo_lo_hi_lo_hi_1 = {{2{maskSplit_1_2[11]}}, {2{maskSplit_1_2[10]}}};
  wire [7:0]         maskSplit_byteMask_lo_lo_hi_lo_1 = {maskSplit_byteMask_lo_lo_hi_lo_hi_1, maskSplit_byteMask_lo_lo_hi_lo_lo_1};
  wire [3:0]         maskSplit_byteMask_lo_lo_hi_hi_lo_1 = {{2{maskSplit_1_2[13]}}, {2{maskSplit_1_2[12]}}};
  wire [3:0]         maskSplit_byteMask_lo_lo_hi_hi_hi_1 = {{2{maskSplit_1_2[15]}}, {2{maskSplit_1_2[14]}}};
  wire [7:0]         maskSplit_byteMask_lo_lo_hi_hi_1 = {maskSplit_byteMask_lo_lo_hi_hi_hi_1, maskSplit_byteMask_lo_lo_hi_hi_lo_1};
  wire [15:0]        maskSplit_byteMask_lo_lo_hi_1 = {maskSplit_byteMask_lo_lo_hi_hi_1, maskSplit_byteMask_lo_lo_hi_lo_1};
  wire [31:0]        maskSplit_byteMask_lo_lo_1 = {maskSplit_byteMask_lo_lo_hi_1, maskSplit_byteMask_lo_lo_lo_1};
  wire [3:0]         maskSplit_byteMask_lo_hi_lo_lo_lo_1 = {{2{maskSplit_1_2[17]}}, {2{maskSplit_1_2[16]}}};
  wire [3:0]         maskSplit_byteMask_lo_hi_lo_lo_hi_1 = {{2{maskSplit_1_2[19]}}, {2{maskSplit_1_2[18]}}};
  wire [7:0]         maskSplit_byteMask_lo_hi_lo_lo_1 = {maskSplit_byteMask_lo_hi_lo_lo_hi_1, maskSplit_byteMask_lo_hi_lo_lo_lo_1};
  wire [3:0]         maskSplit_byteMask_lo_hi_lo_hi_lo_1 = {{2{maskSplit_1_2[21]}}, {2{maskSplit_1_2[20]}}};
  wire [3:0]         maskSplit_byteMask_lo_hi_lo_hi_hi_1 = {{2{maskSplit_1_2[23]}}, {2{maskSplit_1_2[22]}}};
  wire [7:0]         maskSplit_byteMask_lo_hi_lo_hi_1 = {maskSplit_byteMask_lo_hi_lo_hi_hi_1, maskSplit_byteMask_lo_hi_lo_hi_lo_1};
  wire [15:0]        maskSplit_byteMask_lo_hi_lo_1 = {maskSplit_byteMask_lo_hi_lo_hi_1, maskSplit_byteMask_lo_hi_lo_lo_1};
  wire [3:0]         maskSplit_byteMask_lo_hi_hi_lo_lo_1 = {{2{maskSplit_1_2[25]}}, {2{maskSplit_1_2[24]}}};
  wire [3:0]         maskSplit_byteMask_lo_hi_hi_lo_hi_1 = {{2{maskSplit_1_2[27]}}, {2{maskSplit_1_2[26]}}};
  wire [7:0]         maskSplit_byteMask_lo_hi_hi_lo_1 = {maskSplit_byteMask_lo_hi_hi_lo_hi_1, maskSplit_byteMask_lo_hi_hi_lo_lo_1};
  wire [3:0]         maskSplit_byteMask_lo_hi_hi_hi_lo_1 = {{2{maskSplit_1_2[29]}}, {2{maskSplit_1_2[28]}}};
  wire [3:0]         maskSplit_byteMask_lo_hi_hi_hi_hi_1 = {{2{maskSplit_1_2[31]}}, {2{maskSplit_1_2[30]}}};
  wire [7:0]         maskSplit_byteMask_lo_hi_hi_hi_1 = {maskSplit_byteMask_lo_hi_hi_hi_hi_1, maskSplit_byteMask_lo_hi_hi_hi_lo_1};
  wire [15:0]        maskSplit_byteMask_lo_hi_hi_1 = {maskSplit_byteMask_lo_hi_hi_hi_1, maskSplit_byteMask_lo_hi_hi_lo_1};
  wire [31:0]        maskSplit_byteMask_lo_hi_1 = {maskSplit_byteMask_lo_hi_hi_1, maskSplit_byteMask_lo_hi_lo_1};
  wire [63:0]        maskSplit_byteMask_lo_1 = {maskSplit_byteMask_lo_hi_1, maskSplit_byteMask_lo_lo_1};
  wire [3:0]         maskSplit_byteMask_hi_lo_lo_lo_lo_1 = {{2{maskSplit_1_2[33]}}, {2{maskSplit_1_2[32]}}};
  wire [3:0]         maskSplit_byteMask_hi_lo_lo_lo_hi_1 = {{2{maskSplit_1_2[35]}}, {2{maskSplit_1_2[34]}}};
  wire [7:0]         maskSplit_byteMask_hi_lo_lo_lo_1 = {maskSplit_byteMask_hi_lo_lo_lo_hi_1, maskSplit_byteMask_hi_lo_lo_lo_lo_1};
  wire [3:0]         maskSplit_byteMask_hi_lo_lo_hi_lo_1 = {{2{maskSplit_1_2[37]}}, {2{maskSplit_1_2[36]}}};
  wire [3:0]         maskSplit_byteMask_hi_lo_lo_hi_hi_1 = {{2{maskSplit_1_2[39]}}, {2{maskSplit_1_2[38]}}};
  wire [7:0]         maskSplit_byteMask_hi_lo_lo_hi_1 = {maskSplit_byteMask_hi_lo_lo_hi_hi_1, maskSplit_byteMask_hi_lo_lo_hi_lo_1};
  wire [15:0]        maskSplit_byteMask_hi_lo_lo_1 = {maskSplit_byteMask_hi_lo_lo_hi_1, maskSplit_byteMask_hi_lo_lo_lo_1};
  wire [3:0]         maskSplit_byteMask_hi_lo_hi_lo_lo_1 = {{2{maskSplit_1_2[41]}}, {2{maskSplit_1_2[40]}}};
  wire [3:0]         maskSplit_byteMask_hi_lo_hi_lo_hi_1 = {{2{maskSplit_1_2[43]}}, {2{maskSplit_1_2[42]}}};
  wire [7:0]         maskSplit_byteMask_hi_lo_hi_lo_1 = {maskSplit_byteMask_hi_lo_hi_lo_hi_1, maskSplit_byteMask_hi_lo_hi_lo_lo_1};
  wire [3:0]         maskSplit_byteMask_hi_lo_hi_hi_lo_1 = {{2{maskSplit_1_2[45]}}, {2{maskSplit_1_2[44]}}};
  wire [3:0]         maskSplit_byteMask_hi_lo_hi_hi_hi_1 = {{2{maskSplit_1_2[47]}}, {2{maskSplit_1_2[46]}}};
  wire [7:0]         maskSplit_byteMask_hi_lo_hi_hi_1 = {maskSplit_byteMask_hi_lo_hi_hi_hi_1, maskSplit_byteMask_hi_lo_hi_hi_lo_1};
  wire [15:0]        maskSplit_byteMask_hi_lo_hi_1 = {maskSplit_byteMask_hi_lo_hi_hi_1, maskSplit_byteMask_hi_lo_hi_lo_1};
  wire [31:0]        maskSplit_byteMask_hi_lo_1 = {maskSplit_byteMask_hi_lo_hi_1, maskSplit_byteMask_hi_lo_lo_1};
  wire [3:0]         maskSplit_byteMask_hi_hi_lo_lo_lo_1 = {{2{maskSplit_1_2[49]}}, {2{maskSplit_1_2[48]}}};
  wire [3:0]         maskSplit_byteMask_hi_hi_lo_lo_hi_1 = {{2{maskSplit_1_2[51]}}, {2{maskSplit_1_2[50]}}};
  wire [7:0]         maskSplit_byteMask_hi_hi_lo_lo_1 = {maskSplit_byteMask_hi_hi_lo_lo_hi_1, maskSplit_byteMask_hi_hi_lo_lo_lo_1};
  wire [3:0]         maskSplit_byteMask_hi_hi_lo_hi_lo_1 = {{2{maskSplit_1_2[53]}}, {2{maskSplit_1_2[52]}}};
  wire [3:0]         maskSplit_byteMask_hi_hi_lo_hi_hi_1 = {{2{maskSplit_1_2[55]}}, {2{maskSplit_1_2[54]}}};
  wire [7:0]         maskSplit_byteMask_hi_hi_lo_hi_1 = {maskSplit_byteMask_hi_hi_lo_hi_hi_1, maskSplit_byteMask_hi_hi_lo_hi_lo_1};
  wire [15:0]        maskSplit_byteMask_hi_hi_lo_1 = {maskSplit_byteMask_hi_hi_lo_hi_1, maskSplit_byteMask_hi_hi_lo_lo_1};
  wire [3:0]         maskSplit_byteMask_hi_hi_hi_lo_lo_1 = {{2{maskSplit_1_2[57]}}, {2{maskSplit_1_2[56]}}};
  wire [3:0]         maskSplit_byteMask_hi_hi_hi_lo_hi_1 = {{2{maskSplit_1_2[59]}}, {2{maskSplit_1_2[58]}}};
  wire [7:0]         maskSplit_byteMask_hi_hi_hi_lo_1 = {maskSplit_byteMask_hi_hi_hi_lo_hi_1, maskSplit_byteMask_hi_hi_hi_lo_lo_1};
  wire [3:0]         maskSplit_byteMask_hi_hi_hi_hi_lo_1 = {{2{maskSplit_1_2[61]}}, {2{maskSplit_1_2[60]}}};
  wire [3:0]         maskSplit_byteMask_hi_hi_hi_hi_hi_1 = {{2{maskSplit_1_2[63]}}, {2{maskSplit_1_2[62]}}};
  wire [7:0]         maskSplit_byteMask_hi_hi_hi_hi_1 = {maskSplit_byteMask_hi_hi_hi_hi_hi_1, maskSplit_byteMask_hi_hi_hi_hi_lo_1};
  wire [15:0]        maskSplit_byteMask_hi_hi_hi_1 = {maskSplit_byteMask_hi_hi_hi_hi_1, maskSplit_byteMask_hi_hi_hi_lo_1};
  wire [31:0]        maskSplit_byteMask_hi_hi_1 = {maskSplit_byteMask_hi_hi_hi_1, maskSplit_byteMask_hi_hi_lo_1};
  wire [63:0]        maskSplit_byteMask_hi_1 = {maskSplit_byteMask_hi_hi_1, maskSplit_byteMask_hi_lo_1};
  wire [127:0]       maskSplit_1_1 = {maskSplit_byteMask_hi_1, maskSplit_byteMask_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_lo_2 = {maskSplit_maskSelect_lo_lo_lo_lo_hi_2, maskSplit_maskSelect_lo_lo_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_hi_2 = {maskSplit_maskSelect_lo_lo_lo_hi_hi_2, maskSplit_maskSelect_lo_lo_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_lo_lo_2 = {maskSplit_maskSelect_lo_lo_lo_hi_2, maskSplit_maskSelect_lo_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_lo_2 = {maskSplit_maskSelect_lo_lo_hi_lo_hi_2, maskSplit_maskSelect_lo_lo_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_hi_2 = {maskSplit_maskSelect_lo_lo_hi_hi_hi_2, maskSplit_maskSelect_lo_lo_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_lo_hi_2 = {maskSplit_maskSelect_lo_lo_hi_hi_2, maskSplit_maskSelect_lo_lo_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_lo_lo_2 = {maskSplit_maskSelect_lo_lo_hi_2, maskSplit_maskSelect_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_lo_2 = {maskSplit_maskSelect_lo_hi_lo_lo_hi_2, maskSplit_maskSelect_lo_hi_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_hi_2 = {maskSplit_maskSelect_lo_hi_lo_hi_hi_2, maskSplit_maskSelect_lo_hi_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_hi_lo_2 = {maskSplit_maskSelect_lo_hi_lo_hi_2, maskSplit_maskSelect_lo_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_lo_2 = {maskSplit_maskSelect_lo_hi_hi_lo_hi_2, maskSplit_maskSelect_lo_hi_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_hi_2 = {maskSplit_maskSelect_lo_hi_hi_hi_hi_2, maskSplit_maskSelect_lo_hi_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_hi_hi_2 = {maskSplit_maskSelect_lo_hi_hi_hi_2, maskSplit_maskSelect_lo_hi_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_lo_hi_2 = {maskSplit_maskSelect_lo_hi_hi_2, maskSplit_maskSelect_lo_hi_lo_2};
  wire [1023:0]      maskSplit_maskSelect_lo_2 = {maskSplit_maskSelect_lo_hi_2, maskSplit_maskSelect_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_lo_2 = {maskSplit_maskSelect_hi_lo_lo_lo_hi_2, maskSplit_maskSelect_hi_lo_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_hi_2 = {maskSplit_maskSelect_hi_lo_lo_hi_hi_2, maskSplit_maskSelect_hi_lo_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_lo_lo_2 = {maskSplit_maskSelect_hi_lo_lo_hi_2, maskSplit_maskSelect_hi_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_lo_2 = {maskSplit_maskSelect_hi_lo_hi_lo_hi_2, maskSplit_maskSelect_hi_lo_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_hi_2 = {maskSplit_maskSelect_hi_lo_hi_hi_hi_2, maskSplit_maskSelect_hi_lo_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_lo_hi_2 = {maskSplit_maskSelect_hi_lo_hi_hi_2, maskSplit_maskSelect_hi_lo_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_hi_lo_2 = {maskSplit_maskSelect_hi_lo_hi_2, maskSplit_maskSelect_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_lo_2 = {maskSplit_maskSelect_hi_hi_lo_lo_hi_2, maskSplit_maskSelect_hi_hi_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_hi_2 = {maskSplit_maskSelect_hi_hi_lo_hi_hi_2, maskSplit_maskSelect_hi_hi_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_hi_lo_2 = {maskSplit_maskSelect_hi_hi_lo_hi_2, maskSplit_maskSelect_hi_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_lo_2 = {maskSplit_maskSelect_hi_hi_hi_lo_hi_2, maskSplit_maskSelect_hi_hi_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_hi_2 = {maskSplit_maskSelect_hi_hi_hi_hi_hi_2, maskSplit_maskSelect_hi_hi_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_hi_hi_2 = {maskSplit_maskSelect_hi_hi_hi_hi_2, maskSplit_maskSelect_hi_hi_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_hi_hi_2 = {maskSplit_maskSelect_hi_hi_hi_2, maskSplit_maskSelect_hi_hi_lo_2};
  wire [1023:0]      maskSplit_maskSelect_hi_2 = {maskSplit_maskSelect_hi_hi_2, maskSplit_maskSelect_hi_lo_2};
  wire               maskSplit_vlMisAlign_2;
  assign maskSplit_vlMisAlign_2 = |(instReg_vl[4:0]);
  wire [6:0]         maskSplit_lastexecuteGroup_2 = instReg_vl[11:5] - {6'h0, ~maskSplit_vlMisAlign_2};
  wire [6:0]         _GEN_70 = {2'h0, executeGroupCounter};
  wire               maskSplit_isVlBoundary_2 = _GEN_70 == maskSplit_lastexecuteGroup_2;
  wire               maskSplit_validExecuteGroup_2 = _GEN_70 <= maskSplit_lastexecuteGroup_2;
  wire [31:0]        _maskSplit_vlBoundaryCorrection_T_58 = _maskSplit_vlBoundaryCorrection_T_55 | {_maskSplit_vlBoundaryCorrection_T_55[30:0], 1'h0};
  wire [31:0]        _maskSplit_vlBoundaryCorrection_T_61 = _maskSplit_vlBoundaryCorrection_T_58 | {_maskSplit_vlBoundaryCorrection_T_58[29:0], 2'h0};
  wire [31:0]        _maskSplit_vlBoundaryCorrection_T_64 = _maskSplit_vlBoundaryCorrection_T_61 | {_maskSplit_vlBoundaryCorrection_T_61[27:0], 4'h0};
  wire [31:0]        _maskSplit_vlBoundaryCorrection_T_67 = _maskSplit_vlBoundaryCorrection_T_64 | {_maskSplit_vlBoundaryCorrection_T_64[23:0], 8'h0};
  wire [31:0]        maskSplit_vlBoundaryCorrection_2 =
    ~({32{maskSplit_vlMisAlign_2 & maskSplit_isVlBoundary_2}} & (_maskSplit_vlBoundaryCorrection_T_67 | {_maskSplit_vlBoundaryCorrection_T_67[15:0], 16'h0})) & {32{maskSplit_validExecuteGroup_2}};
  wire [31:0][31:0]  _GEN_71 =
    {{maskSplit_maskSelect_lo_2[1023:992]},
     {maskSplit_maskSelect_lo_2[991:960]},
     {maskSplit_maskSelect_lo_2[959:928]},
     {maskSplit_maskSelect_lo_2[927:896]},
     {maskSplit_maskSelect_lo_2[895:864]},
     {maskSplit_maskSelect_lo_2[863:832]},
     {maskSplit_maskSelect_lo_2[831:800]},
     {maskSplit_maskSelect_lo_2[799:768]},
     {maskSplit_maskSelect_lo_2[767:736]},
     {maskSplit_maskSelect_lo_2[735:704]},
     {maskSplit_maskSelect_lo_2[703:672]},
     {maskSplit_maskSelect_lo_2[671:640]},
     {maskSplit_maskSelect_lo_2[639:608]},
     {maskSplit_maskSelect_lo_2[607:576]},
     {maskSplit_maskSelect_lo_2[575:544]},
     {maskSplit_maskSelect_lo_2[543:512]},
     {maskSplit_maskSelect_lo_2[511:480]},
     {maskSplit_maskSelect_lo_2[479:448]},
     {maskSplit_maskSelect_lo_2[447:416]},
     {maskSplit_maskSelect_lo_2[415:384]},
     {maskSplit_maskSelect_lo_2[383:352]},
     {maskSplit_maskSelect_lo_2[351:320]},
     {maskSplit_maskSelect_lo_2[319:288]},
     {maskSplit_maskSelect_lo_2[287:256]},
     {maskSplit_maskSelect_lo_2[255:224]},
     {maskSplit_maskSelect_lo_2[223:192]},
     {maskSplit_maskSelect_lo_2[191:160]},
     {maskSplit_maskSelect_lo_2[159:128]},
     {maskSplit_maskSelect_lo_2[127:96]},
     {maskSplit_maskSelect_lo_2[95:64]},
     {maskSplit_maskSelect_lo_2[63:32]},
     {maskSplit_maskSelect_lo_2[31:0]}};
  wire [31:0]        maskSplit_2_2 = (instReg_maskType ? _GEN_71[executeGroupCounter] : 32'hFFFFFFFF) & maskSplit_vlBoundaryCorrection_2;
  wire [7:0]         maskSplit_byteMask_lo_lo_lo_lo_2 = {{4{maskSplit_2_2[1]}}, {4{maskSplit_2_2[0]}}};
  wire [7:0]         maskSplit_byteMask_lo_lo_lo_hi_2 = {{4{maskSplit_2_2[3]}}, {4{maskSplit_2_2[2]}}};
  wire [15:0]        maskSplit_byteMask_lo_lo_lo_2 = {maskSplit_byteMask_lo_lo_lo_hi_2, maskSplit_byteMask_lo_lo_lo_lo_2};
  wire [7:0]         maskSplit_byteMask_lo_lo_hi_lo_2 = {{4{maskSplit_2_2[5]}}, {4{maskSplit_2_2[4]}}};
  wire [7:0]         maskSplit_byteMask_lo_lo_hi_hi_2 = {{4{maskSplit_2_2[7]}}, {4{maskSplit_2_2[6]}}};
  wire [15:0]        maskSplit_byteMask_lo_lo_hi_2 = {maskSplit_byteMask_lo_lo_hi_hi_2, maskSplit_byteMask_lo_lo_hi_lo_2};
  wire [31:0]        maskSplit_byteMask_lo_lo_2 = {maskSplit_byteMask_lo_lo_hi_2, maskSplit_byteMask_lo_lo_lo_2};
  wire [7:0]         maskSplit_byteMask_lo_hi_lo_lo_2 = {{4{maskSplit_2_2[9]}}, {4{maskSplit_2_2[8]}}};
  wire [7:0]         maskSplit_byteMask_lo_hi_lo_hi_2 = {{4{maskSplit_2_2[11]}}, {4{maskSplit_2_2[10]}}};
  wire [15:0]        maskSplit_byteMask_lo_hi_lo_2 = {maskSplit_byteMask_lo_hi_lo_hi_2, maskSplit_byteMask_lo_hi_lo_lo_2};
  wire [7:0]         maskSplit_byteMask_lo_hi_hi_lo_2 = {{4{maskSplit_2_2[13]}}, {4{maskSplit_2_2[12]}}};
  wire [7:0]         maskSplit_byteMask_lo_hi_hi_hi_2 = {{4{maskSplit_2_2[15]}}, {4{maskSplit_2_2[14]}}};
  wire [15:0]        maskSplit_byteMask_lo_hi_hi_2 = {maskSplit_byteMask_lo_hi_hi_hi_2, maskSplit_byteMask_lo_hi_hi_lo_2};
  wire [31:0]        maskSplit_byteMask_lo_hi_2 = {maskSplit_byteMask_lo_hi_hi_2, maskSplit_byteMask_lo_hi_lo_2};
  wire [63:0]        maskSplit_byteMask_lo_2 = {maskSplit_byteMask_lo_hi_2, maskSplit_byteMask_lo_lo_2};
  wire [7:0]         maskSplit_byteMask_hi_lo_lo_lo_2 = {{4{maskSplit_2_2[17]}}, {4{maskSplit_2_2[16]}}};
  wire [7:0]         maskSplit_byteMask_hi_lo_lo_hi_2 = {{4{maskSplit_2_2[19]}}, {4{maskSplit_2_2[18]}}};
  wire [15:0]        maskSplit_byteMask_hi_lo_lo_2 = {maskSplit_byteMask_hi_lo_lo_hi_2, maskSplit_byteMask_hi_lo_lo_lo_2};
  wire [7:0]         maskSplit_byteMask_hi_lo_hi_lo_2 = {{4{maskSplit_2_2[21]}}, {4{maskSplit_2_2[20]}}};
  wire [7:0]         maskSplit_byteMask_hi_lo_hi_hi_2 = {{4{maskSplit_2_2[23]}}, {4{maskSplit_2_2[22]}}};
  wire [15:0]        maskSplit_byteMask_hi_lo_hi_2 = {maskSplit_byteMask_hi_lo_hi_hi_2, maskSplit_byteMask_hi_lo_hi_lo_2};
  wire [31:0]        maskSplit_byteMask_hi_lo_2 = {maskSplit_byteMask_hi_lo_hi_2, maskSplit_byteMask_hi_lo_lo_2};
  wire [7:0]         maskSplit_byteMask_hi_hi_lo_lo_2 = {{4{maskSplit_2_2[25]}}, {4{maskSplit_2_2[24]}}};
  wire [7:0]         maskSplit_byteMask_hi_hi_lo_hi_2 = {{4{maskSplit_2_2[27]}}, {4{maskSplit_2_2[26]}}};
  wire [15:0]        maskSplit_byteMask_hi_hi_lo_2 = {maskSplit_byteMask_hi_hi_lo_hi_2, maskSplit_byteMask_hi_hi_lo_lo_2};
  wire [7:0]         maskSplit_byteMask_hi_hi_hi_lo_2 = {{4{maskSplit_2_2[29]}}, {4{maskSplit_2_2[28]}}};
  wire [7:0]         maskSplit_byteMask_hi_hi_hi_hi_2 = {{4{maskSplit_2_2[31]}}, {4{maskSplit_2_2[30]}}};
  wire [15:0]        maskSplit_byteMask_hi_hi_hi_2 = {maskSplit_byteMask_hi_hi_hi_hi_2, maskSplit_byteMask_hi_hi_hi_lo_2};
  wire [31:0]        maskSplit_byteMask_hi_hi_2 = {maskSplit_byteMask_hi_hi_hi_2, maskSplit_byteMask_hi_hi_lo_2};
  wire [63:0]        maskSplit_byteMask_hi_2 = {maskSplit_byteMask_hi_hi_2, maskSplit_byteMask_hi_lo_2};
  wire [127:0]       maskSplit_2_1 = {maskSplit_byteMask_hi_2, maskSplit_byteMask_lo_2};
  wire [127:0]       executeByteMask = (sew1H[0] ? maskSplit_0_1 : 128'h0) | (sew1H[1] ? maskSplit_1_1 : 128'h0) | (sew1H[2] ? maskSplit_2_1 : 128'h0);
  wire [127:0]       _executeElementMask_T_3 = sew1H[0] ? maskSplit_0_2 : 128'h0;
  wire [63:0]        _GEN_72 = _executeElementMask_T_3[63:0] | (sew1H[1] ? maskSplit_1_2 : 64'h0);
  wire [127:0]       executeElementMask = {_executeElementMask_T_3[127:64], _GEN_72[63:32], _GEN_72[31:0] | (sew1H[2] ? maskSplit_2_2 : 32'h0)};
  wire [127:0]       maskForDestination_lo_lo_lo_lo = {maskForDestination_lo_lo_lo_lo_hi, maskForDestination_lo_lo_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_lo_lo_hi = {maskForDestination_lo_lo_lo_hi_hi, maskForDestination_lo_lo_lo_hi_lo};
  wire [255:0]       maskForDestination_lo_lo_lo = {maskForDestination_lo_lo_lo_hi, maskForDestination_lo_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_lo_hi_lo = {maskForDestination_lo_lo_hi_lo_hi, maskForDestination_lo_lo_hi_lo_lo};
  wire [127:0]       maskForDestination_lo_lo_hi_hi = {maskForDestination_lo_lo_hi_hi_hi, maskForDestination_lo_lo_hi_hi_lo};
  wire [255:0]       maskForDestination_lo_lo_hi = {maskForDestination_lo_lo_hi_hi, maskForDestination_lo_lo_hi_lo};
  wire [511:0]       maskForDestination_lo_lo = {maskForDestination_lo_lo_hi, maskForDestination_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_lo_lo = {maskForDestination_lo_hi_lo_lo_hi, maskForDestination_lo_hi_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_lo_hi = {maskForDestination_lo_hi_lo_hi_hi, maskForDestination_lo_hi_lo_hi_lo};
  wire [255:0]       maskForDestination_lo_hi_lo = {maskForDestination_lo_hi_lo_hi, maskForDestination_lo_hi_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_hi_lo = {maskForDestination_lo_hi_hi_lo_hi, maskForDestination_lo_hi_hi_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_hi_hi = {maskForDestination_lo_hi_hi_hi_hi, maskForDestination_lo_hi_hi_hi_lo};
  wire [255:0]       maskForDestination_lo_hi_hi = {maskForDestination_lo_hi_hi_hi, maskForDestination_lo_hi_hi_lo};
  wire [511:0]       maskForDestination_lo_hi = {maskForDestination_lo_hi_hi, maskForDestination_lo_hi_lo};
  wire [1023:0]      maskForDestination_lo = {maskForDestination_lo_hi, maskForDestination_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_lo_lo = {maskForDestination_hi_lo_lo_lo_hi, maskForDestination_hi_lo_lo_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_lo_hi = {maskForDestination_hi_lo_lo_hi_hi, maskForDestination_hi_lo_lo_hi_lo};
  wire [255:0]       maskForDestination_hi_lo_lo = {maskForDestination_hi_lo_lo_hi, maskForDestination_hi_lo_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_hi_lo = {maskForDestination_hi_lo_hi_lo_hi, maskForDestination_hi_lo_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_hi_hi = {maskForDestination_hi_lo_hi_hi_hi, maskForDestination_hi_lo_hi_hi_lo};
  wire [255:0]       maskForDestination_hi_lo_hi = {maskForDestination_hi_lo_hi_hi, maskForDestination_hi_lo_hi_lo};
  wire [511:0]       maskForDestination_hi_lo = {maskForDestination_hi_lo_hi, maskForDestination_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_lo_lo = {maskForDestination_hi_hi_lo_lo_hi, maskForDestination_hi_hi_lo_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_lo_hi = {maskForDestination_hi_hi_lo_hi_hi, maskForDestination_hi_hi_lo_hi_lo};
  wire [255:0]       maskForDestination_hi_hi_lo = {maskForDestination_hi_hi_lo_hi, maskForDestination_hi_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_hi_lo = {maskForDestination_hi_hi_hi_lo_hi, maskForDestination_hi_hi_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_hi_hi = {maskForDestination_hi_hi_hi_hi_hi, maskForDestination_hi_hi_hi_hi_lo};
  wire [255:0]       maskForDestination_hi_hi_hi = {maskForDestination_hi_hi_hi_hi, maskForDestination_hi_hi_hi_lo};
  wire [511:0]       maskForDestination_hi_hi = {maskForDestination_hi_hi_hi, maskForDestination_hi_hi_lo};
  wire [1023:0]      maskForDestination_hi = {maskForDestination_hi_hi, maskForDestination_hi_lo};
  wire [1023:0]      _lastGroupMask_T = 1024'h1 << elementTailForMaskDestination;
  wire [1022:0]      _GEN_73 = _lastGroupMask_T[1022:0] | _lastGroupMask_T[1023:1];
  wire [1021:0]      _GEN_74 = _GEN_73[1021:0] | {_lastGroupMask_T[1023], _GEN_73[1022:2]};
  wire [1019:0]      _GEN_75 = _GEN_74[1019:0] | {_lastGroupMask_T[1023], _GEN_73[1022], _GEN_74[1021:4]};
  wire [1015:0]      _GEN_76 = _GEN_75[1015:0] | {_lastGroupMask_T[1023], _GEN_73[1022], _GEN_74[1021:1020], _GEN_75[1019:8]};
  wire [1007:0]      _GEN_77 = _GEN_76[1007:0] | {_lastGroupMask_T[1023], _GEN_73[1022], _GEN_74[1021:1020], _GEN_75[1019:1016], _GEN_76[1015:16]};
  wire [991:0]       _GEN_78 = _GEN_77[991:0] | {_lastGroupMask_T[1023], _GEN_73[1022], _GEN_74[1021:1020], _GEN_75[1019:1016], _GEN_76[1015:1008], _GEN_77[1007:32]};
  wire [959:0]       _GEN_79 = _GEN_78[959:0] | {_lastGroupMask_T[1023], _GEN_73[1022], _GEN_74[1021:1020], _GEN_75[1019:1016], _GEN_76[1015:1008], _GEN_77[1007:992], _GEN_78[991:64]};
  wire [895:0]       _GEN_80 = _GEN_79[895:0] | {_lastGroupMask_T[1023], _GEN_73[1022], _GEN_74[1021:1020], _GEN_75[1019:1016], _GEN_76[1015:1008], _GEN_77[1007:992], _GEN_78[991:960], _GEN_79[959:128]};
  wire [767:0]       _GEN_81 = _GEN_80[767:0] | {_lastGroupMask_T[1023], _GEN_73[1022], _GEN_74[1021:1020], _GEN_75[1019:1016], _GEN_76[1015:1008], _GEN_77[1007:992], _GEN_78[991:960], _GEN_79[959:896], _GEN_80[895:256]};
  wire [1023:0]      lastGroupMask =
    {_lastGroupMask_T[1023],
     _GEN_73[1022],
     _GEN_74[1021:1020],
     _GEN_75[1019:1016],
     _GEN_76[1015:1008],
     _GEN_77[1007:992],
     _GEN_78[991:960],
     _GEN_79[959:896],
     _GEN_80[895:768],
     _GEN_81[767:512],
     _GEN_81[511:0] | {_lastGroupMask_T[1023], _GEN_73[1022], _GEN_74[1021:1020], _GEN_75[1019:1016], _GEN_76[1015:1008], _GEN_77[1007:992], _GEN_78[991:960], _GEN_79[959:896], _GEN_80[895:768], _GEN_81[767:512]}};
  wire [1023:0]      currentMaskGroupForDestination =
    (lastGroup
       ? lastGroupMask
       : 1024'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
    & (instReg_maskType & ~instReg_decodeResult_maskSource
         ? (requestCounter[0] ? maskForDestination_hi : maskForDestination_lo)
         : 1024'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF);
  wire [63:0]        _GEN_82 = {exeReqReg_1_bits_source1, exeReqReg_0_bits_source1};
  wire [63:0]        groupSourceData_lo_lo_lo_lo;
  assign groupSourceData_lo_lo_lo_lo = _GEN_82;
  wire [63:0]        source1_lo_lo_lo_lo;
  assign source1_lo_lo_lo_lo = _GEN_82;
  wire [63:0]        _GEN_83 = {exeReqReg_3_bits_source1, exeReqReg_2_bits_source1};
  wire [63:0]        groupSourceData_lo_lo_lo_hi;
  assign groupSourceData_lo_lo_lo_hi = _GEN_83;
  wire [63:0]        source1_lo_lo_lo_hi;
  assign source1_lo_lo_lo_hi = _GEN_83;
  wire [127:0]       groupSourceData_lo_lo_lo = {groupSourceData_lo_lo_lo_hi, groupSourceData_lo_lo_lo_lo};
  wire [63:0]        _GEN_84 = {exeReqReg_5_bits_source1, exeReqReg_4_bits_source1};
  wire [63:0]        groupSourceData_lo_lo_hi_lo;
  assign groupSourceData_lo_lo_hi_lo = _GEN_84;
  wire [63:0]        source1_lo_lo_hi_lo;
  assign source1_lo_lo_hi_lo = _GEN_84;
  wire [63:0]        _GEN_85 = {exeReqReg_7_bits_source1, exeReqReg_6_bits_source1};
  wire [63:0]        groupSourceData_lo_lo_hi_hi;
  assign groupSourceData_lo_lo_hi_hi = _GEN_85;
  wire [63:0]        source1_lo_lo_hi_hi;
  assign source1_lo_lo_hi_hi = _GEN_85;
  wire [127:0]       groupSourceData_lo_lo_hi = {groupSourceData_lo_lo_hi_hi, groupSourceData_lo_lo_hi_lo};
  wire [255:0]       groupSourceData_lo_lo = {groupSourceData_lo_lo_hi, groupSourceData_lo_lo_lo};
  wire [63:0]        _GEN_86 = {exeReqReg_9_bits_source1, exeReqReg_8_bits_source1};
  wire [63:0]        groupSourceData_lo_hi_lo_lo;
  assign groupSourceData_lo_hi_lo_lo = _GEN_86;
  wire [63:0]        source1_lo_hi_lo_lo;
  assign source1_lo_hi_lo_lo = _GEN_86;
  wire [63:0]        _GEN_87 = {exeReqReg_11_bits_source1, exeReqReg_10_bits_source1};
  wire [63:0]        groupSourceData_lo_hi_lo_hi;
  assign groupSourceData_lo_hi_lo_hi = _GEN_87;
  wire [63:0]        source1_lo_hi_lo_hi;
  assign source1_lo_hi_lo_hi = _GEN_87;
  wire [127:0]       groupSourceData_lo_hi_lo = {groupSourceData_lo_hi_lo_hi, groupSourceData_lo_hi_lo_lo};
  wire [63:0]        _GEN_88 = {exeReqReg_13_bits_source1, exeReqReg_12_bits_source1};
  wire [63:0]        groupSourceData_lo_hi_hi_lo;
  assign groupSourceData_lo_hi_hi_lo = _GEN_88;
  wire [63:0]        source1_lo_hi_hi_lo;
  assign source1_lo_hi_hi_lo = _GEN_88;
  wire [63:0]        _GEN_89 = {exeReqReg_15_bits_source1, exeReqReg_14_bits_source1};
  wire [63:0]        groupSourceData_lo_hi_hi_hi;
  assign groupSourceData_lo_hi_hi_hi = _GEN_89;
  wire [63:0]        source1_lo_hi_hi_hi;
  assign source1_lo_hi_hi_hi = _GEN_89;
  wire [127:0]       groupSourceData_lo_hi_hi = {groupSourceData_lo_hi_hi_hi, groupSourceData_lo_hi_hi_lo};
  wire [255:0]       groupSourceData_lo_hi = {groupSourceData_lo_hi_hi, groupSourceData_lo_hi_lo};
  wire [511:0]       groupSourceData_lo = {groupSourceData_lo_hi, groupSourceData_lo_lo};
  wire [63:0]        _GEN_90 = {exeReqReg_17_bits_source1, exeReqReg_16_bits_source1};
  wire [63:0]        groupSourceData_hi_lo_lo_lo;
  assign groupSourceData_hi_lo_lo_lo = _GEN_90;
  wire [63:0]        source1_hi_lo_lo_lo;
  assign source1_hi_lo_lo_lo = _GEN_90;
  wire [63:0]        _GEN_91 = {exeReqReg_19_bits_source1, exeReqReg_18_bits_source1};
  wire [63:0]        groupSourceData_hi_lo_lo_hi;
  assign groupSourceData_hi_lo_lo_hi = _GEN_91;
  wire [63:0]        source1_hi_lo_lo_hi;
  assign source1_hi_lo_lo_hi = _GEN_91;
  wire [127:0]       groupSourceData_hi_lo_lo = {groupSourceData_hi_lo_lo_hi, groupSourceData_hi_lo_lo_lo};
  wire [63:0]        _GEN_92 = {exeReqReg_21_bits_source1, exeReqReg_20_bits_source1};
  wire [63:0]        groupSourceData_hi_lo_hi_lo;
  assign groupSourceData_hi_lo_hi_lo = _GEN_92;
  wire [63:0]        source1_hi_lo_hi_lo;
  assign source1_hi_lo_hi_lo = _GEN_92;
  wire [63:0]        _GEN_93 = {exeReqReg_23_bits_source1, exeReqReg_22_bits_source1};
  wire [63:0]        groupSourceData_hi_lo_hi_hi;
  assign groupSourceData_hi_lo_hi_hi = _GEN_93;
  wire [63:0]        source1_hi_lo_hi_hi;
  assign source1_hi_lo_hi_hi = _GEN_93;
  wire [127:0]       groupSourceData_hi_lo_hi = {groupSourceData_hi_lo_hi_hi, groupSourceData_hi_lo_hi_lo};
  wire [255:0]       groupSourceData_hi_lo = {groupSourceData_hi_lo_hi, groupSourceData_hi_lo_lo};
  wire [63:0]        _GEN_94 = {exeReqReg_25_bits_source1, exeReqReg_24_bits_source1};
  wire [63:0]        groupSourceData_hi_hi_lo_lo;
  assign groupSourceData_hi_hi_lo_lo = _GEN_94;
  wire [63:0]        source1_hi_hi_lo_lo;
  assign source1_hi_hi_lo_lo = _GEN_94;
  wire [63:0]        _GEN_95 = {exeReqReg_27_bits_source1, exeReqReg_26_bits_source1};
  wire [63:0]        groupSourceData_hi_hi_lo_hi;
  assign groupSourceData_hi_hi_lo_hi = _GEN_95;
  wire [63:0]        source1_hi_hi_lo_hi;
  assign source1_hi_hi_lo_hi = _GEN_95;
  wire [127:0]       groupSourceData_hi_hi_lo = {groupSourceData_hi_hi_lo_hi, groupSourceData_hi_hi_lo_lo};
  wire [63:0]        _GEN_96 = {exeReqReg_29_bits_source1, exeReqReg_28_bits_source1};
  wire [63:0]        groupSourceData_hi_hi_hi_lo;
  assign groupSourceData_hi_hi_hi_lo = _GEN_96;
  wire [63:0]        source1_hi_hi_hi_lo;
  assign source1_hi_hi_hi_lo = _GEN_96;
  wire [63:0]        _GEN_97 = {exeReqReg_31_bits_source1, exeReqReg_30_bits_source1};
  wire [63:0]        groupSourceData_hi_hi_hi_hi;
  assign groupSourceData_hi_hi_hi_hi = _GEN_97;
  wire [63:0]        source1_hi_hi_hi_hi;
  assign source1_hi_hi_hi_hi = _GEN_97;
  wire [127:0]       groupSourceData_hi_hi_hi = {groupSourceData_hi_hi_hi_hi, groupSourceData_hi_hi_hi_lo};
  wire [255:0]       groupSourceData_hi_hi = {groupSourceData_hi_hi_hi, groupSourceData_hi_hi_lo};
  wire [511:0]       groupSourceData_hi = {groupSourceData_hi_hi, groupSourceData_hi_lo};
  wire [1023:0]      groupSourceData = {groupSourceData_hi, groupSourceData_lo};
  wire [1:0]         _GEN_98 = {exeReqReg_1_valid, exeReqReg_0_valid};
  wire [1:0]         groupSourceValid_lo_lo_lo_lo;
  assign groupSourceValid_lo_lo_lo_lo = _GEN_98;
  wire [1:0]         view__in_bits_validInput_lo_lo_lo_lo;
  assign view__in_bits_validInput_lo_lo_lo_lo = _GEN_98;
  wire [1:0]         view__in_bits_sourceValid_lo_lo_lo_lo;
  assign view__in_bits_sourceValid_lo_lo_lo_lo = _GEN_98;
  wire [1:0]         _GEN_99 = {exeReqReg_3_valid, exeReqReg_2_valid};
  wire [1:0]         groupSourceValid_lo_lo_lo_hi;
  assign groupSourceValid_lo_lo_lo_hi = _GEN_99;
  wire [1:0]         view__in_bits_validInput_lo_lo_lo_hi;
  assign view__in_bits_validInput_lo_lo_lo_hi = _GEN_99;
  wire [1:0]         view__in_bits_sourceValid_lo_lo_lo_hi;
  assign view__in_bits_sourceValid_lo_lo_lo_hi = _GEN_99;
  wire [3:0]         groupSourceValid_lo_lo_lo = {groupSourceValid_lo_lo_lo_hi, groupSourceValid_lo_lo_lo_lo};
  wire [1:0]         _GEN_100 = {exeReqReg_5_valid, exeReqReg_4_valid};
  wire [1:0]         groupSourceValid_lo_lo_hi_lo;
  assign groupSourceValid_lo_lo_hi_lo = _GEN_100;
  wire [1:0]         view__in_bits_validInput_lo_lo_hi_lo;
  assign view__in_bits_validInput_lo_lo_hi_lo = _GEN_100;
  wire [1:0]         view__in_bits_sourceValid_lo_lo_hi_lo;
  assign view__in_bits_sourceValid_lo_lo_hi_lo = _GEN_100;
  wire [1:0]         _GEN_101 = {exeReqReg_7_valid, exeReqReg_6_valid};
  wire [1:0]         groupSourceValid_lo_lo_hi_hi;
  assign groupSourceValid_lo_lo_hi_hi = _GEN_101;
  wire [1:0]         view__in_bits_validInput_lo_lo_hi_hi;
  assign view__in_bits_validInput_lo_lo_hi_hi = _GEN_101;
  wire [1:0]         view__in_bits_sourceValid_lo_lo_hi_hi;
  assign view__in_bits_sourceValid_lo_lo_hi_hi = _GEN_101;
  wire [3:0]         groupSourceValid_lo_lo_hi = {groupSourceValid_lo_lo_hi_hi, groupSourceValid_lo_lo_hi_lo};
  wire [7:0]         groupSourceValid_lo_lo = {groupSourceValid_lo_lo_hi, groupSourceValid_lo_lo_lo};
  wire [1:0]         _GEN_102 = {exeReqReg_9_valid, exeReqReg_8_valid};
  wire [1:0]         groupSourceValid_lo_hi_lo_lo;
  assign groupSourceValid_lo_hi_lo_lo = _GEN_102;
  wire [1:0]         view__in_bits_validInput_lo_hi_lo_lo;
  assign view__in_bits_validInput_lo_hi_lo_lo = _GEN_102;
  wire [1:0]         view__in_bits_sourceValid_lo_hi_lo_lo;
  assign view__in_bits_sourceValid_lo_hi_lo_lo = _GEN_102;
  wire [1:0]         _GEN_103 = {exeReqReg_11_valid, exeReqReg_10_valid};
  wire [1:0]         groupSourceValid_lo_hi_lo_hi;
  assign groupSourceValid_lo_hi_lo_hi = _GEN_103;
  wire [1:0]         view__in_bits_validInput_lo_hi_lo_hi;
  assign view__in_bits_validInput_lo_hi_lo_hi = _GEN_103;
  wire [1:0]         view__in_bits_sourceValid_lo_hi_lo_hi;
  assign view__in_bits_sourceValid_lo_hi_lo_hi = _GEN_103;
  wire [3:0]         groupSourceValid_lo_hi_lo = {groupSourceValid_lo_hi_lo_hi, groupSourceValid_lo_hi_lo_lo};
  wire [1:0]         _GEN_104 = {exeReqReg_13_valid, exeReqReg_12_valid};
  wire [1:0]         groupSourceValid_lo_hi_hi_lo;
  assign groupSourceValid_lo_hi_hi_lo = _GEN_104;
  wire [1:0]         view__in_bits_validInput_lo_hi_hi_lo;
  assign view__in_bits_validInput_lo_hi_hi_lo = _GEN_104;
  wire [1:0]         view__in_bits_sourceValid_lo_hi_hi_lo;
  assign view__in_bits_sourceValid_lo_hi_hi_lo = _GEN_104;
  wire [1:0]         _GEN_105 = {exeReqReg_15_valid, exeReqReg_14_valid};
  wire [1:0]         groupSourceValid_lo_hi_hi_hi;
  assign groupSourceValid_lo_hi_hi_hi = _GEN_105;
  wire [1:0]         view__in_bits_validInput_lo_hi_hi_hi;
  assign view__in_bits_validInput_lo_hi_hi_hi = _GEN_105;
  wire [1:0]         view__in_bits_sourceValid_lo_hi_hi_hi;
  assign view__in_bits_sourceValid_lo_hi_hi_hi = _GEN_105;
  wire [3:0]         groupSourceValid_lo_hi_hi = {groupSourceValid_lo_hi_hi_hi, groupSourceValid_lo_hi_hi_lo};
  wire [7:0]         groupSourceValid_lo_hi = {groupSourceValid_lo_hi_hi, groupSourceValid_lo_hi_lo};
  wire [15:0]        groupSourceValid_lo = {groupSourceValid_lo_hi, groupSourceValid_lo_lo};
  wire [1:0]         _GEN_106 = {exeReqReg_17_valid, exeReqReg_16_valid};
  wire [1:0]         groupSourceValid_hi_lo_lo_lo;
  assign groupSourceValid_hi_lo_lo_lo = _GEN_106;
  wire [1:0]         view__in_bits_validInput_hi_lo_lo_lo;
  assign view__in_bits_validInput_hi_lo_lo_lo = _GEN_106;
  wire [1:0]         view__in_bits_sourceValid_hi_lo_lo_lo;
  assign view__in_bits_sourceValid_hi_lo_lo_lo = _GEN_106;
  wire [1:0]         _GEN_107 = {exeReqReg_19_valid, exeReqReg_18_valid};
  wire [1:0]         groupSourceValid_hi_lo_lo_hi;
  assign groupSourceValid_hi_lo_lo_hi = _GEN_107;
  wire [1:0]         view__in_bits_validInput_hi_lo_lo_hi;
  assign view__in_bits_validInput_hi_lo_lo_hi = _GEN_107;
  wire [1:0]         view__in_bits_sourceValid_hi_lo_lo_hi;
  assign view__in_bits_sourceValid_hi_lo_lo_hi = _GEN_107;
  wire [3:0]         groupSourceValid_hi_lo_lo = {groupSourceValid_hi_lo_lo_hi, groupSourceValid_hi_lo_lo_lo};
  wire [1:0]         _GEN_108 = {exeReqReg_21_valid, exeReqReg_20_valid};
  wire [1:0]         groupSourceValid_hi_lo_hi_lo;
  assign groupSourceValid_hi_lo_hi_lo = _GEN_108;
  wire [1:0]         view__in_bits_validInput_hi_lo_hi_lo;
  assign view__in_bits_validInput_hi_lo_hi_lo = _GEN_108;
  wire [1:0]         view__in_bits_sourceValid_hi_lo_hi_lo;
  assign view__in_bits_sourceValid_hi_lo_hi_lo = _GEN_108;
  wire [1:0]         _GEN_109 = {exeReqReg_23_valid, exeReqReg_22_valid};
  wire [1:0]         groupSourceValid_hi_lo_hi_hi;
  assign groupSourceValid_hi_lo_hi_hi = _GEN_109;
  wire [1:0]         view__in_bits_validInput_hi_lo_hi_hi;
  assign view__in_bits_validInput_hi_lo_hi_hi = _GEN_109;
  wire [1:0]         view__in_bits_sourceValid_hi_lo_hi_hi;
  assign view__in_bits_sourceValid_hi_lo_hi_hi = _GEN_109;
  wire [3:0]         groupSourceValid_hi_lo_hi = {groupSourceValid_hi_lo_hi_hi, groupSourceValid_hi_lo_hi_lo};
  wire [7:0]         groupSourceValid_hi_lo = {groupSourceValid_hi_lo_hi, groupSourceValid_hi_lo_lo};
  wire [1:0]         _GEN_110 = {exeReqReg_25_valid, exeReqReg_24_valid};
  wire [1:0]         groupSourceValid_hi_hi_lo_lo;
  assign groupSourceValid_hi_hi_lo_lo = _GEN_110;
  wire [1:0]         view__in_bits_validInput_hi_hi_lo_lo;
  assign view__in_bits_validInput_hi_hi_lo_lo = _GEN_110;
  wire [1:0]         view__in_bits_sourceValid_hi_hi_lo_lo;
  assign view__in_bits_sourceValid_hi_hi_lo_lo = _GEN_110;
  wire [1:0]         _GEN_111 = {exeReqReg_27_valid, exeReqReg_26_valid};
  wire [1:0]         groupSourceValid_hi_hi_lo_hi;
  assign groupSourceValid_hi_hi_lo_hi = _GEN_111;
  wire [1:0]         view__in_bits_validInput_hi_hi_lo_hi;
  assign view__in_bits_validInput_hi_hi_lo_hi = _GEN_111;
  wire [1:0]         view__in_bits_sourceValid_hi_hi_lo_hi;
  assign view__in_bits_sourceValid_hi_hi_lo_hi = _GEN_111;
  wire [3:0]         groupSourceValid_hi_hi_lo = {groupSourceValid_hi_hi_lo_hi, groupSourceValid_hi_hi_lo_lo};
  wire [1:0]         _GEN_112 = {exeReqReg_29_valid, exeReqReg_28_valid};
  wire [1:0]         groupSourceValid_hi_hi_hi_lo;
  assign groupSourceValid_hi_hi_hi_lo = _GEN_112;
  wire [1:0]         view__in_bits_validInput_hi_hi_hi_lo;
  assign view__in_bits_validInput_hi_hi_hi_lo = _GEN_112;
  wire [1:0]         view__in_bits_sourceValid_hi_hi_hi_lo;
  assign view__in_bits_sourceValid_hi_hi_hi_lo = _GEN_112;
  wire [1:0]         _GEN_113 = {exeReqReg_31_valid, exeReqReg_30_valid};
  wire [1:0]         groupSourceValid_hi_hi_hi_hi;
  assign groupSourceValid_hi_hi_hi_hi = _GEN_113;
  wire [1:0]         view__in_bits_validInput_hi_hi_hi_hi;
  assign view__in_bits_validInput_hi_hi_hi_hi = _GEN_113;
  wire [1:0]         view__in_bits_sourceValid_hi_hi_hi_hi;
  assign view__in_bits_sourceValid_hi_hi_hi_hi = _GEN_113;
  wire [3:0]         groupSourceValid_hi_hi_hi = {groupSourceValid_hi_hi_hi_hi, groupSourceValid_hi_hi_hi_lo};
  wire [7:0]         groupSourceValid_hi_hi = {groupSourceValid_hi_hi_hi, groupSourceValid_hi_hi_lo};
  wire [15:0]        groupSourceValid_hi = {groupSourceValid_hi_hi, groupSourceValid_hi_lo};
  wire [31:0]        groupSourceValid = {groupSourceValid_hi, groupSourceValid_lo};
  wire [1:0]         shifterSize = (sourceDataEEW1H[0] ? executeIndex : 2'h0) | (sourceDataEEW1H[1] ? {executeIndex[1], 1'h0} : 2'h0);
  wire [3:0]         _shifterSource_T = 4'h1 << shifterSize;
  wire [1023:0]      _shifterSource_T_8 = _shifterSource_T[0] ? groupSourceData : 1024'h0;
  wire [767:0]       _GEN_114 = _shifterSource_T_8[767:0] | (_shifterSource_T[1] ? groupSourceData[1023:256] : 768'h0);
  wire [511:0]       _GEN_115 = _GEN_114[511:0] | (_shifterSource_T[2] ? groupSourceData[1023:512] : 512'h0);
  wire [1023:0]      shifterSource = {_shifterSource_T_8[1023:768], _GEN_114[767:512], _GEN_115[511:256], _GEN_115[255:0] | (_shifterSource_T[3] ? groupSourceData[1023:768] : 256'h0)};
  wire [7:0]         selectValid_lo_lo_lo_lo = {{4{groupSourceValid[1]}}, {4{groupSourceValid[0]}}};
  wire [7:0]         selectValid_lo_lo_lo_hi = {{4{groupSourceValid[3]}}, {4{groupSourceValid[2]}}};
  wire [15:0]        selectValid_lo_lo_lo = {selectValid_lo_lo_lo_hi, selectValid_lo_lo_lo_lo};
  wire [7:0]         selectValid_lo_lo_hi_lo = {{4{groupSourceValid[5]}}, {4{groupSourceValid[4]}}};
  wire [7:0]         selectValid_lo_lo_hi_hi = {{4{groupSourceValid[7]}}, {4{groupSourceValid[6]}}};
  wire [15:0]        selectValid_lo_lo_hi = {selectValid_lo_lo_hi_hi, selectValid_lo_lo_hi_lo};
  wire [31:0]        selectValid_lo_lo = {selectValid_lo_lo_hi, selectValid_lo_lo_lo};
  wire [7:0]         selectValid_lo_hi_lo_lo = {{4{groupSourceValid[9]}}, {4{groupSourceValid[8]}}};
  wire [7:0]         selectValid_lo_hi_lo_hi = {{4{groupSourceValid[11]}}, {4{groupSourceValid[10]}}};
  wire [15:0]        selectValid_lo_hi_lo = {selectValid_lo_hi_lo_hi, selectValid_lo_hi_lo_lo};
  wire [7:0]         selectValid_lo_hi_hi_lo = {{4{groupSourceValid[13]}}, {4{groupSourceValid[12]}}};
  wire [7:0]         selectValid_lo_hi_hi_hi = {{4{groupSourceValid[15]}}, {4{groupSourceValid[14]}}};
  wire [15:0]        selectValid_lo_hi_hi = {selectValid_lo_hi_hi_hi, selectValid_lo_hi_hi_lo};
  wire [31:0]        selectValid_lo_hi = {selectValid_lo_hi_hi, selectValid_lo_hi_lo};
  wire [63:0]        selectValid_lo = {selectValid_lo_hi, selectValid_lo_lo};
  wire [7:0]         selectValid_hi_lo_lo_lo = {{4{groupSourceValid[17]}}, {4{groupSourceValid[16]}}};
  wire [7:0]         selectValid_hi_lo_lo_hi = {{4{groupSourceValid[19]}}, {4{groupSourceValid[18]}}};
  wire [15:0]        selectValid_hi_lo_lo = {selectValid_hi_lo_lo_hi, selectValid_hi_lo_lo_lo};
  wire [7:0]         selectValid_hi_lo_hi_lo = {{4{groupSourceValid[21]}}, {4{groupSourceValid[20]}}};
  wire [7:0]         selectValid_hi_lo_hi_hi = {{4{groupSourceValid[23]}}, {4{groupSourceValid[22]}}};
  wire [15:0]        selectValid_hi_lo_hi = {selectValid_hi_lo_hi_hi, selectValid_hi_lo_hi_lo};
  wire [31:0]        selectValid_hi_lo = {selectValid_hi_lo_hi, selectValid_hi_lo_lo};
  wire [7:0]         selectValid_hi_hi_lo_lo = {{4{groupSourceValid[25]}}, {4{groupSourceValid[24]}}};
  wire [7:0]         selectValid_hi_hi_lo_hi = {{4{groupSourceValid[27]}}, {4{groupSourceValid[26]}}};
  wire [15:0]        selectValid_hi_hi_lo = {selectValid_hi_hi_lo_hi, selectValid_hi_hi_lo_lo};
  wire [7:0]         selectValid_hi_hi_hi_lo = {{4{groupSourceValid[29]}}, {4{groupSourceValid[28]}}};
  wire [7:0]         selectValid_hi_hi_hi_hi = {{4{groupSourceValid[31]}}, {4{groupSourceValid[30]}}};
  wire [15:0]        selectValid_hi_hi_hi = {selectValid_hi_hi_hi_hi, selectValid_hi_hi_hi_lo};
  wire [31:0]        selectValid_hi_hi = {selectValid_hi_hi_hi, selectValid_hi_hi_lo};
  wire [63:0]        selectValid_hi = {selectValid_hi_hi, selectValid_hi_lo};
  wire [3:0]         selectValid_lo_lo_lo_lo_1 = {{2{groupSourceValid[1]}}, {2{groupSourceValid[0]}}};
  wire [3:0]         selectValid_lo_lo_lo_hi_1 = {{2{groupSourceValid[3]}}, {2{groupSourceValid[2]}}};
  wire [7:0]         selectValid_lo_lo_lo_1 = {selectValid_lo_lo_lo_hi_1, selectValid_lo_lo_lo_lo_1};
  wire [3:0]         selectValid_lo_lo_hi_lo_1 = {{2{groupSourceValid[5]}}, {2{groupSourceValid[4]}}};
  wire [3:0]         selectValid_lo_lo_hi_hi_1 = {{2{groupSourceValid[7]}}, {2{groupSourceValid[6]}}};
  wire [7:0]         selectValid_lo_lo_hi_1 = {selectValid_lo_lo_hi_hi_1, selectValid_lo_lo_hi_lo_1};
  wire [15:0]        selectValid_lo_lo_1 = {selectValid_lo_lo_hi_1, selectValid_lo_lo_lo_1};
  wire [3:0]         selectValid_lo_hi_lo_lo_1 = {{2{groupSourceValid[9]}}, {2{groupSourceValid[8]}}};
  wire [3:0]         selectValid_lo_hi_lo_hi_1 = {{2{groupSourceValid[11]}}, {2{groupSourceValid[10]}}};
  wire [7:0]         selectValid_lo_hi_lo_1 = {selectValid_lo_hi_lo_hi_1, selectValid_lo_hi_lo_lo_1};
  wire [3:0]         selectValid_lo_hi_hi_lo_1 = {{2{groupSourceValid[13]}}, {2{groupSourceValid[12]}}};
  wire [3:0]         selectValid_lo_hi_hi_hi_1 = {{2{groupSourceValid[15]}}, {2{groupSourceValid[14]}}};
  wire [7:0]         selectValid_lo_hi_hi_1 = {selectValid_lo_hi_hi_hi_1, selectValid_lo_hi_hi_lo_1};
  wire [15:0]        selectValid_lo_hi_1 = {selectValid_lo_hi_hi_1, selectValid_lo_hi_lo_1};
  wire [31:0]        selectValid_lo_1 = {selectValid_lo_hi_1, selectValid_lo_lo_1};
  wire [3:0]         selectValid_hi_lo_lo_lo_1 = {{2{groupSourceValid[17]}}, {2{groupSourceValid[16]}}};
  wire [3:0]         selectValid_hi_lo_lo_hi_1 = {{2{groupSourceValid[19]}}, {2{groupSourceValid[18]}}};
  wire [7:0]         selectValid_hi_lo_lo_1 = {selectValid_hi_lo_lo_hi_1, selectValid_hi_lo_lo_lo_1};
  wire [3:0]         selectValid_hi_lo_hi_lo_1 = {{2{groupSourceValid[21]}}, {2{groupSourceValid[20]}}};
  wire [3:0]         selectValid_hi_lo_hi_hi_1 = {{2{groupSourceValid[23]}}, {2{groupSourceValid[22]}}};
  wire [7:0]         selectValid_hi_lo_hi_1 = {selectValid_hi_lo_hi_hi_1, selectValid_hi_lo_hi_lo_1};
  wire [15:0]        selectValid_hi_lo_1 = {selectValid_hi_lo_hi_1, selectValid_hi_lo_lo_1};
  wire [3:0]         selectValid_hi_hi_lo_lo_1 = {{2{groupSourceValid[25]}}, {2{groupSourceValid[24]}}};
  wire [3:0]         selectValid_hi_hi_lo_hi_1 = {{2{groupSourceValid[27]}}, {2{groupSourceValid[26]}}};
  wire [7:0]         selectValid_hi_hi_lo_1 = {selectValid_hi_hi_lo_hi_1, selectValid_hi_hi_lo_lo_1};
  wire [3:0]         selectValid_hi_hi_hi_lo_1 = {{2{groupSourceValid[29]}}, {2{groupSourceValid[28]}}};
  wire [3:0]         selectValid_hi_hi_hi_hi_1 = {{2{groupSourceValid[31]}}, {2{groupSourceValid[30]}}};
  wire [7:0]         selectValid_hi_hi_hi_1 = {selectValid_hi_hi_hi_hi_1, selectValid_hi_hi_hi_lo_1};
  wire [15:0]        selectValid_hi_hi_1 = {selectValid_hi_hi_hi_1, selectValid_hi_hi_lo_1};
  wire [31:0]        selectValid_hi_1 = {selectValid_hi_hi_1, selectValid_hi_lo_1};
  wire [3:0][31:0]   _GEN_116 = {{selectValid_hi[63:32]}, {selectValid_hi[31:0]}, {selectValid_lo[63:32]}, {selectValid_lo[31:0]}};
  wire [31:0]        selectValid = (sourceDataEEW1H[0] ? _GEN_116[executeIndex] : 32'h0) | (sourceDataEEW1H[1] ? (executeIndex[1] ? selectValid_hi_1 : selectValid_lo_1) : 32'h0) | (sourceDataEEW1H[2] ? groupSourceValid : 32'h0);
  wire [31:0]        source_0 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[7:0] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[15:0] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[31:0] : 32'h0);
  wire [31:0]        source_1 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[15:8] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[31:16] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[63:32] : 32'h0);
  wire [31:0]        source_2 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[23:16] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[47:32] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[95:64] : 32'h0);
  wire [31:0]        source_3 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[31:24] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[63:48] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[127:96] : 32'h0);
  wire [31:0]        source_4 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[39:32] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[79:64] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[159:128] : 32'h0);
  wire [31:0]        source_5 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[47:40] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[95:80] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[191:160] : 32'h0);
  wire [31:0]        source_6 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[55:48] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[111:96] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[223:192] : 32'h0);
  wire [31:0]        source_7 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[63:56] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[127:112] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[255:224] : 32'h0);
  wire [31:0]        source_8 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[71:64] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[143:128] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[287:256] : 32'h0);
  wire [31:0]        source_9 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[79:72] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[159:144] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[319:288] : 32'h0);
  wire [31:0]        source_10 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[87:80] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[175:160] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[351:320] : 32'h0);
  wire [31:0]        source_11 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[95:88] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[191:176] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[383:352] : 32'h0);
  wire [31:0]        source_12 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[103:96] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[207:192] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[415:384] : 32'h0);
  wire [31:0]        source_13 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[111:104] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[223:208] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[447:416] : 32'h0);
  wire [31:0]        source_14 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[119:112] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[239:224] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[479:448] : 32'h0);
  wire [31:0]        source_15 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[127:120] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[255:240] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[511:480] : 32'h0);
  wire [31:0]        source_16 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[135:128] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[271:256] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[543:512] : 32'h0);
  wire [31:0]        source_17 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[143:136] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[287:272] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[575:544] : 32'h0);
  wire [31:0]        source_18 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[151:144] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[303:288] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[607:576] : 32'h0);
  wire [31:0]        source_19 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[159:152] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[319:304] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[639:608] : 32'h0);
  wire [31:0]        source_20 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[167:160] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[335:320] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[671:640] : 32'h0);
  wire [31:0]        source_21 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[175:168] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[351:336] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[703:672] : 32'h0);
  wire [31:0]        source_22 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[183:176] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[367:352] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[735:704] : 32'h0);
  wire [31:0]        source_23 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[191:184] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[383:368] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[767:736] : 32'h0);
  wire [31:0]        source_24 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[199:192] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[399:384] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[799:768] : 32'h0);
  wire [31:0]        source_25 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[207:200] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[415:400] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[831:800] : 32'h0);
  wire [31:0]        source_26 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[215:208] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[431:416] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[863:832] : 32'h0);
  wire [31:0]        source_27 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[223:216] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[447:432] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[895:864] : 32'h0);
  wire [31:0]        source_28 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[231:224] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[463:448] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[927:896] : 32'h0);
  wire [31:0]        source_29 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[239:232] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[479:464] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[959:928] : 32'h0);
  wire [31:0]        source_30 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[247:240] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[495:480] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[991:960] : 32'h0);
  wire [31:0]        source_31 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[255:248] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[511:496] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[1023:992] : 32'h0);
  wire [31:0]        _GEN_117 = selectValid & readMaskCorrection;
  wire [31:0]        checkVec_validVec;
  assign checkVec_validVec = _GEN_117;
  wire [31:0]        checkVec_validVec_1;
  assign checkVec_validVec_1 = _GEN_117;
  wire [31:0]        checkVec_validVec_2;
  assign checkVec_validVec_2 = _GEN_117;
  wire               checkVec_checkResultVec_0_6 = checkVec_validVec[0];
  wire [3:0]         _GEN_118 = 4'h1 << instReg_vlmul[1:0];
  wire [3:0]         checkVec_checkResultVec_intLMULInput;
  assign checkVec_checkResultVec_intLMULInput = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_1;
  assign checkVec_checkResultVec_intLMULInput_1 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_2;
  assign checkVec_checkResultVec_intLMULInput_2 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_3;
  assign checkVec_checkResultVec_intLMULInput_3 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_4;
  assign checkVec_checkResultVec_intLMULInput_4 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_5;
  assign checkVec_checkResultVec_intLMULInput_5 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_6;
  assign checkVec_checkResultVec_intLMULInput_6 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_7;
  assign checkVec_checkResultVec_intLMULInput_7 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_8;
  assign checkVec_checkResultVec_intLMULInput_8 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_9;
  assign checkVec_checkResultVec_intLMULInput_9 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_10;
  assign checkVec_checkResultVec_intLMULInput_10 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_11;
  assign checkVec_checkResultVec_intLMULInput_11 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_12;
  assign checkVec_checkResultVec_intLMULInput_12 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_13;
  assign checkVec_checkResultVec_intLMULInput_13 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_14;
  assign checkVec_checkResultVec_intLMULInput_14 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_15;
  assign checkVec_checkResultVec_intLMULInput_15 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_16;
  assign checkVec_checkResultVec_intLMULInput_16 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_17;
  assign checkVec_checkResultVec_intLMULInput_17 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_18;
  assign checkVec_checkResultVec_intLMULInput_18 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_19;
  assign checkVec_checkResultVec_intLMULInput_19 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_20;
  assign checkVec_checkResultVec_intLMULInput_20 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_21;
  assign checkVec_checkResultVec_intLMULInput_21 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_22;
  assign checkVec_checkResultVec_intLMULInput_22 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_23;
  assign checkVec_checkResultVec_intLMULInput_23 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_24;
  assign checkVec_checkResultVec_intLMULInput_24 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_25;
  assign checkVec_checkResultVec_intLMULInput_25 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_26;
  assign checkVec_checkResultVec_intLMULInput_26 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_27;
  assign checkVec_checkResultVec_intLMULInput_27 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_28;
  assign checkVec_checkResultVec_intLMULInput_28 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_29;
  assign checkVec_checkResultVec_intLMULInput_29 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_30;
  assign checkVec_checkResultVec_intLMULInput_30 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_31;
  assign checkVec_checkResultVec_intLMULInput_31 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_32;
  assign checkVec_checkResultVec_intLMULInput_32 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_33;
  assign checkVec_checkResultVec_intLMULInput_33 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_34;
  assign checkVec_checkResultVec_intLMULInput_34 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_35;
  assign checkVec_checkResultVec_intLMULInput_35 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_36;
  assign checkVec_checkResultVec_intLMULInput_36 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_37;
  assign checkVec_checkResultVec_intLMULInput_37 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_38;
  assign checkVec_checkResultVec_intLMULInput_38 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_39;
  assign checkVec_checkResultVec_intLMULInput_39 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_40;
  assign checkVec_checkResultVec_intLMULInput_40 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_41;
  assign checkVec_checkResultVec_intLMULInput_41 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_42;
  assign checkVec_checkResultVec_intLMULInput_42 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_43;
  assign checkVec_checkResultVec_intLMULInput_43 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_44;
  assign checkVec_checkResultVec_intLMULInput_44 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_45;
  assign checkVec_checkResultVec_intLMULInput_45 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_46;
  assign checkVec_checkResultVec_intLMULInput_46 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_47;
  assign checkVec_checkResultVec_intLMULInput_47 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_48;
  assign checkVec_checkResultVec_intLMULInput_48 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_49;
  assign checkVec_checkResultVec_intLMULInput_49 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_50;
  assign checkVec_checkResultVec_intLMULInput_50 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_51;
  assign checkVec_checkResultVec_intLMULInput_51 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_52;
  assign checkVec_checkResultVec_intLMULInput_52 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_53;
  assign checkVec_checkResultVec_intLMULInput_53 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_54;
  assign checkVec_checkResultVec_intLMULInput_54 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_55;
  assign checkVec_checkResultVec_intLMULInput_55 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_56;
  assign checkVec_checkResultVec_intLMULInput_56 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_57;
  assign checkVec_checkResultVec_intLMULInput_57 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_58;
  assign checkVec_checkResultVec_intLMULInput_58 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_59;
  assign checkVec_checkResultVec_intLMULInput_59 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_60;
  assign checkVec_checkResultVec_intLMULInput_60 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_61;
  assign checkVec_checkResultVec_intLMULInput_61 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_62;
  assign checkVec_checkResultVec_intLMULInput_62 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_63;
  assign checkVec_checkResultVec_intLMULInput_63 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_64;
  assign checkVec_checkResultVec_intLMULInput_64 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_65;
  assign checkVec_checkResultVec_intLMULInput_65 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_66;
  assign checkVec_checkResultVec_intLMULInput_66 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_67;
  assign checkVec_checkResultVec_intLMULInput_67 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_68;
  assign checkVec_checkResultVec_intLMULInput_68 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_69;
  assign checkVec_checkResultVec_intLMULInput_69 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_70;
  assign checkVec_checkResultVec_intLMULInput_70 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_71;
  assign checkVec_checkResultVec_intLMULInput_71 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_72;
  assign checkVec_checkResultVec_intLMULInput_72 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_73;
  assign checkVec_checkResultVec_intLMULInput_73 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_74;
  assign checkVec_checkResultVec_intLMULInput_74 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_75;
  assign checkVec_checkResultVec_intLMULInput_75 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_76;
  assign checkVec_checkResultVec_intLMULInput_76 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_77;
  assign checkVec_checkResultVec_intLMULInput_77 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_78;
  assign checkVec_checkResultVec_intLMULInput_78 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_79;
  assign checkVec_checkResultVec_intLMULInput_79 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_80;
  assign checkVec_checkResultVec_intLMULInput_80 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_81;
  assign checkVec_checkResultVec_intLMULInput_81 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_82;
  assign checkVec_checkResultVec_intLMULInput_82 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_83;
  assign checkVec_checkResultVec_intLMULInput_83 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_84;
  assign checkVec_checkResultVec_intLMULInput_84 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_85;
  assign checkVec_checkResultVec_intLMULInput_85 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_86;
  assign checkVec_checkResultVec_intLMULInput_86 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_87;
  assign checkVec_checkResultVec_intLMULInput_87 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_88;
  assign checkVec_checkResultVec_intLMULInput_88 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_89;
  assign checkVec_checkResultVec_intLMULInput_89 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_90;
  assign checkVec_checkResultVec_intLMULInput_90 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_91;
  assign checkVec_checkResultVec_intLMULInput_91 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_92;
  assign checkVec_checkResultVec_intLMULInput_92 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_93;
  assign checkVec_checkResultVec_intLMULInput_93 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_94;
  assign checkVec_checkResultVec_intLMULInput_94 = _GEN_118;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_95;
  assign checkVec_checkResultVec_intLMULInput_95 = _GEN_118;
  wire [10:0]        checkVec_checkResultVec_dataPosition = source_0[10:0];
  wire [3:0]         checkVec_checkResultVec_0_0 = 4'h1 << checkVec_checkResultVec_dataPosition[1:0];
  wire [1:0]         checkVec_checkResultVec_0_1 = checkVec_checkResultVec_dataPosition[1:0];
  wire [4:0]         checkVec_checkResultVec_0_2 = checkVec_checkResultVec_dataPosition[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup = checkVec_checkResultVec_dataPosition[10:7];
  wire               checkVec_checkResultVec_0_3 = checkVec_checkResultVec_dataGroup[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth = checkVec_checkResultVec_dataGroup[3:1];
  wire [2:0]         checkVec_checkResultVec_0_4 = checkVec_checkResultVec_accessRegGrowth;
  wire [5:0]         checkVec_checkResultVec_decimalProportion = {checkVec_checkResultVec_0_3, checkVec_checkResultVec_0_2};
  wire [2:0]         checkVec_checkResultVec_decimal = checkVec_checkResultVec_decimalProportion[5:3];
  wire               checkVec_checkResultVec_overlap =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal >= checkVec_checkResultVec_intLMULInput[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth} >= checkVec_checkResultVec_intLMULInput, source_0[31:11]};
  wire               checkVec_checkResultVec_0_5 = checkVec_checkResultVec_overlap | ~checkVec_checkResultVec_0_6;
  wire               checkVec_checkResultVec_1_6 = checkVec_validVec[1];
  wire [10:0]        checkVec_checkResultVec_dataPosition_1 = source_1[10:0];
  wire [3:0]         checkVec_checkResultVec_1_0 = 4'h1 << checkVec_checkResultVec_dataPosition_1[1:0];
  wire [1:0]         checkVec_checkResultVec_1_1 = checkVec_checkResultVec_dataPosition_1[1:0];
  wire [4:0]         checkVec_checkResultVec_1_2 = checkVec_checkResultVec_dataPosition_1[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_1 = checkVec_checkResultVec_dataPosition_1[10:7];
  wire               checkVec_checkResultVec_1_3 = checkVec_checkResultVec_dataGroup_1[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_1 = checkVec_checkResultVec_dataGroup_1[3:1];
  wire [2:0]         checkVec_checkResultVec_1_4 = checkVec_checkResultVec_accessRegGrowth_1;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_1 = {checkVec_checkResultVec_1_3, checkVec_checkResultVec_1_2};
  wire [2:0]         checkVec_checkResultVec_decimal_1 = checkVec_checkResultVec_decimalProportion_1[5:3];
  wire               checkVec_checkResultVec_overlap_1 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_1 >= checkVec_checkResultVec_intLMULInput_1[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_1} >= checkVec_checkResultVec_intLMULInput_1, source_1[31:11]};
  wire               checkVec_checkResultVec_1_5 = checkVec_checkResultVec_overlap_1 | ~checkVec_checkResultVec_1_6;
  wire               checkVec_checkResultVec_2_6 = checkVec_validVec[2];
  wire [10:0]        checkVec_checkResultVec_dataPosition_2 = source_2[10:0];
  wire [3:0]         checkVec_checkResultVec_2_0 = 4'h1 << checkVec_checkResultVec_dataPosition_2[1:0];
  wire [1:0]         checkVec_checkResultVec_2_1 = checkVec_checkResultVec_dataPosition_2[1:0];
  wire [4:0]         checkVec_checkResultVec_2_2 = checkVec_checkResultVec_dataPosition_2[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_2 = checkVec_checkResultVec_dataPosition_2[10:7];
  wire               checkVec_checkResultVec_2_3 = checkVec_checkResultVec_dataGroup_2[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_2 = checkVec_checkResultVec_dataGroup_2[3:1];
  wire [2:0]         checkVec_checkResultVec_2_4 = checkVec_checkResultVec_accessRegGrowth_2;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_2 = {checkVec_checkResultVec_2_3, checkVec_checkResultVec_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_2 = checkVec_checkResultVec_decimalProportion_2[5:3];
  wire               checkVec_checkResultVec_overlap_2 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_2 >= checkVec_checkResultVec_intLMULInput_2[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_2} >= checkVec_checkResultVec_intLMULInput_2, source_2[31:11]};
  wire               checkVec_checkResultVec_2_5 = checkVec_checkResultVec_overlap_2 | ~checkVec_checkResultVec_2_6;
  wire               checkVec_checkResultVec_3_6 = checkVec_validVec[3];
  wire [10:0]        checkVec_checkResultVec_dataPosition_3 = source_3[10:0];
  wire [3:0]         checkVec_checkResultVec_3_0 = 4'h1 << checkVec_checkResultVec_dataPosition_3[1:0];
  wire [1:0]         checkVec_checkResultVec_3_1 = checkVec_checkResultVec_dataPosition_3[1:0];
  wire [4:0]         checkVec_checkResultVec_3_2 = checkVec_checkResultVec_dataPosition_3[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_3 = checkVec_checkResultVec_dataPosition_3[10:7];
  wire               checkVec_checkResultVec_3_3 = checkVec_checkResultVec_dataGroup_3[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_3 = checkVec_checkResultVec_dataGroup_3[3:1];
  wire [2:0]         checkVec_checkResultVec_3_4 = checkVec_checkResultVec_accessRegGrowth_3;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_3 = {checkVec_checkResultVec_3_3, checkVec_checkResultVec_3_2};
  wire [2:0]         checkVec_checkResultVec_decimal_3 = checkVec_checkResultVec_decimalProportion_3[5:3];
  wire               checkVec_checkResultVec_overlap_3 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_3 >= checkVec_checkResultVec_intLMULInput_3[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_3} >= checkVec_checkResultVec_intLMULInput_3, source_3[31:11]};
  wire               checkVec_checkResultVec_3_5 = checkVec_checkResultVec_overlap_3 | ~checkVec_checkResultVec_3_6;
  wire               checkVec_checkResultVec_4_6 = checkVec_validVec[4];
  wire [10:0]        checkVec_checkResultVec_dataPosition_4 = source_4[10:0];
  wire [3:0]         checkVec_checkResultVec_4_0 = 4'h1 << checkVec_checkResultVec_dataPosition_4[1:0];
  wire [1:0]         checkVec_checkResultVec_4_1 = checkVec_checkResultVec_dataPosition_4[1:0];
  wire [4:0]         checkVec_checkResultVec_4_2 = checkVec_checkResultVec_dataPosition_4[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_4 = checkVec_checkResultVec_dataPosition_4[10:7];
  wire               checkVec_checkResultVec_4_3 = checkVec_checkResultVec_dataGroup_4[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_4 = checkVec_checkResultVec_dataGroup_4[3:1];
  wire [2:0]         checkVec_checkResultVec_4_4 = checkVec_checkResultVec_accessRegGrowth_4;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_4 = {checkVec_checkResultVec_4_3, checkVec_checkResultVec_4_2};
  wire [2:0]         checkVec_checkResultVec_decimal_4 = checkVec_checkResultVec_decimalProportion_4[5:3];
  wire               checkVec_checkResultVec_overlap_4 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_4 >= checkVec_checkResultVec_intLMULInput_4[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_4} >= checkVec_checkResultVec_intLMULInput_4, source_4[31:11]};
  wire               checkVec_checkResultVec_4_5 = checkVec_checkResultVec_overlap_4 | ~checkVec_checkResultVec_4_6;
  wire               checkVec_checkResultVec_5_6 = checkVec_validVec[5];
  wire [10:0]        checkVec_checkResultVec_dataPosition_5 = source_5[10:0];
  wire [3:0]         checkVec_checkResultVec_5_0 = 4'h1 << checkVec_checkResultVec_dataPosition_5[1:0];
  wire [1:0]         checkVec_checkResultVec_5_1 = checkVec_checkResultVec_dataPosition_5[1:0];
  wire [4:0]         checkVec_checkResultVec_5_2 = checkVec_checkResultVec_dataPosition_5[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_5 = checkVec_checkResultVec_dataPosition_5[10:7];
  wire               checkVec_checkResultVec_5_3 = checkVec_checkResultVec_dataGroup_5[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_5 = checkVec_checkResultVec_dataGroup_5[3:1];
  wire [2:0]         checkVec_checkResultVec_5_4 = checkVec_checkResultVec_accessRegGrowth_5;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_5 = {checkVec_checkResultVec_5_3, checkVec_checkResultVec_5_2};
  wire [2:0]         checkVec_checkResultVec_decimal_5 = checkVec_checkResultVec_decimalProportion_5[5:3];
  wire               checkVec_checkResultVec_overlap_5 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_5 >= checkVec_checkResultVec_intLMULInput_5[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_5} >= checkVec_checkResultVec_intLMULInput_5, source_5[31:11]};
  wire               checkVec_checkResultVec_5_5 = checkVec_checkResultVec_overlap_5 | ~checkVec_checkResultVec_5_6;
  wire               checkVec_checkResultVec_6_6 = checkVec_validVec[6];
  wire [10:0]        checkVec_checkResultVec_dataPosition_6 = source_6[10:0];
  wire [3:0]         checkVec_checkResultVec_6_0 = 4'h1 << checkVec_checkResultVec_dataPosition_6[1:0];
  wire [1:0]         checkVec_checkResultVec_6_1 = checkVec_checkResultVec_dataPosition_6[1:0];
  wire [4:0]         checkVec_checkResultVec_6_2 = checkVec_checkResultVec_dataPosition_6[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_6 = checkVec_checkResultVec_dataPosition_6[10:7];
  wire               checkVec_checkResultVec_6_3 = checkVec_checkResultVec_dataGroup_6[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_6 = checkVec_checkResultVec_dataGroup_6[3:1];
  wire [2:0]         checkVec_checkResultVec_6_4 = checkVec_checkResultVec_accessRegGrowth_6;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_6 = {checkVec_checkResultVec_6_3, checkVec_checkResultVec_6_2};
  wire [2:0]         checkVec_checkResultVec_decimal_6 = checkVec_checkResultVec_decimalProportion_6[5:3];
  wire               checkVec_checkResultVec_overlap_6 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_6 >= checkVec_checkResultVec_intLMULInput_6[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_6} >= checkVec_checkResultVec_intLMULInput_6, source_6[31:11]};
  wire               checkVec_checkResultVec_6_5 = checkVec_checkResultVec_overlap_6 | ~checkVec_checkResultVec_6_6;
  wire               checkVec_checkResultVec_7_6 = checkVec_validVec[7];
  wire [10:0]        checkVec_checkResultVec_dataPosition_7 = source_7[10:0];
  wire [3:0]         checkVec_checkResultVec_7_0 = 4'h1 << checkVec_checkResultVec_dataPosition_7[1:0];
  wire [1:0]         checkVec_checkResultVec_7_1 = checkVec_checkResultVec_dataPosition_7[1:0];
  wire [4:0]         checkVec_checkResultVec_7_2 = checkVec_checkResultVec_dataPosition_7[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_7 = checkVec_checkResultVec_dataPosition_7[10:7];
  wire               checkVec_checkResultVec_7_3 = checkVec_checkResultVec_dataGroup_7[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_7 = checkVec_checkResultVec_dataGroup_7[3:1];
  wire [2:0]         checkVec_checkResultVec_7_4 = checkVec_checkResultVec_accessRegGrowth_7;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_7 = {checkVec_checkResultVec_7_3, checkVec_checkResultVec_7_2};
  wire [2:0]         checkVec_checkResultVec_decimal_7 = checkVec_checkResultVec_decimalProportion_7[5:3];
  wire               checkVec_checkResultVec_overlap_7 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_7 >= checkVec_checkResultVec_intLMULInput_7[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_7} >= checkVec_checkResultVec_intLMULInput_7, source_7[31:11]};
  wire               checkVec_checkResultVec_7_5 = checkVec_checkResultVec_overlap_7 | ~checkVec_checkResultVec_7_6;
  wire               checkVec_checkResultVec_8_6 = checkVec_validVec[8];
  wire [10:0]        checkVec_checkResultVec_dataPosition_8 = source_8[10:0];
  wire [3:0]         checkVec_checkResultVec_8_0 = 4'h1 << checkVec_checkResultVec_dataPosition_8[1:0];
  wire [1:0]         checkVec_checkResultVec_8_1 = checkVec_checkResultVec_dataPosition_8[1:0];
  wire [4:0]         checkVec_checkResultVec_8_2 = checkVec_checkResultVec_dataPosition_8[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_8 = checkVec_checkResultVec_dataPosition_8[10:7];
  wire               checkVec_checkResultVec_8_3 = checkVec_checkResultVec_dataGroup_8[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_8 = checkVec_checkResultVec_dataGroup_8[3:1];
  wire [2:0]         checkVec_checkResultVec_8_4 = checkVec_checkResultVec_accessRegGrowth_8;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_8 = {checkVec_checkResultVec_8_3, checkVec_checkResultVec_8_2};
  wire [2:0]         checkVec_checkResultVec_decimal_8 = checkVec_checkResultVec_decimalProportion_8[5:3];
  wire               checkVec_checkResultVec_overlap_8 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_8 >= checkVec_checkResultVec_intLMULInput_8[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_8} >= checkVec_checkResultVec_intLMULInput_8, source_8[31:11]};
  wire               checkVec_checkResultVec_8_5 = checkVec_checkResultVec_overlap_8 | ~checkVec_checkResultVec_8_6;
  wire               checkVec_checkResultVec_9_6 = checkVec_validVec[9];
  wire [10:0]        checkVec_checkResultVec_dataPosition_9 = source_9[10:0];
  wire [3:0]         checkVec_checkResultVec_9_0 = 4'h1 << checkVec_checkResultVec_dataPosition_9[1:0];
  wire [1:0]         checkVec_checkResultVec_9_1 = checkVec_checkResultVec_dataPosition_9[1:0];
  wire [4:0]         checkVec_checkResultVec_9_2 = checkVec_checkResultVec_dataPosition_9[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_9 = checkVec_checkResultVec_dataPosition_9[10:7];
  wire               checkVec_checkResultVec_9_3 = checkVec_checkResultVec_dataGroup_9[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_9 = checkVec_checkResultVec_dataGroup_9[3:1];
  wire [2:0]         checkVec_checkResultVec_9_4 = checkVec_checkResultVec_accessRegGrowth_9;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_9 = {checkVec_checkResultVec_9_3, checkVec_checkResultVec_9_2};
  wire [2:0]         checkVec_checkResultVec_decimal_9 = checkVec_checkResultVec_decimalProportion_9[5:3];
  wire               checkVec_checkResultVec_overlap_9 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_9 >= checkVec_checkResultVec_intLMULInput_9[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_9} >= checkVec_checkResultVec_intLMULInput_9, source_9[31:11]};
  wire               checkVec_checkResultVec_9_5 = checkVec_checkResultVec_overlap_9 | ~checkVec_checkResultVec_9_6;
  wire               checkVec_checkResultVec_10_6 = checkVec_validVec[10];
  wire [10:0]        checkVec_checkResultVec_dataPosition_10 = source_10[10:0];
  wire [3:0]         checkVec_checkResultVec_10_0 = 4'h1 << checkVec_checkResultVec_dataPosition_10[1:0];
  wire [1:0]         checkVec_checkResultVec_10_1 = checkVec_checkResultVec_dataPosition_10[1:0];
  wire [4:0]         checkVec_checkResultVec_10_2 = checkVec_checkResultVec_dataPosition_10[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_10 = checkVec_checkResultVec_dataPosition_10[10:7];
  wire               checkVec_checkResultVec_10_3 = checkVec_checkResultVec_dataGroup_10[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_10 = checkVec_checkResultVec_dataGroup_10[3:1];
  wire [2:0]         checkVec_checkResultVec_10_4 = checkVec_checkResultVec_accessRegGrowth_10;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_10 = {checkVec_checkResultVec_10_3, checkVec_checkResultVec_10_2};
  wire [2:0]         checkVec_checkResultVec_decimal_10 = checkVec_checkResultVec_decimalProportion_10[5:3];
  wire               checkVec_checkResultVec_overlap_10 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_10 >= checkVec_checkResultVec_intLMULInput_10[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_10} >= checkVec_checkResultVec_intLMULInput_10,
      source_10[31:11]};
  wire               checkVec_checkResultVec_10_5 = checkVec_checkResultVec_overlap_10 | ~checkVec_checkResultVec_10_6;
  wire               checkVec_checkResultVec_11_6 = checkVec_validVec[11];
  wire [10:0]        checkVec_checkResultVec_dataPosition_11 = source_11[10:0];
  wire [3:0]         checkVec_checkResultVec_11_0 = 4'h1 << checkVec_checkResultVec_dataPosition_11[1:0];
  wire [1:0]         checkVec_checkResultVec_11_1 = checkVec_checkResultVec_dataPosition_11[1:0];
  wire [4:0]         checkVec_checkResultVec_11_2 = checkVec_checkResultVec_dataPosition_11[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_11 = checkVec_checkResultVec_dataPosition_11[10:7];
  wire               checkVec_checkResultVec_11_3 = checkVec_checkResultVec_dataGroup_11[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_11 = checkVec_checkResultVec_dataGroup_11[3:1];
  wire [2:0]         checkVec_checkResultVec_11_4 = checkVec_checkResultVec_accessRegGrowth_11;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_11 = {checkVec_checkResultVec_11_3, checkVec_checkResultVec_11_2};
  wire [2:0]         checkVec_checkResultVec_decimal_11 = checkVec_checkResultVec_decimalProportion_11[5:3];
  wire               checkVec_checkResultVec_overlap_11 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_11 >= checkVec_checkResultVec_intLMULInput_11[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_11} >= checkVec_checkResultVec_intLMULInput_11,
      source_11[31:11]};
  wire               checkVec_checkResultVec_11_5 = checkVec_checkResultVec_overlap_11 | ~checkVec_checkResultVec_11_6;
  wire               checkVec_checkResultVec_12_6 = checkVec_validVec[12];
  wire [10:0]        checkVec_checkResultVec_dataPosition_12 = source_12[10:0];
  wire [3:0]         checkVec_checkResultVec_12_0 = 4'h1 << checkVec_checkResultVec_dataPosition_12[1:0];
  wire [1:0]         checkVec_checkResultVec_12_1 = checkVec_checkResultVec_dataPosition_12[1:0];
  wire [4:0]         checkVec_checkResultVec_12_2 = checkVec_checkResultVec_dataPosition_12[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_12 = checkVec_checkResultVec_dataPosition_12[10:7];
  wire               checkVec_checkResultVec_12_3 = checkVec_checkResultVec_dataGroup_12[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_12 = checkVec_checkResultVec_dataGroup_12[3:1];
  wire [2:0]         checkVec_checkResultVec_12_4 = checkVec_checkResultVec_accessRegGrowth_12;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_12 = {checkVec_checkResultVec_12_3, checkVec_checkResultVec_12_2};
  wire [2:0]         checkVec_checkResultVec_decimal_12 = checkVec_checkResultVec_decimalProportion_12[5:3];
  wire               checkVec_checkResultVec_overlap_12 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_12 >= checkVec_checkResultVec_intLMULInput_12[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_12} >= checkVec_checkResultVec_intLMULInput_12,
      source_12[31:11]};
  wire               checkVec_checkResultVec_12_5 = checkVec_checkResultVec_overlap_12 | ~checkVec_checkResultVec_12_6;
  wire               checkVec_checkResultVec_13_6 = checkVec_validVec[13];
  wire [10:0]        checkVec_checkResultVec_dataPosition_13 = source_13[10:0];
  wire [3:0]         checkVec_checkResultVec_13_0 = 4'h1 << checkVec_checkResultVec_dataPosition_13[1:0];
  wire [1:0]         checkVec_checkResultVec_13_1 = checkVec_checkResultVec_dataPosition_13[1:0];
  wire [4:0]         checkVec_checkResultVec_13_2 = checkVec_checkResultVec_dataPosition_13[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_13 = checkVec_checkResultVec_dataPosition_13[10:7];
  wire               checkVec_checkResultVec_13_3 = checkVec_checkResultVec_dataGroup_13[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_13 = checkVec_checkResultVec_dataGroup_13[3:1];
  wire [2:0]         checkVec_checkResultVec_13_4 = checkVec_checkResultVec_accessRegGrowth_13;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_13 = {checkVec_checkResultVec_13_3, checkVec_checkResultVec_13_2};
  wire [2:0]         checkVec_checkResultVec_decimal_13 = checkVec_checkResultVec_decimalProportion_13[5:3];
  wire               checkVec_checkResultVec_overlap_13 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_13 >= checkVec_checkResultVec_intLMULInput_13[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_13} >= checkVec_checkResultVec_intLMULInput_13,
      source_13[31:11]};
  wire               checkVec_checkResultVec_13_5 = checkVec_checkResultVec_overlap_13 | ~checkVec_checkResultVec_13_6;
  wire               checkVec_checkResultVec_14_6 = checkVec_validVec[14];
  wire [10:0]        checkVec_checkResultVec_dataPosition_14 = source_14[10:0];
  wire [3:0]         checkVec_checkResultVec_14_0 = 4'h1 << checkVec_checkResultVec_dataPosition_14[1:0];
  wire [1:0]         checkVec_checkResultVec_14_1 = checkVec_checkResultVec_dataPosition_14[1:0];
  wire [4:0]         checkVec_checkResultVec_14_2 = checkVec_checkResultVec_dataPosition_14[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_14 = checkVec_checkResultVec_dataPosition_14[10:7];
  wire               checkVec_checkResultVec_14_3 = checkVec_checkResultVec_dataGroup_14[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_14 = checkVec_checkResultVec_dataGroup_14[3:1];
  wire [2:0]         checkVec_checkResultVec_14_4 = checkVec_checkResultVec_accessRegGrowth_14;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_14 = {checkVec_checkResultVec_14_3, checkVec_checkResultVec_14_2};
  wire [2:0]         checkVec_checkResultVec_decimal_14 = checkVec_checkResultVec_decimalProportion_14[5:3];
  wire               checkVec_checkResultVec_overlap_14 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_14 >= checkVec_checkResultVec_intLMULInput_14[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_14} >= checkVec_checkResultVec_intLMULInput_14,
      source_14[31:11]};
  wire               checkVec_checkResultVec_14_5 = checkVec_checkResultVec_overlap_14 | ~checkVec_checkResultVec_14_6;
  wire               checkVec_checkResultVec_15_6 = checkVec_validVec[15];
  wire [10:0]        checkVec_checkResultVec_dataPosition_15 = source_15[10:0];
  wire [3:0]         checkVec_checkResultVec_15_0 = 4'h1 << checkVec_checkResultVec_dataPosition_15[1:0];
  wire [1:0]         checkVec_checkResultVec_15_1 = checkVec_checkResultVec_dataPosition_15[1:0];
  wire [4:0]         checkVec_checkResultVec_15_2 = checkVec_checkResultVec_dataPosition_15[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_15 = checkVec_checkResultVec_dataPosition_15[10:7];
  wire               checkVec_checkResultVec_15_3 = checkVec_checkResultVec_dataGroup_15[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_15 = checkVec_checkResultVec_dataGroup_15[3:1];
  wire [2:0]         checkVec_checkResultVec_15_4 = checkVec_checkResultVec_accessRegGrowth_15;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_15 = {checkVec_checkResultVec_15_3, checkVec_checkResultVec_15_2};
  wire [2:0]         checkVec_checkResultVec_decimal_15 = checkVec_checkResultVec_decimalProportion_15[5:3];
  wire               checkVec_checkResultVec_overlap_15 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_15 >= checkVec_checkResultVec_intLMULInput_15[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_15} >= checkVec_checkResultVec_intLMULInput_15,
      source_15[31:11]};
  wire               checkVec_checkResultVec_15_5 = checkVec_checkResultVec_overlap_15 | ~checkVec_checkResultVec_15_6;
  wire               checkVec_checkResultVec_16_6 = checkVec_validVec[16];
  wire [10:0]        checkVec_checkResultVec_dataPosition_16 = source_16[10:0];
  wire [3:0]         checkVec_checkResultVec_16_0 = 4'h1 << checkVec_checkResultVec_dataPosition_16[1:0];
  wire [1:0]         checkVec_checkResultVec_16_1 = checkVec_checkResultVec_dataPosition_16[1:0];
  wire [4:0]         checkVec_checkResultVec_16_2 = checkVec_checkResultVec_dataPosition_16[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_16 = checkVec_checkResultVec_dataPosition_16[10:7];
  wire               checkVec_checkResultVec_16_3 = checkVec_checkResultVec_dataGroup_16[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_16 = checkVec_checkResultVec_dataGroup_16[3:1];
  wire [2:0]         checkVec_checkResultVec_16_4 = checkVec_checkResultVec_accessRegGrowth_16;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_16 = {checkVec_checkResultVec_16_3, checkVec_checkResultVec_16_2};
  wire [2:0]         checkVec_checkResultVec_decimal_16 = checkVec_checkResultVec_decimalProportion_16[5:3];
  wire               checkVec_checkResultVec_overlap_16 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_16 >= checkVec_checkResultVec_intLMULInput_16[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_16} >= checkVec_checkResultVec_intLMULInput_16,
      source_16[31:11]};
  wire               checkVec_checkResultVec_16_5 = checkVec_checkResultVec_overlap_16 | ~checkVec_checkResultVec_16_6;
  wire               checkVec_checkResultVec_17_6 = checkVec_validVec[17];
  wire [10:0]        checkVec_checkResultVec_dataPosition_17 = source_17[10:0];
  wire [3:0]         checkVec_checkResultVec_17_0 = 4'h1 << checkVec_checkResultVec_dataPosition_17[1:0];
  wire [1:0]         checkVec_checkResultVec_17_1 = checkVec_checkResultVec_dataPosition_17[1:0];
  wire [4:0]         checkVec_checkResultVec_17_2 = checkVec_checkResultVec_dataPosition_17[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_17 = checkVec_checkResultVec_dataPosition_17[10:7];
  wire               checkVec_checkResultVec_17_3 = checkVec_checkResultVec_dataGroup_17[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_17 = checkVec_checkResultVec_dataGroup_17[3:1];
  wire [2:0]         checkVec_checkResultVec_17_4 = checkVec_checkResultVec_accessRegGrowth_17;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_17 = {checkVec_checkResultVec_17_3, checkVec_checkResultVec_17_2};
  wire [2:0]         checkVec_checkResultVec_decimal_17 = checkVec_checkResultVec_decimalProportion_17[5:3];
  wire               checkVec_checkResultVec_overlap_17 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_17 >= checkVec_checkResultVec_intLMULInput_17[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_17} >= checkVec_checkResultVec_intLMULInput_17,
      source_17[31:11]};
  wire               checkVec_checkResultVec_17_5 = checkVec_checkResultVec_overlap_17 | ~checkVec_checkResultVec_17_6;
  wire               checkVec_checkResultVec_18_6 = checkVec_validVec[18];
  wire [10:0]        checkVec_checkResultVec_dataPosition_18 = source_18[10:0];
  wire [3:0]         checkVec_checkResultVec_18_0 = 4'h1 << checkVec_checkResultVec_dataPosition_18[1:0];
  wire [1:0]         checkVec_checkResultVec_18_1 = checkVec_checkResultVec_dataPosition_18[1:0];
  wire [4:0]         checkVec_checkResultVec_18_2 = checkVec_checkResultVec_dataPosition_18[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_18 = checkVec_checkResultVec_dataPosition_18[10:7];
  wire               checkVec_checkResultVec_18_3 = checkVec_checkResultVec_dataGroup_18[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_18 = checkVec_checkResultVec_dataGroup_18[3:1];
  wire [2:0]         checkVec_checkResultVec_18_4 = checkVec_checkResultVec_accessRegGrowth_18;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_18 = {checkVec_checkResultVec_18_3, checkVec_checkResultVec_18_2};
  wire [2:0]         checkVec_checkResultVec_decimal_18 = checkVec_checkResultVec_decimalProportion_18[5:3];
  wire               checkVec_checkResultVec_overlap_18 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_18 >= checkVec_checkResultVec_intLMULInput_18[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_18} >= checkVec_checkResultVec_intLMULInput_18,
      source_18[31:11]};
  wire               checkVec_checkResultVec_18_5 = checkVec_checkResultVec_overlap_18 | ~checkVec_checkResultVec_18_6;
  wire               checkVec_checkResultVec_19_6 = checkVec_validVec[19];
  wire [10:0]        checkVec_checkResultVec_dataPosition_19 = source_19[10:0];
  wire [3:0]         checkVec_checkResultVec_19_0 = 4'h1 << checkVec_checkResultVec_dataPosition_19[1:0];
  wire [1:0]         checkVec_checkResultVec_19_1 = checkVec_checkResultVec_dataPosition_19[1:0];
  wire [4:0]         checkVec_checkResultVec_19_2 = checkVec_checkResultVec_dataPosition_19[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_19 = checkVec_checkResultVec_dataPosition_19[10:7];
  wire               checkVec_checkResultVec_19_3 = checkVec_checkResultVec_dataGroup_19[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_19 = checkVec_checkResultVec_dataGroup_19[3:1];
  wire [2:0]         checkVec_checkResultVec_19_4 = checkVec_checkResultVec_accessRegGrowth_19;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_19 = {checkVec_checkResultVec_19_3, checkVec_checkResultVec_19_2};
  wire [2:0]         checkVec_checkResultVec_decimal_19 = checkVec_checkResultVec_decimalProportion_19[5:3];
  wire               checkVec_checkResultVec_overlap_19 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_19 >= checkVec_checkResultVec_intLMULInput_19[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_19} >= checkVec_checkResultVec_intLMULInput_19,
      source_19[31:11]};
  wire               checkVec_checkResultVec_19_5 = checkVec_checkResultVec_overlap_19 | ~checkVec_checkResultVec_19_6;
  wire               checkVec_checkResultVec_20_6 = checkVec_validVec[20];
  wire [10:0]        checkVec_checkResultVec_dataPosition_20 = source_20[10:0];
  wire [3:0]         checkVec_checkResultVec_20_0 = 4'h1 << checkVec_checkResultVec_dataPosition_20[1:0];
  wire [1:0]         checkVec_checkResultVec_20_1 = checkVec_checkResultVec_dataPosition_20[1:0];
  wire [4:0]         checkVec_checkResultVec_20_2 = checkVec_checkResultVec_dataPosition_20[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_20 = checkVec_checkResultVec_dataPosition_20[10:7];
  wire               checkVec_checkResultVec_20_3 = checkVec_checkResultVec_dataGroup_20[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_20 = checkVec_checkResultVec_dataGroup_20[3:1];
  wire [2:0]         checkVec_checkResultVec_20_4 = checkVec_checkResultVec_accessRegGrowth_20;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_20 = {checkVec_checkResultVec_20_3, checkVec_checkResultVec_20_2};
  wire [2:0]         checkVec_checkResultVec_decimal_20 = checkVec_checkResultVec_decimalProportion_20[5:3];
  wire               checkVec_checkResultVec_overlap_20 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_20 >= checkVec_checkResultVec_intLMULInput_20[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_20} >= checkVec_checkResultVec_intLMULInput_20,
      source_20[31:11]};
  wire               checkVec_checkResultVec_20_5 = checkVec_checkResultVec_overlap_20 | ~checkVec_checkResultVec_20_6;
  wire               checkVec_checkResultVec_21_6 = checkVec_validVec[21];
  wire [10:0]        checkVec_checkResultVec_dataPosition_21 = source_21[10:0];
  wire [3:0]         checkVec_checkResultVec_21_0 = 4'h1 << checkVec_checkResultVec_dataPosition_21[1:0];
  wire [1:0]         checkVec_checkResultVec_21_1 = checkVec_checkResultVec_dataPosition_21[1:0];
  wire [4:0]         checkVec_checkResultVec_21_2 = checkVec_checkResultVec_dataPosition_21[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_21 = checkVec_checkResultVec_dataPosition_21[10:7];
  wire               checkVec_checkResultVec_21_3 = checkVec_checkResultVec_dataGroup_21[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_21 = checkVec_checkResultVec_dataGroup_21[3:1];
  wire [2:0]         checkVec_checkResultVec_21_4 = checkVec_checkResultVec_accessRegGrowth_21;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_21 = {checkVec_checkResultVec_21_3, checkVec_checkResultVec_21_2};
  wire [2:0]         checkVec_checkResultVec_decimal_21 = checkVec_checkResultVec_decimalProportion_21[5:3];
  wire               checkVec_checkResultVec_overlap_21 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_21 >= checkVec_checkResultVec_intLMULInput_21[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_21} >= checkVec_checkResultVec_intLMULInput_21,
      source_21[31:11]};
  wire               checkVec_checkResultVec_21_5 = checkVec_checkResultVec_overlap_21 | ~checkVec_checkResultVec_21_6;
  wire               checkVec_checkResultVec_22_6 = checkVec_validVec[22];
  wire [10:0]        checkVec_checkResultVec_dataPosition_22 = source_22[10:0];
  wire [3:0]         checkVec_checkResultVec_22_0 = 4'h1 << checkVec_checkResultVec_dataPosition_22[1:0];
  wire [1:0]         checkVec_checkResultVec_22_1 = checkVec_checkResultVec_dataPosition_22[1:0];
  wire [4:0]         checkVec_checkResultVec_22_2 = checkVec_checkResultVec_dataPosition_22[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_22 = checkVec_checkResultVec_dataPosition_22[10:7];
  wire               checkVec_checkResultVec_22_3 = checkVec_checkResultVec_dataGroup_22[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_22 = checkVec_checkResultVec_dataGroup_22[3:1];
  wire [2:0]         checkVec_checkResultVec_22_4 = checkVec_checkResultVec_accessRegGrowth_22;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_22 = {checkVec_checkResultVec_22_3, checkVec_checkResultVec_22_2};
  wire [2:0]         checkVec_checkResultVec_decimal_22 = checkVec_checkResultVec_decimalProportion_22[5:3];
  wire               checkVec_checkResultVec_overlap_22 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_22 >= checkVec_checkResultVec_intLMULInput_22[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_22} >= checkVec_checkResultVec_intLMULInput_22,
      source_22[31:11]};
  wire               checkVec_checkResultVec_22_5 = checkVec_checkResultVec_overlap_22 | ~checkVec_checkResultVec_22_6;
  wire               checkVec_checkResultVec_23_6 = checkVec_validVec[23];
  wire [10:0]        checkVec_checkResultVec_dataPosition_23 = source_23[10:0];
  wire [3:0]         checkVec_checkResultVec_23_0 = 4'h1 << checkVec_checkResultVec_dataPosition_23[1:0];
  wire [1:0]         checkVec_checkResultVec_23_1 = checkVec_checkResultVec_dataPosition_23[1:0];
  wire [4:0]         checkVec_checkResultVec_23_2 = checkVec_checkResultVec_dataPosition_23[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_23 = checkVec_checkResultVec_dataPosition_23[10:7];
  wire               checkVec_checkResultVec_23_3 = checkVec_checkResultVec_dataGroup_23[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_23 = checkVec_checkResultVec_dataGroup_23[3:1];
  wire [2:0]         checkVec_checkResultVec_23_4 = checkVec_checkResultVec_accessRegGrowth_23;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_23 = {checkVec_checkResultVec_23_3, checkVec_checkResultVec_23_2};
  wire [2:0]         checkVec_checkResultVec_decimal_23 = checkVec_checkResultVec_decimalProportion_23[5:3];
  wire               checkVec_checkResultVec_overlap_23 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_23 >= checkVec_checkResultVec_intLMULInput_23[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_23} >= checkVec_checkResultVec_intLMULInput_23,
      source_23[31:11]};
  wire               checkVec_checkResultVec_23_5 = checkVec_checkResultVec_overlap_23 | ~checkVec_checkResultVec_23_6;
  wire               checkVec_checkResultVec_24_6 = checkVec_validVec[24];
  wire [10:0]        checkVec_checkResultVec_dataPosition_24 = source_24[10:0];
  wire [3:0]         checkVec_checkResultVec_24_0 = 4'h1 << checkVec_checkResultVec_dataPosition_24[1:0];
  wire [1:0]         checkVec_checkResultVec_24_1 = checkVec_checkResultVec_dataPosition_24[1:0];
  wire [4:0]         checkVec_checkResultVec_24_2 = checkVec_checkResultVec_dataPosition_24[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_24 = checkVec_checkResultVec_dataPosition_24[10:7];
  wire               checkVec_checkResultVec_24_3 = checkVec_checkResultVec_dataGroup_24[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_24 = checkVec_checkResultVec_dataGroup_24[3:1];
  wire [2:0]         checkVec_checkResultVec_24_4 = checkVec_checkResultVec_accessRegGrowth_24;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_24 = {checkVec_checkResultVec_24_3, checkVec_checkResultVec_24_2};
  wire [2:0]         checkVec_checkResultVec_decimal_24 = checkVec_checkResultVec_decimalProportion_24[5:3];
  wire               checkVec_checkResultVec_overlap_24 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_24 >= checkVec_checkResultVec_intLMULInput_24[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_24} >= checkVec_checkResultVec_intLMULInput_24,
      source_24[31:11]};
  wire               checkVec_checkResultVec_24_5 = checkVec_checkResultVec_overlap_24 | ~checkVec_checkResultVec_24_6;
  wire               checkVec_checkResultVec_25_6 = checkVec_validVec[25];
  wire [10:0]        checkVec_checkResultVec_dataPosition_25 = source_25[10:0];
  wire [3:0]         checkVec_checkResultVec_25_0 = 4'h1 << checkVec_checkResultVec_dataPosition_25[1:0];
  wire [1:0]         checkVec_checkResultVec_25_1 = checkVec_checkResultVec_dataPosition_25[1:0];
  wire [4:0]         checkVec_checkResultVec_25_2 = checkVec_checkResultVec_dataPosition_25[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_25 = checkVec_checkResultVec_dataPosition_25[10:7];
  wire               checkVec_checkResultVec_25_3 = checkVec_checkResultVec_dataGroup_25[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_25 = checkVec_checkResultVec_dataGroup_25[3:1];
  wire [2:0]         checkVec_checkResultVec_25_4 = checkVec_checkResultVec_accessRegGrowth_25;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_25 = {checkVec_checkResultVec_25_3, checkVec_checkResultVec_25_2};
  wire [2:0]         checkVec_checkResultVec_decimal_25 = checkVec_checkResultVec_decimalProportion_25[5:3];
  wire               checkVec_checkResultVec_overlap_25 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_25 >= checkVec_checkResultVec_intLMULInput_25[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_25} >= checkVec_checkResultVec_intLMULInput_25,
      source_25[31:11]};
  wire               checkVec_checkResultVec_25_5 = checkVec_checkResultVec_overlap_25 | ~checkVec_checkResultVec_25_6;
  wire               checkVec_checkResultVec_26_6 = checkVec_validVec[26];
  wire [10:0]        checkVec_checkResultVec_dataPosition_26 = source_26[10:0];
  wire [3:0]         checkVec_checkResultVec_26_0 = 4'h1 << checkVec_checkResultVec_dataPosition_26[1:0];
  wire [1:0]         checkVec_checkResultVec_26_1 = checkVec_checkResultVec_dataPosition_26[1:0];
  wire [4:0]         checkVec_checkResultVec_26_2 = checkVec_checkResultVec_dataPosition_26[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_26 = checkVec_checkResultVec_dataPosition_26[10:7];
  wire               checkVec_checkResultVec_26_3 = checkVec_checkResultVec_dataGroup_26[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_26 = checkVec_checkResultVec_dataGroup_26[3:1];
  wire [2:0]         checkVec_checkResultVec_26_4 = checkVec_checkResultVec_accessRegGrowth_26;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_26 = {checkVec_checkResultVec_26_3, checkVec_checkResultVec_26_2};
  wire [2:0]         checkVec_checkResultVec_decimal_26 = checkVec_checkResultVec_decimalProportion_26[5:3];
  wire               checkVec_checkResultVec_overlap_26 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_26 >= checkVec_checkResultVec_intLMULInput_26[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_26} >= checkVec_checkResultVec_intLMULInput_26,
      source_26[31:11]};
  wire               checkVec_checkResultVec_26_5 = checkVec_checkResultVec_overlap_26 | ~checkVec_checkResultVec_26_6;
  wire               checkVec_checkResultVec_27_6 = checkVec_validVec[27];
  wire [10:0]        checkVec_checkResultVec_dataPosition_27 = source_27[10:0];
  wire [3:0]         checkVec_checkResultVec_27_0 = 4'h1 << checkVec_checkResultVec_dataPosition_27[1:0];
  wire [1:0]         checkVec_checkResultVec_27_1 = checkVec_checkResultVec_dataPosition_27[1:0];
  wire [4:0]         checkVec_checkResultVec_27_2 = checkVec_checkResultVec_dataPosition_27[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_27 = checkVec_checkResultVec_dataPosition_27[10:7];
  wire               checkVec_checkResultVec_27_3 = checkVec_checkResultVec_dataGroup_27[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_27 = checkVec_checkResultVec_dataGroup_27[3:1];
  wire [2:0]         checkVec_checkResultVec_27_4 = checkVec_checkResultVec_accessRegGrowth_27;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_27 = {checkVec_checkResultVec_27_3, checkVec_checkResultVec_27_2};
  wire [2:0]         checkVec_checkResultVec_decimal_27 = checkVec_checkResultVec_decimalProportion_27[5:3];
  wire               checkVec_checkResultVec_overlap_27 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_27 >= checkVec_checkResultVec_intLMULInput_27[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_27} >= checkVec_checkResultVec_intLMULInput_27,
      source_27[31:11]};
  wire               checkVec_checkResultVec_27_5 = checkVec_checkResultVec_overlap_27 | ~checkVec_checkResultVec_27_6;
  wire               checkVec_checkResultVec_28_6 = checkVec_validVec[28];
  wire [10:0]        checkVec_checkResultVec_dataPosition_28 = source_28[10:0];
  wire [3:0]         checkVec_checkResultVec_28_0 = 4'h1 << checkVec_checkResultVec_dataPosition_28[1:0];
  wire [1:0]         checkVec_checkResultVec_28_1 = checkVec_checkResultVec_dataPosition_28[1:0];
  wire [4:0]         checkVec_checkResultVec_28_2 = checkVec_checkResultVec_dataPosition_28[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_28 = checkVec_checkResultVec_dataPosition_28[10:7];
  wire               checkVec_checkResultVec_28_3 = checkVec_checkResultVec_dataGroup_28[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_28 = checkVec_checkResultVec_dataGroup_28[3:1];
  wire [2:0]         checkVec_checkResultVec_28_4 = checkVec_checkResultVec_accessRegGrowth_28;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_28 = {checkVec_checkResultVec_28_3, checkVec_checkResultVec_28_2};
  wire [2:0]         checkVec_checkResultVec_decimal_28 = checkVec_checkResultVec_decimalProportion_28[5:3];
  wire               checkVec_checkResultVec_overlap_28 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_28 >= checkVec_checkResultVec_intLMULInput_28[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_28} >= checkVec_checkResultVec_intLMULInput_28,
      source_28[31:11]};
  wire               checkVec_checkResultVec_28_5 = checkVec_checkResultVec_overlap_28 | ~checkVec_checkResultVec_28_6;
  wire               checkVec_checkResultVec_29_6 = checkVec_validVec[29];
  wire [10:0]        checkVec_checkResultVec_dataPosition_29 = source_29[10:0];
  wire [3:0]         checkVec_checkResultVec_29_0 = 4'h1 << checkVec_checkResultVec_dataPosition_29[1:0];
  wire [1:0]         checkVec_checkResultVec_29_1 = checkVec_checkResultVec_dataPosition_29[1:0];
  wire [4:0]         checkVec_checkResultVec_29_2 = checkVec_checkResultVec_dataPosition_29[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_29 = checkVec_checkResultVec_dataPosition_29[10:7];
  wire               checkVec_checkResultVec_29_3 = checkVec_checkResultVec_dataGroup_29[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_29 = checkVec_checkResultVec_dataGroup_29[3:1];
  wire [2:0]         checkVec_checkResultVec_29_4 = checkVec_checkResultVec_accessRegGrowth_29;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_29 = {checkVec_checkResultVec_29_3, checkVec_checkResultVec_29_2};
  wire [2:0]         checkVec_checkResultVec_decimal_29 = checkVec_checkResultVec_decimalProportion_29[5:3];
  wire               checkVec_checkResultVec_overlap_29 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_29 >= checkVec_checkResultVec_intLMULInput_29[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_29} >= checkVec_checkResultVec_intLMULInput_29,
      source_29[31:11]};
  wire               checkVec_checkResultVec_29_5 = checkVec_checkResultVec_overlap_29 | ~checkVec_checkResultVec_29_6;
  wire               checkVec_checkResultVec_30_6 = checkVec_validVec[30];
  wire [10:0]        checkVec_checkResultVec_dataPosition_30 = source_30[10:0];
  wire [3:0]         checkVec_checkResultVec_30_0 = 4'h1 << checkVec_checkResultVec_dataPosition_30[1:0];
  wire [1:0]         checkVec_checkResultVec_30_1 = checkVec_checkResultVec_dataPosition_30[1:0];
  wire [4:0]         checkVec_checkResultVec_30_2 = checkVec_checkResultVec_dataPosition_30[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_30 = checkVec_checkResultVec_dataPosition_30[10:7];
  wire               checkVec_checkResultVec_30_3 = checkVec_checkResultVec_dataGroup_30[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_30 = checkVec_checkResultVec_dataGroup_30[3:1];
  wire [2:0]         checkVec_checkResultVec_30_4 = checkVec_checkResultVec_accessRegGrowth_30;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_30 = {checkVec_checkResultVec_30_3, checkVec_checkResultVec_30_2};
  wire [2:0]         checkVec_checkResultVec_decimal_30 = checkVec_checkResultVec_decimalProportion_30[5:3];
  wire               checkVec_checkResultVec_overlap_30 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_30 >= checkVec_checkResultVec_intLMULInput_30[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_30} >= checkVec_checkResultVec_intLMULInput_30,
      source_30[31:11]};
  wire               checkVec_checkResultVec_30_5 = checkVec_checkResultVec_overlap_30 | ~checkVec_checkResultVec_30_6;
  wire               checkVec_checkResultVec_31_6 = checkVec_validVec[31];
  wire [10:0]        checkVec_checkResultVec_dataPosition_31 = source_31[10:0];
  wire [3:0]         checkVec_checkResultVec_31_0 = 4'h1 << checkVec_checkResultVec_dataPosition_31[1:0];
  wire [1:0]         checkVec_checkResultVec_31_1 = checkVec_checkResultVec_dataPosition_31[1:0];
  wire [4:0]         checkVec_checkResultVec_31_2 = checkVec_checkResultVec_dataPosition_31[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_31 = checkVec_checkResultVec_dataPosition_31[10:7];
  wire               checkVec_checkResultVec_31_3 = checkVec_checkResultVec_dataGroup_31[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_31 = checkVec_checkResultVec_dataGroup_31[3:1];
  wire [2:0]         checkVec_checkResultVec_31_4 = checkVec_checkResultVec_accessRegGrowth_31;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_31 = {checkVec_checkResultVec_31_3, checkVec_checkResultVec_31_2};
  wire [2:0]         checkVec_checkResultVec_decimal_31 = checkVec_checkResultVec_decimalProportion_31[5:3];
  wire               checkVec_checkResultVec_overlap_31 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_31 >= checkVec_checkResultVec_intLMULInput_31[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_31} >= checkVec_checkResultVec_intLMULInput_31,
      source_31[31:11]};
  wire               checkVec_checkResultVec_31_5 = checkVec_checkResultVec_overlap_31 | ~checkVec_checkResultVec_31_6;
  wire [7:0]         checkVec_checkResult_lo_lo_lo_lo = {checkVec_checkResultVec_1_0, checkVec_checkResultVec_0_0};
  wire [7:0]         checkVec_checkResult_lo_lo_lo_hi = {checkVec_checkResultVec_3_0, checkVec_checkResultVec_2_0};
  wire [15:0]        checkVec_checkResult_lo_lo_lo = {checkVec_checkResult_lo_lo_lo_hi, checkVec_checkResult_lo_lo_lo_lo};
  wire [7:0]         checkVec_checkResult_lo_lo_hi_lo = {checkVec_checkResultVec_5_0, checkVec_checkResultVec_4_0};
  wire [7:0]         checkVec_checkResult_lo_lo_hi_hi = {checkVec_checkResultVec_7_0, checkVec_checkResultVec_6_0};
  wire [15:0]        checkVec_checkResult_lo_lo_hi = {checkVec_checkResult_lo_lo_hi_hi, checkVec_checkResult_lo_lo_hi_lo};
  wire [31:0]        checkVec_checkResult_lo_lo = {checkVec_checkResult_lo_lo_hi, checkVec_checkResult_lo_lo_lo};
  wire [7:0]         checkVec_checkResult_lo_hi_lo_lo = {checkVec_checkResultVec_9_0, checkVec_checkResultVec_8_0};
  wire [7:0]         checkVec_checkResult_lo_hi_lo_hi = {checkVec_checkResultVec_11_0, checkVec_checkResultVec_10_0};
  wire [15:0]        checkVec_checkResult_lo_hi_lo = {checkVec_checkResult_lo_hi_lo_hi, checkVec_checkResult_lo_hi_lo_lo};
  wire [7:0]         checkVec_checkResult_lo_hi_hi_lo = {checkVec_checkResultVec_13_0, checkVec_checkResultVec_12_0};
  wire [7:0]         checkVec_checkResult_lo_hi_hi_hi = {checkVec_checkResultVec_15_0, checkVec_checkResultVec_14_0};
  wire [15:0]        checkVec_checkResult_lo_hi_hi = {checkVec_checkResult_lo_hi_hi_hi, checkVec_checkResult_lo_hi_hi_lo};
  wire [31:0]        checkVec_checkResult_lo_hi = {checkVec_checkResult_lo_hi_hi, checkVec_checkResult_lo_hi_lo};
  wire [63:0]        checkVec_checkResult_lo = {checkVec_checkResult_lo_hi, checkVec_checkResult_lo_lo};
  wire [7:0]         checkVec_checkResult_hi_lo_lo_lo = {checkVec_checkResultVec_17_0, checkVec_checkResultVec_16_0};
  wire [7:0]         checkVec_checkResult_hi_lo_lo_hi = {checkVec_checkResultVec_19_0, checkVec_checkResultVec_18_0};
  wire [15:0]        checkVec_checkResult_hi_lo_lo = {checkVec_checkResult_hi_lo_lo_hi, checkVec_checkResult_hi_lo_lo_lo};
  wire [7:0]         checkVec_checkResult_hi_lo_hi_lo = {checkVec_checkResultVec_21_0, checkVec_checkResultVec_20_0};
  wire [7:0]         checkVec_checkResult_hi_lo_hi_hi = {checkVec_checkResultVec_23_0, checkVec_checkResultVec_22_0};
  wire [15:0]        checkVec_checkResult_hi_lo_hi = {checkVec_checkResult_hi_lo_hi_hi, checkVec_checkResult_hi_lo_hi_lo};
  wire [31:0]        checkVec_checkResult_hi_lo = {checkVec_checkResult_hi_lo_hi, checkVec_checkResult_hi_lo_lo};
  wire [7:0]         checkVec_checkResult_hi_hi_lo_lo = {checkVec_checkResultVec_25_0, checkVec_checkResultVec_24_0};
  wire [7:0]         checkVec_checkResult_hi_hi_lo_hi = {checkVec_checkResultVec_27_0, checkVec_checkResultVec_26_0};
  wire [15:0]        checkVec_checkResult_hi_hi_lo = {checkVec_checkResult_hi_hi_lo_hi, checkVec_checkResult_hi_hi_lo_lo};
  wire [7:0]         checkVec_checkResult_hi_hi_hi_lo = {checkVec_checkResultVec_29_0, checkVec_checkResultVec_28_0};
  wire [7:0]         checkVec_checkResult_hi_hi_hi_hi = {checkVec_checkResultVec_31_0, checkVec_checkResultVec_30_0};
  wire [15:0]        checkVec_checkResult_hi_hi_hi = {checkVec_checkResult_hi_hi_hi_hi, checkVec_checkResult_hi_hi_hi_lo};
  wire [31:0]        checkVec_checkResult_hi_hi = {checkVec_checkResult_hi_hi_hi, checkVec_checkResult_hi_hi_lo};
  wire [63:0]        checkVec_checkResult_hi = {checkVec_checkResult_hi_hi, checkVec_checkResult_hi_lo};
  wire [127:0]       checkVec_0_0 = {checkVec_checkResult_hi, checkVec_checkResult_lo};
  wire [3:0]         checkVec_checkResult_lo_lo_lo_lo_1 = {checkVec_checkResultVec_1_1, checkVec_checkResultVec_0_1};
  wire [3:0]         checkVec_checkResult_lo_lo_lo_hi_1 = {checkVec_checkResultVec_3_1, checkVec_checkResultVec_2_1};
  wire [7:0]         checkVec_checkResult_lo_lo_lo_1 = {checkVec_checkResult_lo_lo_lo_hi_1, checkVec_checkResult_lo_lo_lo_lo_1};
  wire [3:0]         checkVec_checkResult_lo_lo_hi_lo_1 = {checkVec_checkResultVec_5_1, checkVec_checkResultVec_4_1};
  wire [3:0]         checkVec_checkResult_lo_lo_hi_hi_1 = {checkVec_checkResultVec_7_1, checkVec_checkResultVec_6_1};
  wire [7:0]         checkVec_checkResult_lo_lo_hi_1 = {checkVec_checkResult_lo_lo_hi_hi_1, checkVec_checkResult_lo_lo_hi_lo_1};
  wire [15:0]        checkVec_checkResult_lo_lo_1 = {checkVec_checkResult_lo_lo_hi_1, checkVec_checkResult_lo_lo_lo_1};
  wire [3:0]         checkVec_checkResult_lo_hi_lo_lo_1 = {checkVec_checkResultVec_9_1, checkVec_checkResultVec_8_1};
  wire [3:0]         checkVec_checkResult_lo_hi_lo_hi_1 = {checkVec_checkResultVec_11_1, checkVec_checkResultVec_10_1};
  wire [7:0]         checkVec_checkResult_lo_hi_lo_1 = {checkVec_checkResult_lo_hi_lo_hi_1, checkVec_checkResult_lo_hi_lo_lo_1};
  wire [3:0]         checkVec_checkResult_lo_hi_hi_lo_1 = {checkVec_checkResultVec_13_1, checkVec_checkResultVec_12_1};
  wire [3:0]         checkVec_checkResult_lo_hi_hi_hi_1 = {checkVec_checkResultVec_15_1, checkVec_checkResultVec_14_1};
  wire [7:0]         checkVec_checkResult_lo_hi_hi_1 = {checkVec_checkResult_lo_hi_hi_hi_1, checkVec_checkResult_lo_hi_hi_lo_1};
  wire [15:0]        checkVec_checkResult_lo_hi_1 = {checkVec_checkResult_lo_hi_hi_1, checkVec_checkResult_lo_hi_lo_1};
  wire [31:0]        checkVec_checkResult_lo_1 = {checkVec_checkResult_lo_hi_1, checkVec_checkResult_lo_lo_1};
  wire [3:0]         checkVec_checkResult_hi_lo_lo_lo_1 = {checkVec_checkResultVec_17_1, checkVec_checkResultVec_16_1};
  wire [3:0]         checkVec_checkResult_hi_lo_lo_hi_1 = {checkVec_checkResultVec_19_1, checkVec_checkResultVec_18_1};
  wire [7:0]         checkVec_checkResult_hi_lo_lo_1 = {checkVec_checkResult_hi_lo_lo_hi_1, checkVec_checkResult_hi_lo_lo_lo_1};
  wire [3:0]         checkVec_checkResult_hi_lo_hi_lo_1 = {checkVec_checkResultVec_21_1, checkVec_checkResultVec_20_1};
  wire [3:0]         checkVec_checkResult_hi_lo_hi_hi_1 = {checkVec_checkResultVec_23_1, checkVec_checkResultVec_22_1};
  wire [7:0]         checkVec_checkResult_hi_lo_hi_1 = {checkVec_checkResult_hi_lo_hi_hi_1, checkVec_checkResult_hi_lo_hi_lo_1};
  wire [15:0]        checkVec_checkResult_hi_lo_1 = {checkVec_checkResult_hi_lo_hi_1, checkVec_checkResult_hi_lo_lo_1};
  wire [3:0]         checkVec_checkResult_hi_hi_lo_lo_1 = {checkVec_checkResultVec_25_1, checkVec_checkResultVec_24_1};
  wire [3:0]         checkVec_checkResult_hi_hi_lo_hi_1 = {checkVec_checkResultVec_27_1, checkVec_checkResultVec_26_1};
  wire [7:0]         checkVec_checkResult_hi_hi_lo_1 = {checkVec_checkResult_hi_hi_lo_hi_1, checkVec_checkResult_hi_hi_lo_lo_1};
  wire [3:0]         checkVec_checkResult_hi_hi_hi_lo_1 = {checkVec_checkResultVec_29_1, checkVec_checkResultVec_28_1};
  wire [3:0]         checkVec_checkResult_hi_hi_hi_hi_1 = {checkVec_checkResultVec_31_1, checkVec_checkResultVec_30_1};
  wire [7:0]         checkVec_checkResult_hi_hi_hi_1 = {checkVec_checkResult_hi_hi_hi_hi_1, checkVec_checkResult_hi_hi_hi_lo_1};
  wire [15:0]        checkVec_checkResult_hi_hi_1 = {checkVec_checkResult_hi_hi_hi_1, checkVec_checkResult_hi_hi_lo_1};
  wire [31:0]        checkVec_checkResult_hi_1 = {checkVec_checkResult_hi_hi_1, checkVec_checkResult_hi_lo_1};
  wire [63:0]        checkVec_0_1 = {checkVec_checkResult_hi_1, checkVec_checkResult_lo_1};
  wire [9:0]         checkVec_checkResult_lo_lo_lo_lo_2 = {checkVec_checkResultVec_1_2, checkVec_checkResultVec_0_2};
  wire [9:0]         checkVec_checkResult_lo_lo_lo_hi_2 = {checkVec_checkResultVec_3_2, checkVec_checkResultVec_2_2};
  wire [19:0]        checkVec_checkResult_lo_lo_lo_2 = {checkVec_checkResult_lo_lo_lo_hi_2, checkVec_checkResult_lo_lo_lo_lo_2};
  wire [9:0]         checkVec_checkResult_lo_lo_hi_lo_2 = {checkVec_checkResultVec_5_2, checkVec_checkResultVec_4_2};
  wire [9:0]         checkVec_checkResult_lo_lo_hi_hi_2 = {checkVec_checkResultVec_7_2, checkVec_checkResultVec_6_2};
  wire [19:0]        checkVec_checkResult_lo_lo_hi_2 = {checkVec_checkResult_lo_lo_hi_hi_2, checkVec_checkResult_lo_lo_hi_lo_2};
  wire [39:0]        checkVec_checkResult_lo_lo_2 = {checkVec_checkResult_lo_lo_hi_2, checkVec_checkResult_lo_lo_lo_2};
  wire [9:0]         checkVec_checkResult_lo_hi_lo_lo_2 = {checkVec_checkResultVec_9_2, checkVec_checkResultVec_8_2};
  wire [9:0]         checkVec_checkResult_lo_hi_lo_hi_2 = {checkVec_checkResultVec_11_2, checkVec_checkResultVec_10_2};
  wire [19:0]        checkVec_checkResult_lo_hi_lo_2 = {checkVec_checkResult_lo_hi_lo_hi_2, checkVec_checkResult_lo_hi_lo_lo_2};
  wire [9:0]         checkVec_checkResult_lo_hi_hi_lo_2 = {checkVec_checkResultVec_13_2, checkVec_checkResultVec_12_2};
  wire [9:0]         checkVec_checkResult_lo_hi_hi_hi_2 = {checkVec_checkResultVec_15_2, checkVec_checkResultVec_14_2};
  wire [19:0]        checkVec_checkResult_lo_hi_hi_2 = {checkVec_checkResult_lo_hi_hi_hi_2, checkVec_checkResult_lo_hi_hi_lo_2};
  wire [39:0]        checkVec_checkResult_lo_hi_2 = {checkVec_checkResult_lo_hi_hi_2, checkVec_checkResult_lo_hi_lo_2};
  wire [79:0]        checkVec_checkResult_lo_2 = {checkVec_checkResult_lo_hi_2, checkVec_checkResult_lo_lo_2};
  wire [9:0]         checkVec_checkResult_hi_lo_lo_lo_2 = {checkVec_checkResultVec_17_2, checkVec_checkResultVec_16_2};
  wire [9:0]         checkVec_checkResult_hi_lo_lo_hi_2 = {checkVec_checkResultVec_19_2, checkVec_checkResultVec_18_2};
  wire [19:0]        checkVec_checkResult_hi_lo_lo_2 = {checkVec_checkResult_hi_lo_lo_hi_2, checkVec_checkResult_hi_lo_lo_lo_2};
  wire [9:0]         checkVec_checkResult_hi_lo_hi_lo_2 = {checkVec_checkResultVec_21_2, checkVec_checkResultVec_20_2};
  wire [9:0]         checkVec_checkResult_hi_lo_hi_hi_2 = {checkVec_checkResultVec_23_2, checkVec_checkResultVec_22_2};
  wire [19:0]        checkVec_checkResult_hi_lo_hi_2 = {checkVec_checkResult_hi_lo_hi_hi_2, checkVec_checkResult_hi_lo_hi_lo_2};
  wire [39:0]        checkVec_checkResult_hi_lo_2 = {checkVec_checkResult_hi_lo_hi_2, checkVec_checkResult_hi_lo_lo_2};
  wire [9:0]         checkVec_checkResult_hi_hi_lo_lo_2 = {checkVec_checkResultVec_25_2, checkVec_checkResultVec_24_2};
  wire [9:0]         checkVec_checkResult_hi_hi_lo_hi_2 = {checkVec_checkResultVec_27_2, checkVec_checkResultVec_26_2};
  wire [19:0]        checkVec_checkResult_hi_hi_lo_2 = {checkVec_checkResult_hi_hi_lo_hi_2, checkVec_checkResult_hi_hi_lo_lo_2};
  wire [9:0]         checkVec_checkResult_hi_hi_hi_lo_2 = {checkVec_checkResultVec_29_2, checkVec_checkResultVec_28_2};
  wire [9:0]         checkVec_checkResult_hi_hi_hi_hi_2 = {checkVec_checkResultVec_31_2, checkVec_checkResultVec_30_2};
  wire [19:0]        checkVec_checkResult_hi_hi_hi_2 = {checkVec_checkResult_hi_hi_hi_hi_2, checkVec_checkResult_hi_hi_hi_lo_2};
  wire [39:0]        checkVec_checkResult_hi_hi_2 = {checkVec_checkResult_hi_hi_hi_2, checkVec_checkResult_hi_hi_lo_2};
  wire [79:0]        checkVec_checkResult_hi_2 = {checkVec_checkResult_hi_hi_2, checkVec_checkResult_hi_lo_2};
  wire [159:0]       checkVec_0_2 = {checkVec_checkResult_hi_2, checkVec_checkResult_lo_2};
  wire [1:0]         checkVec_checkResult_lo_lo_lo_lo_3 = {checkVec_checkResultVec_1_3, checkVec_checkResultVec_0_3};
  wire [1:0]         checkVec_checkResult_lo_lo_lo_hi_3 = {checkVec_checkResultVec_3_3, checkVec_checkResultVec_2_3};
  wire [3:0]         checkVec_checkResult_lo_lo_lo_3 = {checkVec_checkResult_lo_lo_lo_hi_3, checkVec_checkResult_lo_lo_lo_lo_3};
  wire [1:0]         checkVec_checkResult_lo_lo_hi_lo_3 = {checkVec_checkResultVec_5_3, checkVec_checkResultVec_4_3};
  wire [1:0]         checkVec_checkResult_lo_lo_hi_hi_3 = {checkVec_checkResultVec_7_3, checkVec_checkResultVec_6_3};
  wire [3:0]         checkVec_checkResult_lo_lo_hi_3 = {checkVec_checkResult_lo_lo_hi_hi_3, checkVec_checkResult_lo_lo_hi_lo_3};
  wire [7:0]         checkVec_checkResult_lo_lo_3 = {checkVec_checkResult_lo_lo_hi_3, checkVec_checkResult_lo_lo_lo_3};
  wire [1:0]         checkVec_checkResult_lo_hi_lo_lo_3 = {checkVec_checkResultVec_9_3, checkVec_checkResultVec_8_3};
  wire [1:0]         checkVec_checkResult_lo_hi_lo_hi_3 = {checkVec_checkResultVec_11_3, checkVec_checkResultVec_10_3};
  wire [3:0]         checkVec_checkResult_lo_hi_lo_3 = {checkVec_checkResult_lo_hi_lo_hi_3, checkVec_checkResult_lo_hi_lo_lo_3};
  wire [1:0]         checkVec_checkResult_lo_hi_hi_lo_3 = {checkVec_checkResultVec_13_3, checkVec_checkResultVec_12_3};
  wire [1:0]         checkVec_checkResult_lo_hi_hi_hi_3 = {checkVec_checkResultVec_15_3, checkVec_checkResultVec_14_3};
  wire [3:0]         checkVec_checkResult_lo_hi_hi_3 = {checkVec_checkResult_lo_hi_hi_hi_3, checkVec_checkResult_lo_hi_hi_lo_3};
  wire [7:0]         checkVec_checkResult_lo_hi_3 = {checkVec_checkResult_lo_hi_hi_3, checkVec_checkResult_lo_hi_lo_3};
  wire [15:0]        checkVec_checkResult_lo_3 = {checkVec_checkResult_lo_hi_3, checkVec_checkResult_lo_lo_3};
  wire [1:0]         checkVec_checkResult_hi_lo_lo_lo_3 = {checkVec_checkResultVec_17_3, checkVec_checkResultVec_16_3};
  wire [1:0]         checkVec_checkResult_hi_lo_lo_hi_3 = {checkVec_checkResultVec_19_3, checkVec_checkResultVec_18_3};
  wire [3:0]         checkVec_checkResult_hi_lo_lo_3 = {checkVec_checkResult_hi_lo_lo_hi_3, checkVec_checkResult_hi_lo_lo_lo_3};
  wire [1:0]         checkVec_checkResult_hi_lo_hi_lo_3 = {checkVec_checkResultVec_21_3, checkVec_checkResultVec_20_3};
  wire [1:0]         checkVec_checkResult_hi_lo_hi_hi_3 = {checkVec_checkResultVec_23_3, checkVec_checkResultVec_22_3};
  wire [3:0]         checkVec_checkResult_hi_lo_hi_3 = {checkVec_checkResult_hi_lo_hi_hi_3, checkVec_checkResult_hi_lo_hi_lo_3};
  wire [7:0]         checkVec_checkResult_hi_lo_3 = {checkVec_checkResult_hi_lo_hi_3, checkVec_checkResult_hi_lo_lo_3};
  wire [1:0]         checkVec_checkResult_hi_hi_lo_lo_3 = {checkVec_checkResultVec_25_3, checkVec_checkResultVec_24_3};
  wire [1:0]         checkVec_checkResult_hi_hi_lo_hi_3 = {checkVec_checkResultVec_27_3, checkVec_checkResultVec_26_3};
  wire [3:0]         checkVec_checkResult_hi_hi_lo_3 = {checkVec_checkResult_hi_hi_lo_hi_3, checkVec_checkResult_hi_hi_lo_lo_3};
  wire [1:0]         checkVec_checkResult_hi_hi_hi_lo_3 = {checkVec_checkResultVec_29_3, checkVec_checkResultVec_28_3};
  wire [1:0]         checkVec_checkResult_hi_hi_hi_hi_3 = {checkVec_checkResultVec_31_3, checkVec_checkResultVec_30_3};
  wire [3:0]         checkVec_checkResult_hi_hi_hi_3 = {checkVec_checkResult_hi_hi_hi_hi_3, checkVec_checkResult_hi_hi_hi_lo_3};
  wire [7:0]         checkVec_checkResult_hi_hi_3 = {checkVec_checkResult_hi_hi_hi_3, checkVec_checkResult_hi_hi_lo_3};
  wire [15:0]        checkVec_checkResult_hi_3 = {checkVec_checkResult_hi_hi_3, checkVec_checkResult_hi_lo_3};
  wire [31:0]        checkVec_0_3 = {checkVec_checkResult_hi_3, checkVec_checkResult_lo_3};
  wire [5:0]         checkVec_checkResult_lo_lo_lo_lo_4 = {checkVec_checkResultVec_1_4, checkVec_checkResultVec_0_4};
  wire [5:0]         checkVec_checkResult_lo_lo_lo_hi_4 = {checkVec_checkResultVec_3_4, checkVec_checkResultVec_2_4};
  wire [11:0]        checkVec_checkResult_lo_lo_lo_4 = {checkVec_checkResult_lo_lo_lo_hi_4, checkVec_checkResult_lo_lo_lo_lo_4};
  wire [5:0]         checkVec_checkResult_lo_lo_hi_lo_4 = {checkVec_checkResultVec_5_4, checkVec_checkResultVec_4_4};
  wire [5:0]         checkVec_checkResult_lo_lo_hi_hi_4 = {checkVec_checkResultVec_7_4, checkVec_checkResultVec_6_4};
  wire [11:0]        checkVec_checkResult_lo_lo_hi_4 = {checkVec_checkResult_lo_lo_hi_hi_4, checkVec_checkResult_lo_lo_hi_lo_4};
  wire [23:0]        checkVec_checkResult_lo_lo_4 = {checkVec_checkResult_lo_lo_hi_4, checkVec_checkResult_lo_lo_lo_4};
  wire [5:0]         checkVec_checkResult_lo_hi_lo_lo_4 = {checkVec_checkResultVec_9_4, checkVec_checkResultVec_8_4};
  wire [5:0]         checkVec_checkResult_lo_hi_lo_hi_4 = {checkVec_checkResultVec_11_4, checkVec_checkResultVec_10_4};
  wire [11:0]        checkVec_checkResult_lo_hi_lo_4 = {checkVec_checkResult_lo_hi_lo_hi_4, checkVec_checkResult_lo_hi_lo_lo_4};
  wire [5:0]         checkVec_checkResult_lo_hi_hi_lo_4 = {checkVec_checkResultVec_13_4, checkVec_checkResultVec_12_4};
  wire [5:0]         checkVec_checkResult_lo_hi_hi_hi_4 = {checkVec_checkResultVec_15_4, checkVec_checkResultVec_14_4};
  wire [11:0]        checkVec_checkResult_lo_hi_hi_4 = {checkVec_checkResult_lo_hi_hi_hi_4, checkVec_checkResult_lo_hi_hi_lo_4};
  wire [23:0]        checkVec_checkResult_lo_hi_4 = {checkVec_checkResult_lo_hi_hi_4, checkVec_checkResult_lo_hi_lo_4};
  wire [47:0]        checkVec_checkResult_lo_4 = {checkVec_checkResult_lo_hi_4, checkVec_checkResult_lo_lo_4};
  wire [5:0]         checkVec_checkResult_hi_lo_lo_lo_4 = {checkVec_checkResultVec_17_4, checkVec_checkResultVec_16_4};
  wire [5:0]         checkVec_checkResult_hi_lo_lo_hi_4 = {checkVec_checkResultVec_19_4, checkVec_checkResultVec_18_4};
  wire [11:0]        checkVec_checkResult_hi_lo_lo_4 = {checkVec_checkResult_hi_lo_lo_hi_4, checkVec_checkResult_hi_lo_lo_lo_4};
  wire [5:0]         checkVec_checkResult_hi_lo_hi_lo_4 = {checkVec_checkResultVec_21_4, checkVec_checkResultVec_20_4};
  wire [5:0]         checkVec_checkResult_hi_lo_hi_hi_4 = {checkVec_checkResultVec_23_4, checkVec_checkResultVec_22_4};
  wire [11:0]        checkVec_checkResult_hi_lo_hi_4 = {checkVec_checkResult_hi_lo_hi_hi_4, checkVec_checkResult_hi_lo_hi_lo_4};
  wire [23:0]        checkVec_checkResult_hi_lo_4 = {checkVec_checkResult_hi_lo_hi_4, checkVec_checkResult_hi_lo_lo_4};
  wire [5:0]         checkVec_checkResult_hi_hi_lo_lo_4 = {checkVec_checkResultVec_25_4, checkVec_checkResultVec_24_4};
  wire [5:0]         checkVec_checkResult_hi_hi_lo_hi_4 = {checkVec_checkResultVec_27_4, checkVec_checkResultVec_26_4};
  wire [11:0]        checkVec_checkResult_hi_hi_lo_4 = {checkVec_checkResult_hi_hi_lo_hi_4, checkVec_checkResult_hi_hi_lo_lo_4};
  wire [5:0]         checkVec_checkResult_hi_hi_hi_lo_4 = {checkVec_checkResultVec_29_4, checkVec_checkResultVec_28_4};
  wire [5:0]         checkVec_checkResult_hi_hi_hi_hi_4 = {checkVec_checkResultVec_31_4, checkVec_checkResultVec_30_4};
  wire [11:0]        checkVec_checkResult_hi_hi_hi_4 = {checkVec_checkResult_hi_hi_hi_hi_4, checkVec_checkResult_hi_hi_hi_lo_4};
  wire [23:0]        checkVec_checkResult_hi_hi_4 = {checkVec_checkResult_hi_hi_hi_4, checkVec_checkResult_hi_hi_lo_4};
  wire [47:0]        checkVec_checkResult_hi_4 = {checkVec_checkResult_hi_hi_4, checkVec_checkResult_hi_lo_4};
  wire [95:0]        checkVec_0_4 = {checkVec_checkResult_hi_4, checkVec_checkResult_lo_4};
  wire [1:0]         checkVec_checkResult_lo_lo_lo_lo_5 = {checkVec_checkResultVec_1_5, checkVec_checkResultVec_0_5};
  wire [1:0]         checkVec_checkResult_lo_lo_lo_hi_5 = {checkVec_checkResultVec_3_5, checkVec_checkResultVec_2_5};
  wire [3:0]         checkVec_checkResult_lo_lo_lo_5 = {checkVec_checkResult_lo_lo_lo_hi_5, checkVec_checkResult_lo_lo_lo_lo_5};
  wire [1:0]         checkVec_checkResult_lo_lo_hi_lo_5 = {checkVec_checkResultVec_5_5, checkVec_checkResultVec_4_5};
  wire [1:0]         checkVec_checkResult_lo_lo_hi_hi_5 = {checkVec_checkResultVec_7_5, checkVec_checkResultVec_6_5};
  wire [3:0]         checkVec_checkResult_lo_lo_hi_5 = {checkVec_checkResult_lo_lo_hi_hi_5, checkVec_checkResult_lo_lo_hi_lo_5};
  wire [7:0]         checkVec_checkResult_lo_lo_5 = {checkVec_checkResult_lo_lo_hi_5, checkVec_checkResult_lo_lo_lo_5};
  wire [1:0]         checkVec_checkResult_lo_hi_lo_lo_5 = {checkVec_checkResultVec_9_5, checkVec_checkResultVec_8_5};
  wire [1:0]         checkVec_checkResult_lo_hi_lo_hi_5 = {checkVec_checkResultVec_11_5, checkVec_checkResultVec_10_5};
  wire [3:0]         checkVec_checkResult_lo_hi_lo_5 = {checkVec_checkResult_lo_hi_lo_hi_5, checkVec_checkResult_lo_hi_lo_lo_5};
  wire [1:0]         checkVec_checkResult_lo_hi_hi_lo_5 = {checkVec_checkResultVec_13_5, checkVec_checkResultVec_12_5};
  wire [1:0]         checkVec_checkResult_lo_hi_hi_hi_5 = {checkVec_checkResultVec_15_5, checkVec_checkResultVec_14_5};
  wire [3:0]         checkVec_checkResult_lo_hi_hi_5 = {checkVec_checkResult_lo_hi_hi_hi_5, checkVec_checkResult_lo_hi_hi_lo_5};
  wire [7:0]         checkVec_checkResult_lo_hi_5 = {checkVec_checkResult_lo_hi_hi_5, checkVec_checkResult_lo_hi_lo_5};
  wire [15:0]        checkVec_checkResult_lo_5 = {checkVec_checkResult_lo_hi_5, checkVec_checkResult_lo_lo_5};
  wire [1:0]         checkVec_checkResult_hi_lo_lo_lo_5 = {checkVec_checkResultVec_17_5, checkVec_checkResultVec_16_5};
  wire [1:0]         checkVec_checkResult_hi_lo_lo_hi_5 = {checkVec_checkResultVec_19_5, checkVec_checkResultVec_18_5};
  wire [3:0]         checkVec_checkResult_hi_lo_lo_5 = {checkVec_checkResult_hi_lo_lo_hi_5, checkVec_checkResult_hi_lo_lo_lo_5};
  wire [1:0]         checkVec_checkResult_hi_lo_hi_lo_5 = {checkVec_checkResultVec_21_5, checkVec_checkResultVec_20_5};
  wire [1:0]         checkVec_checkResult_hi_lo_hi_hi_5 = {checkVec_checkResultVec_23_5, checkVec_checkResultVec_22_5};
  wire [3:0]         checkVec_checkResult_hi_lo_hi_5 = {checkVec_checkResult_hi_lo_hi_hi_5, checkVec_checkResult_hi_lo_hi_lo_5};
  wire [7:0]         checkVec_checkResult_hi_lo_5 = {checkVec_checkResult_hi_lo_hi_5, checkVec_checkResult_hi_lo_lo_5};
  wire [1:0]         checkVec_checkResult_hi_hi_lo_lo_5 = {checkVec_checkResultVec_25_5, checkVec_checkResultVec_24_5};
  wire [1:0]         checkVec_checkResult_hi_hi_lo_hi_5 = {checkVec_checkResultVec_27_5, checkVec_checkResultVec_26_5};
  wire [3:0]         checkVec_checkResult_hi_hi_lo_5 = {checkVec_checkResult_hi_hi_lo_hi_5, checkVec_checkResult_hi_hi_lo_lo_5};
  wire [1:0]         checkVec_checkResult_hi_hi_hi_lo_5 = {checkVec_checkResultVec_29_5, checkVec_checkResultVec_28_5};
  wire [1:0]         checkVec_checkResult_hi_hi_hi_hi_5 = {checkVec_checkResultVec_31_5, checkVec_checkResultVec_30_5};
  wire [3:0]         checkVec_checkResult_hi_hi_hi_5 = {checkVec_checkResult_hi_hi_hi_hi_5, checkVec_checkResult_hi_hi_hi_lo_5};
  wire [7:0]         checkVec_checkResult_hi_hi_5 = {checkVec_checkResult_hi_hi_hi_5, checkVec_checkResult_hi_hi_lo_5};
  wire [15:0]        checkVec_checkResult_hi_5 = {checkVec_checkResult_hi_hi_5, checkVec_checkResult_hi_lo_5};
  wire [31:0]        checkVec_0_5 = {checkVec_checkResult_hi_5, checkVec_checkResult_lo_5};
  wire [1:0]         checkVec_checkResult_lo_lo_lo_lo_6 = {checkVec_checkResultVec_1_6, checkVec_checkResultVec_0_6};
  wire [1:0]         checkVec_checkResult_lo_lo_lo_hi_6 = {checkVec_checkResultVec_3_6, checkVec_checkResultVec_2_6};
  wire [3:0]         checkVec_checkResult_lo_lo_lo_6 = {checkVec_checkResult_lo_lo_lo_hi_6, checkVec_checkResult_lo_lo_lo_lo_6};
  wire [1:0]         checkVec_checkResult_lo_lo_hi_lo_6 = {checkVec_checkResultVec_5_6, checkVec_checkResultVec_4_6};
  wire [1:0]         checkVec_checkResult_lo_lo_hi_hi_6 = {checkVec_checkResultVec_7_6, checkVec_checkResultVec_6_6};
  wire [3:0]         checkVec_checkResult_lo_lo_hi_6 = {checkVec_checkResult_lo_lo_hi_hi_6, checkVec_checkResult_lo_lo_hi_lo_6};
  wire [7:0]         checkVec_checkResult_lo_lo_6 = {checkVec_checkResult_lo_lo_hi_6, checkVec_checkResult_lo_lo_lo_6};
  wire [1:0]         checkVec_checkResult_lo_hi_lo_lo_6 = {checkVec_checkResultVec_9_6, checkVec_checkResultVec_8_6};
  wire [1:0]         checkVec_checkResult_lo_hi_lo_hi_6 = {checkVec_checkResultVec_11_6, checkVec_checkResultVec_10_6};
  wire [3:0]         checkVec_checkResult_lo_hi_lo_6 = {checkVec_checkResult_lo_hi_lo_hi_6, checkVec_checkResult_lo_hi_lo_lo_6};
  wire [1:0]         checkVec_checkResult_lo_hi_hi_lo_6 = {checkVec_checkResultVec_13_6, checkVec_checkResultVec_12_6};
  wire [1:0]         checkVec_checkResult_lo_hi_hi_hi_6 = {checkVec_checkResultVec_15_6, checkVec_checkResultVec_14_6};
  wire [3:0]         checkVec_checkResult_lo_hi_hi_6 = {checkVec_checkResult_lo_hi_hi_hi_6, checkVec_checkResult_lo_hi_hi_lo_6};
  wire [7:0]         checkVec_checkResult_lo_hi_6 = {checkVec_checkResult_lo_hi_hi_6, checkVec_checkResult_lo_hi_lo_6};
  wire [15:0]        checkVec_checkResult_lo_6 = {checkVec_checkResult_lo_hi_6, checkVec_checkResult_lo_lo_6};
  wire [1:0]         checkVec_checkResult_hi_lo_lo_lo_6 = {checkVec_checkResultVec_17_6, checkVec_checkResultVec_16_6};
  wire [1:0]         checkVec_checkResult_hi_lo_lo_hi_6 = {checkVec_checkResultVec_19_6, checkVec_checkResultVec_18_6};
  wire [3:0]         checkVec_checkResult_hi_lo_lo_6 = {checkVec_checkResult_hi_lo_lo_hi_6, checkVec_checkResult_hi_lo_lo_lo_6};
  wire [1:0]         checkVec_checkResult_hi_lo_hi_lo_6 = {checkVec_checkResultVec_21_6, checkVec_checkResultVec_20_6};
  wire [1:0]         checkVec_checkResult_hi_lo_hi_hi_6 = {checkVec_checkResultVec_23_6, checkVec_checkResultVec_22_6};
  wire [3:0]         checkVec_checkResult_hi_lo_hi_6 = {checkVec_checkResult_hi_lo_hi_hi_6, checkVec_checkResult_hi_lo_hi_lo_6};
  wire [7:0]         checkVec_checkResult_hi_lo_6 = {checkVec_checkResult_hi_lo_hi_6, checkVec_checkResult_hi_lo_lo_6};
  wire [1:0]         checkVec_checkResult_hi_hi_lo_lo_6 = {checkVec_checkResultVec_25_6, checkVec_checkResultVec_24_6};
  wire [1:0]         checkVec_checkResult_hi_hi_lo_hi_6 = {checkVec_checkResultVec_27_6, checkVec_checkResultVec_26_6};
  wire [3:0]         checkVec_checkResult_hi_hi_lo_6 = {checkVec_checkResult_hi_hi_lo_hi_6, checkVec_checkResult_hi_hi_lo_lo_6};
  wire [1:0]         checkVec_checkResult_hi_hi_hi_lo_6 = {checkVec_checkResultVec_29_6, checkVec_checkResultVec_28_6};
  wire [1:0]         checkVec_checkResult_hi_hi_hi_hi_6 = {checkVec_checkResultVec_31_6, checkVec_checkResultVec_30_6};
  wire [3:0]         checkVec_checkResult_hi_hi_hi_6 = {checkVec_checkResult_hi_hi_hi_hi_6, checkVec_checkResult_hi_hi_hi_lo_6};
  wire [7:0]         checkVec_checkResult_hi_hi_6 = {checkVec_checkResult_hi_hi_hi_6, checkVec_checkResult_hi_hi_lo_6};
  wire [15:0]        checkVec_checkResult_hi_6 = {checkVec_checkResult_hi_hi_6, checkVec_checkResult_hi_lo_6};
  wire [31:0]        checkVec_0_6 = {checkVec_checkResult_hi_6, checkVec_checkResult_lo_6};
  wire               checkVec_checkResultVec_0_6_1 = checkVec_validVec_1[0];
  wire [10:0]        checkVec_checkResultVec_dataPosition_32 = {source_0[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_259 = 2'h1 << checkVec_checkResultVec_dataPosition_32[1];
  wire [3:0]         checkVec_checkResultVec_0_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_259[1]}}, {2{_checkVec_checkResultVec_accessMask_T_259[0]}}};
  wire [1:0]         checkVec_checkResultVec_0_1_1 = {checkVec_checkResultVec_dataPosition_32[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_0_2_1 = checkVec_checkResultVec_dataPosition_32[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_32 = checkVec_checkResultVec_dataPosition_32[10:7];
  wire               checkVec_checkResultVec_0_3_1 = checkVec_checkResultVec_dataGroup_32[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_32 = checkVec_checkResultVec_dataGroup_32[3:1];
  wire [2:0]         checkVec_checkResultVec_0_4_1 = checkVec_checkResultVec_accessRegGrowth_32;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_32 = {checkVec_checkResultVec_0_3_1, checkVec_checkResultVec_0_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_32 = checkVec_checkResultVec_decimalProportion_32[5:3];
  wire               checkVec_checkResultVec_overlap_32 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_32 >= checkVec_checkResultVec_intLMULInput_32[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_32} >= checkVec_checkResultVec_intLMULInput_32,
      source_0[31:11]};
  wire               checkVec_checkResultVec_0_5_1 = checkVec_checkResultVec_overlap_32 | ~checkVec_checkResultVec_0_6_1;
  wire               checkVec_checkResultVec_1_6_1 = checkVec_validVec_1[1];
  wire [10:0]        checkVec_checkResultVec_dataPosition_33 = {source_1[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_267 = 2'h1 << checkVec_checkResultVec_dataPosition_33[1];
  wire [3:0]         checkVec_checkResultVec_1_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_267[1]}}, {2{_checkVec_checkResultVec_accessMask_T_267[0]}}};
  wire [1:0]         checkVec_checkResultVec_1_1_1 = {checkVec_checkResultVec_dataPosition_33[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_1_2_1 = checkVec_checkResultVec_dataPosition_33[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_33 = checkVec_checkResultVec_dataPosition_33[10:7];
  wire               checkVec_checkResultVec_1_3_1 = checkVec_checkResultVec_dataGroup_33[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_33 = checkVec_checkResultVec_dataGroup_33[3:1];
  wire [2:0]         checkVec_checkResultVec_1_4_1 = checkVec_checkResultVec_accessRegGrowth_33;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_33 = {checkVec_checkResultVec_1_3_1, checkVec_checkResultVec_1_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_33 = checkVec_checkResultVec_decimalProportion_33[5:3];
  wire               checkVec_checkResultVec_overlap_33 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_33 >= checkVec_checkResultVec_intLMULInput_33[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_33} >= checkVec_checkResultVec_intLMULInput_33,
      source_1[31:11]};
  wire               checkVec_checkResultVec_1_5_1 = checkVec_checkResultVec_overlap_33 | ~checkVec_checkResultVec_1_6_1;
  wire               checkVec_checkResultVec_2_6_1 = checkVec_validVec_1[2];
  wire [10:0]        checkVec_checkResultVec_dataPosition_34 = {source_2[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_275 = 2'h1 << checkVec_checkResultVec_dataPosition_34[1];
  wire [3:0]         checkVec_checkResultVec_2_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_275[1]}}, {2{_checkVec_checkResultVec_accessMask_T_275[0]}}};
  wire [1:0]         checkVec_checkResultVec_2_1_1 = {checkVec_checkResultVec_dataPosition_34[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_2_2_1 = checkVec_checkResultVec_dataPosition_34[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_34 = checkVec_checkResultVec_dataPosition_34[10:7];
  wire               checkVec_checkResultVec_2_3_1 = checkVec_checkResultVec_dataGroup_34[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_34 = checkVec_checkResultVec_dataGroup_34[3:1];
  wire [2:0]         checkVec_checkResultVec_2_4_1 = checkVec_checkResultVec_accessRegGrowth_34;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_34 = {checkVec_checkResultVec_2_3_1, checkVec_checkResultVec_2_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_34 = checkVec_checkResultVec_decimalProportion_34[5:3];
  wire               checkVec_checkResultVec_overlap_34 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_34 >= checkVec_checkResultVec_intLMULInput_34[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_34} >= checkVec_checkResultVec_intLMULInput_34,
      source_2[31:11]};
  wire               checkVec_checkResultVec_2_5_1 = checkVec_checkResultVec_overlap_34 | ~checkVec_checkResultVec_2_6_1;
  wire               checkVec_checkResultVec_3_6_1 = checkVec_validVec_1[3];
  wire [10:0]        checkVec_checkResultVec_dataPosition_35 = {source_3[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_283 = 2'h1 << checkVec_checkResultVec_dataPosition_35[1];
  wire [3:0]         checkVec_checkResultVec_3_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_283[1]}}, {2{_checkVec_checkResultVec_accessMask_T_283[0]}}};
  wire [1:0]         checkVec_checkResultVec_3_1_1 = {checkVec_checkResultVec_dataPosition_35[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_3_2_1 = checkVec_checkResultVec_dataPosition_35[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_35 = checkVec_checkResultVec_dataPosition_35[10:7];
  wire               checkVec_checkResultVec_3_3_1 = checkVec_checkResultVec_dataGroup_35[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_35 = checkVec_checkResultVec_dataGroup_35[3:1];
  wire [2:0]         checkVec_checkResultVec_3_4_1 = checkVec_checkResultVec_accessRegGrowth_35;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_35 = {checkVec_checkResultVec_3_3_1, checkVec_checkResultVec_3_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_35 = checkVec_checkResultVec_decimalProportion_35[5:3];
  wire               checkVec_checkResultVec_overlap_35 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_35 >= checkVec_checkResultVec_intLMULInput_35[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_35} >= checkVec_checkResultVec_intLMULInput_35,
      source_3[31:11]};
  wire               checkVec_checkResultVec_3_5_1 = checkVec_checkResultVec_overlap_35 | ~checkVec_checkResultVec_3_6_1;
  wire               checkVec_checkResultVec_4_6_1 = checkVec_validVec_1[4];
  wire [10:0]        checkVec_checkResultVec_dataPosition_36 = {source_4[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_291 = 2'h1 << checkVec_checkResultVec_dataPosition_36[1];
  wire [3:0]         checkVec_checkResultVec_4_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_291[1]}}, {2{_checkVec_checkResultVec_accessMask_T_291[0]}}};
  wire [1:0]         checkVec_checkResultVec_4_1_1 = {checkVec_checkResultVec_dataPosition_36[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_4_2_1 = checkVec_checkResultVec_dataPosition_36[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_36 = checkVec_checkResultVec_dataPosition_36[10:7];
  wire               checkVec_checkResultVec_4_3_1 = checkVec_checkResultVec_dataGroup_36[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_36 = checkVec_checkResultVec_dataGroup_36[3:1];
  wire [2:0]         checkVec_checkResultVec_4_4_1 = checkVec_checkResultVec_accessRegGrowth_36;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_36 = {checkVec_checkResultVec_4_3_1, checkVec_checkResultVec_4_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_36 = checkVec_checkResultVec_decimalProportion_36[5:3];
  wire               checkVec_checkResultVec_overlap_36 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_36 >= checkVec_checkResultVec_intLMULInput_36[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_36} >= checkVec_checkResultVec_intLMULInput_36,
      source_4[31:11]};
  wire               checkVec_checkResultVec_4_5_1 = checkVec_checkResultVec_overlap_36 | ~checkVec_checkResultVec_4_6_1;
  wire               checkVec_checkResultVec_5_6_1 = checkVec_validVec_1[5];
  wire [10:0]        checkVec_checkResultVec_dataPosition_37 = {source_5[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_299 = 2'h1 << checkVec_checkResultVec_dataPosition_37[1];
  wire [3:0]         checkVec_checkResultVec_5_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_299[1]}}, {2{_checkVec_checkResultVec_accessMask_T_299[0]}}};
  wire [1:0]         checkVec_checkResultVec_5_1_1 = {checkVec_checkResultVec_dataPosition_37[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_5_2_1 = checkVec_checkResultVec_dataPosition_37[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_37 = checkVec_checkResultVec_dataPosition_37[10:7];
  wire               checkVec_checkResultVec_5_3_1 = checkVec_checkResultVec_dataGroup_37[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_37 = checkVec_checkResultVec_dataGroup_37[3:1];
  wire [2:0]         checkVec_checkResultVec_5_4_1 = checkVec_checkResultVec_accessRegGrowth_37;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_37 = {checkVec_checkResultVec_5_3_1, checkVec_checkResultVec_5_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_37 = checkVec_checkResultVec_decimalProportion_37[5:3];
  wire               checkVec_checkResultVec_overlap_37 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_37 >= checkVec_checkResultVec_intLMULInput_37[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_37} >= checkVec_checkResultVec_intLMULInput_37,
      source_5[31:11]};
  wire               checkVec_checkResultVec_5_5_1 = checkVec_checkResultVec_overlap_37 | ~checkVec_checkResultVec_5_6_1;
  wire               checkVec_checkResultVec_6_6_1 = checkVec_validVec_1[6];
  wire [10:0]        checkVec_checkResultVec_dataPosition_38 = {source_6[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_307 = 2'h1 << checkVec_checkResultVec_dataPosition_38[1];
  wire [3:0]         checkVec_checkResultVec_6_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_307[1]}}, {2{_checkVec_checkResultVec_accessMask_T_307[0]}}};
  wire [1:0]         checkVec_checkResultVec_6_1_1 = {checkVec_checkResultVec_dataPosition_38[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_6_2_1 = checkVec_checkResultVec_dataPosition_38[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_38 = checkVec_checkResultVec_dataPosition_38[10:7];
  wire               checkVec_checkResultVec_6_3_1 = checkVec_checkResultVec_dataGroup_38[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_38 = checkVec_checkResultVec_dataGroup_38[3:1];
  wire [2:0]         checkVec_checkResultVec_6_4_1 = checkVec_checkResultVec_accessRegGrowth_38;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_38 = {checkVec_checkResultVec_6_3_1, checkVec_checkResultVec_6_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_38 = checkVec_checkResultVec_decimalProportion_38[5:3];
  wire               checkVec_checkResultVec_overlap_38 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_38 >= checkVec_checkResultVec_intLMULInput_38[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_38} >= checkVec_checkResultVec_intLMULInput_38,
      source_6[31:11]};
  wire               checkVec_checkResultVec_6_5_1 = checkVec_checkResultVec_overlap_38 | ~checkVec_checkResultVec_6_6_1;
  wire               checkVec_checkResultVec_7_6_1 = checkVec_validVec_1[7];
  wire [10:0]        checkVec_checkResultVec_dataPosition_39 = {source_7[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_315 = 2'h1 << checkVec_checkResultVec_dataPosition_39[1];
  wire [3:0]         checkVec_checkResultVec_7_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_315[1]}}, {2{_checkVec_checkResultVec_accessMask_T_315[0]}}};
  wire [1:0]         checkVec_checkResultVec_7_1_1 = {checkVec_checkResultVec_dataPosition_39[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_7_2_1 = checkVec_checkResultVec_dataPosition_39[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_39 = checkVec_checkResultVec_dataPosition_39[10:7];
  wire               checkVec_checkResultVec_7_3_1 = checkVec_checkResultVec_dataGroup_39[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_39 = checkVec_checkResultVec_dataGroup_39[3:1];
  wire [2:0]         checkVec_checkResultVec_7_4_1 = checkVec_checkResultVec_accessRegGrowth_39;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_39 = {checkVec_checkResultVec_7_3_1, checkVec_checkResultVec_7_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_39 = checkVec_checkResultVec_decimalProportion_39[5:3];
  wire               checkVec_checkResultVec_overlap_39 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_39 >= checkVec_checkResultVec_intLMULInput_39[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_39} >= checkVec_checkResultVec_intLMULInput_39,
      source_7[31:11]};
  wire               checkVec_checkResultVec_7_5_1 = checkVec_checkResultVec_overlap_39 | ~checkVec_checkResultVec_7_6_1;
  wire               checkVec_checkResultVec_8_6_1 = checkVec_validVec_1[8];
  wire [10:0]        checkVec_checkResultVec_dataPosition_40 = {source_8[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_323 = 2'h1 << checkVec_checkResultVec_dataPosition_40[1];
  wire [3:0]         checkVec_checkResultVec_8_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_323[1]}}, {2{_checkVec_checkResultVec_accessMask_T_323[0]}}};
  wire [1:0]         checkVec_checkResultVec_8_1_1 = {checkVec_checkResultVec_dataPosition_40[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_8_2_1 = checkVec_checkResultVec_dataPosition_40[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_40 = checkVec_checkResultVec_dataPosition_40[10:7];
  wire               checkVec_checkResultVec_8_3_1 = checkVec_checkResultVec_dataGroup_40[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_40 = checkVec_checkResultVec_dataGroup_40[3:1];
  wire [2:0]         checkVec_checkResultVec_8_4_1 = checkVec_checkResultVec_accessRegGrowth_40;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_40 = {checkVec_checkResultVec_8_3_1, checkVec_checkResultVec_8_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_40 = checkVec_checkResultVec_decimalProportion_40[5:3];
  wire               checkVec_checkResultVec_overlap_40 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_40 >= checkVec_checkResultVec_intLMULInput_40[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_40} >= checkVec_checkResultVec_intLMULInput_40,
      source_8[31:11]};
  wire               checkVec_checkResultVec_8_5_1 = checkVec_checkResultVec_overlap_40 | ~checkVec_checkResultVec_8_6_1;
  wire               checkVec_checkResultVec_9_6_1 = checkVec_validVec_1[9];
  wire [10:0]        checkVec_checkResultVec_dataPosition_41 = {source_9[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_331 = 2'h1 << checkVec_checkResultVec_dataPosition_41[1];
  wire [3:0]         checkVec_checkResultVec_9_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_331[1]}}, {2{_checkVec_checkResultVec_accessMask_T_331[0]}}};
  wire [1:0]         checkVec_checkResultVec_9_1_1 = {checkVec_checkResultVec_dataPosition_41[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_9_2_1 = checkVec_checkResultVec_dataPosition_41[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_41 = checkVec_checkResultVec_dataPosition_41[10:7];
  wire               checkVec_checkResultVec_9_3_1 = checkVec_checkResultVec_dataGroup_41[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_41 = checkVec_checkResultVec_dataGroup_41[3:1];
  wire [2:0]         checkVec_checkResultVec_9_4_1 = checkVec_checkResultVec_accessRegGrowth_41;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_41 = {checkVec_checkResultVec_9_3_1, checkVec_checkResultVec_9_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_41 = checkVec_checkResultVec_decimalProportion_41[5:3];
  wire               checkVec_checkResultVec_overlap_41 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_41 >= checkVec_checkResultVec_intLMULInput_41[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_41} >= checkVec_checkResultVec_intLMULInput_41,
      source_9[31:11]};
  wire               checkVec_checkResultVec_9_5_1 = checkVec_checkResultVec_overlap_41 | ~checkVec_checkResultVec_9_6_1;
  wire               checkVec_checkResultVec_10_6_1 = checkVec_validVec_1[10];
  wire [10:0]        checkVec_checkResultVec_dataPosition_42 = {source_10[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_339 = 2'h1 << checkVec_checkResultVec_dataPosition_42[1];
  wire [3:0]         checkVec_checkResultVec_10_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_339[1]}}, {2{_checkVec_checkResultVec_accessMask_T_339[0]}}};
  wire [1:0]         checkVec_checkResultVec_10_1_1 = {checkVec_checkResultVec_dataPosition_42[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_10_2_1 = checkVec_checkResultVec_dataPosition_42[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_42 = checkVec_checkResultVec_dataPosition_42[10:7];
  wire               checkVec_checkResultVec_10_3_1 = checkVec_checkResultVec_dataGroup_42[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_42 = checkVec_checkResultVec_dataGroup_42[3:1];
  wire [2:0]         checkVec_checkResultVec_10_4_1 = checkVec_checkResultVec_accessRegGrowth_42;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_42 = {checkVec_checkResultVec_10_3_1, checkVec_checkResultVec_10_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_42 = checkVec_checkResultVec_decimalProportion_42[5:3];
  wire               checkVec_checkResultVec_overlap_42 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_42 >= checkVec_checkResultVec_intLMULInput_42[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_42} >= checkVec_checkResultVec_intLMULInput_42,
      source_10[31:11]};
  wire               checkVec_checkResultVec_10_5_1 = checkVec_checkResultVec_overlap_42 | ~checkVec_checkResultVec_10_6_1;
  wire               checkVec_checkResultVec_11_6_1 = checkVec_validVec_1[11];
  wire [10:0]        checkVec_checkResultVec_dataPosition_43 = {source_11[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_347 = 2'h1 << checkVec_checkResultVec_dataPosition_43[1];
  wire [3:0]         checkVec_checkResultVec_11_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_347[1]}}, {2{_checkVec_checkResultVec_accessMask_T_347[0]}}};
  wire [1:0]         checkVec_checkResultVec_11_1_1 = {checkVec_checkResultVec_dataPosition_43[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_11_2_1 = checkVec_checkResultVec_dataPosition_43[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_43 = checkVec_checkResultVec_dataPosition_43[10:7];
  wire               checkVec_checkResultVec_11_3_1 = checkVec_checkResultVec_dataGroup_43[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_43 = checkVec_checkResultVec_dataGroup_43[3:1];
  wire [2:0]         checkVec_checkResultVec_11_4_1 = checkVec_checkResultVec_accessRegGrowth_43;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_43 = {checkVec_checkResultVec_11_3_1, checkVec_checkResultVec_11_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_43 = checkVec_checkResultVec_decimalProportion_43[5:3];
  wire               checkVec_checkResultVec_overlap_43 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_43 >= checkVec_checkResultVec_intLMULInput_43[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_43} >= checkVec_checkResultVec_intLMULInput_43,
      source_11[31:11]};
  wire               checkVec_checkResultVec_11_5_1 = checkVec_checkResultVec_overlap_43 | ~checkVec_checkResultVec_11_6_1;
  wire               checkVec_checkResultVec_12_6_1 = checkVec_validVec_1[12];
  wire [10:0]        checkVec_checkResultVec_dataPosition_44 = {source_12[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_355 = 2'h1 << checkVec_checkResultVec_dataPosition_44[1];
  wire [3:0]         checkVec_checkResultVec_12_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_355[1]}}, {2{_checkVec_checkResultVec_accessMask_T_355[0]}}};
  wire [1:0]         checkVec_checkResultVec_12_1_1 = {checkVec_checkResultVec_dataPosition_44[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_12_2_1 = checkVec_checkResultVec_dataPosition_44[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_44 = checkVec_checkResultVec_dataPosition_44[10:7];
  wire               checkVec_checkResultVec_12_3_1 = checkVec_checkResultVec_dataGroup_44[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_44 = checkVec_checkResultVec_dataGroup_44[3:1];
  wire [2:0]         checkVec_checkResultVec_12_4_1 = checkVec_checkResultVec_accessRegGrowth_44;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_44 = {checkVec_checkResultVec_12_3_1, checkVec_checkResultVec_12_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_44 = checkVec_checkResultVec_decimalProportion_44[5:3];
  wire               checkVec_checkResultVec_overlap_44 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_44 >= checkVec_checkResultVec_intLMULInput_44[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_44} >= checkVec_checkResultVec_intLMULInput_44,
      source_12[31:11]};
  wire               checkVec_checkResultVec_12_5_1 = checkVec_checkResultVec_overlap_44 | ~checkVec_checkResultVec_12_6_1;
  wire               checkVec_checkResultVec_13_6_1 = checkVec_validVec_1[13];
  wire [10:0]        checkVec_checkResultVec_dataPosition_45 = {source_13[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_363 = 2'h1 << checkVec_checkResultVec_dataPosition_45[1];
  wire [3:0]         checkVec_checkResultVec_13_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_363[1]}}, {2{_checkVec_checkResultVec_accessMask_T_363[0]}}};
  wire [1:0]         checkVec_checkResultVec_13_1_1 = {checkVec_checkResultVec_dataPosition_45[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_13_2_1 = checkVec_checkResultVec_dataPosition_45[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_45 = checkVec_checkResultVec_dataPosition_45[10:7];
  wire               checkVec_checkResultVec_13_3_1 = checkVec_checkResultVec_dataGroup_45[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_45 = checkVec_checkResultVec_dataGroup_45[3:1];
  wire [2:0]         checkVec_checkResultVec_13_4_1 = checkVec_checkResultVec_accessRegGrowth_45;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_45 = {checkVec_checkResultVec_13_3_1, checkVec_checkResultVec_13_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_45 = checkVec_checkResultVec_decimalProportion_45[5:3];
  wire               checkVec_checkResultVec_overlap_45 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_45 >= checkVec_checkResultVec_intLMULInput_45[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_45} >= checkVec_checkResultVec_intLMULInput_45,
      source_13[31:11]};
  wire               checkVec_checkResultVec_13_5_1 = checkVec_checkResultVec_overlap_45 | ~checkVec_checkResultVec_13_6_1;
  wire               checkVec_checkResultVec_14_6_1 = checkVec_validVec_1[14];
  wire [10:0]        checkVec_checkResultVec_dataPosition_46 = {source_14[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_371 = 2'h1 << checkVec_checkResultVec_dataPosition_46[1];
  wire [3:0]         checkVec_checkResultVec_14_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_371[1]}}, {2{_checkVec_checkResultVec_accessMask_T_371[0]}}};
  wire [1:0]         checkVec_checkResultVec_14_1_1 = {checkVec_checkResultVec_dataPosition_46[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_14_2_1 = checkVec_checkResultVec_dataPosition_46[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_46 = checkVec_checkResultVec_dataPosition_46[10:7];
  wire               checkVec_checkResultVec_14_3_1 = checkVec_checkResultVec_dataGroup_46[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_46 = checkVec_checkResultVec_dataGroup_46[3:1];
  wire [2:0]         checkVec_checkResultVec_14_4_1 = checkVec_checkResultVec_accessRegGrowth_46;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_46 = {checkVec_checkResultVec_14_3_1, checkVec_checkResultVec_14_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_46 = checkVec_checkResultVec_decimalProportion_46[5:3];
  wire               checkVec_checkResultVec_overlap_46 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_46 >= checkVec_checkResultVec_intLMULInput_46[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_46} >= checkVec_checkResultVec_intLMULInput_46,
      source_14[31:11]};
  wire               checkVec_checkResultVec_14_5_1 = checkVec_checkResultVec_overlap_46 | ~checkVec_checkResultVec_14_6_1;
  wire               checkVec_checkResultVec_15_6_1 = checkVec_validVec_1[15];
  wire [10:0]        checkVec_checkResultVec_dataPosition_47 = {source_15[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_379 = 2'h1 << checkVec_checkResultVec_dataPosition_47[1];
  wire [3:0]         checkVec_checkResultVec_15_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_379[1]}}, {2{_checkVec_checkResultVec_accessMask_T_379[0]}}};
  wire [1:0]         checkVec_checkResultVec_15_1_1 = {checkVec_checkResultVec_dataPosition_47[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_15_2_1 = checkVec_checkResultVec_dataPosition_47[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_47 = checkVec_checkResultVec_dataPosition_47[10:7];
  wire               checkVec_checkResultVec_15_3_1 = checkVec_checkResultVec_dataGroup_47[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_47 = checkVec_checkResultVec_dataGroup_47[3:1];
  wire [2:0]         checkVec_checkResultVec_15_4_1 = checkVec_checkResultVec_accessRegGrowth_47;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_47 = {checkVec_checkResultVec_15_3_1, checkVec_checkResultVec_15_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_47 = checkVec_checkResultVec_decimalProportion_47[5:3];
  wire               checkVec_checkResultVec_overlap_47 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_47 >= checkVec_checkResultVec_intLMULInput_47[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_47} >= checkVec_checkResultVec_intLMULInput_47,
      source_15[31:11]};
  wire               checkVec_checkResultVec_15_5_1 = checkVec_checkResultVec_overlap_47 | ~checkVec_checkResultVec_15_6_1;
  wire               checkVec_checkResultVec_16_6_1 = checkVec_validVec_1[16];
  wire [10:0]        checkVec_checkResultVec_dataPosition_48 = {source_16[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_387 = 2'h1 << checkVec_checkResultVec_dataPosition_48[1];
  wire [3:0]         checkVec_checkResultVec_16_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_387[1]}}, {2{_checkVec_checkResultVec_accessMask_T_387[0]}}};
  wire [1:0]         checkVec_checkResultVec_16_1_1 = {checkVec_checkResultVec_dataPosition_48[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_16_2_1 = checkVec_checkResultVec_dataPosition_48[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_48 = checkVec_checkResultVec_dataPosition_48[10:7];
  wire               checkVec_checkResultVec_16_3_1 = checkVec_checkResultVec_dataGroup_48[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_48 = checkVec_checkResultVec_dataGroup_48[3:1];
  wire [2:0]         checkVec_checkResultVec_16_4_1 = checkVec_checkResultVec_accessRegGrowth_48;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_48 = {checkVec_checkResultVec_16_3_1, checkVec_checkResultVec_16_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_48 = checkVec_checkResultVec_decimalProportion_48[5:3];
  wire               checkVec_checkResultVec_overlap_48 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_48 >= checkVec_checkResultVec_intLMULInput_48[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_48} >= checkVec_checkResultVec_intLMULInput_48,
      source_16[31:11]};
  wire               checkVec_checkResultVec_16_5_1 = checkVec_checkResultVec_overlap_48 | ~checkVec_checkResultVec_16_6_1;
  wire               checkVec_checkResultVec_17_6_1 = checkVec_validVec_1[17];
  wire [10:0]        checkVec_checkResultVec_dataPosition_49 = {source_17[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_395 = 2'h1 << checkVec_checkResultVec_dataPosition_49[1];
  wire [3:0]         checkVec_checkResultVec_17_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_395[1]}}, {2{_checkVec_checkResultVec_accessMask_T_395[0]}}};
  wire [1:0]         checkVec_checkResultVec_17_1_1 = {checkVec_checkResultVec_dataPosition_49[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_17_2_1 = checkVec_checkResultVec_dataPosition_49[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_49 = checkVec_checkResultVec_dataPosition_49[10:7];
  wire               checkVec_checkResultVec_17_3_1 = checkVec_checkResultVec_dataGroup_49[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_49 = checkVec_checkResultVec_dataGroup_49[3:1];
  wire [2:0]         checkVec_checkResultVec_17_4_1 = checkVec_checkResultVec_accessRegGrowth_49;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_49 = {checkVec_checkResultVec_17_3_1, checkVec_checkResultVec_17_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_49 = checkVec_checkResultVec_decimalProportion_49[5:3];
  wire               checkVec_checkResultVec_overlap_49 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_49 >= checkVec_checkResultVec_intLMULInput_49[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_49} >= checkVec_checkResultVec_intLMULInput_49,
      source_17[31:11]};
  wire               checkVec_checkResultVec_17_5_1 = checkVec_checkResultVec_overlap_49 | ~checkVec_checkResultVec_17_6_1;
  wire               checkVec_checkResultVec_18_6_1 = checkVec_validVec_1[18];
  wire [10:0]        checkVec_checkResultVec_dataPosition_50 = {source_18[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_403 = 2'h1 << checkVec_checkResultVec_dataPosition_50[1];
  wire [3:0]         checkVec_checkResultVec_18_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_403[1]}}, {2{_checkVec_checkResultVec_accessMask_T_403[0]}}};
  wire [1:0]         checkVec_checkResultVec_18_1_1 = {checkVec_checkResultVec_dataPosition_50[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_18_2_1 = checkVec_checkResultVec_dataPosition_50[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_50 = checkVec_checkResultVec_dataPosition_50[10:7];
  wire               checkVec_checkResultVec_18_3_1 = checkVec_checkResultVec_dataGroup_50[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_50 = checkVec_checkResultVec_dataGroup_50[3:1];
  wire [2:0]         checkVec_checkResultVec_18_4_1 = checkVec_checkResultVec_accessRegGrowth_50;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_50 = {checkVec_checkResultVec_18_3_1, checkVec_checkResultVec_18_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_50 = checkVec_checkResultVec_decimalProportion_50[5:3];
  wire               checkVec_checkResultVec_overlap_50 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_50 >= checkVec_checkResultVec_intLMULInput_50[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_50} >= checkVec_checkResultVec_intLMULInput_50,
      source_18[31:11]};
  wire               checkVec_checkResultVec_18_5_1 = checkVec_checkResultVec_overlap_50 | ~checkVec_checkResultVec_18_6_1;
  wire               checkVec_checkResultVec_19_6_1 = checkVec_validVec_1[19];
  wire [10:0]        checkVec_checkResultVec_dataPosition_51 = {source_19[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_411 = 2'h1 << checkVec_checkResultVec_dataPosition_51[1];
  wire [3:0]         checkVec_checkResultVec_19_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_411[1]}}, {2{_checkVec_checkResultVec_accessMask_T_411[0]}}};
  wire [1:0]         checkVec_checkResultVec_19_1_1 = {checkVec_checkResultVec_dataPosition_51[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_19_2_1 = checkVec_checkResultVec_dataPosition_51[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_51 = checkVec_checkResultVec_dataPosition_51[10:7];
  wire               checkVec_checkResultVec_19_3_1 = checkVec_checkResultVec_dataGroup_51[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_51 = checkVec_checkResultVec_dataGroup_51[3:1];
  wire [2:0]         checkVec_checkResultVec_19_4_1 = checkVec_checkResultVec_accessRegGrowth_51;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_51 = {checkVec_checkResultVec_19_3_1, checkVec_checkResultVec_19_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_51 = checkVec_checkResultVec_decimalProportion_51[5:3];
  wire               checkVec_checkResultVec_overlap_51 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_51 >= checkVec_checkResultVec_intLMULInput_51[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_51} >= checkVec_checkResultVec_intLMULInput_51,
      source_19[31:11]};
  wire               checkVec_checkResultVec_19_5_1 = checkVec_checkResultVec_overlap_51 | ~checkVec_checkResultVec_19_6_1;
  wire               checkVec_checkResultVec_20_6_1 = checkVec_validVec_1[20];
  wire [10:0]        checkVec_checkResultVec_dataPosition_52 = {source_20[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_419 = 2'h1 << checkVec_checkResultVec_dataPosition_52[1];
  wire [3:0]         checkVec_checkResultVec_20_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_419[1]}}, {2{_checkVec_checkResultVec_accessMask_T_419[0]}}};
  wire [1:0]         checkVec_checkResultVec_20_1_1 = {checkVec_checkResultVec_dataPosition_52[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_20_2_1 = checkVec_checkResultVec_dataPosition_52[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_52 = checkVec_checkResultVec_dataPosition_52[10:7];
  wire               checkVec_checkResultVec_20_3_1 = checkVec_checkResultVec_dataGroup_52[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_52 = checkVec_checkResultVec_dataGroup_52[3:1];
  wire [2:0]         checkVec_checkResultVec_20_4_1 = checkVec_checkResultVec_accessRegGrowth_52;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_52 = {checkVec_checkResultVec_20_3_1, checkVec_checkResultVec_20_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_52 = checkVec_checkResultVec_decimalProportion_52[5:3];
  wire               checkVec_checkResultVec_overlap_52 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_52 >= checkVec_checkResultVec_intLMULInput_52[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_52} >= checkVec_checkResultVec_intLMULInput_52,
      source_20[31:11]};
  wire               checkVec_checkResultVec_20_5_1 = checkVec_checkResultVec_overlap_52 | ~checkVec_checkResultVec_20_6_1;
  wire               checkVec_checkResultVec_21_6_1 = checkVec_validVec_1[21];
  wire [10:0]        checkVec_checkResultVec_dataPosition_53 = {source_21[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_427 = 2'h1 << checkVec_checkResultVec_dataPosition_53[1];
  wire [3:0]         checkVec_checkResultVec_21_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_427[1]}}, {2{_checkVec_checkResultVec_accessMask_T_427[0]}}};
  wire [1:0]         checkVec_checkResultVec_21_1_1 = {checkVec_checkResultVec_dataPosition_53[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_21_2_1 = checkVec_checkResultVec_dataPosition_53[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_53 = checkVec_checkResultVec_dataPosition_53[10:7];
  wire               checkVec_checkResultVec_21_3_1 = checkVec_checkResultVec_dataGroup_53[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_53 = checkVec_checkResultVec_dataGroup_53[3:1];
  wire [2:0]         checkVec_checkResultVec_21_4_1 = checkVec_checkResultVec_accessRegGrowth_53;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_53 = {checkVec_checkResultVec_21_3_1, checkVec_checkResultVec_21_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_53 = checkVec_checkResultVec_decimalProportion_53[5:3];
  wire               checkVec_checkResultVec_overlap_53 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_53 >= checkVec_checkResultVec_intLMULInput_53[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_53} >= checkVec_checkResultVec_intLMULInput_53,
      source_21[31:11]};
  wire               checkVec_checkResultVec_21_5_1 = checkVec_checkResultVec_overlap_53 | ~checkVec_checkResultVec_21_6_1;
  wire               checkVec_checkResultVec_22_6_1 = checkVec_validVec_1[22];
  wire [10:0]        checkVec_checkResultVec_dataPosition_54 = {source_22[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_435 = 2'h1 << checkVec_checkResultVec_dataPosition_54[1];
  wire [3:0]         checkVec_checkResultVec_22_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_435[1]}}, {2{_checkVec_checkResultVec_accessMask_T_435[0]}}};
  wire [1:0]         checkVec_checkResultVec_22_1_1 = {checkVec_checkResultVec_dataPosition_54[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_22_2_1 = checkVec_checkResultVec_dataPosition_54[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_54 = checkVec_checkResultVec_dataPosition_54[10:7];
  wire               checkVec_checkResultVec_22_3_1 = checkVec_checkResultVec_dataGroup_54[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_54 = checkVec_checkResultVec_dataGroup_54[3:1];
  wire [2:0]         checkVec_checkResultVec_22_4_1 = checkVec_checkResultVec_accessRegGrowth_54;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_54 = {checkVec_checkResultVec_22_3_1, checkVec_checkResultVec_22_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_54 = checkVec_checkResultVec_decimalProportion_54[5:3];
  wire               checkVec_checkResultVec_overlap_54 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_54 >= checkVec_checkResultVec_intLMULInput_54[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_54} >= checkVec_checkResultVec_intLMULInput_54,
      source_22[31:11]};
  wire               checkVec_checkResultVec_22_5_1 = checkVec_checkResultVec_overlap_54 | ~checkVec_checkResultVec_22_6_1;
  wire               checkVec_checkResultVec_23_6_1 = checkVec_validVec_1[23];
  wire [10:0]        checkVec_checkResultVec_dataPosition_55 = {source_23[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_443 = 2'h1 << checkVec_checkResultVec_dataPosition_55[1];
  wire [3:0]         checkVec_checkResultVec_23_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_443[1]}}, {2{_checkVec_checkResultVec_accessMask_T_443[0]}}};
  wire [1:0]         checkVec_checkResultVec_23_1_1 = {checkVec_checkResultVec_dataPosition_55[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_23_2_1 = checkVec_checkResultVec_dataPosition_55[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_55 = checkVec_checkResultVec_dataPosition_55[10:7];
  wire               checkVec_checkResultVec_23_3_1 = checkVec_checkResultVec_dataGroup_55[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_55 = checkVec_checkResultVec_dataGroup_55[3:1];
  wire [2:0]         checkVec_checkResultVec_23_4_1 = checkVec_checkResultVec_accessRegGrowth_55;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_55 = {checkVec_checkResultVec_23_3_1, checkVec_checkResultVec_23_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_55 = checkVec_checkResultVec_decimalProportion_55[5:3];
  wire               checkVec_checkResultVec_overlap_55 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_55 >= checkVec_checkResultVec_intLMULInput_55[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_55} >= checkVec_checkResultVec_intLMULInput_55,
      source_23[31:11]};
  wire               checkVec_checkResultVec_23_5_1 = checkVec_checkResultVec_overlap_55 | ~checkVec_checkResultVec_23_6_1;
  wire               checkVec_checkResultVec_24_6_1 = checkVec_validVec_1[24];
  wire [10:0]        checkVec_checkResultVec_dataPosition_56 = {source_24[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_451 = 2'h1 << checkVec_checkResultVec_dataPosition_56[1];
  wire [3:0]         checkVec_checkResultVec_24_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_451[1]}}, {2{_checkVec_checkResultVec_accessMask_T_451[0]}}};
  wire [1:0]         checkVec_checkResultVec_24_1_1 = {checkVec_checkResultVec_dataPosition_56[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_24_2_1 = checkVec_checkResultVec_dataPosition_56[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_56 = checkVec_checkResultVec_dataPosition_56[10:7];
  wire               checkVec_checkResultVec_24_3_1 = checkVec_checkResultVec_dataGroup_56[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_56 = checkVec_checkResultVec_dataGroup_56[3:1];
  wire [2:0]         checkVec_checkResultVec_24_4_1 = checkVec_checkResultVec_accessRegGrowth_56;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_56 = {checkVec_checkResultVec_24_3_1, checkVec_checkResultVec_24_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_56 = checkVec_checkResultVec_decimalProportion_56[5:3];
  wire               checkVec_checkResultVec_overlap_56 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_56 >= checkVec_checkResultVec_intLMULInput_56[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_56} >= checkVec_checkResultVec_intLMULInput_56,
      source_24[31:11]};
  wire               checkVec_checkResultVec_24_5_1 = checkVec_checkResultVec_overlap_56 | ~checkVec_checkResultVec_24_6_1;
  wire               checkVec_checkResultVec_25_6_1 = checkVec_validVec_1[25];
  wire [10:0]        checkVec_checkResultVec_dataPosition_57 = {source_25[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_459 = 2'h1 << checkVec_checkResultVec_dataPosition_57[1];
  wire [3:0]         checkVec_checkResultVec_25_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_459[1]}}, {2{_checkVec_checkResultVec_accessMask_T_459[0]}}};
  wire [1:0]         checkVec_checkResultVec_25_1_1 = {checkVec_checkResultVec_dataPosition_57[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_25_2_1 = checkVec_checkResultVec_dataPosition_57[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_57 = checkVec_checkResultVec_dataPosition_57[10:7];
  wire               checkVec_checkResultVec_25_3_1 = checkVec_checkResultVec_dataGroup_57[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_57 = checkVec_checkResultVec_dataGroup_57[3:1];
  wire [2:0]         checkVec_checkResultVec_25_4_1 = checkVec_checkResultVec_accessRegGrowth_57;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_57 = {checkVec_checkResultVec_25_3_1, checkVec_checkResultVec_25_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_57 = checkVec_checkResultVec_decimalProportion_57[5:3];
  wire               checkVec_checkResultVec_overlap_57 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_57 >= checkVec_checkResultVec_intLMULInput_57[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_57} >= checkVec_checkResultVec_intLMULInput_57,
      source_25[31:11]};
  wire               checkVec_checkResultVec_25_5_1 = checkVec_checkResultVec_overlap_57 | ~checkVec_checkResultVec_25_6_1;
  wire               checkVec_checkResultVec_26_6_1 = checkVec_validVec_1[26];
  wire [10:0]        checkVec_checkResultVec_dataPosition_58 = {source_26[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_467 = 2'h1 << checkVec_checkResultVec_dataPosition_58[1];
  wire [3:0]         checkVec_checkResultVec_26_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_467[1]}}, {2{_checkVec_checkResultVec_accessMask_T_467[0]}}};
  wire [1:0]         checkVec_checkResultVec_26_1_1 = {checkVec_checkResultVec_dataPosition_58[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_26_2_1 = checkVec_checkResultVec_dataPosition_58[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_58 = checkVec_checkResultVec_dataPosition_58[10:7];
  wire               checkVec_checkResultVec_26_3_1 = checkVec_checkResultVec_dataGroup_58[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_58 = checkVec_checkResultVec_dataGroup_58[3:1];
  wire [2:0]         checkVec_checkResultVec_26_4_1 = checkVec_checkResultVec_accessRegGrowth_58;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_58 = {checkVec_checkResultVec_26_3_1, checkVec_checkResultVec_26_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_58 = checkVec_checkResultVec_decimalProportion_58[5:3];
  wire               checkVec_checkResultVec_overlap_58 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_58 >= checkVec_checkResultVec_intLMULInput_58[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_58} >= checkVec_checkResultVec_intLMULInput_58,
      source_26[31:11]};
  wire               checkVec_checkResultVec_26_5_1 = checkVec_checkResultVec_overlap_58 | ~checkVec_checkResultVec_26_6_1;
  wire               checkVec_checkResultVec_27_6_1 = checkVec_validVec_1[27];
  wire [10:0]        checkVec_checkResultVec_dataPosition_59 = {source_27[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_475 = 2'h1 << checkVec_checkResultVec_dataPosition_59[1];
  wire [3:0]         checkVec_checkResultVec_27_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_475[1]}}, {2{_checkVec_checkResultVec_accessMask_T_475[0]}}};
  wire [1:0]         checkVec_checkResultVec_27_1_1 = {checkVec_checkResultVec_dataPosition_59[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_27_2_1 = checkVec_checkResultVec_dataPosition_59[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_59 = checkVec_checkResultVec_dataPosition_59[10:7];
  wire               checkVec_checkResultVec_27_3_1 = checkVec_checkResultVec_dataGroup_59[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_59 = checkVec_checkResultVec_dataGroup_59[3:1];
  wire [2:0]         checkVec_checkResultVec_27_4_1 = checkVec_checkResultVec_accessRegGrowth_59;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_59 = {checkVec_checkResultVec_27_3_1, checkVec_checkResultVec_27_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_59 = checkVec_checkResultVec_decimalProportion_59[5:3];
  wire               checkVec_checkResultVec_overlap_59 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_59 >= checkVec_checkResultVec_intLMULInput_59[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_59} >= checkVec_checkResultVec_intLMULInput_59,
      source_27[31:11]};
  wire               checkVec_checkResultVec_27_5_1 = checkVec_checkResultVec_overlap_59 | ~checkVec_checkResultVec_27_6_1;
  wire               checkVec_checkResultVec_28_6_1 = checkVec_validVec_1[28];
  wire [10:0]        checkVec_checkResultVec_dataPosition_60 = {source_28[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_483 = 2'h1 << checkVec_checkResultVec_dataPosition_60[1];
  wire [3:0]         checkVec_checkResultVec_28_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_483[1]}}, {2{_checkVec_checkResultVec_accessMask_T_483[0]}}};
  wire [1:0]         checkVec_checkResultVec_28_1_1 = {checkVec_checkResultVec_dataPosition_60[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_28_2_1 = checkVec_checkResultVec_dataPosition_60[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_60 = checkVec_checkResultVec_dataPosition_60[10:7];
  wire               checkVec_checkResultVec_28_3_1 = checkVec_checkResultVec_dataGroup_60[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_60 = checkVec_checkResultVec_dataGroup_60[3:1];
  wire [2:0]         checkVec_checkResultVec_28_4_1 = checkVec_checkResultVec_accessRegGrowth_60;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_60 = {checkVec_checkResultVec_28_3_1, checkVec_checkResultVec_28_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_60 = checkVec_checkResultVec_decimalProportion_60[5:3];
  wire               checkVec_checkResultVec_overlap_60 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_60 >= checkVec_checkResultVec_intLMULInput_60[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_60} >= checkVec_checkResultVec_intLMULInput_60,
      source_28[31:11]};
  wire               checkVec_checkResultVec_28_5_1 = checkVec_checkResultVec_overlap_60 | ~checkVec_checkResultVec_28_6_1;
  wire               checkVec_checkResultVec_29_6_1 = checkVec_validVec_1[29];
  wire [10:0]        checkVec_checkResultVec_dataPosition_61 = {source_29[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_491 = 2'h1 << checkVec_checkResultVec_dataPosition_61[1];
  wire [3:0]         checkVec_checkResultVec_29_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_491[1]}}, {2{_checkVec_checkResultVec_accessMask_T_491[0]}}};
  wire [1:0]         checkVec_checkResultVec_29_1_1 = {checkVec_checkResultVec_dataPosition_61[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_29_2_1 = checkVec_checkResultVec_dataPosition_61[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_61 = checkVec_checkResultVec_dataPosition_61[10:7];
  wire               checkVec_checkResultVec_29_3_1 = checkVec_checkResultVec_dataGroup_61[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_61 = checkVec_checkResultVec_dataGroup_61[3:1];
  wire [2:0]         checkVec_checkResultVec_29_4_1 = checkVec_checkResultVec_accessRegGrowth_61;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_61 = {checkVec_checkResultVec_29_3_1, checkVec_checkResultVec_29_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_61 = checkVec_checkResultVec_decimalProportion_61[5:3];
  wire               checkVec_checkResultVec_overlap_61 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_61 >= checkVec_checkResultVec_intLMULInput_61[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_61} >= checkVec_checkResultVec_intLMULInput_61,
      source_29[31:11]};
  wire               checkVec_checkResultVec_29_5_1 = checkVec_checkResultVec_overlap_61 | ~checkVec_checkResultVec_29_6_1;
  wire               checkVec_checkResultVec_30_6_1 = checkVec_validVec_1[30];
  wire [10:0]        checkVec_checkResultVec_dataPosition_62 = {source_30[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_499 = 2'h1 << checkVec_checkResultVec_dataPosition_62[1];
  wire [3:0]         checkVec_checkResultVec_30_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_499[1]}}, {2{_checkVec_checkResultVec_accessMask_T_499[0]}}};
  wire [1:0]         checkVec_checkResultVec_30_1_1 = {checkVec_checkResultVec_dataPosition_62[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_30_2_1 = checkVec_checkResultVec_dataPosition_62[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_62 = checkVec_checkResultVec_dataPosition_62[10:7];
  wire               checkVec_checkResultVec_30_3_1 = checkVec_checkResultVec_dataGroup_62[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_62 = checkVec_checkResultVec_dataGroup_62[3:1];
  wire [2:0]         checkVec_checkResultVec_30_4_1 = checkVec_checkResultVec_accessRegGrowth_62;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_62 = {checkVec_checkResultVec_30_3_1, checkVec_checkResultVec_30_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_62 = checkVec_checkResultVec_decimalProportion_62[5:3];
  wire               checkVec_checkResultVec_overlap_62 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_62 >= checkVec_checkResultVec_intLMULInput_62[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_62} >= checkVec_checkResultVec_intLMULInput_62,
      source_30[31:11]};
  wire               checkVec_checkResultVec_30_5_1 = checkVec_checkResultVec_overlap_62 | ~checkVec_checkResultVec_30_6_1;
  wire               checkVec_checkResultVec_31_6_1 = checkVec_validVec_1[31];
  wire [10:0]        checkVec_checkResultVec_dataPosition_63 = {source_31[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_507 = 2'h1 << checkVec_checkResultVec_dataPosition_63[1];
  wire [3:0]         checkVec_checkResultVec_31_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_507[1]}}, {2{_checkVec_checkResultVec_accessMask_T_507[0]}}};
  wire [1:0]         checkVec_checkResultVec_31_1_1 = {checkVec_checkResultVec_dataPosition_63[1], 1'h0};
  wire [4:0]         checkVec_checkResultVec_31_2_1 = checkVec_checkResultVec_dataPosition_63[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_63 = checkVec_checkResultVec_dataPosition_63[10:7];
  wire               checkVec_checkResultVec_31_3_1 = checkVec_checkResultVec_dataGroup_63[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_63 = checkVec_checkResultVec_dataGroup_63[3:1];
  wire [2:0]         checkVec_checkResultVec_31_4_1 = checkVec_checkResultVec_accessRegGrowth_63;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_63 = {checkVec_checkResultVec_31_3_1, checkVec_checkResultVec_31_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_63 = checkVec_checkResultVec_decimalProportion_63[5:3];
  wire               checkVec_checkResultVec_overlap_63 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_63 >= checkVec_checkResultVec_intLMULInput_63[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_63} >= checkVec_checkResultVec_intLMULInput_63,
      source_31[31:11]};
  wire               checkVec_checkResultVec_31_5_1 = checkVec_checkResultVec_overlap_63 | ~checkVec_checkResultVec_31_6_1;
  wire [7:0]         checkVec_checkResult_lo_lo_lo_lo_7 = {checkVec_checkResultVec_1_0_1, checkVec_checkResultVec_0_0_1};
  wire [7:0]         checkVec_checkResult_lo_lo_lo_hi_7 = {checkVec_checkResultVec_3_0_1, checkVec_checkResultVec_2_0_1};
  wire [15:0]        checkVec_checkResult_lo_lo_lo_7 = {checkVec_checkResult_lo_lo_lo_hi_7, checkVec_checkResult_lo_lo_lo_lo_7};
  wire [7:0]         checkVec_checkResult_lo_lo_hi_lo_7 = {checkVec_checkResultVec_5_0_1, checkVec_checkResultVec_4_0_1};
  wire [7:0]         checkVec_checkResult_lo_lo_hi_hi_7 = {checkVec_checkResultVec_7_0_1, checkVec_checkResultVec_6_0_1};
  wire [15:0]        checkVec_checkResult_lo_lo_hi_7 = {checkVec_checkResult_lo_lo_hi_hi_7, checkVec_checkResult_lo_lo_hi_lo_7};
  wire [31:0]        checkVec_checkResult_lo_lo_7 = {checkVec_checkResult_lo_lo_hi_7, checkVec_checkResult_lo_lo_lo_7};
  wire [7:0]         checkVec_checkResult_lo_hi_lo_lo_7 = {checkVec_checkResultVec_9_0_1, checkVec_checkResultVec_8_0_1};
  wire [7:0]         checkVec_checkResult_lo_hi_lo_hi_7 = {checkVec_checkResultVec_11_0_1, checkVec_checkResultVec_10_0_1};
  wire [15:0]        checkVec_checkResult_lo_hi_lo_7 = {checkVec_checkResult_lo_hi_lo_hi_7, checkVec_checkResult_lo_hi_lo_lo_7};
  wire [7:0]         checkVec_checkResult_lo_hi_hi_lo_7 = {checkVec_checkResultVec_13_0_1, checkVec_checkResultVec_12_0_1};
  wire [7:0]         checkVec_checkResult_lo_hi_hi_hi_7 = {checkVec_checkResultVec_15_0_1, checkVec_checkResultVec_14_0_1};
  wire [15:0]        checkVec_checkResult_lo_hi_hi_7 = {checkVec_checkResult_lo_hi_hi_hi_7, checkVec_checkResult_lo_hi_hi_lo_7};
  wire [31:0]        checkVec_checkResult_lo_hi_7 = {checkVec_checkResult_lo_hi_hi_7, checkVec_checkResult_lo_hi_lo_7};
  wire [63:0]        checkVec_checkResult_lo_7 = {checkVec_checkResult_lo_hi_7, checkVec_checkResult_lo_lo_7};
  wire [7:0]         checkVec_checkResult_hi_lo_lo_lo_7 = {checkVec_checkResultVec_17_0_1, checkVec_checkResultVec_16_0_1};
  wire [7:0]         checkVec_checkResult_hi_lo_lo_hi_7 = {checkVec_checkResultVec_19_0_1, checkVec_checkResultVec_18_0_1};
  wire [15:0]        checkVec_checkResult_hi_lo_lo_7 = {checkVec_checkResult_hi_lo_lo_hi_7, checkVec_checkResult_hi_lo_lo_lo_7};
  wire [7:0]         checkVec_checkResult_hi_lo_hi_lo_7 = {checkVec_checkResultVec_21_0_1, checkVec_checkResultVec_20_0_1};
  wire [7:0]         checkVec_checkResult_hi_lo_hi_hi_7 = {checkVec_checkResultVec_23_0_1, checkVec_checkResultVec_22_0_1};
  wire [15:0]        checkVec_checkResult_hi_lo_hi_7 = {checkVec_checkResult_hi_lo_hi_hi_7, checkVec_checkResult_hi_lo_hi_lo_7};
  wire [31:0]        checkVec_checkResult_hi_lo_7 = {checkVec_checkResult_hi_lo_hi_7, checkVec_checkResult_hi_lo_lo_7};
  wire [7:0]         checkVec_checkResult_hi_hi_lo_lo_7 = {checkVec_checkResultVec_25_0_1, checkVec_checkResultVec_24_0_1};
  wire [7:0]         checkVec_checkResult_hi_hi_lo_hi_7 = {checkVec_checkResultVec_27_0_1, checkVec_checkResultVec_26_0_1};
  wire [15:0]        checkVec_checkResult_hi_hi_lo_7 = {checkVec_checkResult_hi_hi_lo_hi_7, checkVec_checkResult_hi_hi_lo_lo_7};
  wire [7:0]         checkVec_checkResult_hi_hi_hi_lo_7 = {checkVec_checkResultVec_29_0_1, checkVec_checkResultVec_28_0_1};
  wire [7:0]         checkVec_checkResult_hi_hi_hi_hi_7 = {checkVec_checkResultVec_31_0_1, checkVec_checkResultVec_30_0_1};
  wire [15:0]        checkVec_checkResult_hi_hi_hi_7 = {checkVec_checkResult_hi_hi_hi_hi_7, checkVec_checkResult_hi_hi_hi_lo_7};
  wire [31:0]        checkVec_checkResult_hi_hi_7 = {checkVec_checkResult_hi_hi_hi_7, checkVec_checkResult_hi_hi_lo_7};
  wire [63:0]        checkVec_checkResult_hi_7 = {checkVec_checkResult_hi_hi_7, checkVec_checkResult_hi_lo_7};
  wire [127:0]       checkVec_1_0 = {checkVec_checkResult_hi_7, checkVec_checkResult_lo_7};
  wire [3:0]         checkVec_checkResult_lo_lo_lo_lo_8 = {checkVec_checkResultVec_1_1_1, checkVec_checkResultVec_0_1_1};
  wire [3:0]         checkVec_checkResult_lo_lo_lo_hi_8 = {checkVec_checkResultVec_3_1_1, checkVec_checkResultVec_2_1_1};
  wire [7:0]         checkVec_checkResult_lo_lo_lo_8 = {checkVec_checkResult_lo_lo_lo_hi_8, checkVec_checkResult_lo_lo_lo_lo_8};
  wire [3:0]         checkVec_checkResult_lo_lo_hi_lo_8 = {checkVec_checkResultVec_5_1_1, checkVec_checkResultVec_4_1_1};
  wire [3:0]         checkVec_checkResult_lo_lo_hi_hi_8 = {checkVec_checkResultVec_7_1_1, checkVec_checkResultVec_6_1_1};
  wire [7:0]         checkVec_checkResult_lo_lo_hi_8 = {checkVec_checkResult_lo_lo_hi_hi_8, checkVec_checkResult_lo_lo_hi_lo_8};
  wire [15:0]        checkVec_checkResult_lo_lo_8 = {checkVec_checkResult_lo_lo_hi_8, checkVec_checkResult_lo_lo_lo_8};
  wire [3:0]         checkVec_checkResult_lo_hi_lo_lo_8 = {checkVec_checkResultVec_9_1_1, checkVec_checkResultVec_8_1_1};
  wire [3:0]         checkVec_checkResult_lo_hi_lo_hi_8 = {checkVec_checkResultVec_11_1_1, checkVec_checkResultVec_10_1_1};
  wire [7:0]         checkVec_checkResult_lo_hi_lo_8 = {checkVec_checkResult_lo_hi_lo_hi_8, checkVec_checkResult_lo_hi_lo_lo_8};
  wire [3:0]         checkVec_checkResult_lo_hi_hi_lo_8 = {checkVec_checkResultVec_13_1_1, checkVec_checkResultVec_12_1_1};
  wire [3:0]         checkVec_checkResult_lo_hi_hi_hi_8 = {checkVec_checkResultVec_15_1_1, checkVec_checkResultVec_14_1_1};
  wire [7:0]         checkVec_checkResult_lo_hi_hi_8 = {checkVec_checkResult_lo_hi_hi_hi_8, checkVec_checkResult_lo_hi_hi_lo_8};
  wire [15:0]        checkVec_checkResult_lo_hi_8 = {checkVec_checkResult_lo_hi_hi_8, checkVec_checkResult_lo_hi_lo_8};
  wire [31:0]        checkVec_checkResult_lo_8 = {checkVec_checkResult_lo_hi_8, checkVec_checkResult_lo_lo_8};
  wire [3:0]         checkVec_checkResult_hi_lo_lo_lo_8 = {checkVec_checkResultVec_17_1_1, checkVec_checkResultVec_16_1_1};
  wire [3:0]         checkVec_checkResult_hi_lo_lo_hi_8 = {checkVec_checkResultVec_19_1_1, checkVec_checkResultVec_18_1_1};
  wire [7:0]         checkVec_checkResult_hi_lo_lo_8 = {checkVec_checkResult_hi_lo_lo_hi_8, checkVec_checkResult_hi_lo_lo_lo_8};
  wire [3:0]         checkVec_checkResult_hi_lo_hi_lo_8 = {checkVec_checkResultVec_21_1_1, checkVec_checkResultVec_20_1_1};
  wire [3:0]         checkVec_checkResult_hi_lo_hi_hi_8 = {checkVec_checkResultVec_23_1_1, checkVec_checkResultVec_22_1_1};
  wire [7:0]         checkVec_checkResult_hi_lo_hi_8 = {checkVec_checkResult_hi_lo_hi_hi_8, checkVec_checkResult_hi_lo_hi_lo_8};
  wire [15:0]        checkVec_checkResult_hi_lo_8 = {checkVec_checkResult_hi_lo_hi_8, checkVec_checkResult_hi_lo_lo_8};
  wire [3:0]         checkVec_checkResult_hi_hi_lo_lo_8 = {checkVec_checkResultVec_25_1_1, checkVec_checkResultVec_24_1_1};
  wire [3:0]         checkVec_checkResult_hi_hi_lo_hi_8 = {checkVec_checkResultVec_27_1_1, checkVec_checkResultVec_26_1_1};
  wire [7:0]         checkVec_checkResult_hi_hi_lo_8 = {checkVec_checkResult_hi_hi_lo_hi_8, checkVec_checkResult_hi_hi_lo_lo_8};
  wire [3:0]         checkVec_checkResult_hi_hi_hi_lo_8 = {checkVec_checkResultVec_29_1_1, checkVec_checkResultVec_28_1_1};
  wire [3:0]         checkVec_checkResult_hi_hi_hi_hi_8 = {checkVec_checkResultVec_31_1_1, checkVec_checkResultVec_30_1_1};
  wire [7:0]         checkVec_checkResult_hi_hi_hi_8 = {checkVec_checkResult_hi_hi_hi_hi_8, checkVec_checkResult_hi_hi_hi_lo_8};
  wire [15:0]        checkVec_checkResult_hi_hi_8 = {checkVec_checkResult_hi_hi_hi_8, checkVec_checkResult_hi_hi_lo_8};
  wire [31:0]        checkVec_checkResult_hi_8 = {checkVec_checkResult_hi_hi_8, checkVec_checkResult_hi_lo_8};
  wire [63:0]        checkVec_1_1 = {checkVec_checkResult_hi_8, checkVec_checkResult_lo_8};
  wire [9:0]         checkVec_checkResult_lo_lo_lo_lo_9 = {checkVec_checkResultVec_1_2_1, checkVec_checkResultVec_0_2_1};
  wire [9:0]         checkVec_checkResult_lo_lo_lo_hi_9 = {checkVec_checkResultVec_3_2_1, checkVec_checkResultVec_2_2_1};
  wire [19:0]        checkVec_checkResult_lo_lo_lo_9 = {checkVec_checkResult_lo_lo_lo_hi_9, checkVec_checkResult_lo_lo_lo_lo_9};
  wire [9:0]         checkVec_checkResult_lo_lo_hi_lo_9 = {checkVec_checkResultVec_5_2_1, checkVec_checkResultVec_4_2_1};
  wire [9:0]         checkVec_checkResult_lo_lo_hi_hi_9 = {checkVec_checkResultVec_7_2_1, checkVec_checkResultVec_6_2_1};
  wire [19:0]        checkVec_checkResult_lo_lo_hi_9 = {checkVec_checkResult_lo_lo_hi_hi_9, checkVec_checkResult_lo_lo_hi_lo_9};
  wire [39:0]        checkVec_checkResult_lo_lo_9 = {checkVec_checkResult_lo_lo_hi_9, checkVec_checkResult_lo_lo_lo_9};
  wire [9:0]         checkVec_checkResult_lo_hi_lo_lo_9 = {checkVec_checkResultVec_9_2_1, checkVec_checkResultVec_8_2_1};
  wire [9:0]         checkVec_checkResult_lo_hi_lo_hi_9 = {checkVec_checkResultVec_11_2_1, checkVec_checkResultVec_10_2_1};
  wire [19:0]        checkVec_checkResult_lo_hi_lo_9 = {checkVec_checkResult_lo_hi_lo_hi_9, checkVec_checkResult_lo_hi_lo_lo_9};
  wire [9:0]         checkVec_checkResult_lo_hi_hi_lo_9 = {checkVec_checkResultVec_13_2_1, checkVec_checkResultVec_12_2_1};
  wire [9:0]         checkVec_checkResult_lo_hi_hi_hi_9 = {checkVec_checkResultVec_15_2_1, checkVec_checkResultVec_14_2_1};
  wire [19:0]        checkVec_checkResult_lo_hi_hi_9 = {checkVec_checkResult_lo_hi_hi_hi_9, checkVec_checkResult_lo_hi_hi_lo_9};
  wire [39:0]        checkVec_checkResult_lo_hi_9 = {checkVec_checkResult_lo_hi_hi_9, checkVec_checkResult_lo_hi_lo_9};
  wire [79:0]        checkVec_checkResult_lo_9 = {checkVec_checkResult_lo_hi_9, checkVec_checkResult_lo_lo_9};
  wire [9:0]         checkVec_checkResult_hi_lo_lo_lo_9 = {checkVec_checkResultVec_17_2_1, checkVec_checkResultVec_16_2_1};
  wire [9:0]         checkVec_checkResult_hi_lo_lo_hi_9 = {checkVec_checkResultVec_19_2_1, checkVec_checkResultVec_18_2_1};
  wire [19:0]        checkVec_checkResult_hi_lo_lo_9 = {checkVec_checkResult_hi_lo_lo_hi_9, checkVec_checkResult_hi_lo_lo_lo_9};
  wire [9:0]         checkVec_checkResult_hi_lo_hi_lo_9 = {checkVec_checkResultVec_21_2_1, checkVec_checkResultVec_20_2_1};
  wire [9:0]         checkVec_checkResult_hi_lo_hi_hi_9 = {checkVec_checkResultVec_23_2_1, checkVec_checkResultVec_22_2_1};
  wire [19:0]        checkVec_checkResult_hi_lo_hi_9 = {checkVec_checkResult_hi_lo_hi_hi_9, checkVec_checkResult_hi_lo_hi_lo_9};
  wire [39:0]        checkVec_checkResult_hi_lo_9 = {checkVec_checkResult_hi_lo_hi_9, checkVec_checkResult_hi_lo_lo_9};
  wire [9:0]         checkVec_checkResult_hi_hi_lo_lo_9 = {checkVec_checkResultVec_25_2_1, checkVec_checkResultVec_24_2_1};
  wire [9:0]         checkVec_checkResult_hi_hi_lo_hi_9 = {checkVec_checkResultVec_27_2_1, checkVec_checkResultVec_26_2_1};
  wire [19:0]        checkVec_checkResult_hi_hi_lo_9 = {checkVec_checkResult_hi_hi_lo_hi_9, checkVec_checkResult_hi_hi_lo_lo_9};
  wire [9:0]         checkVec_checkResult_hi_hi_hi_lo_9 = {checkVec_checkResultVec_29_2_1, checkVec_checkResultVec_28_2_1};
  wire [9:0]         checkVec_checkResult_hi_hi_hi_hi_9 = {checkVec_checkResultVec_31_2_1, checkVec_checkResultVec_30_2_1};
  wire [19:0]        checkVec_checkResult_hi_hi_hi_9 = {checkVec_checkResult_hi_hi_hi_hi_9, checkVec_checkResult_hi_hi_hi_lo_9};
  wire [39:0]        checkVec_checkResult_hi_hi_9 = {checkVec_checkResult_hi_hi_hi_9, checkVec_checkResult_hi_hi_lo_9};
  wire [79:0]        checkVec_checkResult_hi_9 = {checkVec_checkResult_hi_hi_9, checkVec_checkResult_hi_lo_9};
  wire [159:0]       checkVec_1_2 = {checkVec_checkResult_hi_9, checkVec_checkResult_lo_9};
  wire [1:0]         checkVec_checkResult_lo_lo_lo_lo_10 = {checkVec_checkResultVec_1_3_1, checkVec_checkResultVec_0_3_1};
  wire [1:0]         checkVec_checkResult_lo_lo_lo_hi_10 = {checkVec_checkResultVec_3_3_1, checkVec_checkResultVec_2_3_1};
  wire [3:0]         checkVec_checkResult_lo_lo_lo_10 = {checkVec_checkResult_lo_lo_lo_hi_10, checkVec_checkResult_lo_lo_lo_lo_10};
  wire [1:0]         checkVec_checkResult_lo_lo_hi_lo_10 = {checkVec_checkResultVec_5_3_1, checkVec_checkResultVec_4_3_1};
  wire [1:0]         checkVec_checkResult_lo_lo_hi_hi_10 = {checkVec_checkResultVec_7_3_1, checkVec_checkResultVec_6_3_1};
  wire [3:0]         checkVec_checkResult_lo_lo_hi_10 = {checkVec_checkResult_lo_lo_hi_hi_10, checkVec_checkResult_lo_lo_hi_lo_10};
  wire [7:0]         checkVec_checkResult_lo_lo_10 = {checkVec_checkResult_lo_lo_hi_10, checkVec_checkResult_lo_lo_lo_10};
  wire [1:0]         checkVec_checkResult_lo_hi_lo_lo_10 = {checkVec_checkResultVec_9_3_1, checkVec_checkResultVec_8_3_1};
  wire [1:0]         checkVec_checkResult_lo_hi_lo_hi_10 = {checkVec_checkResultVec_11_3_1, checkVec_checkResultVec_10_3_1};
  wire [3:0]         checkVec_checkResult_lo_hi_lo_10 = {checkVec_checkResult_lo_hi_lo_hi_10, checkVec_checkResult_lo_hi_lo_lo_10};
  wire [1:0]         checkVec_checkResult_lo_hi_hi_lo_10 = {checkVec_checkResultVec_13_3_1, checkVec_checkResultVec_12_3_1};
  wire [1:0]         checkVec_checkResult_lo_hi_hi_hi_10 = {checkVec_checkResultVec_15_3_1, checkVec_checkResultVec_14_3_1};
  wire [3:0]         checkVec_checkResult_lo_hi_hi_10 = {checkVec_checkResult_lo_hi_hi_hi_10, checkVec_checkResult_lo_hi_hi_lo_10};
  wire [7:0]         checkVec_checkResult_lo_hi_10 = {checkVec_checkResult_lo_hi_hi_10, checkVec_checkResult_lo_hi_lo_10};
  wire [15:0]        checkVec_checkResult_lo_10 = {checkVec_checkResult_lo_hi_10, checkVec_checkResult_lo_lo_10};
  wire [1:0]         checkVec_checkResult_hi_lo_lo_lo_10 = {checkVec_checkResultVec_17_3_1, checkVec_checkResultVec_16_3_1};
  wire [1:0]         checkVec_checkResult_hi_lo_lo_hi_10 = {checkVec_checkResultVec_19_3_1, checkVec_checkResultVec_18_3_1};
  wire [3:0]         checkVec_checkResult_hi_lo_lo_10 = {checkVec_checkResult_hi_lo_lo_hi_10, checkVec_checkResult_hi_lo_lo_lo_10};
  wire [1:0]         checkVec_checkResult_hi_lo_hi_lo_10 = {checkVec_checkResultVec_21_3_1, checkVec_checkResultVec_20_3_1};
  wire [1:0]         checkVec_checkResult_hi_lo_hi_hi_10 = {checkVec_checkResultVec_23_3_1, checkVec_checkResultVec_22_3_1};
  wire [3:0]         checkVec_checkResult_hi_lo_hi_10 = {checkVec_checkResult_hi_lo_hi_hi_10, checkVec_checkResult_hi_lo_hi_lo_10};
  wire [7:0]         checkVec_checkResult_hi_lo_10 = {checkVec_checkResult_hi_lo_hi_10, checkVec_checkResult_hi_lo_lo_10};
  wire [1:0]         checkVec_checkResult_hi_hi_lo_lo_10 = {checkVec_checkResultVec_25_3_1, checkVec_checkResultVec_24_3_1};
  wire [1:0]         checkVec_checkResult_hi_hi_lo_hi_10 = {checkVec_checkResultVec_27_3_1, checkVec_checkResultVec_26_3_1};
  wire [3:0]         checkVec_checkResult_hi_hi_lo_10 = {checkVec_checkResult_hi_hi_lo_hi_10, checkVec_checkResult_hi_hi_lo_lo_10};
  wire [1:0]         checkVec_checkResult_hi_hi_hi_lo_10 = {checkVec_checkResultVec_29_3_1, checkVec_checkResultVec_28_3_1};
  wire [1:0]         checkVec_checkResult_hi_hi_hi_hi_10 = {checkVec_checkResultVec_31_3_1, checkVec_checkResultVec_30_3_1};
  wire [3:0]         checkVec_checkResult_hi_hi_hi_10 = {checkVec_checkResult_hi_hi_hi_hi_10, checkVec_checkResult_hi_hi_hi_lo_10};
  wire [7:0]         checkVec_checkResult_hi_hi_10 = {checkVec_checkResult_hi_hi_hi_10, checkVec_checkResult_hi_hi_lo_10};
  wire [15:0]        checkVec_checkResult_hi_10 = {checkVec_checkResult_hi_hi_10, checkVec_checkResult_hi_lo_10};
  wire [31:0]        checkVec_1_3 = {checkVec_checkResult_hi_10, checkVec_checkResult_lo_10};
  wire [5:0]         checkVec_checkResult_lo_lo_lo_lo_11 = {checkVec_checkResultVec_1_4_1, checkVec_checkResultVec_0_4_1};
  wire [5:0]         checkVec_checkResult_lo_lo_lo_hi_11 = {checkVec_checkResultVec_3_4_1, checkVec_checkResultVec_2_4_1};
  wire [11:0]        checkVec_checkResult_lo_lo_lo_11 = {checkVec_checkResult_lo_lo_lo_hi_11, checkVec_checkResult_lo_lo_lo_lo_11};
  wire [5:0]         checkVec_checkResult_lo_lo_hi_lo_11 = {checkVec_checkResultVec_5_4_1, checkVec_checkResultVec_4_4_1};
  wire [5:0]         checkVec_checkResult_lo_lo_hi_hi_11 = {checkVec_checkResultVec_7_4_1, checkVec_checkResultVec_6_4_1};
  wire [11:0]        checkVec_checkResult_lo_lo_hi_11 = {checkVec_checkResult_lo_lo_hi_hi_11, checkVec_checkResult_lo_lo_hi_lo_11};
  wire [23:0]        checkVec_checkResult_lo_lo_11 = {checkVec_checkResult_lo_lo_hi_11, checkVec_checkResult_lo_lo_lo_11};
  wire [5:0]         checkVec_checkResult_lo_hi_lo_lo_11 = {checkVec_checkResultVec_9_4_1, checkVec_checkResultVec_8_4_1};
  wire [5:0]         checkVec_checkResult_lo_hi_lo_hi_11 = {checkVec_checkResultVec_11_4_1, checkVec_checkResultVec_10_4_1};
  wire [11:0]        checkVec_checkResult_lo_hi_lo_11 = {checkVec_checkResult_lo_hi_lo_hi_11, checkVec_checkResult_lo_hi_lo_lo_11};
  wire [5:0]         checkVec_checkResult_lo_hi_hi_lo_11 = {checkVec_checkResultVec_13_4_1, checkVec_checkResultVec_12_4_1};
  wire [5:0]         checkVec_checkResult_lo_hi_hi_hi_11 = {checkVec_checkResultVec_15_4_1, checkVec_checkResultVec_14_4_1};
  wire [11:0]        checkVec_checkResult_lo_hi_hi_11 = {checkVec_checkResult_lo_hi_hi_hi_11, checkVec_checkResult_lo_hi_hi_lo_11};
  wire [23:0]        checkVec_checkResult_lo_hi_11 = {checkVec_checkResult_lo_hi_hi_11, checkVec_checkResult_lo_hi_lo_11};
  wire [47:0]        checkVec_checkResult_lo_11 = {checkVec_checkResult_lo_hi_11, checkVec_checkResult_lo_lo_11};
  wire [5:0]         checkVec_checkResult_hi_lo_lo_lo_11 = {checkVec_checkResultVec_17_4_1, checkVec_checkResultVec_16_4_1};
  wire [5:0]         checkVec_checkResult_hi_lo_lo_hi_11 = {checkVec_checkResultVec_19_4_1, checkVec_checkResultVec_18_4_1};
  wire [11:0]        checkVec_checkResult_hi_lo_lo_11 = {checkVec_checkResult_hi_lo_lo_hi_11, checkVec_checkResult_hi_lo_lo_lo_11};
  wire [5:0]         checkVec_checkResult_hi_lo_hi_lo_11 = {checkVec_checkResultVec_21_4_1, checkVec_checkResultVec_20_4_1};
  wire [5:0]         checkVec_checkResult_hi_lo_hi_hi_11 = {checkVec_checkResultVec_23_4_1, checkVec_checkResultVec_22_4_1};
  wire [11:0]        checkVec_checkResult_hi_lo_hi_11 = {checkVec_checkResult_hi_lo_hi_hi_11, checkVec_checkResult_hi_lo_hi_lo_11};
  wire [23:0]        checkVec_checkResult_hi_lo_11 = {checkVec_checkResult_hi_lo_hi_11, checkVec_checkResult_hi_lo_lo_11};
  wire [5:0]         checkVec_checkResult_hi_hi_lo_lo_11 = {checkVec_checkResultVec_25_4_1, checkVec_checkResultVec_24_4_1};
  wire [5:0]         checkVec_checkResult_hi_hi_lo_hi_11 = {checkVec_checkResultVec_27_4_1, checkVec_checkResultVec_26_4_1};
  wire [11:0]        checkVec_checkResult_hi_hi_lo_11 = {checkVec_checkResult_hi_hi_lo_hi_11, checkVec_checkResult_hi_hi_lo_lo_11};
  wire [5:0]         checkVec_checkResult_hi_hi_hi_lo_11 = {checkVec_checkResultVec_29_4_1, checkVec_checkResultVec_28_4_1};
  wire [5:0]         checkVec_checkResult_hi_hi_hi_hi_11 = {checkVec_checkResultVec_31_4_1, checkVec_checkResultVec_30_4_1};
  wire [11:0]        checkVec_checkResult_hi_hi_hi_11 = {checkVec_checkResult_hi_hi_hi_hi_11, checkVec_checkResult_hi_hi_hi_lo_11};
  wire [23:0]        checkVec_checkResult_hi_hi_11 = {checkVec_checkResult_hi_hi_hi_11, checkVec_checkResult_hi_hi_lo_11};
  wire [47:0]        checkVec_checkResult_hi_11 = {checkVec_checkResult_hi_hi_11, checkVec_checkResult_hi_lo_11};
  wire [95:0]        checkVec_1_4 = {checkVec_checkResult_hi_11, checkVec_checkResult_lo_11};
  wire [1:0]         checkVec_checkResult_lo_lo_lo_lo_12 = {checkVec_checkResultVec_1_5_1, checkVec_checkResultVec_0_5_1};
  wire [1:0]         checkVec_checkResult_lo_lo_lo_hi_12 = {checkVec_checkResultVec_3_5_1, checkVec_checkResultVec_2_5_1};
  wire [3:0]         checkVec_checkResult_lo_lo_lo_12 = {checkVec_checkResult_lo_lo_lo_hi_12, checkVec_checkResult_lo_lo_lo_lo_12};
  wire [1:0]         checkVec_checkResult_lo_lo_hi_lo_12 = {checkVec_checkResultVec_5_5_1, checkVec_checkResultVec_4_5_1};
  wire [1:0]         checkVec_checkResult_lo_lo_hi_hi_12 = {checkVec_checkResultVec_7_5_1, checkVec_checkResultVec_6_5_1};
  wire [3:0]         checkVec_checkResult_lo_lo_hi_12 = {checkVec_checkResult_lo_lo_hi_hi_12, checkVec_checkResult_lo_lo_hi_lo_12};
  wire [7:0]         checkVec_checkResult_lo_lo_12 = {checkVec_checkResult_lo_lo_hi_12, checkVec_checkResult_lo_lo_lo_12};
  wire [1:0]         checkVec_checkResult_lo_hi_lo_lo_12 = {checkVec_checkResultVec_9_5_1, checkVec_checkResultVec_8_5_1};
  wire [1:0]         checkVec_checkResult_lo_hi_lo_hi_12 = {checkVec_checkResultVec_11_5_1, checkVec_checkResultVec_10_5_1};
  wire [3:0]         checkVec_checkResult_lo_hi_lo_12 = {checkVec_checkResult_lo_hi_lo_hi_12, checkVec_checkResult_lo_hi_lo_lo_12};
  wire [1:0]         checkVec_checkResult_lo_hi_hi_lo_12 = {checkVec_checkResultVec_13_5_1, checkVec_checkResultVec_12_5_1};
  wire [1:0]         checkVec_checkResult_lo_hi_hi_hi_12 = {checkVec_checkResultVec_15_5_1, checkVec_checkResultVec_14_5_1};
  wire [3:0]         checkVec_checkResult_lo_hi_hi_12 = {checkVec_checkResult_lo_hi_hi_hi_12, checkVec_checkResult_lo_hi_hi_lo_12};
  wire [7:0]         checkVec_checkResult_lo_hi_12 = {checkVec_checkResult_lo_hi_hi_12, checkVec_checkResult_lo_hi_lo_12};
  wire [15:0]        checkVec_checkResult_lo_12 = {checkVec_checkResult_lo_hi_12, checkVec_checkResult_lo_lo_12};
  wire [1:0]         checkVec_checkResult_hi_lo_lo_lo_12 = {checkVec_checkResultVec_17_5_1, checkVec_checkResultVec_16_5_1};
  wire [1:0]         checkVec_checkResult_hi_lo_lo_hi_12 = {checkVec_checkResultVec_19_5_1, checkVec_checkResultVec_18_5_1};
  wire [3:0]         checkVec_checkResult_hi_lo_lo_12 = {checkVec_checkResult_hi_lo_lo_hi_12, checkVec_checkResult_hi_lo_lo_lo_12};
  wire [1:0]         checkVec_checkResult_hi_lo_hi_lo_12 = {checkVec_checkResultVec_21_5_1, checkVec_checkResultVec_20_5_1};
  wire [1:0]         checkVec_checkResult_hi_lo_hi_hi_12 = {checkVec_checkResultVec_23_5_1, checkVec_checkResultVec_22_5_1};
  wire [3:0]         checkVec_checkResult_hi_lo_hi_12 = {checkVec_checkResult_hi_lo_hi_hi_12, checkVec_checkResult_hi_lo_hi_lo_12};
  wire [7:0]         checkVec_checkResult_hi_lo_12 = {checkVec_checkResult_hi_lo_hi_12, checkVec_checkResult_hi_lo_lo_12};
  wire [1:0]         checkVec_checkResult_hi_hi_lo_lo_12 = {checkVec_checkResultVec_25_5_1, checkVec_checkResultVec_24_5_1};
  wire [1:0]         checkVec_checkResult_hi_hi_lo_hi_12 = {checkVec_checkResultVec_27_5_1, checkVec_checkResultVec_26_5_1};
  wire [3:0]         checkVec_checkResult_hi_hi_lo_12 = {checkVec_checkResult_hi_hi_lo_hi_12, checkVec_checkResult_hi_hi_lo_lo_12};
  wire [1:0]         checkVec_checkResult_hi_hi_hi_lo_12 = {checkVec_checkResultVec_29_5_1, checkVec_checkResultVec_28_5_1};
  wire [1:0]         checkVec_checkResult_hi_hi_hi_hi_12 = {checkVec_checkResultVec_31_5_1, checkVec_checkResultVec_30_5_1};
  wire [3:0]         checkVec_checkResult_hi_hi_hi_12 = {checkVec_checkResult_hi_hi_hi_hi_12, checkVec_checkResult_hi_hi_hi_lo_12};
  wire [7:0]         checkVec_checkResult_hi_hi_12 = {checkVec_checkResult_hi_hi_hi_12, checkVec_checkResult_hi_hi_lo_12};
  wire [15:0]        checkVec_checkResult_hi_12 = {checkVec_checkResult_hi_hi_12, checkVec_checkResult_hi_lo_12};
  wire [31:0]        checkVec_1_5 = {checkVec_checkResult_hi_12, checkVec_checkResult_lo_12};
  wire [1:0]         checkVec_checkResult_lo_lo_lo_lo_13 = {checkVec_checkResultVec_1_6_1, checkVec_checkResultVec_0_6_1};
  wire [1:0]         checkVec_checkResult_lo_lo_lo_hi_13 = {checkVec_checkResultVec_3_6_1, checkVec_checkResultVec_2_6_1};
  wire [3:0]         checkVec_checkResult_lo_lo_lo_13 = {checkVec_checkResult_lo_lo_lo_hi_13, checkVec_checkResult_lo_lo_lo_lo_13};
  wire [1:0]         checkVec_checkResult_lo_lo_hi_lo_13 = {checkVec_checkResultVec_5_6_1, checkVec_checkResultVec_4_6_1};
  wire [1:0]         checkVec_checkResult_lo_lo_hi_hi_13 = {checkVec_checkResultVec_7_6_1, checkVec_checkResultVec_6_6_1};
  wire [3:0]         checkVec_checkResult_lo_lo_hi_13 = {checkVec_checkResult_lo_lo_hi_hi_13, checkVec_checkResult_lo_lo_hi_lo_13};
  wire [7:0]         checkVec_checkResult_lo_lo_13 = {checkVec_checkResult_lo_lo_hi_13, checkVec_checkResult_lo_lo_lo_13};
  wire [1:0]         checkVec_checkResult_lo_hi_lo_lo_13 = {checkVec_checkResultVec_9_6_1, checkVec_checkResultVec_8_6_1};
  wire [1:0]         checkVec_checkResult_lo_hi_lo_hi_13 = {checkVec_checkResultVec_11_6_1, checkVec_checkResultVec_10_6_1};
  wire [3:0]         checkVec_checkResult_lo_hi_lo_13 = {checkVec_checkResult_lo_hi_lo_hi_13, checkVec_checkResult_lo_hi_lo_lo_13};
  wire [1:0]         checkVec_checkResult_lo_hi_hi_lo_13 = {checkVec_checkResultVec_13_6_1, checkVec_checkResultVec_12_6_1};
  wire [1:0]         checkVec_checkResult_lo_hi_hi_hi_13 = {checkVec_checkResultVec_15_6_1, checkVec_checkResultVec_14_6_1};
  wire [3:0]         checkVec_checkResult_lo_hi_hi_13 = {checkVec_checkResult_lo_hi_hi_hi_13, checkVec_checkResult_lo_hi_hi_lo_13};
  wire [7:0]         checkVec_checkResult_lo_hi_13 = {checkVec_checkResult_lo_hi_hi_13, checkVec_checkResult_lo_hi_lo_13};
  wire [15:0]        checkVec_checkResult_lo_13 = {checkVec_checkResult_lo_hi_13, checkVec_checkResult_lo_lo_13};
  wire [1:0]         checkVec_checkResult_hi_lo_lo_lo_13 = {checkVec_checkResultVec_17_6_1, checkVec_checkResultVec_16_6_1};
  wire [1:0]         checkVec_checkResult_hi_lo_lo_hi_13 = {checkVec_checkResultVec_19_6_1, checkVec_checkResultVec_18_6_1};
  wire [3:0]         checkVec_checkResult_hi_lo_lo_13 = {checkVec_checkResult_hi_lo_lo_hi_13, checkVec_checkResult_hi_lo_lo_lo_13};
  wire [1:0]         checkVec_checkResult_hi_lo_hi_lo_13 = {checkVec_checkResultVec_21_6_1, checkVec_checkResultVec_20_6_1};
  wire [1:0]         checkVec_checkResult_hi_lo_hi_hi_13 = {checkVec_checkResultVec_23_6_1, checkVec_checkResultVec_22_6_1};
  wire [3:0]         checkVec_checkResult_hi_lo_hi_13 = {checkVec_checkResult_hi_lo_hi_hi_13, checkVec_checkResult_hi_lo_hi_lo_13};
  wire [7:0]         checkVec_checkResult_hi_lo_13 = {checkVec_checkResult_hi_lo_hi_13, checkVec_checkResult_hi_lo_lo_13};
  wire [1:0]         checkVec_checkResult_hi_hi_lo_lo_13 = {checkVec_checkResultVec_25_6_1, checkVec_checkResultVec_24_6_1};
  wire [1:0]         checkVec_checkResult_hi_hi_lo_hi_13 = {checkVec_checkResultVec_27_6_1, checkVec_checkResultVec_26_6_1};
  wire [3:0]         checkVec_checkResult_hi_hi_lo_13 = {checkVec_checkResult_hi_hi_lo_hi_13, checkVec_checkResult_hi_hi_lo_lo_13};
  wire [1:0]         checkVec_checkResult_hi_hi_hi_lo_13 = {checkVec_checkResultVec_29_6_1, checkVec_checkResultVec_28_6_1};
  wire [1:0]         checkVec_checkResult_hi_hi_hi_hi_13 = {checkVec_checkResultVec_31_6_1, checkVec_checkResultVec_30_6_1};
  wire [3:0]         checkVec_checkResult_hi_hi_hi_13 = {checkVec_checkResult_hi_hi_hi_hi_13, checkVec_checkResult_hi_hi_hi_lo_13};
  wire [7:0]         checkVec_checkResult_hi_hi_13 = {checkVec_checkResult_hi_hi_hi_13, checkVec_checkResult_hi_hi_lo_13};
  wire [15:0]        checkVec_checkResult_hi_13 = {checkVec_checkResult_hi_hi_13, checkVec_checkResult_hi_lo_13};
  wire [31:0]        checkVec_1_6 = {checkVec_checkResult_hi_13, checkVec_checkResult_lo_13};
  wire               checkVec_checkResultVec_0_6_2 = checkVec_validVec_2[0];
  wire [10:0]        checkVec_checkResultVec_dataPosition_64 = {source_0[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_0_2_2 = checkVec_checkResultVec_dataPosition_64[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_64 = checkVec_checkResultVec_dataPosition_64[10:7];
  wire               checkVec_checkResultVec_0_3_2 = checkVec_checkResultVec_dataGroup_64[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_64 = checkVec_checkResultVec_dataGroup_64[3:1];
  wire [2:0]         checkVec_checkResultVec_0_4_2 = checkVec_checkResultVec_accessRegGrowth_64;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_64 = {checkVec_checkResultVec_0_3_2, checkVec_checkResultVec_0_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_64 = checkVec_checkResultVec_decimalProportion_64[5:3];
  wire               checkVec_checkResultVec_overlap_64 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_64 >= checkVec_checkResultVec_intLMULInput_64[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_64} >= checkVec_checkResultVec_intLMULInput_64,
      source_0[31:11]};
  wire               checkVec_checkResultVec_0_5_2 = checkVec_checkResultVec_overlap_64 | ~checkVec_checkResultVec_0_6_2;
  wire               checkVec_checkResultVec_1_6_2 = checkVec_validVec_2[1];
  wire [10:0]        checkVec_checkResultVec_dataPosition_65 = {source_1[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_1_2_2 = checkVec_checkResultVec_dataPosition_65[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_65 = checkVec_checkResultVec_dataPosition_65[10:7];
  wire               checkVec_checkResultVec_1_3_2 = checkVec_checkResultVec_dataGroup_65[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_65 = checkVec_checkResultVec_dataGroup_65[3:1];
  wire [2:0]         checkVec_checkResultVec_1_4_2 = checkVec_checkResultVec_accessRegGrowth_65;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_65 = {checkVec_checkResultVec_1_3_2, checkVec_checkResultVec_1_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_65 = checkVec_checkResultVec_decimalProportion_65[5:3];
  wire               checkVec_checkResultVec_overlap_65 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_65 >= checkVec_checkResultVec_intLMULInput_65[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_65} >= checkVec_checkResultVec_intLMULInput_65,
      source_1[31:11]};
  wire               checkVec_checkResultVec_1_5_2 = checkVec_checkResultVec_overlap_65 | ~checkVec_checkResultVec_1_6_2;
  wire               checkVec_checkResultVec_2_6_2 = checkVec_validVec_2[2];
  wire [10:0]        checkVec_checkResultVec_dataPosition_66 = {source_2[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_2_2_2 = checkVec_checkResultVec_dataPosition_66[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_66 = checkVec_checkResultVec_dataPosition_66[10:7];
  wire               checkVec_checkResultVec_2_3_2 = checkVec_checkResultVec_dataGroup_66[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_66 = checkVec_checkResultVec_dataGroup_66[3:1];
  wire [2:0]         checkVec_checkResultVec_2_4_2 = checkVec_checkResultVec_accessRegGrowth_66;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_66 = {checkVec_checkResultVec_2_3_2, checkVec_checkResultVec_2_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_66 = checkVec_checkResultVec_decimalProportion_66[5:3];
  wire               checkVec_checkResultVec_overlap_66 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_66 >= checkVec_checkResultVec_intLMULInput_66[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_66} >= checkVec_checkResultVec_intLMULInput_66,
      source_2[31:11]};
  wire               checkVec_checkResultVec_2_5_2 = checkVec_checkResultVec_overlap_66 | ~checkVec_checkResultVec_2_6_2;
  wire               checkVec_checkResultVec_3_6_2 = checkVec_validVec_2[3];
  wire [10:0]        checkVec_checkResultVec_dataPosition_67 = {source_3[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_3_2_2 = checkVec_checkResultVec_dataPosition_67[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_67 = checkVec_checkResultVec_dataPosition_67[10:7];
  wire               checkVec_checkResultVec_3_3_2 = checkVec_checkResultVec_dataGroup_67[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_67 = checkVec_checkResultVec_dataGroup_67[3:1];
  wire [2:0]         checkVec_checkResultVec_3_4_2 = checkVec_checkResultVec_accessRegGrowth_67;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_67 = {checkVec_checkResultVec_3_3_2, checkVec_checkResultVec_3_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_67 = checkVec_checkResultVec_decimalProportion_67[5:3];
  wire               checkVec_checkResultVec_overlap_67 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_67 >= checkVec_checkResultVec_intLMULInput_67[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_67} >= checkVec_checkResultVec_intLMULInput_67,
      source_3[31:11]};
  wire               checkVec_checkResultVec_3_5_2 = checkVec_checkResultVec_overlap_67 | ~checkVec_checkResultVec_3_6_2;
  wire               checkVec_checkResultVec_4_6_2 = checkVec_validVec_2[4];
  wire [10:0]        checkVec_checkResultVec_dataPosition_68 = {source_4[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_4_2_2 = checkVec_checkResultVec_dataPosition_68[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_68 = checkVec_checkResultVec_dataPosition_68[10:7];
  wire               checkVec_checkResultVec_4_3_2 = checkVec_checkResultVec_dataGroup_68[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_68 = checkVec_checkResultVec_dataGroup_68[3:1];
  wire [2:0]         checkVec_checkResultVec_4_4_2 = checkVec_checkResultVec_accessRegGrowth_68;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_68 = {checkVec_checkResultVec_4_3_2, checkVec_checkResultVec_4_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_68 = checkVec_checkResultVec_decimalProportion_68[5:3];
  wire               checkVec_checkResultVec_overlap_68 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_68 >= checkVec_checkResultVec_intLMULInput_68[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_68} >= checkVec_checkResultVec_intLMULInput_68,
      source_4[31:11]};
  wire               checkVec_checkResultVec_4_5_2 = checkVec_checkResultVec_overlap_68 | ~checkVec_checkResultVec_4_6_2;
  wire               checkVec_checkResultVec_5_6_2 = checkVec_validVec_2[5];
  wire [10:0]        checkVec_checkResultVec_dataPosition_69 = {source_5[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_5_2_2 = checkVec_checkResultVec_dataPosition_69[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_69 = checkVec_checkResultVec_dataPosition_69[10:7];
  wire               checkVec_checkResultVec_5_3_2 = checkVec_checkResultVec_dataGroup_69[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_69 = checkVec_checkResultVec_dataGroup_69[3:1];
  wire [2:0]         checkVec_checkResultVec_5_4_2 = checkVec_checkResultVec_accessRegGrowth_69;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_69 = {checkVec_checkResultVec_5_3_2, checkVec_checkResultVec_5_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_69 = checkVec_checkResultVec_decimalProportion_69[5:3];
  wire               checkVec_checkResultVec_overlap_69 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_69 >= checkVec_checkResultVec_intLMULInput_69[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_69} >= checkVec_checkResultVec_intLMULInput_69,
      source_5[31:11]};
  wire               checkVec_checkResultVec_5_5_2 = checkVec_checkResultVec_overlap_69 | ~checkVec_checkResultVec_5_6_2;
  wire               checkVec_checkResultVec_6_6_2 = checkVec_validVec_2[6];
  wire [10:0]        checkVec_checkResultVec_dataPosition_70 = {source_6[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_6_2_2 = checkVec_checkResultVec_dataPosition_70[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_70 = checkVec_checkResultVec_dataPosition_70[10:7];
  wire               checkVec_checkResultVec_6_3_2 = checkVec_checkResultVec_dataGroup_70[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_70 = checkVec_checkResultVec_dataGroup_70[3:1];
  wire [2:0]         checkVec_checkResultVec_6_4_2 = checkVec_checkResultVec_accessRegGrowth_70;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_70 = {checkVec_checkResultVec_6_3_2, checkVec_checkResultVec_6_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_70 = checkVec_checkResultVec_decimalProportion_70[5:3];
  wire               checkVec_checkResultVec_overlap_70 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_70 >= checkVec_checkResultVec_intLMULInput_70[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_70} >= checkVec_checkResultVec_intLMULInput_70,
      source_6[31:11]};
  wire               checkVec_checkResultVec_6_5_2 = checkVec_checkResultVec_overlap_70 | ~checkVec_checkResultVec_6_6_2;
  wire               checkVec_checkResultVec_7_6_2 = checkVec_validVec_2[7];
  wire [10:0]        checkVec_checkResultVec_dataPosition_71 = {source_7[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_7_2_2 = checkVec_checkResultVec_dataPosition_71[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_71 = checkVec_checkResultVec_dataPosition_71[10:7];
  wire               checkVec_checkResultVec_7_3_2 = checkVec_checkResultVec_dataGroup_71[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_71 = checkVec_checkResultVec_dataGroup_71[3:1];
  wire [2:0]         checkVec_checkResultVec_7_4_2 = checkVec_checkResultVec_accessRegGrowth_71;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_71 = {checkVec_checkResultVec_7_3_2, checkVec_checkResultVec_7_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_71 = checkVec_checkResultVec_decimalProportion_71[5:3];
  wire               checkVec_checkResultVec_overlap_71 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_71 >= checkVec_checkResultVec_intLMULInput_71[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_71} >= checkVec_checkResultVec_intLMULInput_71,
      source_7[31:11]};
  wire               checkVec_checkResultVec_7_5_2 = checkVec_checkResultVec_overlap_71 | ~checkVec_checkResultVec_7_6_2;
  wire               checkVec_checkResultVec_8_6_2 = checkVec_validVec_2[8];
  wire [10:0]        checkVec_checkResultVec_dataPosition_72 = {source_8[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_8_2_2 = checkVec_checkResultVec_dataPosition_72[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_72 = checkVec_checkResultVec_dataPosition_72[10:7];
  wire               checkVec_checkResultVec_8_3_2 = checkVec_checkResultVec_dataGroup_72[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_72 = checkVec_checkResultVec_dataGroup_72[3:1];
  wire [2:0]         checkVec_checkResultVec_8_4_2 = checkVec_checkResultVec_accessRegGrowth_72;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_72 = {checkVec_checkResultVec_8_3_2, checkVec_checkResultVec_8_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_72 = checkVec_checkResultVec_decimalProportion_72[5:3];
  wire               checkVec_checkResultVec_overlap_72 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_72 >= checkVec_checkResultVec_intLMULInput_72[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_72} >= checkVec_checkResultVec_intLMULInput_72,
      source_8[31:11]};
  wire               checkVec_checkResultVec_8_5_2 = checkVec_checkResultVec_overlap_72 | ~checkVec_checkResultVec_8_6_2;
  wire               checkVec_checkResultVec_9_6_2 = checkVec_validVec_2[9];
  wire [10:0]        checkVec_checkResultVec_dataPosition_73 = {source_9[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_9_2_2 = checkVec_checkResultVec_dataPosition_73[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_73 = checkVec_checkResultVec_dataPosition_73[10:7];
  wire               checkVec_checkResultVec_9_3_2 = checkVec_checkResultVec_dataGroup_73[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_73 = checkVec_checkResultVec_dataGroup_73[3:1];
  wire [2:0]         checkVec_checkResultVec_9_4_2 = checkVec_checkResultVec_accessRegGrowth_73;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_73 = {checkVec_checkResultVec_9_3_2, checkVec_checkResultVec_9_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_73 = checkVec_checkResultVec_decimalProportion_73[5:3];
  wire               checkVec_checkResultVec_overlap_73 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_73 >= checkVec_checkResultVec_intLMULInput_73[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_73} >= checkVec_checkResultVec_intLMULInput_73,
      source_9[31:11]};
  wire               checkVec_checkResultVec_9_5_2 = checkVec_checkResultVec_overlap_73 | ~checkVec_checkResultVec_9_6_2;
  wire               checkVec_checkResultVec_10_6_2 = checkVec_validVec_2[10];
  wire [10:0]        checkVec_checkResultVec_dataPosition_74 = {source_10[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_10_2_2 = checkVec_checkResultVec_dataPosition_74[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_74 = checkVec_checkResultVec_dataPosition_74[10:7];
  wire               checkVec_checkResultVec_10_3_2 = checkVec_checkResultVec_dataGroup_74[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_74 = checkVec_checkResultVec_dataGroup_74[3:1];
  wire [2:0]         checkVec_checkResultVec_10_4_2 = checkVec_checkResultVec_accessRegGrowth_74;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_74 = {checkVec_checkResultVec_10_3_2, checkVec_checkResultVec_10_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_74 = checkVec_checkResultVec_decimalProportion_74[5:3];
  wire               checkVec_checkResultVec_overlap_74 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_74 >= checkVec_checkResultVec_intLMULInput_74[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_74} >= checkVec_checkResultVec_intLMULInput_74,
      source_10[31:11]};
  wire               checkVec_checkResultVec_10_5_2 = checkVec_checkResultVec_overlap_74 | ~checkVec_checkResultVec_10_6_2;
  wire               checkVec_checkResultVec_11_6_2 = checkVec_validVec_2[11];
  wire [10:0]        checkVec_checkResultVec_dataPosition_75 = {source_11[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_11_2_2 = checkVec_checkResultVec_dataPosition_75[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_75 = checkVec_checkResultVec_dataPosition_75[10:7];
  wire               checkVec_checkResultVec_11_3_2 = checkVec_checkResultVec_dataGroup_75[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_75 = checkVec_checkResultVec_dataGroup_75[3:1];
  wire [2:0]         checkVec_checkResultVec_11_4_2 = checkVec_checkResultVec_accessRegGrowth_75;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_75 = {checkVec_checkResultVec_11_3_2, checkVec_checkResultVec_11_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_75 = checkVec_checkResultVec_decimalProportion_75[5:3];
  wire               checkVec_checkResultVec_overlap_75 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_75 >= checkVec_checkResultVec_intLMULInput_75[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_75} >= checkVec_checkResultVec_intLMULInput_75,
      source_11[31:11]};
  wire               checkVec_checkResultVec_11_5_2 = checkVec_checkResultVec_overlap_75 | ~checkVec_checkResultVec_11_6_2;
  wire               checkVec_checkResultVec_12_6_2 = checkVec_validVec_2[12];
  wire [10:0]        checkVec_checkResultVec_dataPosition_76 = {source_12[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_12_2_2 = checkVec_checkResultVec_dataPosition_76[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_76 = checkVec_checkResultVec_dataPosition_76[10:7];
  wire               checkVec_checkResultVec_12_3_2 = checkVec_checkResultVec_dataGroup_76[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_76 = checkVec_checkResultVec_dataGroup_76[3:1];
  wire [2:0]         checkVec_checkResultVec_12_4_2 = checkVec_checkResultVec_accessRegGrowth_76;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_76 = {checkVec_checkResultVec_12_3_2, checkVec_checkResultVec_12_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_76 = checkVec_checkResultVec_decimalProportion_76[5:3];
  wire               checkVec_checkResultVec_overlap_76 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_76 >= checkVec_checkResultVec_intLMULInput_76[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_76} >= checkVec_checkResultVec_intLMULInput_76,
      source_12[31:11]};
  wire               checkVec_checkResultVec_12_5_2 = checkVec_checkResultVec_overlap_76 | ~checkVec_checkResultVec_12_6_2;
  wire               checkVec_checkResultVec_13_6_2 = checkVec_validVec_2[13];
  wire [10:0]        checkVec_checkResultVec_dataPosition_77 = {source_13[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_13_2_2 = checkVec_checkResultVec_dataPosition_77[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_77 = checkVec_checkResultVec_dataPosition_77[10:7];
  wire               checkVec_checkResultVec_13_3_2 = checkVec_checkResultVec_dataGroup_77[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_77 = checkVec_checkResultVec_dataGroup_77[3:1];
  wire [2:0]         checkVec_checkResultVec_13_4_2 = checkVec_checkResultVec_accessRegGrowth_77;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_77 = {checkVec_checkResultVec_13_3_2, checkVec_checkResultVec_13_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_77 = checkVec_checkResultVec_decimalProportion_77[5:3];
  wire               checkVec_checkResultVec_overlap_77 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_77 >= checkVec_checkResultVec_intLMULInput_77[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_77} >= checkVec_checkResultVec_intLMULInput_77,
      source_13[31:11]};
  wire               checkVec_checkResultVec_13_5_2 = checkVec_checkResultVec_overlap_77 | ~checkVec_checkResultVec_13_6_2;
  wire               checkVec_checkResultVec_14_6_2 = checkVec_validVec_2[14];
  wire [10:0]        checkVec_checkResultVec_dataPosition_78 = {source_14[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_14_2_2 = checkVec_checkResultVec_dataPosition_78[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_78 = checkVec_checkResultVec_dataPosition_78[10:7];
  wire               checkVec_checkResultVec_14_3_2 = checkVec_checkResultVec_dataGroup_78[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_78 = checkVec_checkResultVec_dataGroup_78[3:1];
  wire [2:0]         checkVec_checkResultVec_14_4_2 = checkVec_checkResultVec_accessRegGrowth_78;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_78 = {checkVec_checkResultVec_14_3_2, checkVec_checkResultVec_14_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_78 = checkVec_checkResultVec_decimalProportion_78[5:3];
  wire               checkVec_checkResultVec_overlap_78 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_78 >= checkVec_checkResultVec_intLMULInput_78[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_78} >= checkVec_checkResultVec_intLMULInput_78,
      source_14[31:11]};
  wire               checkVec_checkResultVec_14_5_2 = checkVec_checkResultVec_overlap_78 | ~checkVec_checkResultVec_14_6_2;
  wire               checkVec_checkResultVec_15_6_2 = checkVec_validVec_2[15];
  wire [10:0]        checkVec_checkResultVec_dataPosition_79 = {source_15[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_15_2_2 = checkVec_checkResultVec_dataPosition_79[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_79 = checkVec_checkResultVec_dataPosition_79[10:7];
  wire               checkVec_checkResultVec_15_3_2 = checkVec_checkResultVec_dataGroup_79[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_79 = checkVec_checkResultVec_dataGroup_79[3:1];
  wire [2:0]         checkVec_checkResultVec_15_4_2 = checkVec_checkResultVec_accessRegGrowth_79;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_79 = {checkVec_checkResultVec_15_3_2, checkVec_checkResultVec_15_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_79 = checkVec_checkResultVec_decimalProportion_79[5:3];
  wire               checkVec_checkResultVec_overlap_79 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_79 >= checkVec_checkResultVec_intLMULInput_79[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_79} >= checkVec_checkResultVec_intLMULInput_79,
      source_15[31:11]};
  wire               checkVec_checkResultVec_15_5_2 = checkVec_checkResultVec_overlap_79 | ~checkVec_checkResultVec_15_6_2;
  wire               checkVec_checkResultVec_16_6_2 = checkVec_validVec_2[16];
  wire [10:0]        checkVec_checkResultVec_dataPosition_80 = {source_16[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_16_2_2 = checkVec_checkResultVec_dataPosition_80[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_80 = checkVec_checkResultVec_dataPosition_80[10:7];
  wire               checkVec_checkResultVec_16_3_2 = checkVec_checkResultVec_dataGroup_80[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_80 = checkVec_checkResultVec_dataGroup_80[3:1];
  wire [2:0]         checkVec_checkResultVec_16_4_2 = checkVec_checkResultVec_accessRegGrowth_80;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_80 = {checkVec_checkResultVec_16_3_2, checkVec_checkResultVec_16_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_80 = checkVec_checkResultVec_decimalProportion_80[5:3];
  wire               checkVec_checkResultVec_overlap_80 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_80 >= checkVec_checkResultVec_intLMULInput_80[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_80} >= checkVec_checkResultVec_intLMULInput_80,
      source_16[31:11]};
  wire               checkVec_checkResultVec_16_5_2 = checkVec_checkResultVec_overlap_80 | ~checkVec_checkResultVec_16_6_2;
  wire               checkVec_checkResultVec_17_6_2 = checkVec_validVec_2[17];
  wire [10:0]        checkVec_checkResultVec_dataPosition_81 = {source_17[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_17_2_2 = checkVec_checkResultVec_dataPosition_81[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_81 = checkVec_checkResultVec_dataPosition_81[10:7];
  wire               checkVec_checkResultVec_17_3_2 = checkVec_checkResultVec_dataGroup_81[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_81 = checkVec_checkResultVec_dataGroup_81[3:1];
  wire [2:0]         checkVec_checkResultVec_17_4_2 = checkVec_checkResultVec_accessRegGrowth_81;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_81 = {checkVec_checkResultVec_17_3_2, checkVec_checkResultVec_17_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_81 = checkVec_checkResultVec_decimalProportion_81[5:3];
  wire               checkVec_checkResultVec_overlap_81 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_81 >= checkVec_checkResultVec_intLMULInput_81[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_81} >= checkVec_checkResultVec_intLMULInput_81,
      source_17[31:11]};
  wire               checkVec_checkResultVec_17_5_2 = checkVec_checkResultVec_overlap_81 | ~checkVec_checkResultVec_17_6_2;
  wire               checkVec_checkResultVec_18_6_2 = checkVec_validVec_2[18];
  wire [10:0]        checkVec_checkResultVec_dataPosition_82 = {source_18[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_18_2_2 = checkVec_checkResultVec_dataPosition_82[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_82 = checkVec_checkResultVec_dataPosition_82[10:7];
  wire               checkVec_checkResultVec_18_3_2 = checkVec_checkResultVec_dataGroup_82[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_82 = checkVec_checkResultVec_dataGroup_82[3:1];
  wire [2:0]         checkVec_checkResultVec_18_4_2 = checkVec_checkResultVec_accessRegGrowth_82;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_82 = {checkVec_checkResultVec_18_3_2, checkVec_checkResultVec_18_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_82 = checkVec_checkResultVec_decimalProportion_82[5:3];
  wire               checkVec_checkResultVec_overlap_82 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_82 >= checkVec_checkResultVec_intLMULInput_82[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_82} >= checkVec_checkResultVec_intLMULInput_82,
      source_18[31:11]};
  wire               checkVec_checkResultVec_18_5_2 = checkVec_checkResultVec_overlap_82 | ~checkVec_checkResultVec_18_6_2;
  wire               checkVec_checkResultVec_19_6_2 = checkVec_validVec_2[19];
  wire [10:0]        checkVec_checkResultVec_dataPosition_83 = {source_19[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_19_2_2 = checkVec_checkResultVec_dataPosition_83[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_83 = checkVec_checkResultVec_dataPosition_83[10:7];
  wire               checkVec_checkResultVec_19_3_2 = checkVec_checkResultVec_dataGroup_83[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_83 = checkVec_checkResultVec_dataGroup_83[3:1];
  wire [2:0]         checkVec_checkResultVec_19_4_2 = checkVec_checkResultVec_accessRegGrowth_83;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_83 = {checkVec_checkResultVec_19_3_2, checkVec_checkResultVec_19_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_83 = checkVec_checkResultVec_decimalProportion_83[5:3];
  wire               checkVec_checkResultVec_overlap_83 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_83 >= checkVec_checkResultVec_intLMULInput_83[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_83} >= checkVec_checkResultVec_intLMULInput_83,
      source_19[31:11]};
  wire               checkVec_checkResultVec_19_5_2 = checkVec_checkResultVec_overlap_83 | ~checkVec_checkResultVec_19_6_2;
  wire               checkVec_checkResultVec_20_6_2 = checkVec_validVec_2[20];
  wire [10:0]        checkVec_checkResultVec_dataPosition_84 = {source_20[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_20_2_2 = checkVec_checkResultVec_dataPosition_84[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_84 = checkVec_checkResultVec_dataPosition_84[10:7];
  wire               checkVec_checkResultVec_20_3_2 = checkVec_checkResultVec_dataGroup_84[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_84 = checkVec_checkResultVec_dataGroup_84[3:1];
  wire [2:0]         checkVec_checkResultVec_20_4_2 = checkVec_checkResultVec_accessRegGrowth_84;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_84 = {checkVec_checkResultVec_20_3_2, checkVec_checkResultVec_20_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_84 = checkVec_checkResultVec_decimalProportion_84[5:3];
  wire               checkVec_checkResultVec_overlap_84 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_84 >= checkVec_checkResultVec_intLMULInput_84[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_84} >= checkVec_checkResultVec_intLMULInput_84,
      source_20[31:11]};
  wire               checkVec_checkResultVec_20_5_2 = checkVec_checkResultVec_overlap_84 | ~checkVec_checkResultVec_20_6_2;
  wire               checkVec_checkResultVec_21_6_2 = checkVec_validVec_2[21];
  wire [10:0]        checkVec_checkResultVec_dataPosition_85 = {source_21[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_21_2_2 = checkVec_checkResultVec_dataPosition_85[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_85 = checkVec_checkResultVec_dataPosition_85[10:7];
  wire               checkVec_checkResultVec_21_3_2 = checkVec_checkResultVec_dataGroup_85[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_85 = checkVec_checkResultVec_dataGroup_85[3:1];
  wire [2:0]         checkVec_checkResultVec_21_4_2 = checkVec_checkResultVec_accessRegGrowth_85;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_85 = {checkVec_checkResultVec_21_3_2, checkVec_checkResultVec_21_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_85 = checkVec_checkResultVec_decimalProportion_85[5:3];
  wire               checkVec_checkResultVec_overlap_85 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_85 >= checkVec_checkResultVec_intLMULInput_85[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_85} >= checkVec_checkResultVec_intLMULInput_85,
      source_21[31:11]};
  wire               checkVec_checkResultVec_21_5_2 = checkVec_checkResultVec_overlap_85 | ~checkVec_checkResultVec_21_6_2;
  wire               checkVec_checkResultVec_22_6_2 = checkVec_validVec_2[22];
  wire [10:0]        checkVec_checkResultVec_dataPosition_86 = {source_22[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_22_2_2 = checkVec_checkResultVec_dataPosition_86[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_86 = checkVec_checkResultVec_dataPosition_86[10:7];
  wire               checkVec_checkResultVec_22_3_2 = checkVec_checkResultVec_dataGroup_86[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_86 = checkVec_checkResultVec_dataGroup_86[3:1];
  wire [2:0]         checkVec_checkResultVec_22_4_2 = checkVec_checkResultVec_accessRegGrowth_86;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_86 = {checkVec_checkResultVec_22_3_2, checkVec_checkResultVec_22_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_86 = checkVec_checkResultVec_decimalProportion_86[5:3];
  wire               checkVec_checkResultVec_overlap_86 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_86 >= checkVec_checkResultVec_intLMULInput_86[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_86} >= checkVec_checkResultVec_intLMULInput_86,
      source_22[31:11]};
  wire               checkVec_checkResultVec_22_5_2 = checkVec_checkResultVec_overlap_86 | ~checkVec_checkResultVec_22_6_2;
  wire               checkVec_checkResultVec_23_6_2 = checkVec_validVec_2[23];
  wire [10:0]        checkVec_checkResultVec_dataPosition_87 = {source_23[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_23_2_2 = checkVec_checkResultVec_dataPosition_87[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_87 = checkVec_checkResultVec_dataPosition_87[10:7];
  wire               checkVec_checkResultVec_23_3_2 = checkVec_checkResultVec_dataGroup_87[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_87 = checkVec_checkResultVec_dataGroup_87[3:1];
  wire [2:0]         checkVec_checkResultVec_23_4_2 = checkVec_checkResultVec_accessRegGrowth_87;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_87 = {checkVec_checkResultVec_23_3_2, checkVec_checkResultVec_23_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_87 = checkVec_checkResultVec_decimalProportion_87[5:3];
  wire               checkVec_checkResultVec_overlap_87 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_87 >= checkVec_checkResultVec_intLMULInput_87[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_87} >= checkVec_checkResultVec_intLMULInput_87,
      source_23[31:11]};
  wire               checkVec_checkResultVec_23_5_2 = checkVec_checkResultVec_overlap_87 | ~checkVec_checkResultVec_23_6_2;
  wire               checkVec_checkResultVec_24_6_2 = checkVec_validVec_2[24];
  wire [10:0]        checkVec_checkResultVec_dataPosition_88 = {source_24[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_24_2_2 = checkVec_checkResultVec_dataPosition_88[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_88 = checkVec_checkResultVec_dataPosition_88[10:7];
  wire               checkVec_checkResultVec_24_3_2 = checkVec_checkResultVec_dataGroup_88[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_88 = checkVec_checkResultVec_dataGroup_88[3:1];
  wire [2:0]         checkVec_checkResultVec_24_4_2 = checkVec_checkResultVec_accessRegGrowth_88;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_88 = {checkVec_checkResultVec_24_3_2, checkVec_checkResultVec_24_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_88 = checkVec_checkResultVec_decimalProportion_88[5:3];
  wire               checkVec_checkResultVec_overlap_88 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_88 >= checkVec_checkResultVec_intLMULInput_88[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_88} >= checkVec_checkResultVec_intLMULInput_88,
      source_24[31:11]};
  wire               checkVec_checkResultVec_24_5_2 = checkVec_checkResultVec_overlap_88 | ~checkVec_checkResultVec_24_6_2;
  wire               checkVec_checkResultVec_25_6_2 = checkVec_validVec_2[25];
  wire [10:0]        checkVec_checkResultVec_dataPosition_89 = {source_25[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_25_2_2 = checkVec_checkResultVec_dataPosition_89[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_89 = checkVec_checkResultVec_dataPosition_89[10:7];
  wire               checkVec_checkResultVec_25_3_2 = checkVec_checkResultVec_dataGroup_89[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_89 = checkVec_checkResultVec_dataGroup_89[3:1];
  wire [2:0]         checkVec_checkResultVec_25_4_2 = checkVec_checkResultVec_accessRegGrowth_89;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_89 = {checkVec_checkResultVec_25_3_2, checkVec_checkResultVec_25_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_89 = checkVec_checkResultVec_decimalProportion_89[5:3];
  wire               checkVec_checkResultVec_overlap_89 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_89 >= checkVec_checkResultVec_intLMULInput_89[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_89} >= checkVec_checkResultVec_intLMULInput_89,
      source_25[31:11]};
  wire               checkVec_checkResultVec_25_5_2 = checkVec_checkResultVec_overlap_89 | ~checkVec_checkResultVec_25_6_2;
  wire               checkVec_checkResultVec_26_6_2 = checkVec_validVec_2[26];
  wire [10:0]        checkVec_checkResultVec_dataPosition_90 = {source_26[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_26_2_2 = checkVec_checkResultVec_dataPosition_90[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_90 = checkVec_checkResultVec_dataPosition_90[10:7];
  wire               checkVec_checkResultVec_26_3_2 = checkVec_checkResultVec_dataGroup_90[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_90 = checkVec_checkResultVec_dataGroup_90[3:1];
  wire [2:0]         checkVec_checkResultVec_26_4_2 = checkVec_checkResultVec_accessRegGrowth_90;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_90 = {checkVec_checkResultVec_26_3_2, checkVec_checkResultVec_26_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_90 = checkVec_checkResultVec_decimalProportion_90[5:3];
  wire               checkVec_checkResultVec_overlap_90 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_90 >= checkVec_checkResultVec_intLMULInput_90[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_90} >= checkVec_checkResultVec_intLMULInput_90,
      source_26[31:11]};
  wire               checkVec_checkResultVec_26_5_2 = checkVec_checkResultVec_overlap_90 | ~checkVec_checkResultVec_26_6_2;
  wire               checkVec_checkResultVec_27_6_2 = checkVec_validVec_2[27];
  wire [10:0]        checkVec_checkResultVec_dataPosition_91 = {source_27[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_27_2_2 = checkVec_checkResultVec_dataPosition_91[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_91 = checkVec_checkResultVec_dataPosition_91[10:7];
  wire               checkVec_checkResultVec_27_3_2 = checkVec_checkResultVec_dataGroup_91[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_91 = checkVec_checkResultVec_dataGroup_91[3:1];
  wire [2:0]         checkVec_checkResultVec_27_4_2 = checkVec_checkResultVec_accessRegGrowth_91;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_91 = {checkVec_checkResultVec_27_3_2, checkVec_checkResultVec_27_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_91 = checkVec_checkResultVec_decimalProportion_91[5:3];
  wire               checkVec_checkResultVec_overlap_91 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_91 >= checkVec_checkResultVec_intLMULInput_91[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_91} >= checkVec_checkResultVec_intLMULInput_91,
      source_27[31:11]};
  wire               checkVec_checkResultVec_27_5_2 = checkVec_checkResultVec_overlap_91 | ~checkVec_checkResultVec_27_6_2;
  wire               checkVec_checkResultVec_28_6_2 = checkVec_validVec_2[28];
  wire [10:0]        checkVec_checkResultVec_dataPosition_92 = {source_28[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_28_2_2 = checkVec_checkResultVec_dataPosition_92[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_92 = checkVec_checkResultVec_dataPosition_92[10:7];
  wire               checkVec_checkResultVec_28_3_2 = checkVec_checkResultVec_dataGroup_92[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_92 = checkVec_checkResultVec_dataGroup_92[3:1];
  wire [2:0]         checkVec_checkResultVec_28_4_2 = checkVec_checkResultVec_accessRegGrowth_92;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_92 = {checkVec_checkResultVec_28_3_2, checkVec_checkResultVec_28_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_92 = checkVec_checkResultVec_decimalProportion_92[5:3];
  wire               checkVec_checkResultVec_overlap_92 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_92 >= checkVec_checkResultVec_intLMULInput_92[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_92} >= checkVec_checkResultVec_intLMULInput_92,
      source_28[31:11]};
  wire               checkVec_checkResultVec_28_5_2 = checkVec_checkResultVec_overlap_92 | ~checkVec_checkResultVec_28_6_2;
  wire               checkVec_checkResultVec_29_6_2 = checkVec_validVec_2[29];
  wire [10:0]        checkVec_checkResultVec_dataPosition_93 = {source_29[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_29_2_2 = checkVec_checkResultVec_dataPosition_93[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_93 = checkVec_checkResultVec_dataPosition_93[10:7];
  wire               checkVec_checkResultVec_29_3_2 = checkVec_checkResultVec_dataGroup_93[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_93 = checkVec_checkResultVec_dataGroup_93[3:1];
  wire [2:0]         checkVec_checkResultVec_29_4_2 = checkVec_checkResultVec_accessRegGrowth_93;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_93 = {checkVec_checkResultVec_29_3_2, checkVec_checkResultVec_29_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_93 = checkVec_checkResultVec_decimalProportion_93[5:3];
  wire               checkVec_checkResultVec_overlap_93 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_93 >= checkVec_checkResultVec_intLMULInput_93[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_93} >= checkVec_checkResultVec_intLMULInput_93,
      source_29[31:11]};
  wire               checkVec_checkResultVec_29_5_2 = checkVec_checkResultVec_overlap_93 | ~checkVec_checkResultVec_29_6_2;
  wire               checkVec_checkResultVec_30_6_2 = checkVec_validVec_2[30];
  wire [10:0]        checkVec_checkResultVec_dataPosition_94 = {source_30[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_30_2_2 = checkVec_checkResultVec_dataPosition_94[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_94 = checkVec_checkResultVec_dataPosition_94[10:7];
  wire               checkVec_checkResultVec_30_3_2 = checkVec_checkResultVec_dataGroup_94[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_94 = checkVec_checkResultVec_dataGroup_94[3:1];
  wire [2:0]         checkVec_checkResultVec_30_4_2 = checkVec_checkResultVec_accessRegGrowth_94;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_94 = {checkVec_checkResultVec_30_3_2, checkVec_checkResultVec_30_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_94 = checkVec_checkResultVec_decimalProportion_94[5:3];
  wire               checkVec_checkResultVec_overlap_94 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_94 >= checkVec_checkResultVec_intLMULInput_94[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_94} >= checkVec_checkResultVec_intLMULInput_94,
      source_30[31:11]};
  wire               checkVec_checkResultVec_30_5_2 = checkVec_checkResultVec_overlap_94 | ~checkVec_checkResultVec_30_6_2;
  wire               checkVec_checkResultVec_31_6_2 = checkVec_validVec_2[31];
  wire [10:0]        checkVec_checkResultVec_dataPosition_95 = {source_31[8:0], 2'h0};
  wire [4:0]         checkVec_checkResultVec_31_2_2 = checkVec_checkResultVec_dataPosition_95[6:2];
  wire [3:0]         checkVec_checkResultVec_dataGroup_95 = checkVec_checkResultVec_dataPosition_95[10:7];
  wire               checkVec_checkResultVec_31_3_2 = checkVec_checkResultVec_dataGroup_95[0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_95 = checkVec_checkResultVec_dataGroup_95[3:1];
  wire [2:0]         checkVec_checkResultVec_31_4_2 = checkVec_checkResultVec_accessRegGrowth_95;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_95 = {checkVec_checkResultVec_31_3_2, checkVec_checkResultVec_31_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_95 = checkVec_checkResultVec_decimalProportion_95[5:3];
  wire               checkVec_checkResultVec_overlap_95 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_95 >= checkVec_checkResultVec_intLMULInput_95[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_95} >= checkVec_checkResultVec_intLMULInput_95,
      source_31[31:11]};
  wire               checkVec_checkResultVec_31_5_2 = checkVec_checkResultVec_overlap_95 | ~checkVec_checkResultVec_31_6_2;
  wire [9:0]         checkVec_checkResult_lo_lo_lo_lo_16 = {checkVec_checkResultVec_1_2_2, checkVec_checkResultVec_0_2_2};
  wire [9:0]         checkVec_checkResult_lo_lo_lo_hi_16 = {checkVec_checkResultVec_3_2_2, checkVec_checkResultVec_2_2_2};
  wire [19:0]        checkVec_checkResult_lo_lo_lo_16 = {checkVec_checkResult_lo_lo_lo_hi_16, checkVec_checkResult_lo_lo_lo_lo_16};
  wire [9:0]         checkVec_checkResult_lo_lo_hi_lo_16 = {checkVec_checkResultVec_5_2_2, checkVec_checkResultVec_4_2_2};
  wire [9:0]         checkVec_checkResult_lo_lo_hi_hi_16 = {checkVec_checkResultVec_7_2_2, checkVec_checkResultVec_6_2_2};
  wire [19:0]        checkVec_checkResult_lo_lo_hi_16 = {checkVec_checkResult_lo_lo_hi_hi_16, checkVec_checkResult_lo_lo_hi_lo_16};
  wire [39:0]        checkVec_checkResult_lo_lo_16 = {checkVec_checkResult_lo_lo_hi_16, checkVec_checkResult_lo_lo_lo_16};
  wire [9:0]         checkVec_checkResult_lo_hi_lo_lo_16 = {checkVec_checkResultVec_9_2_2, checkVec_checkResultVec_8_2_2};
  wire [9:0]         checkVec_checkResult_lo_hi_lo_hi_16 = {checkVec_checkResultVec_11_2_2, checkVec_checkResultVec_10_2_2};
  wire [19:0]        checkVec_checkResult_lo_hi_lo_16 = {checkVec_checkResult_lo_hi_lo_hi_16, checkVec_checkResult_lo_hi_lo_lo_16};
  wire [9:0]         checkVec_checkResult_lo_hi_hi_lo_16 = {checkVec_checkResultVec_13_2_2, checkVec_checkResultVec_12_2_2};
  wire [9:0]         checkVec_checkResult_lo_hi_hi_hi_16 = {checkVec_checkResultVec_15_2_2, checkVec_checkResultVec_14_2_2};
  wire [19:0]        checkVec_checkResult_lo_hi_hi_16 = {checkVec_checkResult_lo_hi_hi_hi_16, checkVec_checkResult_lo_hi_hi_lo_16};
  wire [39:0]        checkVec_checkResult_lo_hi_16 = {checkVec_checkResult_lo_hi_hi_16, checkVec_checkResult_lo_hi_lo_16};
  wire [79:0]        checkVec_checkResult_lo_16 = {checkVec_checkResult_lo_hi_16, checkVec_checkResult_lo_lo_16};
  wire [9:0]         checkVec_checkResult_hi_lo_lo_lo_16 = {checkVec_checkResultVec_17_2_2, checkVec_checkResultVec_16_2_2};
  wire [9:0]         checkVec_checkResult_hi_lo_lo_hi_16 = {checkVec_checkResultVec_19_2_2, checkVec_checkResultVec_18_2_2};
  wire [19:0]        checkVec_checkResult_hi_lo_lo_16 = {checkVec_checkResult_hi_lo_lo_hi_16, checkVec_checkResult_hi_lo_lo_lo_16};
  wire [9:0]         checkVec_checkResult_hi_lo_hi_lo_16 = {checkVec_checkResultVec_21_2_2, checkVec_checkResultVec_20_2_2};
  wire [9:0]         checkVec_checkResult_hi_lo_hi_hi_16 = {checkVec_checkResultVec_23_2_2, checkVec_checkResultVec_22_2_2};
  wire [19:0]        checkVec_checkResult_hi_lo_hi_16 = {checkVec_checkResult_hi_lo_hi_hi_16, checkVec_checkResult_hi_lo_hi_lo_16};
  wire [39:0]        checkVec_checkResult_hi_lo_16 = {checkVec_checkResult_hi_lo_hi_16, checkVec_checkResult_hi_lo_lo_16};
  wire [9:0]         checkVec_checkResult_hi_hi_lo_lo_16 = {checkVec_checkResultVec_25_2_2, checkVec_checkResultVec_24_2_2};
  wire [9:0]         checkVec_checkResult_hi_hi_lo_hi_16 = {checkVec_checkResultVec_27_2_2, checkVec_checkResultVec_26_2_2};
  wire [19:0]        checkVec_checkResult_hi_hi_lo_16 = {checkVec_checkResult_hi_hi_lo_hi_16, checkVec_checkResult_hi_hi_lo_lo_16};
  wire [9:0]         checkVec_checkResult_hi_hi_hi_lo_16 = {checkVec_checkResultVec_29_2_2, checkVec_checkResultVec_28_2_2};
  wire [9:0]         checkVec_checkResult_hi_hi_hi_hi_16 = {checkVec_checkResultVec_31_2_2, checkVec_checkResultVec_30_2_2};
  wire [19:0]        checkVec_checkResult_hi_hi_hi_16 = {checkVec_checkResult_hi_hi_hi_hi_16, checkVec_checkResult_hi_hi_hi_lo_16};
  wire [39:0]        checkVec_checkResult_hi_hi_16 = {checkVec_checkResult_hi_hi_hi_16, checkVec_checkResult_hi_hi_lo_16};
  wire [79:0]        checkVec_checkResult_hi_16 = {checkVec_checkResult_hi_hi_16, checkVec_checkResult_hi_lo_16};
  wire [159:0]       checkVec_2_2 = {checkVec_checkResult_hi_16, checkVec_checkResult_lo_16};
  wire [1:0]         checkVec_checkResult_lo_lo_lo_lo_17 = {checkVec_checkResultVec_1_3_2, checkVec_checkResultVec_0_3_2};
  wire [1:0]         checkVec_checkResult_lo_lo_lo_hi_17 = {checkVec_checkResultVec_3_3_2, checkVec_checkResultVec_2_3_2};
  wire [3:0]         checkVec_checkResult_lo_lo_lo_17 = {checkVec_checkResult_lo_lo_lo_hi_17, checkVec_checkResult_lo_lo_lo_lo_17};
  wire [1:0]         checkVec_checkResult_lo_lo_hi_lo_17 = {checkVec_checkResultVec_5_3_2, checkVec_checkResultVec_4_3_2};
  wire [1:0]         checkVec_checkResult_lo_lo_hi_hi_17 = {checkVec_checkResultVec_7_3_2, checkVec_checkResultVec_6_3_2};
  wire [3:0]         checkVec_checkResult_lo_lo_hi_17 = {checkVec_checkResult_lo_lo_hi_hi_17, checkVec_checkResult_lo_lo_hi_lo_17};
  wire [7:0]         checkVec_checkResult_lo_lo_17 = {checkVec_checkResult_lo_lo_hi_17, checkVec_checkResult_lo_lo_lo_17};
  wire [1:0]         checkVec_checkResult_lo_hi_lo_lo_17 = {checkVec_checkResultVec_9_3_2, checkVec_checkResultVec_8_3_2};
  wire [1:0]         checkVec_checkResult_lo_hi_lo_hi_17 = {checkVec_checkResultVec_11_3_2, checkVec_checkResultVec_10_3_2};
  wire [3:0]         checkVec_checkResult_lo_hi_lo_17 = {checkVec_checkResult_lo_hi_lo_hi_17, checkVec_checkResult_lo_hi_lo_lo_17};
  wire [1:0]         checkVec_checkResult_lo_hi_hi_lo_17 = {checkVec_checkResultVec_13_3_2, checkVec_checkResultVec_12_3_2};
  wire [1:0]         checkVec_checkResult_lo_hi_hi_hi_17 = {checkVec_checkResultVec_15_3_2, checkVec_checkResultVec_14_3_2};
  wire [3:0]         checkVec_checkResult_lo_hi_hi_17 = {checkVec_checkResult_lo_hi_hi_hi_17, checkVec_checkResult_lo_hi_hi_lo_17};
  wire [7:0]         checkVec_checkResult_lo_hi_17 = {checkVec_checkResult_lo_hi_hi_17, checkVec_checkResult_lo_hi_lo_17};
  wire [15:0]        checkVec_checkResult_lo_17 = {checkVec_checkResult_lo_hi_17, checkVec_checkResult_lo_lo_17};
  wire [1:0]         checkVec_checkResult_hi_lo_lo_lo_17 = {checkVec_checkResultVec_17_3_2, checkVec_checkResultVec_16_3_2};
  wire [1:0]         checkVec_checkResult_hi_lo_lo_hi_17 = {checkVec_checkResultVec_19_3_2, checkVec_checkResultVec_18_3_2};
  wire [3:0]         checkVec_checkResult_hi_lo_lo_17 = {checkVec_checkResult_hi_lo_lo_hi_17, checkVec_checkResult_hi_lo_lo_lo_17};
  wire [1:0]         checkVec_checkResult_hi_lo_hi_lo_17 = {checkVec_checkResultVec_21_3_2, checkVec_checkResultVec_20_3_2};
  wire [1:0]         checkVec_checkResult_hi_lo_hi_hi_17 = {checkVec_checkResultVec_23_3_2, checkVec_checkResultVec_22_3_2};
  wire [3:0]         checkVec_checkResult_hi_lo_hi_17 = {checkVec_checkResult_hi_lo_hi_hi_17, checkVec_checkResult_hi_lo_hi_lo_17};
  wire [7:0]         checkVec_checkResult_hi_lo_17 = {checkVec_checkResult_hi_lo_hi_17, checkVec_checkResult_hi_lo_lo_17};
  wire [1:0]         checkVec_checkResult_hi_hi_lo_lo_17 = {checkVec_checkResultVec_25_3_2, checkVec_checkResultVec_24_3_2};
  wire [1:0]         checkVec_checkResult_hi_hi_lo_hi_17 = {checkVec_checkResultVec_27_3_2, checkVec_checkResultVec_26_3_2};
  wire [3:0]         checkVec_checkResult_hi_hi_lo_17 = {checkVec_checkResult_hi_hi_lo_hi_17, checkVec_checkResult_hi_hi_lo_lo_17};
  wire [1:0]         checkVec_checkResult_hi_hi_hi_lo_17 = {checkVec_checkResultVec_29_3_2, checkVec_checkResultVec_28_3_2};
  wire [1:0]         checkVec_checkResult_hi_hi_hi_hi_17 = {checkVec_checkResultVec_31_3_2, checkVec_checkResultVec_30_3_2};
  wire [3:0]         checkVec_checkResult_hi_hi_hi_17 = {checkVec_checkResult_hi_hi_hi_hi_17, checkVec_checkResult_hi_hi_hi_lo_17};
  wire [7:0]         checkVec_checkResult_hi_hi_17 = {checkVec_checkResult_hi_hi_hi_17, checkVec_checkResult_hi_hi_lo_17};
  wire [15:0]        checkVec_checkResult_hi_17 = {checkVec_checkResult_hi_hi_17, checkVec_checkResult_hi_lo_17};
  wire [31:0]        checkVec_2_3 = {checkVec_checkResult_hi_17, checkVec_checkResult_lo_17};
  wire [5:0]         checkVec_checkResult_lo_lo_lo_lo_18 = {checkVec_checkResultVec_1_4_2, checkVec_checkResultVec_0_4_2};
  wire [5:0]         checkVec_checkResult_lo_lo_lo_hi_18 = {checkVec_checkResultVec_3_4_2, checkVec_checkResultVec_2_4_2};
  wire [11:0]        checkVec_checkResult_lo_lo_lo_18 = {checkVec_checkResult_lo_lo_lo_hi_18, checkVec_checkResult_lo_lo_lo_lo_18};
  wire [5:0]         checkVec_checkResult_lo_lo_hi_lo_18 = {checkVec_checkResultVec_5_4_2, checkVec_checkResultVec_4_4_2};
  wire [5:0]         checkVec_checkResult_lo_lo_hi_hi_18 = {checkVec_checkResultVec_7_4_2, checkVec_checkResultVec_6_4_2};
  wire [11:0]        checkVec_checkResult_lo_lo_hi_18 = {checkVec_checkResult_lo_lo_hi_hi_18, checkVec_checkResult_lo_lo_hi_lo_18};
  wire [23:0]        checkVec_checkResult_lo_lo_18 = {checkVec_checkResult_lo_lo_hi_18, checkVec_checkResult_lo_lo_lo_18};
  wire [5:0]         checkVec_checkResult_lo_hi_lo_lo_18 = {checkVec_checkResultVec_9_4_2, checkVec_checkResultVec_8_4_2};
  wire [5:0]         checkVec_checkResult_lo_hi_lo_hi_18 = {checkVec_checkResultVec_11_4_2, checkVec_checkResultVec_10_4_2};
  wire [11:0]        checkVec_checkResult_lo_hi_lo_18 = {checkVec_checkResult_lo_hi_lo_hi_18, checkVec_checkResult_lo_hi_lo_lo_18};
  wire [5:0]         checkVec_checkResult_lo_hi_hi_lo_18 = {checkVec_checkResultVec_13_4_2, checkVec_checkResultVec_12_4_2};
  wire [5:0]         checkVec_checkResult_lo_hi_hi_hi_18 = {checkVec_checkResultVec_15_4_2, checkVec_checkResultVec_14_4_2};
  wire [11:0]        checkVec_checkResult_lo_hi_hi_18 = {checkVec_checkResult_lo_hi_hi_hi_18, checkVec_checkResult_lo_hi_hi_lo_18};
  wire [23:0]        checkVec_checkResult_lo_hi_18 = {checkVec_checkResult_lo_hi_hi_18, checkVec_checkResult_lo_hi_lo_18};
  wire [47:0]        checkVec_checkResult_lo_18 = {checkVec_checkResult_lo_hi_18, checkVec_checkResult_lo_lo_18};
  wire [5:0]         checkVec_checkResult_hi_lo_lo_lo_18 = {checkVec_checkResultVec_17_4_2, checkVec_checkResultVec_16_4_2};
  wire [5:0]         checkVec_checkResult_hi_lo_lo_hi_18 = {checkVec_checkResultVec_19_4_2, checkVec_checkResultVec_18_4_2};
  wire [11:0]        checkVec_checkResult_hi_lo_lo_18 = {checkVec_checkResult_hi_lo_lo_hi_18, checkVec_checkResult_hi_lo_lo_lo_18};
  wire [5:0]         checkVec_checkResult_hi_lo_hi_lo_18 = {checkVec_checkResultVec_21_4_2, checkVec_checkResultVec_20_4_2};
  wire [5:0]         checkVec_checkResult_hi_lo_hi_hi_18 = {checkVec_checkResultVec_23_4_2, checkVec_checkResultVec_22_4_2};
  wire [11:0]        checkVec_checkResult_hi_lo_hi_18 = {checkVec_checkResult_hi_lo_hi_hi_18, checkVec_checkResult_hi_lo_hi_lo_18};
  wire [23:0]        checkVec_checkResult_hi_lo_18 = {checkVec_checkResult_hi_lo_hi_18, checkVec_checkResult_hi_lo_lo_18};
  wire [5:0]         checkVec_checkResult_hi_hi_lo_lo_18 = {checkVec_checkResultVec_25_4_2, checkVec_checkResultVec_24_4_2};
  wire [5:0]         checkVec_checkResult_hi_hi_lo_hi_18 = {checkVec_checkResultVec_27_4_2, checkVec_checkResultVec_26_4_2};
  wire [11:0]        checkVec_checkResult_hi_hi_lo_18 = {checkVec_checkResult_hi_hi_lo_hi_18, checkVec_checkResult_hi_hi_lo_lo_18};
  wire [5:0]         checkVec_checkResult_hi_hi_hi_lo_18 = {checkVec_checkResultVec_29_4_2, checkVec_checkResultVec_28_4_2};
  wire [5:0]         checkVec_checkResult_hi_hi_hi_hi_18 = {checkVec_checkResultVec_31_4_2, checkVec_checkResultVec_30_4_2};
  wire [11:0]        checkVec_checkResult_hi_hi_hi_18 = {checkVec_checkResult_hi_hi_hi_hi_18, checkVec_checkResult_hi_hi_hi_lo_18};
  wire [23:0]        checkVec_checkResult_hi_hi_18 = {checkVec_checkResult_hi_hi_hi_18, checkVec_checkResult_hi_hi_lo_18};
  wire [47:0]        checkVec_checkResult_hi_18 = {checkVec_checkResult_hi_hi_18, checkVec_checkResult_hi_lo_18};
  wire [95:0]        checkVec_2_4 = {checkVec_checkResult_hi_18, checkVec_checkResult_lo_18};
  wire [1:0]         checkVec_checkResult_lo_lo_lo_lo_19 = {checkVec_checkResultVec_1_5_2, checkVec_checkResultVec_0_5_2};
  wire [1:0]         checkVec_checkResult_lo_lo_lo_hi_19 = {checkVec_checkResultVec_3_5_2, checkVec_checkResultVec_2_5_2};
  wire [3:0]         checkVec_checkResult_lo_lo_lo_19 = {checkVec_checkResult_lo_lo_lo_hi_19, checkVec_checkResult_lo_lo_lo_lo_19};
  wire [1:0]         checkVec_checkResult_lo_lo_hi_lo_19 = {checkVec_checkResultVec_5_5_2, checkVec_checkResultVec_4_5_2};
  wire [1:0]         checkVec_checkResult_lo_lo_hi_hi_19 = {checkVec_checkResultVec_7_5_2, checkVec_checkResultVec_6_5_2};
  wire [3:0]         checkVec_checkResult_lo_lo_hi_19 = {checkVec_checkResult_lo_lo_hi_hi_19, checkVec_checkResult_lo_lo_hi_lo_19};
  wire [7:0]         checkVec_checkResult_lo_lo_19 = {checkVec_checkResult_lo_lo_hi_19, checkVec_checkResult_lo_lo_lo_19};
  wire [1:0]         checkVec_checkResult_lo_hi_lo_lo_19 = {checkVec_checkResultVec_9_5_2, checkVec_checkResultVec_8_5_2};
  wire [1:0]         checkVec_checkResult_lo_hi_lo_hi_19 = {checkVec_checkResultVec_11_5_2, checkVec_checkResultVec_10_5_2};
  wire [3:0]         checkVec_checkResult_lo_hi_lo_19 = {checkVec_checkResult_lo_hi_lo_hi_19, checkVec_checkResult_lo_hi_lo_lo_19};
  wire [1:0]         checkVec_checkResult_lo_hi_hi_lo_19 = {checkVec_checkResultVec_13_5_2, checkVec_checkResultVec_12_5_2};
  wire [1:0]         checkVec_checkResult_lo_hi_hi_hi_19 = {checkVec_checkResultVec_15_5_2, checkVec_checkResultVec_14_5_2};
  wire [3:0]         checkVec_checkResult_lo_hi_hi_19 = {checkVec_checkResult_lo_hi_hi_hi_19, checkVec_checkResult_lo_hi_hi_lo_19};
  wire [7:0]         checkVec_checkResult_lo_hi_19 = {checkVec_checkResult_lo_hi_hi_19, checkVec_checkResult_lo_hi_lo_19};
  wire [15:0]        checkVec_checkResult_lo_19 = {checkVec_checkResult_lo_hi_19, checkVec_checkResult_lo_lo_19};
  wire [1:0]         checkVec_checkResult_hi_lo_lo_lo_19 = {checkVec_checkResultVec_17_5_2, checkVec_checkResultVec_16_5_2};
  wire [1:0]         checkVec_checkResult_hi_lo_lo_hi_19 = {checkVec_checkResultVec_19_5_2, checkVec_checkResultVec_18_5_2};
  wire [3:0]         checkVec_checkResult_hi_lo_lo_19 = {checkVec_checkResult_hi_lo_lo_hi_19, checkVec_checkResult_hi_lo_lo_lo_19};
  wire [1:0]         checkVec_checkResult_hi_lo_hi_lo_19 = {checkVec_checkResultVec_21_5_2, checkVec_checkResultVec_20_5_2};
  wire [1:0]         checkVec_checkResult_hi_lo_hi_hi_19 = {checkVec_checkResultVec_23_5_2, checkVec_checkResultVec_22_5_2};
  wire [3:0]         checkVec_checkResult_hi_lo_hi_19 = {checkVec_checkResult_hi_lo_hi_hi_19, checkVec_checkResult_hi_lo_hi_lo_19};
  wire [7:0]         checkVec_checkResult_hi_lo_19 = {checkVec_checkResult_hi_lo_hi_19, checkVec_checkResult_hi_lo_lo_19};
  wire [1:0]         checkVec_checkResult_hi_hi_lo_lo_19 = {checkVec_checkResultVec_25_5_2, checkVec_checkResultVec_24_5_2};
  wire [1:0]         checkVec_checkResult_hi_hi_lo_hi_19 = {checkVec_checkResultVec_27_5_2, checkVec_checkResultVec_26_5_2};
  wire [3:0]         checkVec_checkResult_hi_hi_lo_19 = {checkVec_checkResult_hi_hi_lo_hi_19, checkVec_checkResult_hi_hi_lo_lo_19};
  wire [1:0]         checkVec_checkResult_hi_hi_hi_lo_19 = {checkVec_checkResultVec_29_5_2, checkVec_checkResultVec_28_5_2};
  wire [1:0]         checkVec_checkResult_hi_hi_hi_hi_19 = {checkVec_checkResultVec_31_5_2, checkVec_checkResultVec_30_5_2};
  wire [3:0]         checkVec_checkResult_hi_hi_hi_19 = {checkVec_checkResult_hi_hi_hi_hi_19, checkVec_checkResult_hi_hi_hi_lo_19};
  wire [7:0]         checkVec_checkResult_hi_hi_19 = {checkVec_checkResult_hi_hi_hi_19, checkVec_checkResult_hi_hi_lo_19};
  wire [15:0]        checkVec_checkResult_hi_19 = {checkVec_checkResult_hi_hi_19, checkVec_checkResult_hi_lo_19};
  wire [31:0]        checkVec_2_5 = {checkVec_checkResult_hi_19, checkVec_checkResult_lo_19};
  wire [1:0]         checkVec_checkResult_lo_lo_lo_lo_20 = {checkVec_checkResultVec_1_6_2, checkVec_checkResultVec_0_6_2};
  wire [1:0]         checkVec_checkResult_lo_lo_lo_hi_20 = {checkVec_checkResultVec_3_6_2, checkVec_checkResultVec_2_6_2};
  wire [3:0]         checkVec_checkResult_lo_lo_lo_20 = {checkVec_checkResult_lo_lo_lo_hi_20, checkVec_checkResult_lo_lo_lo_lo_20};
  wire [1:0]         checkVec_checkResult_lo_lo_hi_lo_20 = {checkVec_checkResultVec_5_6_2, checkVec_checkResultVec_4_6_2};
  wire [1:0]         checkVec_checkResult_lo_lo_hi_hi_20 = {checkVec_checkResultVec_7_6_2, checkVec_checkResultVec_6_6_2};
  wire [3:0]         checkVec_checkResult_lo_lo_hi_20 = {checkVec_checkResult_lo_lo_hi_hi_20, checkVec_checkResult_lo_lo_hi_lo_20};
  wire [7:0]         checkVec_checkResult_lo_lo_20 = {checkVec_checkResult_lo_lo_hi_20, checkVec_checkResult_lo_lo_lo_20};
  wire [1:0]         checkVec_checkResult_lo_hi_lo_lo_20 = {checkVec_checkResultVec_9_6_2, checkVec_checkResultVec_8_6_2};
  wire [1:0]         checkVec_checkResult_lo_hi_lo_hi_20 = {checkVec_checkResultVec_11_6_2, checkVec_checkResultVec_10_6_2};
  wire [3:0]         checkVec_checkResult_lo_hi_lo_20 = {checkVec_checkResult_lo_hi_lo_hi_20, checkVec_checkResult_lo_hi_lo_lo_20};
  wire [1:0]         checkVec_checkResult_lo_hi_hi_lo_20 = {checkVec_checkResultVec_13_6_2, checkVec_checkResultVec_12_6_2};
  wire [1:0]         checkVec_checkResult_lo_hi_hi_hi_20 = {checkVec_checkResultVec_15_6_2, checkVec_checkResultVec_14_6_2};
  wire [3:0]         checkVec_checkResult_lo_hi_hi_20 = {checkVec_checkResult_lo_hi_hi_hi_20, checkVec_checkResult_lo_hi_hi_lo_20};
  wire [7:0]         checkVec_checkResult_lo_hi_20 = {checkVec_checkResult_lo_hi_hi_20, checkVec_checkResult_lo_hi_lo_20};
  wire [15:0]        checkVec_checkResult_lo_20 = {checkVec_checkResult_lo_hi_20, checkVec_checkResult_lo_lo_20};
  wire [1:0]         checkVec_checkResult_hi_lo_lo_lo_20 = {checkVec_checkResultVec_17_6_2, checkVec_checkResultVec_16_6_2};
  wire [1:0]         checkVec_checkResult_hi_lo_lo_hi_20 = {checkVec_checkResultVec_19_6_2, checkVec_checkResultVec_18_6_2};
  wire [3:0]         checkVec_checkResult_hi_lo_lo_20 = {checkVec_checkResult_hi_lo_lo_hi_20, checkVec_checkResult_hi_lo_lo_lo_20};
  wire [1:0]         checkVec_checkResult_hi_lo_hi_lo_20 = {checkVec_checkResultVec_21_6_2, checkVec_checkResultVec_20_6_2};
  wire [1:0]         checkVec_checkResult_hi_lo_hi_hi_20 = {checkVec_checkResultVec_23_6_2, checkVec_checkResultVec_22_6_2};
  wire [3:0]         checkVec_checkResult_hi_lo_hi_20 = {checkVec_checkResult_hi_lo_hi_hi_20, checkVec_checkResult_hi_lo_hi_lo_20};
  wire [7:0]         checkVec_checkResult_hi_lo_20 = {checkVec_checkResult_hi_lo_hi_20, checkVec_checkResult_hi_lo_lo_20};
  wire [1:0]         checkVec_checkResult_hi_hi_lo_lo_20 = {checkVec_checkResultVec_25_6_2, checkVec_checkResultVec_24_6_2};
  wire [1:0]         checkVec_checkResult_hi_hi_lo_hi_20 = {checkVec_checkResultVec_27_6_2, checkVec_checkResultVec_26_6_2};
  wire [3:0]         checkVec_checkResult_hi_hi_lo_20 = {checkVec_checkResult_hi_hi_lo_hi_20, checkVec_checkResult_hi_hi_lo_lo_20};
  wire [1:0]         checkVec_checkResult_hi_hi_hi_lo_20 = {checkVec_checkResultVec_29_6_2, checkVec_checkResultVec_28_6_2};
  wire [1:0]         checkVec_checkResult_hi_hi_hi_hi_20 = {checkVec_checkResultVec_31_6_2, checkVec_checkResultVec_30_6_2};
  wire [3:0]         checkVec_checkResult_hi_hi_hi_20 = {checkVec_checkResult_hi_hi_hi_hi_20, checkVec_checkResult_hi_hi_hi_lo_20};
  wire [7:0]         checkVec_checkResult_hi_hi_20 = {checkVec_checkResult_hi_hi_hi_20, checkVec_checkResult_hi_hi_lo_20};
  wire [15:0]        checkVec_checkResult_hi_20 = {checkVec_checkResult_hi_hi_20, checkVec_checkResult_hi_lo_20};
  wire [31:0]        checkVec_2_6 = {checkVec_checkResult_hi_20, checkVec_checkResult_lo_20};
  wire [63:0]        dataOffsetSelect = (sew1H[0] ? checkVec_0_1 : 64'h0) | (sew1H[1] ? checkVec_1_1 : 64'h0);
  wire [159:0]       accessLaneSelect = (sew1H[0] ? checkVec_0_2 : 160'h0) | (sew1H[1] ? checkVec_1_2 : 160'h0) | (sew1H[2] ? checkVec_2_2 : 160'h0);
  wire [31:0]        offsetSelect = (sew1H[0] ? checkVec_0_3 : 32'h0) | (sew1H[1] ? checkVec_1_3 : 32'h0) | (sew1H[2] ? checkVec_2_3 : 32'h0);
  wire [95:0]        growthSelect = (sew1H[0] ? checkVec_0_4 : 96'h0) | (sew1H[1] ? checkVec_1_4 : 96'h0) | (sew1H[2] ? checkVec_2_4 : 96'h0);
  wire [31:0]        notReadSelect = (sew1H[0] ? checkVec_0_5 : 32'h0) | (sew1H[1] ? checkVec_1_5 : 32'h0) | (sew1H[2] ? checkVec_2_5 : 32'h0);
  wire [31:0]        elementValidSelect = (sew1H[0] ? checkVec_0_6 : 32'h0) | (sew1H[1] ? checkVec_1_6 : 32'h0) | (sew1H[2] ? checkVec_2_6 : 32'h0);
  wire               readTypeRequestDeq;
  wire               waiteStageEnqReady;
  wire               readWaitQueue_deq_valid;
  assign readWaitQueue_deq_valid = ~_readWaitQueue_fifo_empty;
  wire [6:0]         readWaitQueue_dataOut_executeGroup;
  wire [31:0]        readWaitQueue_dataOut_sourceValid;
  wire [31:0]        readWaitQueue_dataOut_replaceVs1;
  wire [31:0]        readWaitQueue_dataOut_needRead;
  wire               readWaitQueue_dataOut_last;
  wire [32:0]        readWaitQueue_dataIn_lo = {readWaitQueue_enq_bits_needRead, readWaitQueue_enq_bits_last};
  wire [38:0]        readWaitQueue_dataIn_hi_hi = {readWaitQueue_enq_bits_executeGroup, readWaitQueue_enq_bits_sourceValid};
  wire [70:0]        readWaitQueue_dataIn_hi = {readWaitQueue_dataIn_hi_hi, readWaitQueue_enq_bits_replaceVs1};
  wire [103:0]       readWaitQueue_dataIn = {readWaitQueue_dataIn_hi, readWaitQueue_dataIn_lo};
  assign readWaitQueue_dataOut_last = _readWaitQueue_fifo_data_out[0];
  assign readWaitQueue_dataOut_needRead = _readWaitQueue_fifo_data_out[32:1];
  assign readWaitQueue_dataOut_replaceVs1 = _readWaitQueue_fifo_data_out[64:33];
  assign readWaitQueue_dataOut_sourceValid = _readWaitQueue_fifo_data_out[96:65];
  assign readWaitQueue_dataOut_executeGroup = _readWaitQueue_fifo_data_out[103:97];
  wire [6:0]         readWaitQueue_deq_bits_executeGroup = readWaitQueue_dataOut_executeGroup;
  wire [31:0]        readWaitQueue_deq_bits_sourceValid = readWaitQueue_dataOut_sourceValid;
  wire [31:0]        readWaitQueue_deq_bits_replaceVs1 = readWaitQueue_dataOut_replaceVs1;
  wire [31:0]        readWaitQueue_deq_bits_needRead = readWaitQueue_dataOut_needRead;
  wire               readWaitQueue_deq_bits_last = readWaitQueue_dataOut_last;
  wire               readWaitQueue_enq_ready = ~_readWaitQueue_fifo_full;
  wire               readWaitQueue_enq_valid;
  wire               readWaitQueue_deq_ready;
  wire               _GEN_119 = lastExecuteGroupDeq | viota;
  assign exeRequestQueue_0_deq_ready = ~exeReqReg_0_valid | _GEN_119;
  assign exeRequestQueue_1_deq_ready = ~exeReqReg_1_valid | _GEN_119;
  assign exeRequestQueue_2_deq_ready = ~exeReqReg_2_valid | _GEN_119;
  assign exeRequestQueue_3_deq_ready = ~exeReqReg_3_valid | _GEN_119;
  assign exeRequestQueue_4_deq_ready = ~exeReqReg_4_valid | _GEN_119;
  assign exeRequestQueue_5_deq_ready = ~exeReqReg_5_valid | _GEN_119;
  assign exeRequestQueue_6_deq_ready = ~exeReqReg_6_valid | _GEN_119;
  assign exeRequestQueue_7_deq_ready = ~exeReqReg_7_valid | _GEN_119;
  assign exeRequestQueue_8_deq_ready = ~exeReqReg_8_valid | _GEN_119;
  assign exeRequestQueue_9_deq_ready = ~exeReqReg_9_valid | _GEN_119;
  assign exeRequestQueue_10_deq_ready = ~exeReqReg_10_valid | _GEN_119;
  assign exeRequestQueue_11_deq_ready = ~exeReqReg_11_valid | _GEN_119;
  assign exeRequestQueue_12_deq_ready = ~exeReqReg_12_valid | _GEN_119;
  assign exeRequestQueue_13_deq_ready = ~exeReqReg_13_valid | _GEN_119;
  assign exeRequestQueue_14_deq_ready = ~exeReqReg_14_valid | _GEN_119;
  assign exeRequestQueue_15_deq_ready = ~exeReqReg_15_valid | _GEN_119;
  assign exeRequestQueue_16_deq_ready = ~exeReqReg_16_valid | _GEN_119;
  assign exeRequestQueue_17_deq_ready = ~exeReqReg_17_valid | _GEN_119;
  assign exeRequestQueue_18_deq_ready = ~exeReqReg_18_valid | _GEN_119;
  assign exeRequestQueue_19_deq_ready = ~exeReqReg_19_valid | _GEN_119;
  assign exeRequestQueue_20_deq_ready = ~exeReqReg_20_valid | _GEN_119;
  assign exeRequestQueue_21_deq_ready = ~exeReqReg_21_valid | _GEN_119;
  assign exeRequestQueue_22_deq_ready = ~exeReqReg_22_valid | _GEN_119;
  assign exeRequestQueue_23_deq_ready = ~exeReqReg_23_valid | _GEN_119;
  assign exeRequestQueue_24_deq_ready = ~exeReqReg_24_valid | _GEN_119;
  assign exeRequestQueue_25_deq_ready = ~exeReqReg_25_valid | _GEN_119;
  assign exeRequestQueue_26_deq_ready = ~exeReqReg_26_valid | _GEN_119;
  assign exeRequestQueue_27_deq_ready = ~exeReqReg_27_valid | _GEN_119;
  assign exeRequestQueue_28_deq_ready = ~exeReqReg_28_valid | _GEN_119;
  assign exeRequestQueue_29_deq_ready = ~exeReqReg_29_valid | _GEN_119;
  assign exeRequestQueue_30_deq_ready = ~exeReqReg_30_valid | _GEN_119;
  assign exeRequestQueue_31_deq_ready = ~exeReqReg_31_valid | _GEN_119;
  wire               isLastExecuteGroup = executeIndex == lastExecuteIndex;
  wire               allDataValid =
    (exeReqReg_0_valid | ~(groupDataNeed[0])) & (exeReqReg_1_valid | ~(groupDataNeed[1])) & (exeReqReg_2_valid | ~(groupDataNeed[2])) & (exeReqReg_3_valid | ~(groupDataNeed[3])) & (exeReqReg_4_valid | ~(groupDataNeed[4]))
    & (exeReqReg_5_valid | ~(groupDataNeed[5])) & (exeReqReg_6_valid | ~(groupDataNeed[6])) & (exeReqReg_7_valid | ~(groupDataNeed[7])) & (exeReqReg_8_valid | ~(groupDataNeed[8])) & (exeReqReg_9_valid | ~(groupDataNeed[9]))
    & (exeReqReg_10_valid | ~(groupDataNeed[10])) & (exeReqReg_11_valid | ~(groupDataNeed[11])) & (exeReqReg_12_valid | ~(groupDataNeed[12])) & (exeReqReg_13_valid | ~(groupDataNeed[13])) & (exeReqReg_14_valid | ~(groupDataNeed[14]))
    & (exeReqReg_15_valid | ~(groupDataNeed[15])) & (exeReqReg_16_valid | ~(groupDataNeed[16])) & (exeReqReg_17_valid | ~(groupDataNeed[17])) & (exeReqReg_18_valid | ~(groupDataNeed[18])) & (exeReqReg_19_valid | ~(groupDataNeed[19]))
    & (exeReqReg_20_valid | ~(groupDataNeed[20])) & (exeReqReg_21_valid | ~(groupDataNeed[21])) & (exeReqReg_22_valid | ~(groupDataNeed[22])) & (exeReqReg_23_valid | ~(groupDataNeed[23])) & (exeReqReg_24_valid | ~(groupDataNeed[24]))
    & (exeReqReg_25_valid | ~(groupDataNeed[25])) & (exeReqReg_26_valid | ~(groupDataNeed[26])) & (exeReqReg_27_valid | ~(groupDataNeed[27])) & (exeReqReg_28_valid | ~(groupDataNeed[28])) & (exeReqReg_29_valid | ~(groupDataNeed[29]))
    & (exeReqReg_30_valid | ~(groupDataNeed[30])) & (exeReqReg_31_valid | ~(groupDataNeed[31]));
  wire               anyDataValid =
    exeReqReg_0_valid | exeReqReg_1_valid | exeReqReg_2_valid | exeReqReg_3_valid | exeReqReg_4_valid | exeReqReg_5_valid | exeReqReg_6_valid | exeReqReg_7_valid | exeReqReg_8_valid | exeReqReg_9_valid | exeReqReg_10_valid
    | exeReqReg_11_valid | exeReqReg_12_valid | exeReqReg_13_valid | exeReqReg_14_valid | exeReqReg_15_valid | exeReqReg_16_valid | exeReqReg_17_valid | exeReqReg_18_valid | exeReqReg_19_valid | exeReqReg_20_valid | exeReqReg_21_valid
    | exeReqReg_22_valid | exeReqReg_23_valid | exeReqReg_24_valid | exeReqReg_25_valid | exeReqReg_26_valid | exeReqReg_27_valid | exeReqReg_28_valid | exeReqReg_29_valid | exeReqReg_30_valid | exeReqReg_31_valid;
  wire               _GEN_120 = compress | mvRd;
  wire               readVs1Valid = (unitType[2] | _GEN_120) & ~readVS1Reg_requestSend | gatherSRead;
  wire               _GEN_121 = compress | ~gatherSRead;
  wire [4:0]         readVS1Req_vs = _GEN_121 ? instReg_vs1 : instReg_vs1 + {2'h0, gatherGrowth};
  wire               readVS1Req_offset = ~compress & gatherSRead & gatherOffset;
  wire [4:0]         readVS1Req_readLane = compress ? {1'h0, readVS1Reg_readIndex} : gatherSRead ? gatherLane : 5'h0;
  wire [1:0]         readVS1Req_dataOffset = _GEN_121 ? 2'h0 : gatherDatOffset;
  wire               selectExecuteReq_1_bits_offset = readIssueStageState_readOffset[1];
  wire               selectExecuteReq_2_bits_offset = readIssueStageState_readOffset[2];
  wire               selectExecuteReq_3_bits_offset = readIssueStageState_readOffset[3];
  wire               selectExecuteReq_4_bits_offset = readIssueStageState_readOffset[4];
  wire               selectExecuteReq_5_bits_offset = readIssueStageState_readOffset[5];
  wire               selectExecuteReq_6_bits_offset = readIssueStageState_readOffset[6];
  wire               selectExecuteReq_7_bits_offset = readIssueStageState_readOffset[7];
  wire               selectExecuteReq_8_bits_offset = readIssueStageState_readOffset[8];
  wire               selectExecuteReq_9_bits_offset = readIssueStageState_readOffset[9];
  wire               selectExecuteReq_10_bits_offset = readIssueStageState_readOffset[10];
  wire               selectExecuteReq_11_bits_offset = readIssueStageState_readOffset[11];
  wire               selectExecuteReq_12_bits_offset = readIssueStageState_readOffset[12];
  wire               selectExecuteReq_13_bits_offset = readIssueStageState_readOffset[13];
  wire               selectExecuteReq_14_bits_offset = readIssueStageState_readOffset[14];
  wire               selectExecuteReq_15_bits_offset = readIssueStageState_readOffset[15];
  wire               selectExecuteReq_16_bits_offset = readIssueStageState_readOffset[16];
  wire               selectExecuteReq_17_bits_offset = readIssueStageState_readOffset[17];
  wire               selectExecuteReq_18_bits_offset = readIssueStageState_readOffset[18];
  wire               selectExecuteReq_19_bits_offset = readIssueStageState_readOffset[19];
  wire               selectExecuteReq_20_bits_offset = readIssueStageState_readOffset[20];
  wire               selectExecuteReq_21_bits_offset = readIssueStageState_readOffset[21];
  wire               selectExecuteReq_22_bits_offset = readIssueStageState_readOffset[22];
  wire               selectExecuteReq_23_bits_offset = readIssueStageState_readOffset[23];
  wire               selectExecuteReq_24_bits_offset = readIssueStageState_readOffset[24];
  wire               selectExecuteReq_25_bits_offset = readIssueStageState_readOffset[25];
  wire               selectExecuteReq_26_bits_offset = readIssueStageState_readOffset[26];
  wire               selectExecuteReq_27_bits_offset = readIssueStageState_readOffset[27];
  wire               selectExecuteReq_28_bits_offset = readIssueStageState_readOffset[28];
  wire               selectExecuteReq_29_bits_offset = readIssueStageState_readOffset[29];
  wire               selectExecuteReq_30_bits_offset = readIssueStageState_readOffset[30];
  wire               selectExecuteReq_31_bits_offset = readIssueStageState_readOffset[31];
  wire [1:0]         selectExecuteReq_1_bits_dataOffset = readIssueStageState_readDataOffset[3:2];
  wire [1:0]         selectExecuteReq_2_bits_dataOffset = readIssueStageState_readDataOffset[5:4];
  wire [1:0]         selectExecuteReq_3_bits_dataOffset = readIssueStageState_readDataOffset[7:6];
  wire [1:0]         selectExecuteReq_4_bits_dataOffset = readIssueStageState_readDataOffset[9:8];
  wire [1:0]         selectExecuteReq_5_bits_dataOffset = readIssueStageState_readDataOffset[11:10];
  wire [1:0]         selectExecuteReq_6_bits_dataOffset = readIssueStageState_readDataOffset[13:12];
  wire [1:0]         selectExecuteReq_7_bits_dataOffset = readIssueStageState_readDataOffset[15:14];
  wire [1:0]         selectExecuteReq_8_bits_dataOffset = readIssueStageState_readDataOffset[17:16];
  wire [1:0]         selectExecuteReq_9_bits_dataOffset = readIssueStageState_readDataOffset[19:18];
  wire [1:0]         selectExecuteReq_10_bits_dataOffset = readIssueStageState_readDataOffset[21:20];
  wire [1:0]         selectExecuteReq_11_bits_dataOffset = readIssueStageState_readDataOffset[23:22];
  wire [1:0]         selectExecuteReq_12_bits_dataOffset = readIssueStageState_readDataOffset[25:24];
  wire [1:0]         selectExecuteReq_13_bits_dataOffset = readIssueStageState_readDataOffset[27:26];
  wire [1:0]         selectExecuteReq_14_bits_dataOffset = readIssueStageState_readDataOffset[29:28];
  wire [1:0]         selectExecuteReq_15_bits_dataOffset = readIssueStageState_readDataOffset[31:30];
  wire [1:0]         selectExecuteReq_16_bits_dataOffset = readIssueStageState_readDataOffset[33:32];
  wire [1:0]         selectExecuteReq_17_bits_dataOffset = readIssueStageState_readDataOffset[35:34];
  wire [1:0]         selectExecuteReq_18_bits_dataOffset = readIssueStageState_readDataOffset[37:36];
  wire [1:0]         selectExecuteReq_19_bits_dataOffset = readIssueStageState_readDataOffset[39:38];
  wire [1:0]         selectExecuteReq_20_bits_dataOffset = readIssueStageState_readDataOffset[41:40];
  wire [1:0]         selectExecuteReq_21_bits_dataOffset = readIssueStageState_readDataOffset[43:42];
  wire [1:0]         selectExecuteReq_22_bits_dataOffset = readIssueStageState_readDataOffset[45:44];
  wire [1:0]         selectExecuteReq_23_bits_dataOffset = readIssueStageState_readDataOffset[47:46];
  wire [1:0]         selectExecuteReq_24_bits_dataOffset = readIssueStageState_readDataOffset[49:48];
  wire [1:0]         selectExecuteReq_25_bits_dataOffset = readIssueStageState_readDataOffset[51:50];
  wire [1:0]         selectExecuteReq_26_bits_dataOffset = readIssueStageState_readDataOffset[53:52];
  wire [1:0]         selectExecuteReq_27_bits_dataOffset = readIssueStageState_readDataOffset[55:54];
  wire [1:0]         selectExecuteReq_28_bits_dataOffset = readIssueStageState_readDataOffset[57:56];
  wire [1:0]         selectExecuteReq_29_bits_dataOffset = readIssueStageState_readDataOffset[59:58];
  wire [1:0]         selectExecuteReq_30_bits_dataOffset = readIssueStageState_readDataOffset[61:60];
  wire [1:0]         selectExecuteReq_31_bits_dataOffset = readIssueStageState_readDataOffset[63:62];
  wire               selectExecuteReq_0_valid = readVs1Valid | readIssueStageValid & ~(readIssueStageState_groupReadState[0]) & readIssueStageState_needRead[0] & readType;
  wire [4:0]         selectExecuteReq_0_bits_vs = readVs1Valid ? readVS1Req_vs : instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_0};
  wire               selectExecuteReq_0_bits_offset = readVs1Valid ? readVS1Req_offset : readIssueStageState_readOffset[0];
  wire [4:0]         selectExecuteReq_0_bits_readLane = readVs1Valid ? readVS1Req_readLane : readIssueStageState_accessLane_0;
  wire [1:0]         selectExecuteReq_0_bits_dataOffset = readVs1Valid ? readVS1Req_dataOffset : readIssueStageState_readDataOffset[1:0];
  wire               _tokenCheck_T = _readCrossBar_input_0_ready & readCrossBar_input_0_valid;
  wire               pipeReadFire_0 = ~readVs1Valid & _tokenCheck_T;
  wire [4:0]         selectExecuteReq_1_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_1};
  wire               selectExecuteReq_1_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[1]) & readIssueStageState_needRead[1] & readType;
  wire               pipeReadFire_1 = _readCrossBar_input_1_ready & readCrossBar_input_1_valid;
  wire [4:0]         selectExecuteReq_2_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_2};
  wire               selectExecuteReq_2_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[2]) & readIssueStageState_needRead[2] & readType;
  wire               pipeReadFire_2 = _readCrossBar_input_2_ready & readCrossBar_input_2_valid;
  wire [4:0]         selectExecuteReq_3_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_3};
  wire               selectExecuteReq_3_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[3]) & readIssueStageState_needRead[3] & readType;
  wire               pipeReadFire_3 = _readCrossBar_input_3_ready & readCrossBar_input_3_valid;
  wire [4:0]         selectExecuteReq_4_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_4};
  wire               selectExecuteReq_4_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[4]) & readIssueStageState_needRead[4] & readType;
  wire               pipeReadFire_4 = _readCrossBar_input_4_ready & readCrossBar_input_4_valid;
  wire [4:0]         selectExecuteReq_5_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_5};
  wire               selectExecuteReq_5_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[5]) & readIssueStageState_needRead[5] & readType;
  wire               pipeReadFire_5 = _readCrossBar_input_5_ready & readCrossBar_input_5_valid;
  wire [4:0]         selectExecuteReq_6_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_6};
  wire               selectExecuteReq_6_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[6]) & readIssueStageState_needRead[6] & readType;
  wire               pipeReadFire_6 = _readCrossBar_input_6_ready & readCrossBar_input_6_valid;
  wire [4:0]         selectExecuteReq_7_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_7};
  wire               selectExecuteReq_7_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[7]) & readIssueStageState_needRead[7] & readType;
  wire               pipeReadFire_7 = _readCrossBar_input_7_ready & readCrossBar_input_7_valid;
  wire [4:0]         selectExecuteReq_8_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_8};
  wire               selectExecuteReq_8_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[8]) & readIssueStageState_needRead[8] & readType;
  wire               pipeReadFire_8 = _readCrossBar_input_8_ready & readCrossBar_input_8_valid;
  wire [4:0]         selectExecuteReq_9_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_9};
  wire               selectExecuteReq_9_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[9]) & readIssueStageState_needRead[9] & readType;
  wire               pipeReadFire_9 = _readCrossBar_input_9_ready & readCrossBar_input_9_valid;
  wire [4:0]         selectExecuteReq_10_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_10};
  wire               selectExecuteReq_10_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[10]) & readIssueStageState_needRead[10] & readType;
  wire               pipeReadFire_10 = _readCrossBar_input_10_ready & readCrossBar_input_10_valid;
  wire [4:0]         selectExecuteReq_11_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_11};
  wire               selectExecuteReq_11_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[11]) & readIssueStageState_needRead[11] & readType;
  wire               pipeReadFire_11 = _readCrossBar_input_11_ready & readCrossBar_input_11_valid;
  wire [4:0]         selectExecuteReq_12_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_12};
  wire               selectExecuteReq_12_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[12]) & readIssueStageState_needRead[12] & readType;
  wire               pipeReadFire_12 = _readCrossBar_input_12_ready & readCrossBar_input_12_valid;
  wire [4:0]         selectExecuteReq_13_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_13};
  wire               selectExecuteReq_13_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[13]) & readIssueStageState_needRead[13] & readType;
  wire               pipeReadFire_13 = _readCrossBar_input_13_ready & readCrossBar_input_13_valid;
  wire [4:0]         selectExecuteReq_14_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_14};
  wire               selectExecuteReq_14_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[14]) & readIssueStageState_needRead[14] & readType;
  wire               pipeReadFire_14 = _readCrossBar_input_14_ready & readCrossBar_input_14_valid;
  wire [4:0]         selectExecuteReq_15_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_15};
  wire               selectExecuteReq_15_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[15]) & readIssueStageState_needRead[15] & readType;
  wire               pipeReadFire_15 = _readCrossBar_input_15_ready & readCrossBar_input_15_valid;
  wire [4:0]         selectExecuteReq_16_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_16};
  wire               selectExecuteReq_16_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[16]) & readIssueStageState_needRead[16] & readType;
  wire               pipeReadFire_16 = _readCrossBar_input_16_ready & readCrossBar_input_16_valid;
  wire [4:0]         selectExecuteReq_17_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_17};
  wire               selectExecuteReq_17_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[17]) & readIssueStageState_needRead[17] & readType;
  wire               pipeReadFire_17 = _readCrossBar_input_17_ready & readCrossBar_input_17_valid;
  wire [4:0]         selectExecuteReq_18_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_18};
  wire               selectExecuteReq_18_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[18]) & readIssueStageState_needRead[18] & readType;
  wire               pipeReadFire_18 = _readCrossBar_input_18_ready & readCrossBar_input_18_valid;
  wire [4:0]         selectExecuteReq_19_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_19};
  wire               selectExecuteReq_19_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[19]) & readIssueStageState_needRead[19] & readType;
  wire               pipeReadFire_19 = _readCrossBar_input_19_ready & readCrossBar_input_19_valid;
  wire [4:0]         selectExecuteReq_20_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_20};
  wire               selectExecuteReq_20_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[20]) & readIssueStageState_needRead[20] & readType;
  wire               pipeReadFire_20 = _readCrossBar_input_20_ready & readCrossBar_input_20_valid;
  wire [4:0]         selectExecuteReq_21_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_21};
  wire               selectExecuteReq_21_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[21]) & readIssueStageState_needRead[21] & readType;
  wire               pipeReadFire_21 = _readCrossBar_input_21_ready & readCrossBar_input_21_valid;
  wire [4:0]         selectExecuteReq_22_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_22};
  wire               selectExecuteReq_22_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[22]) & readIssueStageState_needRead[22] & readType;
  wire               pipeReadFire_22 = _readCrossBar_input_22_ready & readCrossBar_input_22_valid;
  wire [4:0]         selectExecuteReq_23_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_23};
  wire               selectExecuteReq_23_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[23]) & readIssueStageState_needRead[23] & readType;
  wire               pipeReadFire_23 = _readCrossBar_input_23_ready & readCrossBar_input_23_valid;
  wire [4:0]         selectExecuteReq_24_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_24};
  wire               selectExecuteReq_24_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[24]) & readIssueStageState_needRead[24] & readType;
  wire               pipeReadFire_24 = _readCrossBar_input_24_ready & readCrossBar_input_24_valid;
  wire [4:0]         selectExecuteReq_25_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_25};
  wire               selectExecuteReq_25_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[25]) & readIssueStageState_needRead[25] & readType;
  wire               pipeReadFire_25 = _readCrossBar_input_25_ready & readCrossBar_input_25_valid;
  wire [4:0]         selectExecuteReq_26_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_26};
  wire               selectExecuteReq_26_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[26]) & readIssueStageState_needRead[26] & readType;
  wire               pipeReadFire_26 = _readCrossBar_input_26_ready & readCrossBar_input_26_valid;
  wire [4:0]         selectExecuteReq_27_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_27};
  wire               selectExecuteReq_27_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[27]) & readIssueStageState_needRead[27] & readType;
  wire               pipeReadFire_27 = _readCrossBar_input_27_ready & readCrossBar_input_27_valid;
  wire [4:0]         selectExecuteReq_28_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_28};
  wire               selectExecuteReq_28_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[28]) & readIssueStageState_needRead[28] & readType;
  wire               pipeReadFire_28 = _readCrossBar_input_28_ready & readCrossBar_input_28_valid;
  wire [4:0]         selectExecuteReq_29_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_29};
  wire               selectExecuteReq_29_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[29]) & readIssueStageState_needRead[29] & readType;
  wire               pipeReadFire_29 = _readCrossBar_input_29_ready & readCrossBar_input_29_valid;
  wire [4:0]         selectExecuteReq_30_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_30};
  wire               selectExecuteReq_30_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[30]) & readIssueStageState_needRead[30] & readType;
  wire               pipeReadFire_30 = _readCrossBar_input_30_ready & readCrossBar_input_30_valid;
  wire [4:0]         selectExecuteReq_31_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_31};
  wire               selectExecuteReq_31_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[31]) & readIssueStageState_needRead[31] & readType;
  wire               pipeReadFire_31 = _readCrossBar_input_31_ready & readCrossBar_input_31_valid;
  reg  [3:0]         tokenCheck_counter;
  wire [3:0]         tokenCheck_counterChange = _tokenCheck_T ? 4'h1 : 4'hF;
  wire               tokenCheck = ~(tokenCheck_counter[3]);
  assign readCrossBar_input_0_valid = selectExecuteReq_0_valid & tokenCheck;
  reg  [3:0]         tokenCheck_counter_1;
  wire [3:0]         tokenCheck_counterChange_1 = pipeReadFire_1 ? 4'h1 : 4'hF;
  wire               tokenCheck_1 = ~(tokenCheck_counter_1[3]);
  assign readCrossBar_input_1_valid = selectExecuteReq_1_valid & tokenCheck_1;
  reg  [3:0]         tokenCheck_counter_2;
  wire [3:0]         tokenCheck_counterChange_2 = pipeReadFire_2 ? 4'h1 : 4'hF;
  wire               tokenCheck_2 = ~(tokenCheck_counter_2[3]);
  assign readCrossBar_input_2_valid = selectExecuteReq_2_valid & tokenCheck_2;
  reg  [3:0]         tokenCheck_counter_3;
  wire [3:0]         tokenCheck_counterChange_3 = pipeReadFire_3 ? 4'h1 : 4'hF;
  wire               tokenCheck_3 = ~(tokenCheck_counter_3[3]);
  assign readCrossBar_input_3_valid = selectExecuteReq_3_valid & tokenCheck_3;
  reg  [3:0]         tokenCheck_counter_4;
  wire [3:0]         tokenCheck_counterChange_4 = pipeReadFire_4 ? 4'h1 : 4'hF;
  wire               tokenCheck_4 = ~(tokenCheck_counter_4[3]);
  assign readCrossBar_input_4_valid = selectExecuteReq_4_valid & tokenCheck_4;
  reg  [3:0]         tokenCheck_counter_5;
  wire [3:0]         tokenCheck_counterChange_5 = pipeReadFire_5 ? 4'h1 : 4'hF;
  wire               tokenCheck_5 = ~(tokenCheck_counter_5[3]);
  assign readCrossBar_input_5_valid = selectExecuteReq_5_valid & tokenCheck_5;
  reg  [3:0]         tokenCheck_counter_6;
  wire [3:0]         tokenCheck_counterChange_6 = pipeReadFire_6 ? 4'h1 : 4'hF;
  wire               tokenCheck_6 = ~(tokenCheck_counter_6[3]);
  assign readCrossBar_input_6_valid = selectExecuteReq_6_valid & tokenCheck_6;
  reg  [3:0]         tokenCheck_counter_7;
  wire [3:0]         tokenCheck_counterChange_7 = pipeReadFire_7 ? 4'h1 : 4'hF;
  wire               tokenCheck_7 = ~(tokenCheck_counter_7[3]);
  assign readCrossBar_input_7_valid = selectExecuteReq_7_valid & tokenCheck_7;
  reg  [3:0]         tokenCheck_counter_8;
  wire [3:0]         tokenCheck_counterChange_8 = pipeReadFire_8 ? 4'h1 : 4'hF;
  wire               tokenCheck_8 = ~(tokenCheck_counter_8[3]);
  assign readCrossBar_input_8_valid = selectExecuteReq_8_valid & tokenCheck_8;
  reg  [3:0]         tokenCheck_counter_9;
  wire [3:0]         tokenCheck_counterChange_9 = pipeReadFire_9 ? 4'h1 : 4'hF;
  wire               tokenCheck_9 = ~(tokenCheck_counter_9[3]);
  assign readCrossBar_input_9_valid = selectExecuteReq_9_valid & tokenCheck_9;
  reg  [3:0]         tokenCheck_counter_10;
  wire [3:0]         tokenCheck_counterChange_10 = pipeReadFire_10 ? 4'h1 : 4'hF;
  wire               tokenCheck_10 = ~(tokenCheck_counter_10[3]);
  assign readCrossBar_input_10_valid = selectExecuteReq_10_valid & tokenCheck_10;
  reg  [3:0]         tokenCheck_counter_11;
  wire [3:0]         tokenCheck_counterChange_11 = pipeReadFire_11 ? 4'h1 : 4'hF;
  wire               tokenCheck_11 = ~(tokenCheck_counter_11[3]);
  assign readCrossBar_input_11_valid = selectExecuteReq_11_valid & tokenCheck_11;
  reg  [3:0]         tokenCheck_counter_12;
  wire [3:0]         tokenCheck_counterChange_12 = pipeReadFire_12 ? 4'h1 : 4'hF;
  wire               tokenCheck_12 = ~(tokenCheck_counter_12[3]);
  assign readCrossBar_input_12_valid = selectExecuteReq_12_valid & tokenCheck_12;
  reg  [3:0]         tokenCheck_counter_13;
  wire [3:0]         tokenCheck_counterChange_13 = pipeReadFire_13 ? 4'h1 : 4'hF;
  wire               tokenCheck_13 = ~(tokenCheck_counter_13[3]);
  assign readCrossBar_input_13_valid = selectExecuteReq_13_valid & tokenCheck_13;
  reg  [3:0]         tokenCheck_counter_14;
  wire [3:0]         tokenCheck_counterChange_14 = pipeReadFire_14 ? 4'h1 : 4'hF;
  wire               tokenCheck_14 = ~(tokenCheck_counter_14[3]);
  assign readCrossBar_input_14_valid = selectExecuteReq_14_valid & tokenCheck_14;
  reg  [3:0]         tokenCheck_counter_15;
  wire [3:0]         tokenCheck_counterChange_15 = pipeReadFire_15 ? 4'h1 : 4'hF;
  wire               tokenCheck_15 = ~(tokenCheck_counter_15[3]);
  assign readCrossBar_input_15_valid = selectExecuteReq_15_valid & tokenCheck_15;
  reg  [3:0]         tokenCheck_counter_16;
  wire [3:0]         tokenCheck_counterChange_16 = pipeReadFire_16 ? 4'h1 : 4'hF;
  wire               tokenCheck_16 = ~(tokenCheck_counter_16[3]);
  assign readCrossBar_input_16_valid = selectExecuteReq_16_valid & tokenCheck_16;
  reg  [3:0]         tokenCheck_counter_17;
  wire [3:0]         tokenCheck_counterChange_17 = pipeReadFire_17 ? 4'h1 : 4'hF;
  wire               tokenCheck_17 = ~(tokenCheck_counter_17[3]);
  assign readCrossBar_input_17_valid = selectExecuteReq_17_valid & tokenCheck_17;
  reg  [3:0]         tokenCheck_counter_18;
  wire [3:0]         tokenCheck_counterChange_18 = pipeReadFire_18 ? 4'h1 : 4'hF;
  wire               tokenCheck_18 = ~(tokenCheck_counter_18[3]);
  assign readCrossBar_input_18_valid = selectExecuteReq_18_valid & tokenCheck_18;
  reg  [3:0]         tokenCheck_counter_19;
  wire [3:0]         tokenCheck_counterChange_19 = pipeReadFire_19 ? 4'h1 : 4'hF;
  wire               tokenCheck_19 = ~(tokenCheck_counter_19[3]);
  assign readCrossBar_input_19_valid = selectExecuteReq_19_valid & tokenCheck_19;
  reg  [3:0]         tokenCheck_counter_20;
  wire [3:0]         tokenCheck_counterChange_20 = pipeReadFire_20 ? 4'h1 : 4'hF;
  wire               tokenCheck_20 = ~(tokenCheck_counter_20[3]);
  assign readCrossBar_input_20_valid = selectExecuteReq_20_valid & tokenCheck_20;
  reg  [3:0]         tokenCheck_counter_21;
  wire [3:0]         tokenCheck_counterChange_21 = pipeReadFire_21 ? 4'h1 : 4'hF;
  wire               tokenCheck_21 = ~(tokenCheck_counter_21[3]);
  assign readCrossBar_input_21_valid = selectExecuteReq_21_valid & tokenCheck_21;
  reg  [3:0]         tokenCheck_counter_22;
  wire [3:0]         tokenCheck_counterChange_22 = pipeReadFire_22 ? 4'h1 : 4'hF;
  wire               tokenCheck_22 = ~(tokenCheck_counter_22[3]);
  assign readCrossBar_input_22_valid = selectExecuteReq_22_valid & tokenCheck_22;
  reg  [3:0]         tokenCheck_counter_23;
  wire [3:0]         tokenCheck_counterChange_23 = pipeReadFire_23 ? 4'h1 : 4'hF;
  wire               tokenCheck_23 = ~(tokenCheck_counter_23[3]);
  assign readCrossBar_input_23_valid = selectExecuteReq_23_valid & tokenCheck_23;
  reg  [3:0]         tokenCheck_counter_24;
  wire [3:0]         tokenCheck_counterChange_24 = pipeReadFire_24 ? 4'h1 : 4'hF;
  wire               tokenCheck_24 = ~(tokenCheck_counter_24[3]);
  assign readCrossBar_input_24_valid = selectExecuteReq_24_valid & tokenCheck_24;
  reg  [3:0]         tokenCheck_counter_25;
  wire [3:0]         tokenCheck_counterChange_25 = pipeReadFire_25 ? 4'h1 : 4'hF;
  wire               tokenCheck_25 = ~(tokenCheck_counter_25[3]);
  assign readCrossBar_input_25_valid = selectExecuteReq_25_valid & tokenCheck_25;
  reg  [3:0]         tokenCheck_counter_26;
  wire [3:0]         tokenCheck_counterChange_26 = pipeReadFire_26 ? 4'h1 : 4'hF;
  wire               tokenCheck_26 = ~(tokenCheck_counter_26[3]);
  assign readCrossBar_input_26_valid = selectExecuteReq_26_valid & tokenCheck_26;
  reg  [3:0]         tokenCheck_counter_27;
  wire [3:0]         tokenCheck_counterChange_27 = pipeReadFire_27 ? 4'h1 : 4'hF;
  wire               tokenCheck_27 = ~(tokenCheck_counter_27[3]);
  assign readCrossBar_input_27_valid = selectExecuteReq_27_valid & tokenCheck_27;
  reg  [3:0]         tokenCheck_counter_28;
  wire [3:0]         tokenCheck_counterChange_28 = pipeReadFire_28 ? 4'h1 : 4'hF;
  wire               tokenCheck_28 = ~(tokenCheck_counter_28[3]);
  assign readCrossBar_input_28_valid = selectExecuteReq_28_valid & tokenCheck_28;
  reg  [3:0]         tokenCheck_counter_29;
  wire [3:0]         tokenCheck_counterChange_29 = pipeReadFire_29 ? 4'h1 : 4'hF;
  wire               tokenCheck_29 = ~(tokenCheck_counter_29[3]);
  assign readCrossBar_input_29_valid = selectExecuteReq_29_valid & tokenCheck_29;
  reg  [3:0]         tokenCheck_counter_30;
  wire [3:0]         tokenCheck_counterChange_30 = pipeReadFire_30 ? 4'h1 : 4'hF;
  wire               tokenCheck_30 = ~(tokenCheck_counter_30[3]);
  assign readCrossBar_input_30_valid = selectExecuteReq_30_valid & tokenCheck_30;
  reg  [3:0]         tokenCheck_counter_31;
  wire [3:0]         tokenCheck_counterChange_31 = pipeReadFire_31 ? 4'h1 : 4'hF;
  wire               tokenCheck_31 = ~(tokenCheck_counter_31[3]);
  assign readCrossBar_input_31_valid = selectExecuteReq_31_valid & tokenCheck_31;
  wire [1:0]         readFire_lo_lo_lo_lo = {pipeReadFire_1, pipeReadFire_0};
  wire [1:0]         readFire_lo_lo_lo_hi = {pipeReadFire_3, pipeReadFire_2};
  wire [3:0]         readFire_lo_lo_lo = {readFire_lo_lo_lo_hi, readFire_lo_lo_lo_lo};
  wire [1:0]         readFire_lo_lo_hi_lo = {pipeReadFire_5, pipeReadFire_4};
  wire [1:0]         readFire_lo_lo_hi_hi = {pipeReadFire_7, pipeReadFire_6};
  wire [3:0]         readFire_lo_lo_hi = {readFire_lo_lo_hi_hi, readFire_lo_lo_hi_lo};
  wire [7:0]         readFire_lo_lo = {readFire_lo_lo_hi, readFire_lo_lo_lo};
  wire [1:0]         readFire_lo_hi_lo_lo = {pipeReadFire_9, pipeReadFire_8};
  wire [1:0]         readFire_lo_hi_lo_hi = {pipeReadFire_11, pipeReadFire_10};
  wire [3:0]         readFire_lo_hi_lo = {readFire_lo_hi_lo_hi, readFire_lo_hi_lo_lo};
  wire [1:0]         readFire_lo_hi_hi_lo = {pipeReadFire_13, pipeReadFire_12};
  wire [1:0]         readFire_lo_hi_hi_hi = {pipeReadFire_15, pipeReadFire_14};
  wire [3:0]         readFire_lo_hi_hi = {readFire_lo_hi_hi_hi, readFire_lo_hi_hi_lo};
  wire [7:0]         readFire_lo_hi = {readFire_lo_hi_hi, readFire_lo_hi_lo};
  wire [15:0]        readFire_lo = {readFire_lo_hi, readFire_lo_lo};
  wire [1:0]         readFire_hi_lo_lo_lo = {pipeReadFire_17, pipeReadFire_16};
  wire [1:0]         readFire_hi_lo_lo_hi = {pipeReadFire_19, pipeReadFire_18};
  wire [3:0]         readFire_hi_lo_lo = {readFire_hi_lo_lo_hi, readFire_hi_lo_lo_lo};
  wire [1:0]         readFire_hi_lo_hi_lo = {pipeReadFire_21, pipeReadFire_20};
  wire [1:0]         readFire_hi_lo_hi_hi = {pipeReadFire_23, pipeReadFire_22};
  wire [3:0]         readFire_hi_lo_hi = {readFire_hi_lo_hi_hi, readFire_hi_lo_hi_lo};
  wire [7:0]         readFire_hi_lo = {readFire_hi_lo_hi, readFire_hi_lo_lo};
  wire [1:0]         readFire_hi_hi_lo_lo = {pipeReadFire_25, pipeReadFire_24};
  wire [1:0]         readFire_hi_hi_lo_hi = {pipeReadFire_27, pipeReadFire_26};
  wire [3:0]         readFire_hi_hi_lo = {readFire_hi_hi_lo_hi, readFire_hi_hi_lo_lo};
  wire [1:0]         readFire_hi_hi_hi_lo = {pipeReadFire_29, pipeReadFire_28};
  wire [1:0]         readFire_hi_hi_hi_hi = {pipeReadFire_31, pipeReadFire_30};
  wire [3:0]         readFire_hi_hi_hi = {readFire_hi_hi_hi_hi, readFire_hi_hi_hi_lo};
  wire [7:0]         readFire_hi_hi = {readFire_hi_hi_hi, readFire_hi_hi_lo};
  wire [15:0]        readFire_hi = {readFire_hi_hi, readFire_hi_lo};
  wire [31:0]        readFire = {readFire_hi, readFire_lo};
  wire               anyReadFire = |readFire;
  wire [31:0]        readStateUpdate = readFire | readIssueStageState_groupReadState;
  wire               groupReadFinish = readStateUpdate == readIssueStageState_needRead;
  assign readTypeRequestDeq = anyReadFire & groupReadFinish | readIssueStageValid & readIssueStageState_needRead == 32'h0;
  assign readWaitQueue_enq_valid = readTypeRequestDeq;
  wire [31:0]        compressUnitResultQueue_enq_bits_ffoOutput;
  wire               compressUnitResultQueue_enq_bits_compressValid;
  wire [32:0]        compressUnitResultQueue_dataIn_lo = {compressUnitResultQueue_enq_bits_ffoOutput, compressUnitResultQueue_enq_bits_compressValid};
  wire [1023:0]      compressUnitResultQueue_enq_bits_data;
  wire [127:0]       compressUnitResultQueue_enq_bits_mask;
  wire [1151:0]      compressUnitResultQueue_dataIn_hi_hi = {compressUnitResultQueue_enq_bits_data, compressUnitResultQueue_enq_bits_mask};
  wire [4:0]         compressUnitResultQueue_enq_bits_groupCounter;
  wire [1156:0]      compressUnitResultQueue_dataIn_hi = {compressUnitResultQueue_dataIn_hi_hi, compressUnitResultQueue_enq_bits_groupCounter};
  wire [1189:0]      compressUnitResultQueue_dataIn = {compressUnitResultQueue_dataIn_hi, compressUnitResultQueue_dataIn_lo};
  wire               compressUnitResultQueue_dataOut_compressValid = _compressUnitResultQueue_fifo_data_out[0];
  wire [31:0]        compressUnitResultQueue_dataOut_ffoOutput = _compressUnitResultQueue_fifo_data_out[32:1];
  wire [4:0]         compressUnitResultQueue_dataOut_groupCounter = _compressUnitResultQueue_fifo_data_out[37:33];
  wire [127:0]       compressUnitResultQueue_dataOut_mask = _compressUnitResultQueue_fifo_data_out[165:38];
  wire [1023:0]      compressUnitResultQueue_dataOut_data = _compressUnitResultQueue_fifo_data_out[1189:166];
  wire               compressUnitResultQueue_enq_ready = ~_compressUnitResultQueue_fifo_full;
  wire               compressUnitResultQueue_deq_ready;
  wire               compressUnitResultQueue_enq_valid;
  wire               compressUnitResultQueue_deq_valid = ~_compressUnitResultQueue_fifo_empty | compressUnitResultQueue_enq_valid;
  wire [1023:0]      compressUnitResultQueue_deq_bits_data = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_data : compressUnitResultQueue_dataOut_data;
  wire [127:0]       compressUnitResultQueue_deq_bits_mask = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_mask : compressUnitResultQueue_dataOut_mask;
  wire [4:0]         compressUnitResultQueue_deq_bits_groupCounter = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_groupCounter : compressUnitResultQueue_dataOut_groupCounter;
  wire [31:0]        compressUnitResultQueue_deq_bits_ffoOutput = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_ffoOutput : compressUnitResultQueue_dataOut_ffoOutput;
  wire               compressUnitResultQueue_deq_bits_compressValid = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_compressValid : compressUnitResultQueue_dataOut_compressValid;
  wire               noSourceValid = noSource & counterValid & ((|instReg_vl) | mvRd & ~readVS1Reg_sendToExecution);
  wire               vs1DataValid = readVS1Reg_dataValid | ~(unitType[2] | _GEN_120);
  wire [1:0]         _GEN_122 = {_maskedWrite_in_1_ready, _maskedWrite_in_0_ready};
  wire [1:0]         executeDeqReady_lo_lo_lo_lo;
  assign executeDeqReady_lo_lo_lo_lo = _GEN_122;
  wire [1:0]         compressUnitResultQueue_deq_ready_lo_lo_lo_lo;
  assign compressUnitResultQueue_deq_ready_lo_lo_lo_lo = _GEN_122;
  wire [1:0]         _GEN_123 = {_maskedWrite_in_3_ready, _maskedWrite_in_2_ready};
  wire [1:0]         executeDeqReady_lo_lo_lo_hi;
  assign executeDeqReady_lo_lo_lo_hi = _GEN_123;
  wire [1:0]         compressUnitResultQueue_deq_ready_lo_lo_lo_hi;
  assign compressUnitResultQueue_deq_ready_lo_lo_lo_hi = _GEN_123;
  wire [3:0]         executeDeqReady_lo_lo_lo = {executeDeqReady_lo_lo_lo_hi, executeDeqReady_lo_lo_lo_lo};
  wire [1:0]         _GEN_124 = {_maskedWrite_in_5_ready, _maskedWrite_in_4_ready};
  wire [1:0]         executeDeqReady_lo_lo_hi_lo;
  assign executeDeqReady_lo_lo_hi_lo = _GEN_124;
  wire [1:0]         compressUnitResultQueue_deq_ready_lo_lo_hi_lo;
  assign compressUnitResultQueue_deq_ready_lo_lo_hi_lo = _GEN_124;
  wire [1:0]         _GEN_125 = {_maskedWrite_in_7_ready, _maskedWrite_in_6_ready};
  wire [1:0]         executeDeqReady_lo_lo_hi_hi;
  assign executeDeqReady_lo_lo_hi_hi = _GEN_125;
  wire [1:0]         compressUnitResultQueue_deq_ready_lo_lo_hi_hi;
  assign compressUnitResultQueue_deq_ready_lo_lo_hi_hi = _GEN_125;
  wire [3:0]         executeDeqReady_lo_lo_hi = {executeDeqReady_lo_lo_hi_hi, executeDeqReady_lo_lo_hi_lo};
  wire [7:0]         executeDeqReady_lo_lo = {executeDeqReady_lo_lo_hi, executeDeqReady_lo_lo_lo};
  wire [1:0]         _GEN_126 = {_maskedWrite_in_9_ready, _maskedWrite_in_8_ready};
  wire [1:0]         executeDeqReady_lo_hi_lo_lo;
  assign executeDeqReady_lo_hi_lo_lo = _GEN_126;
  wire [1:0]         compressUnitResultQueue_deq_ready_lo_hi_lo_lo;
  assign compressUnitResultQueue_deq_ready_lo_hi_lo_lo = _GEN_126;
  wire [1:0]         _GEN_127 = {_maskedWrite_in_11_ready, _maskedWrite_in_10_ready};
  wire [1:0]         executeDeqReady_lo_hi_lo_hi;
  assign executeDeqReady_lo_hi_lo_hi = _GEN_127;
  wire [1:0]         compressUnitResultQueue_deq_ready_lo_hi_lo_hi;
  assign compressUnitResultQueue_deq_ready_lo_hi_lo_hi = _GEN_127;
  wire [3:0]         executeDeqReady_lo_hi_lo = {executeDeqReady_lo_hi_lo_hi, executeDeqReady_lo_hi_lo_lo};
  wire [1:0]         _GEN_128 = {_maskedWrite_in_13_ready, _maskedWrite_in_12_ready};
  wire [1:0]         executeDeqReady_lo_hi_hi_lo;
  assign executeDeqReady_lo_hi_hi_lo = _GEN_128;
  wire [1:0]         compressUnitResultQueue_deq_ready_lo_hi_hi_lo;
  assign compressUnitResultQueue_deq_ready_lo_hi_hi_lo = _GEN_128;
  wire [1:0]         _GEN_129 = {_maskedWrite_in_15_ready, _maskedWrite_in_14_ready};
  wire [1:0]         executeDeqReady_lo_hi_hi_hi;
  assign executeDeqReady_lo_hi_hi_hi = _GEN_129;
  wire [1:0]         compressUnitResultQueue_deq_ready_lo_hi_hi_hi;
  assign compressUnitResultQueue_deq_ready_lo_hi_hi_hi = _GEN_129;
  wire [3:0]         executeDeqReady_lo_hi_hi = {executeDeqReady_lo_hi_hi_hi, executeDeqReady_lo_hi_hi_lo};
  wire [7:0]         executeDeqReady_lo_hi = {executeDeqReady_lo_hi_hi, executeDeqReady_lo_hi_lo};
  wire [15:0]        executeDeqReady_lo = {executeDeqReady_lo_hi, executeDeqReady_lo_lo};
  wire [1:0]         _GEN_130 = {_maskedWrite_in_17_ready, _maskedWrite_in_16_ready};
  wire [1:0]         executeDeqReady_hi_lo_lo_lo;
  assign executeDeqReady_hi_lo_lo_lo = _GEN_130;
  wire [1:0]         compressUnitResultQueue_deq_ready_hi_lo_lo_lo;
  assign compressUnitResultQueue_deq_ready_hi_lo_lo_lo = _GEN_130;
  wire [1:0]         _GEN_131 = {_maskedWrite_in_19_ready, _maskedWrite_in_18_ready};
  wire [1:0]         executeDeqReady_hi_lo_lo_hi;
  assign executeDeqReady_hi_lo_lo_hi = _GEN_131;
  wire [1:0]         compressUnitResultQueue_deq_ready_hi_lo_lo_hi;
  assign compressUnitResultQueue_deq_ready_hi_lo_lo_hi = _GEN_131;
  wire [3:0]         executeDeqReady_hi_lo_lo = {executeDeqReady_hi_lo_lo_hi, executeDeqReady_hi_lo_lo_lo};
  wire [1:0]         _GEN_132 = {_maskedWrite_in_21_ready, _maskedWrite_in_20_ready};
  wire [1:0]         executeDeqReady_hi_lo_hi_lo;
  assign executeDeqReady_hi_lo_hi_lo = _GEN_132;
  wire [1:0]         compressUnitResultQueue_deq_ready_hi_lo_hi_lo;
  assign compressUnitResultQueue_deq_ready_hi_lo_hi_lo = _GEN_132;
  wire [1:0]         _GEN_133 = {_maskedWrite_in_23_ready, _maskedWrite_in_22_ready};
  wire [1:0]         executeDeqReady_hi_lo_hi_hi;
  assign executeDeqReady_hi_lo_hi_hi = _GEN_133;
  wire [1:0]         compressUnitResultQueue_deq_ready_hi_lo_hi_hi;
  assign compressUnitResultQueue_deq_ready_hi_lo_hi_hi = _GEN_133;
  wire [3:0]         executeDeqReady_hi_lo_hi = {executeDeqReady_hi_lo_hi_hi, executeDeqReady_hi_lo_hi_lo};
  wire [7:0]         executeDeqReady_hi_lo = {executeDeqReady_hi_lo_hi, executeDeqReady_hi_lo_lo};
  wire [1:0]         _GEN_134 = {_maskedWrite_in_25_ready, _maskedWrite_in_24_ready};
  wire [1:0]         executeDeqReady_hi_hi_lo_lo;
  assign executeDeqReady_hi_hi_lo_lo = _GEN_134;
  wire [1:0]         compressUnitResultQueue_deq_ready_hi_hi_lo_lo;
  assign compressUnitResultQueue_deq_ready_hi_hi_lo_lo = _GEN_134;
  wire [1:0]         _GEN_135 = {_maskedWrite_in_27_ready, _maskedWrite_in_26_ready};
  wire [1:0]         executeDeqReady_hi_hi_lo_hi;
  assign executeDeqReady_hi_hi_lo_hi = _GEN_135;
  wire [1:0]         compressUnitResultQueue_deq_ready_hi_hi_lo_hi;
  assign compressUnitResultQueue_deq_ready_hi_hi_lo_hi = _GEN_135;
  wire [3:0]         executeDeqReady_hi_hi_lo = {executeDeqReady_hi_hi_lo_hi, executeDeqReady_hi_hi_lo_lo};
  wire [1:0]         _GEN_136 = {_maskedWrite_in_29_ready, _maskedWrite_in_28_ready};
  wire [1:0]         executeDeqReady_hi_hi_hi_lo;
  assign executeDeqReady_hi_hi_hi_lo = _GEN_136;
  wire [1:0]         compressUnitResultQueue_deq_ready_hi_hi_hi_lo;
  assign compressUnitResultQueue_deq_ready_hi_hi_hi_lo = _GEN_136;
  wire [1:0]         _GEN_137 = {_maskedWrite_in_31_ready, _maskedWrite_in_30_ready};
  wire [1:0]         executeDeqReady_hi_hi_hi_hi;
  assign executeDeqReady_hi_hi_hi_hi = _GEN_137;
  wire [1:0]         compressUnitResultQueue_deq_ready_hi_hi_hi_hi;
  assign compressUnitResultQueue_deq_ready_hi_hi_hi_hi = _GEN_137;
  wire [3:0]         executeDeqReady_hi_hi_hi = {executeDeqReady_hi_hi_hi_hi, executeDeqReady_hi_hi_hi_lo};
  wire [7:0]         executeDeqReady_hi_hi = {executeDeqReady_hi_hi_hi, executeDeqReady_hi_hi_lo};
  wire [15:0]        executeDeqReady_hi = {executeDeqReady_hi_hi, executeDeqReady_hi_lo};
  wire               compressUnitResultQueue_empty;
  wire               executeDeqReady = (&{executeDeqReady_hi, executeDeqReady_lo}) & compressUnitResultQueue_empty;
  wire               otherTypeRequestDeq = (noSource ? noSourceValid : allDataValid) & vs1DataValid & instVlValid & executeDeqReady;
  wire               reorderQueueAllocate;
  wire               _GEN_138 = accessCountQueue_enq_ready & reorderQueueAllocate;
  assign readIssueStageEnq = (allDataValid | _slideAddressGen_indexDeq_valid) & (readTypeRequestDeq | ~readIssueStageValid) & instVlValid & readType & _GEN_138;
  assign accessCountQueue_enq_valid = readIssueStageEnq;
  wire               executeReady;
  wire               requestStageDeq = readType ? readIssueStageEnq : otherTypeRequestDeq & executeReady;
  wire               slideAddressGen_indexDeq_ready = (readTypeRequestDeq | ~readIssueStageValid) & _GEN_138;
  wire               _GEN_139 = slideAddressGen_indexDeq_ready & _slideAddressGen_indexDeq_valid;
  wire               _GEN_140 = readIssueStageEnq & _GEN_139;
  assign accessCountEnq_0 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[22]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[26]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h0 & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h0 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h0 & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h0 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h0 & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h0 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h0 & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h0 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h0 & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h0 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h0 & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h0 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h0 & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h0 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h0 & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h0 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h0 & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h0 & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h0 & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h0 & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h0 & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h0 & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h0 & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h0 & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h0 & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h0 & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h0 & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h0 & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h0 & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h0 & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h0 & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h0 & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h0 & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_1 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[22]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[26]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h1 & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h1 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h1 & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h1 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h1 & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h1 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h1 & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h1 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h1 & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h1 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h1 & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h1 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h1 & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h1 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h1 & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h1 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h1 & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h1 & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h1 & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h1 & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h1 & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h1 & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h1 & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h1 & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h1 & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h1 & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h1 & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h1 & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h1 & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h1 & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h1 & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h1 & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h1 & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_2 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[22]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[26]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h2 & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h2 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h2 & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h2 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h2 & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h2 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h2 & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h2 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h2 & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h2 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h2 & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h2 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h2 & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h2 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h2 & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h2 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h2 & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h2 & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h2 & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h2 & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h2 & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h2 & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h2 & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h2 & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h2 & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h2 & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h2 & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h2 & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h2 & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h2 & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h2 & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h2 & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h2 & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_3 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[22]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[26]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h3 & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h3 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h3 & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h3 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h3 & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h3 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h3 & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h3 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h3 & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h3 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h3 & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h3 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h3 & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h3 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h3 & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h3 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h3 & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h3 & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h3 & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h3 & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h3 & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h3 & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h3 & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h3 & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h3 & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h3 & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h3 & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h3 & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h3 & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h3 & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h3 & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h3 & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h3 & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_4 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[22]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[26]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h4 & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h4 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h4 & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h4 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h4 & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h4 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h4 & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h4 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h4 & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h4 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h4 & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h4 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h4 & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h4 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h4 & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h4 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h4 & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h4 & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h4 & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h4 & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h4 & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h4 & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h4 & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h4 & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h4 & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h4 & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h4 & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h4 & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h4 & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h4 & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h4 & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h4 & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h4 & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_5 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[22]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[26]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h5 & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h5 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h5 & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h5 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h5 & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h5 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h5 & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h5 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h5 & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h5 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h5 & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h5 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h5 & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h5 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h5 & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h5 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h5 & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h5 & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h5 & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h5 & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h5 & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h5 & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h5 & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h5 & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h5 & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h5 & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h5 & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h5 & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h5 & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h5 & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h5 & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h5 & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h5 & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_6 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[22]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[26]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h6 & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h6 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h6 & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h6 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h6 & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h6 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h6 & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h6 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h6 & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h6 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h6 & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h6 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h6 & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h6 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h6 & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h6 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h6 & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h6 & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h6 & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h6 & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h6 & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h6 & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h6 & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h6 & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h6 & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h6 & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h6 & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h6 & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h6 & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h6 & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h6 & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h6 & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h6 & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_7 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[22]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[26]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h7 & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h7 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h7 & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h7 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h7 & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h7 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h7 & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h7 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h7 & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h7 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h7 & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h7 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h7 & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h7 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h7 & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h7 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h7 & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h7 & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h7 & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h7 & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h7 & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h7 & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h7 & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h7 & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h7 & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h7 & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h7 & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h7 & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h7 & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h7 & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h7 & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h7 & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h7 & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_8 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[22]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[26]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h8 & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h8 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h8 & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h8 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h8 & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h8 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h8 & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h8 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h8 & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h8 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h8 & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h8 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h8 & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h8 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h8 & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h8 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h8 & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h8 & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h8 & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h8 & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h8 & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h8 & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h8 & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h8 & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h8 & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h8 & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h8 & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h8 & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h8 & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h8 & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h8 & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h8 & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h8 & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_9 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[22]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[26]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h9 & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h9 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h9 & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h9 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h9 & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h9 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h9 & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h9 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h9 & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h9 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h9 & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h9 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h9 & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h9 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h9 & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h9 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h9 & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h9 & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h9 & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h9 & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h9 & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h9 & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h9 & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h9 & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h9 & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h9 & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h9 & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h9 & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h9 & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h9 & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h9 & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h9 & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h9 & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_10 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[22]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[26]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'hA & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'hA & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'hA & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'hA & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'hA & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'hA & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'hA & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'hA & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'hA & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'hA & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'hA & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'hA & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'hA & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'hA & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'hA & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'hA & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'hA & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'hA & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'hA & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'hA & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'hA & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'hA & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'hA & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'hA & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'hA & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'hA & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'hA & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'hA & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'hA & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'hA & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'hA & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'hA & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'hA & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_11 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[22]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[26]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'hB & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'hB & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'hB & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'hB & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'hB & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'hB & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'hB & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'hB & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'hB & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'hB & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'hB & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'hB & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'hB & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'hB & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'hB & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'hB & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'hB & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'hB & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'hB & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'hB & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'hB & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'hB & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'hB & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'hB & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'hB & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'hB & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'hB & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'hB & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'hB & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'hB & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'hB & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'hB & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'hB & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_12 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[22]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[26]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'hC & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'hC & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'hC & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'hC & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'hC & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'hC & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'hC & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'hC & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'hC & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'hC & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'hC & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'hC & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'hC & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'hC & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'hC & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'hC & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'hC & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'hC & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'hC & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'hC & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'hC & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'hC & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'hC & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'hC & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'hC & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'hC & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'hC & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'hC & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'hC & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'hC & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'hC & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'hC & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'hC & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_13 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[22]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[26]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'hD & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'hD & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'hD & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'hD & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'hD & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'hD & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'hD & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'hD & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'hD & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'hD & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'hD & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'hD & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'hD & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'hD & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'hD & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'hD & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'hD & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'hD & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'hD & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'hD & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'hD & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'hD & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'hD & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'hD & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'hD & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'hD & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'hD & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'hD & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'hD & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'hD & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'hD & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'hD & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'hD & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_14 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[22]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[26]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'hE & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'hE & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'hE & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'hE & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'hE & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'hE & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'hE & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'hE & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'hE & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'hE & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'hE & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'hE & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'hE & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'hE & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'hE & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'hE & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'hE & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'hE & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'hE & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'hE & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'hE & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'hE & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'hE & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'hE & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'hE & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'hE & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'hE & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'hE & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'hE & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'hE & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'hE & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'hE & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'hE & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_15 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[22]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[26]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'hF & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'hF & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'hF & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'hF & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'hF & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'hF & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'hF & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'hF & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'hF & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'hF & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'hF & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'hF & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'hF & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'hF & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'hF & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'hF & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'hF & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'hF & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'hF & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'hF & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'hF & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'hF & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'hF & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'hF & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'hF & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'hF & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'hF & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'hF & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'hF & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'hF & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'hF & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'hF & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'hF & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_16 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[22]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[26]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h10 & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h10 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h10 & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h10 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h10 & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h10 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h10 & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h10 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h10 & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h10 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h10 & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h10 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h10 & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h10 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h10 & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h10 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h10 & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h10 & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h10 & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h10 & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h10 & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h10 & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h10 & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h10 & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h10 & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h10 & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h10 & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h10 & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h10 & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h10 & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h10 & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h10 & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h10 & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_17 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[22]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[26]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h11 & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h11 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h11 & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h11 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h11 & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h11 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h11 & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h11 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h11 & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h11 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h11 & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h11 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h11 & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h11 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h11 & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h11 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h11 & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h11 & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h11 & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h11 & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h11 & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h11 & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h11 & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h11 & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h11 & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h11 & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h11 & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h11 & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h11 & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h11 & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h11 & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h11 & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h11 & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_18 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[22]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[26]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h12 & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h12 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h12 & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h12 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h12 & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h12 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h12 & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h12 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h12 & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h12 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h12 & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h12 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h12 & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h12 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h12 & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h12 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h12 & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h12 & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h12 & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h12 & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h12 & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h12 & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h12 & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h12 & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h12 & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h12 & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h12 & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h12 & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h12 & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h12 & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h12 & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h12 & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h12 & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_19 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[22]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[26]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h13 & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h13 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h13 & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h13 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h13 & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h13 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h13 & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h13 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h13 & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h13 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h13 & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h13 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h13 & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h13 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h13 & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h13 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h13 & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h13 & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h13 & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h13 & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h13 & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h13 & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h13 & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h13 & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h13 & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h13 & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h13 & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h13 & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h13 & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h13 & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h13 & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h13 & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h13 & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_20 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[22]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[26]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h14 & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h14 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h14 & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h14 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h14 & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h14 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h14 & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h14 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h14 & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h14 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h14 & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h14 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h14 & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h14 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h14 & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h14 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h14 & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h14 & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h14 & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h14 & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h14 & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h14 & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h14 & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h14 & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h14 & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h14 & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h14 & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h14 & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h14 & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h14 & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h14 & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h14 & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h14 & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_21 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[22]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[26]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h15 & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h15 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h15 & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h15 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h15 & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h15 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h15 & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h15 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h15 & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h15 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h15 & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h15 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h15 & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h15 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h15 & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h15 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h15 & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h15 & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h15 & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h15 & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h15 & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h15 & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h15 & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h15 & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h15 & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h15 & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h15 & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h15 & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h15 & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h15 & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h15 & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h15 & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h15 & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_22 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[22]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[26]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h16 & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h16 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h16 & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h16 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h16 & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h16 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h16 & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h16 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h16 & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h16 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h16 & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h16 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h16 & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h16 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h16 & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h16 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h16 & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h16 & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h16 & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h16 & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h16 & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h16 & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h16 & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h16 & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h16 & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h16 & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h16 & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h16 & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h16 & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h16 & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h16 & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h16 & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h16 & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_23 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[22]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[26]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h17 & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h17 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h17 & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h17 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h17 & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h17 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h17 & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h17 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h17 & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h17 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h17 & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h17 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h17 & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h17 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h17 & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h17 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h17 & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h17 & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h17 & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h17 & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h17 & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h17 & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h17 & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h17 & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h17 & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h17 & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h17 & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h17 & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h17 & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h17 & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h17 & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h17 & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h17 & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_24 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[22]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[26]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h18 & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h18 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h18 & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h18 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h18 & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h18 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h18 & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h18 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h18 & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h18 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h18 & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h18 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h18 & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h18 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h18 & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h18 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h18 & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h18 & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h18 & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h18 & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h18 & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h18 & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h18 & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h18 & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h18 & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h18 & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h18 & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h18 & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h18 & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h18 & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h18 & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h18 & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h18 & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_25 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[22]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[26]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h19 & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h19 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h19 & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h19 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h19 & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h19 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h19 & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h19 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h19 & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h19 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h19 & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h19 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h19 & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h19 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h19 & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h19 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h19 & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h19 & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h19 & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h19 & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h19 & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h19 & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h19 & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h19 & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h19 & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h19 & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h19 & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h19 & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h19 & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h19 & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h19 & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h19 & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h19 & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_26 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[22]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[26]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h1A & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h1A & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h1A & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h1A & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h1A & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h1A & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h1A & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h1A & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h1A & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h1A & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h1A & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h1A & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h1A & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h1A & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h1A & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h1A & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h1A & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h1A & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h1A & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h1A & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h1A & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h1A & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h1A & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h1A & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h1A & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h1A & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h1A & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h1A & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h1A & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h1A & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h1A & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h1A & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h1A & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_27 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[22]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[26]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h1B & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h1B & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h1B & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h1B & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h1B & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h1B & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h1B & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h1B & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h1B & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h1B & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h1B & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h1B & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h1B & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h1B & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h1B & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h1B & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h1B & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h1B & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h1B & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h1B & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h1B & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h1B & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h1B & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h1B & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h1B & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h1B & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h1B & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h1B & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h1B & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h1B & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h1B & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h1B & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h1B & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_28 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[22]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[26]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h1C & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h1C & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h1C & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h1C & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h1C & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h1C & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h1C & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h1C & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h1C & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h1C & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h1C & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h1C & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h1C & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h1C & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h1C & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h1C & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h1C & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h1C & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h1C & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h1C & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h1C & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h1C & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h1C & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h1C & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h1C & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h1C & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h1C & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h1C & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h1C & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h1C & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h1C & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h1C & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h1C & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_29 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[22]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[26]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h1D & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h1D & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h1D & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h1D & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h1D & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h1D & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h1D & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h1D & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h1D & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h1D & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h1D & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h1D & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h1D & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h1D & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h1D & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h1D & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h1D & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h1D & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h1D & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h1D & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h1D & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h1D & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h1D & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h1D & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h1D & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h1D & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h1D & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h1D & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h1D & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h1D & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h1D & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h1D & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h1D & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_30 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0,
                    {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0,
                        {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[14]}
                          + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_16 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_17 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_18 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_19 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_20 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_21 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_22 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[22]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_23 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0,
                  {1'h0, _slideAddressGen_indexDeq_bits_accessLane_24 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_25 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_26 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[26]}
                        + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_27 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0,
                      {1'h0, _slideAddressGen_indexDeq_bits_accessLane_28 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_29 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, _slideAddressGen_indexDeq_bits_accessLane_30 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[30]}
                            + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_31 == 5'h1E & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, accessLaneSelect[4:0] == 5'h1E & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[9:5] == 5'h1E & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, accessLaneSelect[14:10] == 5'h1E & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[19:15] == 5'h1E & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, accessLaneSelect[24:20] == 5'h1E & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[29:25] == 5'h1E & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, accessLaneSelect[34:30] == 5'h1E & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[39:35] == 5'h1E & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, accessLaneSelect[44:40] == 5'h1E & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[49:45] == 5'h1E & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, accessLaneSelect[54:50] == 5'h1E & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[59:55] == 5'h1E & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, accessLaneSelect[64:60] == 5'h1E & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[69:65] == 5'h1E & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, accessLaneSelect[74:70] == 5'h1E & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[79:75] == 5'h1E & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, accessLaneSelect[84:80] == 5'h1E & ~(notReadSelect[16])} + {1'h0, accessLaneSelect[89:85] == 5'h1E & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, accessLaneSelect[94:90] == 5'h1E & ~(notReadSelect[18])} + {1'h0, accessLaneSelect[99:95] == 5'h1E & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[104:100] == 5'h1E & ~(notReadSelect[20])} + {1'h0, accessLaneSelect[109:105] == 5'h1E & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, accessLaneSelect[114:110] == 5'h1E & ~(notReadSelect[22])} + {1'h0, accessLaneSelect[119:115] == 5'h1E & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, accessLaneSelect[124:120] == 5'h1E & ~(notReadSelect[24])} + {1'h0, accessLaneSelect[129:125] == 5'h1E & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, accessLaneSelect[134:130] == 5'h1E & ~(notReadSelect[26])} + {1'h0, accessLaneSelect[139:135] == 5'h1E & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, accessLaneSelect[144:140] == 5'h1E & ~(notReadSelect[28])} + {1'h0, accessLaneSelect[149:145] == 5'h1E & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, accessLaneSelect[154:150] == 5'h1E & ~(notReadSelect[30])} + {1'h0, accessLaneSelect[159:155] == 5'h1E & ~(notReadSelect[31])}}}}};
  assign accessCountEnq_31 =
    _GEN_140
      ? {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_0) & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_1) & _slideAddressGen_indexDeq_bits_needRead[1]}}
             + {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_2) & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_3) & _slideAddressGen_indexDeq_bits_needRead[3]}}}
            + {1'h0,
               {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_4) & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_5) & _slideAddressGen_indexDeq_bits_needRead[5]}}
                 + {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_6) & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_7) & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_8) & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_9) & _slideAddressGen_indexDeq_bits_needRead[9]}}
                 + {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_10) & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_11) & _slideAddressGen_indexDeq_bits_needRead[11]}}}
                + {1'h0,
                   {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_12) & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_13) & _slideAddressGen_indexDeq_bits_needRead[13]}}
                     + {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_14) & _slideAddressGen_indexDeq_bits_needRead[14]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_15) & _slideAddressGen_indexDeq_bits_needRead[15]}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_16) & _slideAddressGen_indexDeq_bits_needRead[16]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_17) & _slideAddressGen_indexDeq_bits_needRead[17]}}
               + {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_18) & _slideAddressGen_indexDeq_bits_needRead[18]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_19) & _slideAddressGen_indexDeq_bits_needRead[19]}}}
              + {1'h0,
                 {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_20) & _slideAddressGen_indexDeq_bits_needRead[20]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_21) & _slideAddressGen_indexDeq_bits_needRead[21]}}
                   + {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_22) & _slideAddressGen_indexDeq_bits_needRead[22]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_23) & _slideAddressGen_indexDeq_bits_needRead[23]}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_24) & _slideAddressGen_indexDeq_bits_needRead[24]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_25) & _slideAddressGen_indexDeq_bits_needRead[25]}}
                   + {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_26) & _slideAddressGen_indexDeq_bits_needRead[26]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_27) & _slideAddressGen_indexDeq_bits_needRead[27]}}}
                  + {1'h0,
                     {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_28) & _slideAddressGen_indexDeq_bits_needRead[28]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_29) & _slideAddressGen_indexDeq_bits_needRead[29]}}
                       + {1'h0,
                          {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_30) & _slideAddressGen_indexDeq_bits_needRead[30]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_31) & _slideAddressGen_indexDeq_bits_needRead[31]}}}}}
      : {1'h0,
         {1'h0,
          {1'h0,
           {1'h0, {1'h0, (&(accessLaneSelect[4:0])) & ~(notReadSelect[0])} + {1'h0, (&(accessLaneSelect[9:5])) & ~(notReadSelect[1])}}
             + {1'h0, {1'h0, (&(accessLaneSelect[14:10])) & ~(notReadSelect[2])} + {1'h0, (&(accessLaneSelect[19:15])) & ~(notReadSelect[3])}}}
            + {1'h0,
               {1'h0, {1'h0, (&(accessLaneSelect[24:20])) & ~(notReadSelect[4])} + {1'h0, (&(accessLaneSelect[29:25])) & ~(notReadSelect[5])}}
                 + {1'h0, {1'h0, (&(accessLaneSelect[34:30])) & ~(notReadSelect[6])} + {1'h0, (&(accessLaneSelect[39:35])) & ~(notReadSelect[7])}}}}
           + {1'h0,
              {1'h0,
               {1'h0, {1'h0, (&(accessLaneSelect[44:40])) & ~(notReadSelect[8])} + {1'h0, (&(accessLaneSelect[49:45])) & ~(notReadSelect[9])}}
                 + {1'h0, {1'h0, (&(accessLaneSelect[54:50])) & ~(notReadSelect[10])} + {1'h0, (&(accessLaneSelect[59:55])) & ~(notReadSelect[11])}}}
                + {1'h0,
                   {1'h0, {1'h0, (&(accessLaneSelect[64:60])) & ~(notReadSelect[12])} + {1'h0, (&(accessLaneSelect[69:65])) & ~(notReadSelect[13])}}
                     + {1'h0, {1'h0, (&(accessLaneSelect[74:70])) & ~(notReadSelect[14])} + {1'h0, (&(accessLaneSelect[79:75])) & ~(notReadSelect[15])}}}}}
        + {1'h0,
           {1'h0,
            {1'h0,
             {1'h0, {1'h0, (&(accessLaneSelect[84:80])) & ~(notReadSelect[16])} + {1'h0, (&(accessLaneSelect[89:85])) & ~(notReadSelect[17])}}
               + {1'h0, {1'h0, (&(accessLaneSelect[94:90])) & ~(notReadSelect[18])} + {1'h0, (&(accessLaneSelect[99:95])) & ~(notReadSelect[19])}}}
              + {1'h0,
                 {1'h0, {1'h0, (&(accessLaneSelect[104:100])) & ~(notReadSelect[20])} + {1'h0, (&(accessLaneSelect[109:105])) & ~(notReadSelect[21])}}
                   + {1'h0, {1'h0, (&(accessLaneSelect[114:110])) & ~(notReadSelect[22])} + {1'h0, (&(accessLaneSelect[119:115])) & ~(notReadSelect[23])}}}}
             + {1'h0,
                {1'h0,
                 {1'h0, {1'h0, (&(accessLaneSelect[124:120])) & ~(notReadSelect[24])} + {1'h0, (&(accessLaneSelect[129:125])) & ~(notReadSelect[25])}}
                   + {1'h0, {1'h0, (&(accessLaneSelect[134:130])) & ~(notReadSelect[26])} + {1'h0, (&(accessLaneSelect[139:135])) & ~(notReadSelect[27])}}}
                  + {1'h0,
                     {1'h0, {1'h0, (&(accessLaneSelect[144:140])) & ~(notReadSelect[28])} + {1'h0, (&(accessLaneSelect[149:145])) & ~(notReadSelect[29])}}
                       + {1'h0, {1'h0, (&(accessLaneSelect[154:150])) & ~(notReadSelect[30])} + {1'h0, (&(accessLaneSelect[159:155])) & ~(notReadSelect[31])}}}}};
  assign lastExecuteGroupDeq = requestStageDeq & isLastExecuteGroup;
  wire [31:0]        readMessageQueue_deq_bits_readSource;
  wire               deqAllocate;
  wire               reorderQueueVec_0_deq_valid;
  assign reorderQueueVec_0_deq_valid = ~_reorderQueueVec_fifo_empty;
  wire [31:0]        reorderQueueVec_dataOut_data;
  wire [31:0]        reorderQueueVec_dataOut_write1H;
  wire [31:0]        dataAfterReorderCheck_0 = reorderQueueVec_0_deq_bits_data;
  wire [31:0]        reorderQueueVec_0_enq_bits_data;
  wire [31:0]        reorderQueueVec_0_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn = {reorderQueueVec_0_enq_bits_data, reorderQueueVec_0_enq_bits_write1H};
  assign reorderQueueVec_dataOut_write1H = _reorderQueueVec_fifo_data_out[31:0];
  assign reorderQueueVec_dataOut_data = _reorderQueueVec_fifo_data_out[63:32];
  assign reorderQueueVec_0_deq_bits_data = reorderQueueVec_dataOut_data;
  wire [31:0]        reorderQueueVec_0_deq_bits_write1H = reorderQueueVec_dataOut_write1H;
  wire               reorderQueueVec_0_enq_ready = ~_reorderQueueVec_fifo_full;
  wire               reorderQueueVec_0_deq_ready;
  wire [31:0]        readMessageQueue_1_deq_bits_readSource;
  wire               deqAllocate_1;
  wire               reorderQueueVec_1_deq_valid;
  assign reorderQueueVec_1_deq_valid = ~_reorderQueueVec_fifo_1_empty;
  wire [31:0]        reorderQueueVec_dataOut_1_data;
  wire [31:0]        reorderQueueVec_dataOut_1_write1H;
  wire [31:0]        dataAfterReorderCheck_1 = reorderQueueVec_1_deq_bits_data;
  wire [31:0]        reorderQueueVec_1_enq_bits_data;
  wire [31:0]        reorderQueueVec_1_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_1 = {reorderQueueVec_1_enq_bits_data, reorderQueueVec_1_enq_bits_write1H};
  assign reorderQueueVec_dataOut_1_write1H = _reorderQueueVec_fifo_1_data_out[31:0];
  assign reorderQueueVec_dataOut_1_data = _reorderQueueVec_fifo_1_data_out[63:32];
  assign reorderQueueVec_1_deq_bits_data = reorderQueueVec_dataOut_1_data;
  wire [31:0]        reorderQueueVec_1_deq_bits_write1H = reorderQueueVec_dataOut_1_write1H;
  wire               reorderQueueVec_1_enq_ready = ~_reorderQueueVec_fifo_1_full;
  wire               reorderQueueVec_1_deq_ready;
  wire [31:0]        readMessageQueue_2_deq_bits_readSource;
  wire               deqAllocate_2;
  wire               reorderQueueVec_2_deq_valid;
  assign reorderQueueVec_2_deq_valid = ~_reorderQueueVec_fifo_2_empty;
  wire [31:0]        reorderQueueVec_dataOut_2_data;
  wire [31:0]        reorderQueueVec_dataOut_2_write1H;
  wire [31:0]        dataAfterReorderCheck_2 = reorderQueueVec_2_deq_bits_data;
  wire [31:0]        reorderQueueVec_2_enq_bits_data;
  wire [31:0]        reorderQueueVec_2_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_2 = {reorderQueueVec_2_enq_bits_data, reorderQueueVec_2_enq_bits_write1H};
  assign reorderQueueVec_dataOut_2_write1H = _reorderQueueVec_fifo_2_data_out[31:0];
  assign reorderQueueVec_dataOut_2_data = _reorderQueueVec_fifo_2_data_out[63:32];
  assign reorderQueueVec_2_deq_bits_data = reorderQueueVec_dataOut_2_data;
  wire [31:0]        reorderQueueVec_2_deq_bits_write1H = reorderQueueVec_dataOut_2_write1H;
  wire               reorderQueueVec_2_enq_ready = ~_reorderQueueVec_fifo_2_full;
  wire               reorderQueueVec_2_deq_ready;
  wire [31:0]        readMessageQueue_3_deq_bits_readSource;
  wire               deqAllocate_3;
  wire               reorderQueueVec_3_deq_valid;
  assign reorderQueueVec_3_deq_valid = ~_reorderQueueVec_fifo_3_empty;
  wire [31:0]        reorderQueueVec_dataOut_3_data;
  wire [31:0]        reorderQueueVec_dataOut_3_write1H;
  wire [31:0]        dataAfterReorderCheck_3 = reorderQueueVec_3_deq_bits_data;
  wire [31:0]        reorderQueueVec_3_enq_bits_data;
  wire [31:0]        reorderQueueVec_3_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_3 = {reorderQueueVec_3_enq_bits_data, reorderQueueVec_3_enq_bits_write1H};
  assign reorderQueueVec_dataOut_3_write1H = _reorderQueueVec_fifo_3_data_out[31:0];
  assign reorderQueueVec_dataOut_3_data = _reorderQueueVec_fifo_3_data_out[63:32];
  assign reorderQueueVec_3_deq_bits_data = reorderQueueVec_dataOut_3_data;
  wire [31:0]        reorderQueueVec_3_deq_bits_write1H = reorderQueueVec_dataOut_3_write1H;
  wire               reorderQueueVec_3_enq_ready = ~_reorderQueueVec_fifo_3_full;
  wire               reorderQueueVec_3_deq_ready;
  wire [31:0]        readMessageQueue_4_deq_bits_readSource;
  wire               deqAllocate_4;
  wire               reorderQueueVec_4_deq_valid;
  assign reorderQueueVec_4_deq_valid = ~_reorderQueueVec_fifo_4_empty;
  wire [31:0]        reorderQueueVec_dataOut_4_data;
  wire [31:0]        reorderQueueVec_dataOut_4_write1H;
  wire [31:0]        dataAfterReorderCheck_4 = reorderQueueVec_4_deq_bits_data;
  wire [31:0]        reorderQueueVec_4_enq_bits_data;
  wire [31:0]        reorderQueueVec_4_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_4 = {reorderQueueVec_4_enq_bits_data, reorderQueueVec_4_enq_bits_write1H};
  assign reorderQueueVec_dataOut_4_write1H = _reorderQueueVec_fifo_4_data_out[31:0];
  assign reorderQueueVec_dataOut_4_data = _reorderQueueVec_fifo_4_data_out[63:32];
  assign reorderQueueVec_4_deq_bits_data = reorderQueueVec_dataOut_4_data;
  wire [31:0]        reorderQueueVec_4_deq_bits_write1H = reorderQueueVec_dataOut_4_write1H;
  wire               reorderQueueVec_4_enq_ready = ~_reorderQueueVec_fifo_4_full;
  wire               reorderQueueVec_4_deq_ready;
  wire [31:0]        readMessageQueue_5_deq_bits_readSource;
  wire               deqAllocate_5;
  wire               reorderQueueVec_5_deq_valid;
  assign reorderQueueVec_5_deq_valid = ~_reorderQueueVec_fifo_5_empty;
  wire [31:0]        reorderQueueVec_dataOut_5_data;
  wire [31:0]        reorderQueueVec_dataOut_5_write1H;
  wire [31:0]        dataAfterReorderCheck_5 = reorderQueueVec_5_deq_bits_data;
  wire [31:0]        reorderQueueVec_5_enq_bits_data;
  wire [31:0]        reorderQueueVec_5_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_5 = {reorderQueueVec_5_enq_bits_data, reorderQueueVec_5_enq_bits_write1H};
  assign reorderQueueVec_dataOut_5_write1H = _reorderQueueVec_fifo_5_data_out[31:0];
  assign reorderQueueVec_dataOut_5_data = _reorderQueueVec_fifo_5_data_out[63:32];
  assign reorderQueueVec_5_deq_bits_data = reorderQueueVec_dataOut_5_data;
  wire [31:0]        reorderQueueVec_5_deq_bits_write1H = reorderQueueVec_dataOut_5_write1H;
  wire               reorderQueueVec_5_enq_ready = ~_reorderQueueVec_fifo_5_full;
  wire               reorderQueueVec_5_deq_ready;
  wire [31:0]        readMessageQueue_6_deq_bits_readSource;
  wire               deqAllocate_6;
  wire               reorderQueueVec_6_deq_valid;
  assign reorderQueueVec_6_deq_valid = ~_reorderQueueVec_fifo_6_empty;
  wire [31:0]        reorderQueueVec_dataOut_6_data;
  wire [31:0]        reorderQueueVec_dataOut_6_write1H;
  wire [31:0]        dataAfterReorderCheck_6 = reorderQueueVec_6_deq_bits_data;
  wire [31:0]        reorderQueueVec_6_enq_bits_data;
  wire [31:0]        reorderQueueVec_6_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_6 = {reorderQueueVec_6_enq_bits_data, reorderQueueVec_6_enq_bits_write1H};
  assign reorderQueueVec_dataOut_6_write1H = _reorderQueueVec_fifo_6_data_out[31:0];
  assign reorderQueueVec_dataOut_6_data = _reorderQueueVec_fifo_6_data_out[63:32];
  assign reorderQueueVec_6_deq_bits_data = reorderQueueVec_dataOut_6_data;
  wire [31:0]        reorderQueueVec_6_deq_bits_write1H = reorderQueueVec_dataOut_6_write1H;
  wire               reorderQueueVec_6_enq_ready = ~_reorderQueueVec_fifo_6_full;
  wire               reorderQueueVec_6_deq_ready;
  wire [31:0]        readMessageQueue_7_deq_bits_readSource;
  wire               deqAllocate_7;
  wire               reorderQueueVec_7_deq_valid;
  assign reorderQueueVec_7_deq_valid = ~_reorderQueueVec_fifo_7_empty;
  wire [31:0]        reorderQueueVec_dataOut_7_data;
  wire [31:0]        reorderQueueVec_dataOut_7_write1H;
  wire [31:0]        dataAfterReorderCheck_7 = reorderQueueVec_7_deq_bits_data;
  wire [31:0]        reorderQueueVec_7_enq_bits_data;
  wire [31:0]        reorderQueueVec_7_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_7 = {reorderQueueVec_7_enq_bits_data, reorderQueueVec_7_enq_bits_write1H};
  assign reorderQueueVec_dataOut_7_write1H = _reorderQueueVec_fifo_7_data_out[31:0];
  assign reorderQueueVec_dataOut_7_data = _reorderQueueVec_fifo_7_data_out[63:32];
  assign reorderQueueVec_7_deq_bits_data = reorderQueueVec_dataOut_7_data;
  wire [31:0]        reorderQueueVec_7_deq_bits_write1H = reorderQueueVec_dataOut_7_write1H;
  wire               reorderQueueVec_7_enq_ready = ~_reorderQueueVec_fifo_7_full;
  wire               reorderQueueVec_7_deq_ready;
  wire [31:0]        readMessageQueue_8_deq_bits_readSource;
  wire               deqAllocate_8;
  wire               reorderQueueVec_8_deq_valid;
  assign reorderQueueVec_8_deq_valid = ~_reorderQueueVec_fifo_8_empty;
  wire [31:0]        reorderQueueVec_dataOut_8_data;
  wire [31:0]        reorderQueueVec_dataOut_8_write1H;
  wire [31:0]        dataAfterReorderCheck_8 = reorderQueueVec_8_deq_bits_data;
  wire [31:0]        reorderQueueVec_8_enq_bits_data;
  wire [31:0]        reorderQueueVec_8_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_8 = {reorderQueueVec_8_enq_bits_data, reorderQueueVec_8_enq_bits_write1H};
  assign reorderQueueVec_dataOut_8_write1H = _reorderQueueVec_fifo_8_data_out[31:0];
  assign reorderQueueVec_dataOut_8_data = _reorderQueueVec_fifo_8_data_out[63:32];
  assign reorderQueueVec_8_deq_bits_data = reorderQueueVec_dataOut_8_data;
  wire [31:0]        reorderQueueVec_8_deq_bits_write1H = reorderQueueVec_dataOut_8_write1H;
  wire               reorderQueueVec_8_enq_ready = ~_reorderQueueVec_fifo_8_full;
  wire               reorderQueueVec_8_deq_ready;
  wire [31:0]        readMessageQueue_9_deq_bits_readSource;
  wire               deqAllocate_9;
  wire               reorderQueueVec_9_deq_valid;
  assign reorderQueueVec_9_deq_valid = ~_reorderQueueVec_fifo_9_empty;
  wire [31:0]        reorderQueueVec_dataOut_9_data;
  wire [31:0]        reorderQueueVec_dataOut_9_write1H;
  wire [31:0]        dataAfterReorderCheck_9 = reorderQueueVec_9_deq_bits_data;
  wire [31:0]        reorderQueueVec_9_enq_bits_data;
  wire [31:0]        reorderQueueVec_9_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_9 = {reorderQueueVec_9_enq_bits_data, reorderQueueVec_9_enq_bits_write1H};
  assign reorderQueueVec_dataOut_9_write1H = _reorderQueueVec_fifo_9_data_out[31:0];
  assign reorderQueueVec_dataOut_9_data = _reorderQueueVec_fifo_9_data_out[63:32];
  assign reorderQueueVec_9_deq_bits_data = reorderQueueVec_dataOut_9_data;
  wire [31:0]        reorderQueueVec_9_deq_bits_write1H = reorderQueueVec_dataOut_9_write1H;
  wire               reorderQueueVec_9_enq_ready = ~_reorderQueueVec_fifo_9_full;
  wire               reorderQueueVec_9_deq_ready;
  wire [31:0]        readMessageQueue_10_deq_bits_readSource;
  wire               deqAllocate_10;
  wire               reorderQueueVec_10_deq_valid;
  assign reorderQueueVec_10_deq_valid = ~_reorderQueueVec_fifo_10_empty;
  wire [31:0]        reorderQueueVec_dataOut_10_data;
  wire [31:0]        reorderQueueVec_dataOut_10_write1H;
  wire [31:0]        dataAfterReorderCheck_10 = reorderQueueVec_10_deq_bits_data;
  wire [31:0]        reorderQueueVec_10_enq_bits_data;
  wire [31:0]        reorderQueueVec_10_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_10 = {reorderQueueVec_10_enq_bits_data, reorderQueueVec_10_enq_bits_write1H};
  assign reorderQueueVec_dataOut_10_write1H = _reorderQueueVec_fifo_10_data_out[31:0];
  assign reorderQueueVec_dataOut_10_data = _reorderQueueVec_fifo_10_data_out[63:32];
  assign reorderQueueVec_10_deq_bits_data = reorderQueueVec_dataOut_10_data;
  wire [31:0]        reorderQueueVec_10_deq_bits_write1H = reorderQueueVec_dataOut_10_write1H;
  wire               reorderQueueVec_10_enq_ready = ~_reorderQueueVec_fifo_10_full;
  wire               reorderQueueVec_10_deq_ready;
  wire [31:0]        readMessageQueue_11_deq_bits_readSource;
  wire               deqAllocate_11;
  wire               reorderQueueVec_11_deq_valid;
  assign reorderQueueVec_11_deq_valid = ~_reorderQueueVec_fifo_11_empty;
  wire [31:0]        reorderQueueVec_dataOut_11_data;
  wire [31:0]        reorderQueueVec_dataOut_11_write1H;
  wire [31:0]        dataAfterReorderCheck_11 = reorderQueueVec_11_deq_bits_data;
  wire [31:0]        reorderQueueVec_11_enq_bits_data;
  wire [31:0]        reorderQueueVec_11_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_11 = {reorderQueueVec_11_enq_bits_data, reorderQueueVec_11_enq_bits_write1H};
  assign reorderQueueVec_dataOut_11_write1H = _reorderQueueVec_fifo_11_data_out[31:0];
  assign reorderQueueVec_dataOut_11_data = _reorderQueueVec_fifo_11_data_out[63:32];
  assign reorderQueueVec_11_deq_bits_data = reorderQueueVec_dataOut_11_data;
  wire [31:0]        reorderQueueVec_11_deq_bits_write1H = reorderQueueVec_dataOut_11_write1H;
  wire               reorderQueueVec_11_enq_ready = ~_reorderQueueVec_fifo_11_full;
  wire               reorderQueueVec_11_deq_ready;
  wire [31:0]        readMessageQueue_12_deq_bits_readSource;
  wire               deqAllocate_12;
  wire               reorderQueueVec_12_deq_valid;
  assign reorderQueueVec_12_deq_valid = ~_reorderQueueVec_fifo_12_empty;
  wire [31:0]        reorderQueueVec_dataOut_12_data;
  wire [31:0]        reorderQueueVec_dataOut_12_write1H;
  wire [31:0]        dataAfterReorderCheck_12 = reorderQueueVec_12_deq_bits_data;
  wire [31:0]        reorderQueueVec_12_enq_bits_data;
  wire [31:0]        reorderQueueVec_12_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_12 = {reorderQueueVec_12_enq_bits_data, reorderQueueVec_12_enq_bits_write1H};
  assign reorderQueueVec_dataOut_12_write1H = _reorderQueueVec_fifo_12_data_out[31:0];
  assign reorderQueueVec_dataOut_12_data = _reorderQueueVec_fifo_12_data_out[63:32];
  assign reorderQueueVec_12_deq_bits_data = reorderQueueVec_dataOut_12_data;
  wire [31:0]        reorderQueueVec_12_deq_bits_write1H = reorderQueueVec_dataOut_12_write1H;
  wire               reorderQueueVec_12_enq_ready = ~_reorderQueueVec_fifo_12_full;
  wire               reorderQueueVec_12_deq_ready;
  wire [31:0]        readMessageQueue_13_deq_bits_readSource;
  wire               deqAllocate_13;
  wire               reorderQueueVec_13_deq_valid;
  assign reorderQueueVec_13_deq_valid = ~_reorderQueueVec_fifo_13_empty;
  wire [31:0]        reorderQueueVec_dataOut_13_data;
  wire [31:0]        reorderQueueVec_dataOut_13_write1H;
  wire [31:0]        dataAfterReorderCheck_13 = reorderQueueVec_13_deq_bits_data;
  wire [31:0]        reorderQueueVec_13_enq_bits_data;
  wire [31:0]        reorderQueueVec_13_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_13 = {reorderQueueVec_13_enq_bits_data, reorderQueueVec_13_enq_bits_write1H};
  assign reorderQueueVec_dataOut_13_write1H = _reorderQueueVec_fifo_13_data_out[31:0];
  assign reorderQueueVec_dataOut_13_data = _reorderQueueVec_fifo_13_data_out[63:32];
  assign reorderQueueVec_13_deq_bits_data = reorderQueueVec_dataOut_13_data;
  wire [31:0]        reorderQueueVec_13_deq_bits_write1H = reorderQueueVec_dataOut_13_write1H;
  wire               reorderQueueVec_13_enq_ready = ~_reorderQueueVec_fifo_13_full;
  wire               reorderQueueVec_13_deq_ready;
  wire [31:0]        readMessageQueue_14_deq_bits_readSource;
  wire               deqAllocate_14;
  wire               reorderQueueVec_14_deq_valid;
  assign reorderQueueVec_14_deq_valid = ~_reorderQueueVec_fifo_14_empty;
  wire [31:0]        reorderQueueVec_dataOut_14_data;
  wire [31:0]        reorderQueueVec_dataOut_14_write1H;
  wire [31:0]        dataAfterReorderCheck_14 = reorderQueueVec_14_deq_bits_data;
  wire [31:0]        reorderQueueVec_14_enq_bits_data;
  wire [31:0]        reorderQueueVec_14_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_14 = {reorderQueueVec_14_enq_bits_data, reorderQueueVec_14_enq_bits_write1H};
  assign reorderQueueVec_dataOut_14_write1H = _reorderQueueVec_fifo_14_data_out[31:0];
  assign reorderQueueVec_dataOut_14_data = _reorderQueueVec_fifo_14_data_out[63:32];
  assign reorderQueueVec_14_deq_bits_data = reorderQueueVec_dataOut_14_data;
  wire [31:0]        reorderQueueVec_14_deq_bits_write1H = reorderQueueVec_dataOut_14_write1H;
  wire               reorderQueueVec_14_enq_ready = ~_reorderQueueVec_fifo_14_full;
  wire               reorderQueueVec_14_deq_ready;
  wire [31:0]        readMessageQueue_15_deq_bits_readSource;
  wire               deqAllocate_15;
  wire               reorderQueueVec_15_deq_valid;
  assign reorderQueueVec_15_deq_valid = ~_reorderQueueVec_fifo_15_empty;
  wire [31:0]        reorderQueueVec_dataOut_15_data;
  wire [31:0]        reorderQueueVec_dataOut_15_write1H;
  wire [31:0]        dataAfterReorderCheck_15 = reorderQueueVec_15_deq_bits_data;
  wire [31:0]        reorderQueueVec_15_enq_bits_data;
  wire [31:0]        reorderQueueVec_15_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_15 = {reorderQueueVec_15_enq_bits_data, reorderQueueVec_15_enq_bits_write1H};
  assign reorderQueueVec_dataOut_15_write1H = _reorderQueueVec_fifo_15_data_out[31:0];
  assign reorderQueueVec_dataOut_15_data = _reorderQueueVec_fifo_15_data_out[63:32];
  assign reorderQueueVec_15_deq_bits_data = reorderQueueVec_dataOut_15_data;
  wire [31:0]        reorderQueueVec_15_deq_bits_write1H = reorderQueueVec_dataOut_15_write1H;
  wire               reorderQueueVec_15_enq_ready = ~_reorderQueueVec_fifo_15_full;
  wire               reorderQueueVec_15_deq_ready;
  wire [31:0]        readMessageQueue_16_deq_bits_readSource;
  wire               deqAllocate_16;
  wire               reorderQueueVec_16_deq_valid;
  assign reorderQueueVec_16_deq_valid = ~_reorderQueueVec_fifo_16_empty;
  wire [31:0]        reorderQueueVec_dataOut_16_data;
  wire [31:0]        reorderQueueVec_dataOut_16_write1H;
  wire [31:0]        dataAfterReorderCheck_16 = reorderQueueVec_16_deq_bits_data;
  wire [31:0]        reorderQueueVec_16_enq_bits_data;
  wire [31:0]        reorderQueueVec_16_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_16 = {reorderQueueVec_16_enq_bits_data, reorderQueueVec_16_enq_bits_write1H};
  assign reorderQueueVec_dataOut_16_write1H = _reorderQueueVec_fifo_16_data_out[31:0];
  assign reorderQueueVec_dataOut_16_data = _reorderQueueVec_fifo_16_data_out[63:32];
  assign reorderQueueVec_16_deq_bits_data = reorderQueueVec_dataOut_16_data;
  wire [31:0]        reorderQueueVec_16_deq_bits_write1H = reorderQueueVec_dataOut_16_write1H;
  wire               reorderQueueVec_16_enq_ready = ~_reorderQueueVec_fifo_16_full;
  wire               reorderQueueVec_16_deq_ready;
  wire [31:0]        readMessageQueue_17_deq_bits_readSource;
  wire               deqAllocate_17;
  wire               reorderQueueVec_17_deq_valid;
  assign reorderQueueVec_17_deq_valid = ~_reorderQueueVec_fifo_17_empty;
  wire [31:0]        reorderQueueVec_dataOut_17_data;
  wire [31:0]        reorderQueueVec_dataOut_17_write1H;
  wire [31:0]        dataAfterReorderCheck_17 = reorderQueueVec_17_deq_bits_data;
  wire [31:0]        reorderQueueVec_17_enq_bits_data;
  wire [31:0]        reorderQueueVec_17_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_17 = {reorderQueueVec_17_enq_bits_data, reorderQueueVec_17_enq_bits_write1H};
  assign reorderQueueVec_dataOut_17_write1H = _reorderQueueVec_fifo_17_data_out[31:0];
  assign reorderQueueVec_dataOut_17_data = _reorderQueueVec_fifo_17_data_out[63:32];
  assign reorderQueueVec_17_deq_bits_data = reorderQueueVec_dataOut_17_data;
  wire [31:0]        reorderQueueVec_17_deq_bits_write1H = reorderQueueVec_dataOut_17_write1H;
  wire               reorderQueueVec_17_enq_ready = ~_reorderQueueVec_fifo_17_full;
  wire               reorderQueueVec_17_deq_ready;
  wire [31:0]        readMessageQueue_18_deq_bits_readSource;
  wire               deqAllocate_18;
  wire               reorderQueueVec_18_deq_valid;
  assign reorderQueueVec_18_deq_valid = ~_reorderQueueVec_fifo_18_empty;
  wire [31:0]        reorderQueueVec_dataOut_18_data;
  wire [31:0]        reorderQueueVec_dataOut_18_write1H;
  wire [31:0]        dataAfterReorderCheck_18 = reorderQueueVec_18_deq_bits_data;
  wire [31:0]        reorderQueueVec_18_enq_bits_data;
  wire [31:0]        reorderQueueVec_18_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_18 = {reorderQueueVec_18_enq_bits_data, reorderQueueVec_18_enq_bits_write1H};
  assign reorderQueueVec_dataOut_18_write1H = _reorderQueueVec_fifo_18_data_out[31:0];
  assign reorderQueueVec_dataOut_18_data = _reorderQueueVec_fifo_18_data_out[63:32];
  assign reorderQueueVec_18_deq_bits_data = reorderQueueVec_dataOut_18_data;
  wire [31:0]        reorderQueueVec_18_deq_bits_write1H = reorderQueueVec_dataOut_18_write1H;
  wire               reorderQueueVec_18_enq_ready = ~_reorderQueueVec_fifo_18_full;
  wire               reorderQueueVec_18_deq_ready;
  wire [31:0]        readMessageQueue_19_deq_bits_readSource;
  wire               deqAllocate_19;
  wire               reorderQueueVec_19_deq_valid;
  assign reorderQueueVec_19_deq_valid = ~_reorderQueueVec_fifo_19_empty;
  wire [31:0]        reorderQueueVec_dataOut_19_data;
  wire [31:0]        reorderQueueVec_dataOut_19_write1H;
  wire [31:0]        dataAfterReorderCheck_19 = reorderQueueVec_19_deq_bits_data;
  wire [31:0]        reorderQueueVec_19_enq_bits_data;
  wire [31:0]        reorderQueueVec_19_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_19 = {reorderQueueVec_19_enq_bits_data, reorderQueueVec_19_enq_bits_write1H};
  assign reorderQueueVec_dataOut_19_write1H = _reorderQueueVec_fifo_19_data_out[31:0];
  assign reorderQueueVec_dataOut_19_data = _reorderQueueVec_fifo_19_data_out[63:32];
  assign reorderQueueVec_19_deq_bits_data = reorderQueueVec_dataOut_19_data;
  wire [31:0]        reorderQueueVec_19_deq_bits_write1H = reorderQueueVec_dataOut_19_write1H;
  wire               reorderQueueVec_19_enq_ready = ~_reorderQueueVec_fifo_19_full;
  wire               reorderQueueVec_19_deq_ready;
  wire [31:0]        readMessageQueue_20_deq_bits_readSource;
  wire               deqAllocate_20;
  wire               reorderQueueVec_20_deq_valid;
  assign reorderQueueVec_20_deq_valid = ~_reorderQueueVec_fifo_20_empty;
  wire [31:0]        reorderQueueVec_dataOut_20_data;
  wire [31:0]        reorderQueueVec_dataOut_20_write1H;
  wire [31:0]        dataAfterReorderCheck_20 = reorderQueueVec_20_deq_bits_data;
  wire [31:0]        reorderQueueVec_20_enq_bits_data;
  wire [31:0]        reorderQueueVec_20_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_20 = {reorderQueueVec_20_enq_bits_data, reorderQueueVec_20_enq_bits_write1H};
  assign reorderQueueVec_dataOut_20_write1H = _reorderQueueVec_fifo_20_data_out[31:0];
  assign reorderQueueVec_dataOut_20_data = _reorderQueueVec_fifo_20_data_out[63:32];
  assign reorderQueueVec_20_deq_bits_data = reorderQueueVec_dataOut_20_data;
  wire [31:0]        reorderQueueVec_20_deq_bits_write1H = reorderQueueVec_dataOut_20_write1H;
  wire               reorderQueueVec_20_enq_ready = ~_reorderQueueVec_fifo_20_full;
  wire               reorderQueueVec_20_deq_ready;
  wire [31:0]        readMessageQueue_21_deq_bits_readSource;
  wire               deqAllocate_21;
  wire               reorderQueueVec_21_deq_valid;
  assign reorderQueueVec_21_deq_valid = ~_reorderQueueVec_fifo_21_empty;
  wire [31:0]        reorderQueueVec_dataOut_21_data;
  wire [31:0]        reorderQueueVec_dataOut_21_write1H;
  wire [31:0]        dataAfterReorderCheck_21 = reorderQueueVec_21_deq_bits_data;
  wire [31:0]        reorderQueueVec_21_enq_bits_data;
  wire [31:0]        reorderQueueVec_21_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_21 = {reorderQueueVec_21_enq_bits_data, reorderQueueVec_21_enq_bits_write1H};
  assign reorderQueueVec_dataOut_21_write1H = _reorderQueueVec_fifo_21_data_out[31:0];
  assign reorderQueueVec_dataOut_21_data = _reorderQueueVec_fifo_21_data_out[63:32];
  assign reorderQueueVec_21_deq_bits_data = reorderQueueVec_dataOut_21_data;
  wire [31:0]        reorderQueueVec_21_deq_bits_write1H = reorderQueueVec_dataOut_21_write1H;
  wire               reorderQueueVec_21_enq_ready = ~_reorderQueueVec_fifo_21_full;
  wire               reorderQueueVec_21_deq_ready;
  wire [31:0]        readMessageQueue_22_deq_bits_readSource;
  wire               deqAllocate_22;
  wire               reorderQueueVec_22_deq_valid;
  assign reorderQueueVec_22_deq_valid = ~_reorderQueueVec_fifo_22_empty;
  wire [31:0]        reorderQueueVec_dataOut_22_data;
  wire [31:0]        reorderQueueVec_dataOut_22_write1H;
  wire [31:0]        dataAfterReorderCheck_22 = reorderQueueVec_22_deq_bits_data;
  wire [31:0]        reorderQueueVec_22_enq_bits_data;
  wire [31:0]        reorderQueueVec_22_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_22 = {reorderQueueVec_22_enq_bits_data, reorderQueueVec_22_enq_bits_write1H};
  assign reorderQueueVec_dataOut_22_write1H = _reorderQueueVec_fifo_22_data_out[31:0];
  assign reorderQueueVec_dataOut_22_data = _reorderQueueVec_fifo_22_data_out[63:32];
  assign reorderQueueVec_22_deq_bits_data = reorderQueueVec_dataOut_22_data;
  wire [31:0]        reorderQueueVec_22_deq_bits_write1H = reorderQueueVec_dataOut_22_write1H;
  wire               reorderQueueVec_22_enq_ready = ~_reorderQueueVec_fifo_22_full;
  wire               reorderQueueVec_22_deq_ready;
  wire [31:0]        readMessageQueue_23_deq_bits_readSource;
  wire               deqAllocate_23;
  wire               reorderQueueVec_23_deq_valid;
  assign reorderQueueVec_23_deq_valid = ~_reorderQueueVec_fifo_23_empty;
  wire [31:0]        reorderQueueVec_dataOut_23_data;
  wire [31:0]        reorderQueueVec_dataOut_23_write1H;
  wire [31:0]        dataAfterReorderCheck_23 = reorderQueueVec_23_deq_bits_data;
  wire [31:0]        reorderQueueVec_23_enq_bits_data;
  wire [31:0]        reorderQueueVec_23_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_23 = {reorderQueueVec_23_enq_bits_data, reorderQueueVec_23_enq_bits_write1H};
  assign reorderQueueVec_dataOut_23_write1H = _reorderQueueVec_fifo_23_data_out[31:0];
  assign reorderQueueVec_dataOut_23_data = _reorderQueueVec_fifo_23_data_out[63:32];
  assign reorderQueueVec_23_deq_bits_data = reorderQueueVec_dataOut_23_data;
  wire [31:0]        reorderQueueVec_23_deq_bits_write1H = reorderQueueVec_dataOut_23_write1H;
  wire               reorderQueueVec_23_enq_ready = ~_reorderQueueVec_fifo_23_full;
  wire               reorderQueueVec_23_deq_ready;
  wire [31:0]        readMessageQueue_24_deq_bits_readSource;
  wire               deqAllocate_24;
  wire               reorderQueueVec_24_deq_valid;
  assign reorderQueueVec_24_deq_valid = ~_reorderQueueVec_fifo_24_empty;
  wire [31:0]        reorderQueueVec_dataOut_24_data;
  wire [31:0]        reorderQueueVec_dataOut_24_write1H;
  wire [31:0]        dataAfterReorderCheck_24 = reorderQueueVec_24_deq_bits_data;
  wire [31:0]        reorderQueueVec_24_enq_bits_data;
  wire [31:0]        reorderQueueVec_24_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_24 = {reorderQueueVec_24_enq_bits_data, reorderQueueVec_24_enq_bits_write1H};
  assign reorderQueueVec_dataOut_24_write1H = _reorderQueueVec_fifo_24_data_out[31:0];
  assign reorderQueueVec_dataOut_24_data = _reorderQueueVec_fifo_24_data_out[63:32];
  assign reorderQueueVec_24_deq_bits_data = reorderQueueVec_dataOut_24_data;
  wire [31:0]        reorderQueueVec_24_deq_bits_write1H = reorderQueueVec_dataOut_24_write1H;
  wire               reorderQueueVec_24_enq_ready = ~_reorderQueueVec_fifo_24_full;
  wire               reorderQueueVec_24_deq_ready;
  wire [31:0]        readMessageQueue_25_deq_bits_readSource;
  wire               deqAllocate_25;
  wire               reorderQueueVec_25_deq_valid;
  assign reorderQueueVec_25_deq_valid = ~_reorderQueueVec_fifo_25_empty;
  wire [31:0]        reorderQueueVec_dataOut_25_data;
  wire [31:0]        reorderQueueVec_dataOut_25_write1H;
  wire [31:0]        dataAfterReorderCheck_25 = reorderQueueVec_25_deq_bits_data;
  wire [31:0]        reorderQueueVec_25_enq_bits_data;
  wire [31:0]        reorderQueueVec_25_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_25 = {reorderQueueVec_25_enq_bits_data, reorderQueueVec_25_enq_bits_write1H};
  assign reorderQueueVec_dataOut_25_write1H = _reorderQueueVec_fifo_25_data_out[31:0];
  assign reorderQueueVec_dataOut_25_data = _reorderQueueVec_fifo_25_data_out[63:32];
  assign reorderQueueVec_25_deq_bits_data = reorderQueueVec_dataOut_25_data;
  wire [31:0]        reorderQueueVec_25_deq_bits_write1H = reorderQueueVec_dataOut_25_write1H;
  wire               reorderQueueVec_25_enq_ready = ~_reorderQueueVec_fifo_25_full;
  wire               reorderQueueVec_25_deq_ready;
  wire [31:0]        readMessageQueue_26_deq_bits_readSource;
  wire               deqAllocate_26;
  wire               reorderQueueVec_26_deq_valid;
  assign reorderQueueVec_26_deq_valid = ~_reorderQueueVec_fifo_26_empty;
  wire [31:0]        reorderQueueVec_dataOut_26_data;
  wire [31:0]        reorderQueueVec_dataOut_26_write1H;
  wire [31:0]        dataAfterReorderCheck_26 = reorderQueueVec_26_deq_bits_data;
  wire [31:0]        reorderQueueVec_26_enq_bits_data;
  wire [31:0]        reorderQueueVec_26_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_26 = {reorderQueueVec_26_enq_bits_data, reorderQueueVec_26_enq_bits_write1H};
  assign reorderQueueVec_dataOut_26_write1H = _reorderQueueVec_fifo_26_data_out[31:0];
  assign reorderQueueVec_dataOut_26_data = _reorderQueueVec_fifo_26_data_out[63:32];
  assign reorderQueueVec_26_deq_bits_data = reorderQueueVec_dataOut_26_data;
  wire [31:0]        reorderQueueVec_26_deq_bits_write1H = reorderQueueVec_dataOut_26_write1H;
  wire               reorderQueueVec_26_enq_ready = ~_reorderQueueVec_fifo_26_full;
  wire               reorderQueueVec_26_deq_ready;
  wire [31:0]        readMessageQueue_27_deq_bits_readSource;
  wire               deqAllocate_27;
  wire               reorderQueueVec_27_deq_valid;
  assign reorderQueueVec_27_deq_valid = ~_reorderQueueVec_fifo_27_empty;
  wire [31:0]        reorderQueueVec_dataOut_27_data;
  wire [31:0]        reorderQueueVec_dataOut_27_write1H;
  wire [31:0]        dataAfterReorderCheck_27 = reorderQueueVec_27_deq_bits_data;
  wire [31:0]        reorderQueueVec_27_enq_bits_data;
  wire [31:0]        reorderQueueVec_27_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_27 = {reorderQueueVec_27_enq_bits_data, reorderQueueVec_27_enq_bits_write1H};
  assign reorderQueueVec_dataOut_27_write1H = _reorderQueueVec_fifo_27_data_out[31:0];
  assign reorderQueueVec_dataOut_27_data = _reorderQueueVec_fifo_27_data_out[63:32];
  assign reorderQueueVec_27_deq_bits_data = reorderQueueVec_dataOut_27_data;
  wire [31:0]        reorderQueueVec_27_deq_bits_write1H = reorderQueueVec_dataOut_27_write1H;
  wire               reorderQueueVec_27_enq_ready = ~_reorderQueueVec_fifo_27_full;
  wire               reorderQueueVec_27_deq_ready;
  wire [31:0]        readMessageQueue_28_deq_bits_readSource;
  wire               deqAllocate_28;
  wire               reorderQueueVec_28_deq_valid;
  assign reorderQueueVec_28_deq_valid = ~_reorderQueueVec_fifo_28_empty;
  wire [31:0]        reorderQueueVec_dataOut_28_data;
  wire [31:0]        reorderQueueVec_dataOut_28_write1H;
  wire [31:0]        dataAfterReorderCheck_28 = reorderQueueVec_28_deq_bits_data;
  wire [31:0]        reorderQueueVec_28_enq_bits_data;
  wire [31:0]        reorderQueueVec_28_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_28 = {reorderQueueVec_28_enq_bits_data, reorderQueueVec_28_enq_bits_write1H};
  assign reorderQueueVec_dataOut_28_write1H = _reorderQueueVec_fifo_28_data_out[31:0];
  assign reorderQueueVec_dataOut_28_data = _reorderQueueVec_fifo_28_data_out[63:32];
  assign reorderQueueVec_28_deq_bits_data = reorderQueueVec_dataOut_28_data;
  wire [31:0]        reorderQueueVec_28_deq_bits_write1H = reorderQueueVec_dataOut_28_write1H;
  wire               reorderQueueVec_28_enq_ready = ~_reorderQueueVec_fifo_28_full;
  wire               reorderQueueVec_28_deq_ready;
  wire [31:0]        readMessageQueue_29_deq_bits_readSource;
  wire               deqAllocate_29;
  wire               reorderQueueVec_29_deq_valid;
  assign reorderQueueVec_29_deq_valid = ~_reorderQueueVec_fifo_29_empty;
  wire [31:0]        reorderQueueVec_dataOut_29_data;
  wire [31:0]        reorderQueueVec_dataOut_29_write1H;
  wire [31:0]        dataAfterReorderCheck_29 = reorderQueueVec_29_deq_bits_data;
  wire [31:0]        reorderQueueVec_29_enq_bits_data;
  wire [31:0]        reorderQueueVec_29_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_29 = {reorderQueueVec_29_enq_bits_data, reorderQueueVec_29_enq_bits_write1H};
  assign reorderQueueVec_dataOut_29_write1H = _reorderQueueVec_fifo_29_data_out[31:0];
  assign reorderQueueVec_dataOut_29_data = _reorderQueueVec_fifo_29_data_out[63:32];
  assign reorderQueueVec_29_deq_bits_data = reorderQueueVec_dataOut_29_data;
  wire [31:0]        reorderQueueVec_29_deq_bits_write1H = reorderQueueVec_dataOut_29_write1H;
  wire               reorderQueueVec_29_enq_ready = ~_reorderQueueVec_fifo_29_full;
  wire               reorderQueueVec_29_deq_ready;
  wire [31:0]        readMessageQueue_30_deq_bits_readSource;
  wire               deqAllocate_30;
  wire               reorderQueueVec_30_deq_valid;
  assign reorderQueueVec_30_deq_valid = ~_reorderQueueVec_fifo_30_empty;
  wire [31:0]        reorderQueueVec_dataOut_30_data;
  wire [31:0]        reorderQueueVec_dataOut_30_write1H;
  wire [31:0]        dataAfterReorderCheck_30 = reorderQueueVec_30_deq_bits_data;
  wire [31:0]        reorderQueueVec_30_enq_bits_data;
  wire [31:0]        reorderQueueVec_30_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_30 = {reorderQueueVec_30_enq_bits_data, reorderQueueVec_30_enq_bits_write1H};
  assign reorderQueueVec_dataOut_30_write1H = _reorderQueueVec_fifo_30_data_out[31:0];
  assign reorderQueueVec_dataOut_30_data = _reorderQueueVec_fifo_30_data_out[63:32];
  assign reorderQueueVec_30_deq_bits_data = reorderQueueVec_dataOut_30_data;
  wire [31:0]        reorderQueueVec_30_deq_bits_write1H = reorderQueueVec_dataOut_30_write1H;
  wire               reorderQueueVec_30_enq_ready = ~_reorderQueueVec_fifo_30_full;
  wire               reorderQueueVec_30_deq_ready;
  wire [31:0]        readMessageQueue_31_deq_bits_readSource;
  wire               deqAllocate_31;
  wire               reorderQueueVec_31_deq_valid;
  assign reorderQueueVec_31_deq_valid = ~_reorderQueueVec_fifo_31_empty;
  wire [31:0]        reorderQueueVec_dataOut_31_data;
  wire [31:0]        reorderQueueVec_dataOut_31_write1H;
  wire [31:0]        dataAfterReorderCheck_31 = reorderQueueVec_31_deq_bits_data;
  wire [31:0]        reorderQueueVec_31_enq_bits_data;
  wire [31:0]        reorderQueueVec_31_enq_bits_write1H;
  wire [63:0]        reorderQueueVec_dataIn_31 = {reorderQueueVec_31_enq_bits_data, reorderQueueVec_31_enq_bits_write1H};
  assign reorderQueueVec_dataOut_31_write1H = _reorderQueueVec_fifo_31_data_out[31:0];
  assign reorderQueueVec_dataOut_31_data = _reorderQueueVec_fifo_31_data_out[63:32];
  assign reorderQueueVec_31_deq_bits_data = reorderQueueVec_dataOut_31_data;
  wire [31:0]        reorderQueueVec_31_deq_bits_write1H = reorderQueueVec_dataOut_31_write1H;
  wire               reorderQueueVec_31_enq_ready = ~_reorderQueueVec_fifo_31_full;
  wire               reorderQueueVec_31_deq_ready;
  reg  [6:0]         reorderQueueAllocate_counter;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate;
  wire               _write1HPipe_0_T = reorderQueueVec_0_deq_ready & reorderQueueVec_0_deq_valid;
  wire               reorderQueueAllocate_release = _write1HPipe_0_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate = readIssueStageEnq ? accessCountEnq_0 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate = reorderQueueAllocate_counter + {1'h0, reorderQueueAllocate_allocate} - {6'h0, reorderQueueAllocate_release};
  reg  [6:0]         reorderQueueAllocate_counter_1;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_1;
  wire               _write1HPipe_1_T = reorderQueueVec_1_deq_ready & reorderQueueVec_1_deq_valid;
  wire               reorderQueueAllocate_release_1 = _write1HPipe_1_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_1 = readIssueStageEnq ? accessCountEnq_1 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_1 = reorderQueueAllocate_counter_1 + {1'h0, reorderQueueAllocate_allocate_1} - {6'h0, reorderQueueAllocate_release_1};
  reg  [6:0]         reorderQueueAllocate_counter_2;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_2;
  wire               _write1HPipe_2_T = reorderQueueVec_2_deq_ready & reorderQueueVec_2_deq_valid;
  wire               reorderQueueAllocate_release_2 = _write1HPipe_2_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_2 = readIssueStageEnq ? accessCountEnq_2 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_2 = reorderQueueAllocate_counter_2 + {1'h0, reorderQueueAllocate_allocate_2} - {6'h0, reorderQueueAllocate_release_2};
  reg  [6:0]         reorderQueueAllocate_counter_3;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_3;
  wire               _write1HPipe_3_T = reorderQueueVec_3_deq_ready & reorderQueueVec_3_deq_valid;
  wire               reorderQueueAllocate_release_3 = _write1HPipe_3_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_3 = readIssueStageEnq ? accessCountEnq_3 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_3 = reorderQueueAllocate_counter_3 + {1'h0, reorderQueueAllocate_allocate_3} - {6'h0, reorderQueueAllocate_release_3};
  reg  [6:0]         reorderQueueAllocate_counter_4;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_4;
  wire               _write1HPipe_4_T = reorderQueueVec_4_deq_ready & reorderQueueVec_4_deq_valid;
  wire               reorderQueueAllocate_release_4 = _write1HPipe_4_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_4 = readIssueStageEnq ? accessCountEnq_4 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_4 = reorderQueueAllocate_counter_4 + {1'h0, reorderQueueAllocate_allocate_4} - {6'h0, reorderQueueAllocate_release_4};
  reg  [6:0]         reorderQueueAllocate_counter_5;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_5;
  wire               _write1HPipe_5_T = reorderQueueVec_5_deq_ready & reorderQueueVec_5_deq_valid;
  wire               reorderQueueAllocate_release_5 = _write1HPipe_5_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_5 = readIssueStageEnq ? accessCountEnq_5 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_5 = reorderQueueAllocate_counter_5 + {1'h0, reorderQueueAllocate_allocate_5} - {6'h0, reorderQueueAllocate_release_5};
  reg  [6:0]         reorderQueueAllocate_counter_6;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_6;
  wire               _write1HPipe_6_T = reorderQueueVec_6_deq_ready & reorderQueueVec_6_deq_valid;
  wire               reorderQueueAllocate_release_6 = _write1HPipe_6_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_6 = readIssueStageEnq ? accessCountEnq_6 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_6 = reorderQueueAllocate_counter_6 + {1'h0, reorderQueueAllocate_allocate_6} - {6'h0, reorderQueueAllocate_release_6};
  reg  [6:0]         reorderQueueAllocate_counter_7;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_7;
  wire               _write1HPipe_7_T = reorderQueueVec_7_deq_ready & reorderQueueVec_7_deq_valid;
  wire               reorderQueueAllocate_release_7 = _write1HPipe_7_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_7 = readIssueStageEnq ? accessCountEnq_7 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_7 = reorderQueueAllocate_counter_7 + {1'h0, reorderQueueAllocate_allocate_7} - {6'h0, reorderQueueAllocate_release_7};
  reg  [6:0]         reorderQueueAllocate_counter_8;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_8;
  wire               _write1HPipe_8_T = reorderQueueVec_8_deq_ready & reorderQueueVec_8_deq_valid;
  wire               reorderQueueAllocate_release_8 = _write1HPipe_8_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_8 = readIssueStageEnq ? accessCountEnq_8 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_8 = reorderQueueAllocate_counter_8 + {1'h0, reorderQueueAllocate_allocate_8} - {6'h0, reorderQueueAllocate_release_8};
  reg  [6:0]         reorderQueueAllocate_counter_9;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_9;
  wire               _write1HPipe_9_T = reorderQueueVec_9_deq_ready & reorderQueueVec_9_deq_valid;
  wire               reorderQueueAllocate_release_9 = _write1HPipe_9_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_9 = readIssueStageEnq ? accessCountEnq_9 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_9 = reorderQueueAllocate_counter_9 + {1'h0, reorderQueueAllocate_allocate_9} - {6'h0, reorderQueueAllocate_release_9};
  reg  [6:0]         reorderQueueAllocate_counter_10;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_10;
  wire               _write1HPipe_10_T = reorderQueueVec_10_deq_ready & reorderQueueVec_10_deq_valid;
  wire               reorderQueueAllocate_release_10 = _write1HPipe_10_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_10 = readIssueStageEnq ? accessCountEnq_10 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_10 = reorderQueueAllocate_counter_10 + {1'h0, reorderQueueAllocate_allocate_10} - {6'h0, reorderQueueAllocate_release_10};
  reg  [6:0]         reorderQueueAllocate_counter_11;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_11;
  wire               _write1HPipe_11_T = reorderQueueVec_11_deq_ready & reorderQueueVec_11_deq_valid;
  wire               reorderQueueAllocate_release_11 = _write1HPipe_11_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_11 = readIssueStageEnq ? accessCountEnq_11 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_11 = reorderQueueAllocate_counter_11 + {1'h0, reorderQueueAllocate_allocate_11} - {6'h0, reorderQueueAllocate_release_11};
  reg  [6:0]         reorderQueueAllocate_counter_12;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_12;
  wire               _write1HPipe_12_T = reorderQueueVec_12_deq_ready & reorderQueueVec_12_deq_valid;
  wire               reorderQueueAllocate_release_12 = _write1HPipe_12_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_12 = readIssueStageEnq ? accessCountEnq_12 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_12 = reorderQueueAllocate_counter_12 + {1'h0, reorderQueueAllocate_allocate_12} - {6'h0, reorderQueueAllocate_release_12};
  reg  [6:0]         reorderQueueAllocate_counter_13;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_13;
  wire               _write1HPipe_13_T = reorderQueueVec_13_deq_ready & reorderQueueVec_13_deq_valid;
  wire               reorderQueueAllocate_release_13 = _write1HPipe_13_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_13 = readIssueStageEnq ? accessCountEnq_13 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_13 = reorderQueueAllocate_counter_13 + {1'h0, reorderQueueAllocate_allocate_13} - {6'h0, reorderQueueAllocate_release_13};
  reg  [6:0]         reorderQueueAllocate_counter_14;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_14;
  wire               _write1HPipe_14_T = reorderQueueVec_14_deq_ready & reorderQueueVec_14_deq_valid;
  wire               reorderQueueAllocate_release_14 = _write1HPipe_14_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_14 = readIssueStageEnq ? accessCountEnq_14 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_14 = reorderQueueAllocate_counter_14 + {1'h0, reorderQueueAllocate_allocate_14} - {6'h0, reorderQueueAllocate_release_14};
  reg  [6:0]         reorderQueueAllocate_counter_15;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_15;
  wire               _write1HPipe_15_T = reorderQueueVec_15_deq_ready & reorderQueueVec_15_deq_valid;
  wire               reorderQueueAllocate_release_15 = _write1HPipe_15_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_15 = readIssueStageEnq ? accessCountEnq_15 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_15 = reorderQueueAllocate_counter_15 + {1'h0, reorderQueueAllocate_allocate_15} - {6'h0, reorderQueueAllocate_release_15};
  reg  [6:0]         reorderQueueAllocate_counter_16;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_16;
  wire               _write1HPipe_16_T = reorderQueueVec_16_deq_ready & reorderQueueVec_16_deq_valid;
  wire               reorderQueueAllocate_release_16 = _write1HPipe_16_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_16 = readIssueStageEnq ? accessCountEnq_16 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_16 = reorderQueueAllocate_counter_16 + {1'h0, reorderQueueAllocate_allocate_16} - {6'h0, reorderQueueAllocate_release_16};
  reg  [6:0]         reorderQueueAllocate_counter_17;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_17;
  wire               _write1HPipe_17_T = reorderQueueVec_17_deq_ready & reorderQueueVec_17_deq_valid;
  wire               reorderQueueAllocate_release_17 = _write1HPipe_17_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_17 = readIssueStageEnq ? accessCountEnq_17 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_17 = reorderQueueAllocate_counter_17 + {1'h0, reorderQueueAllocate_allocate_17} - {6'h0, reorderQueueAllocate_release_17};
  reg  [6:0]         reorderQueueAllocate_counter_18;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_18;
  wire               _write1HPipe_18_T = reorderQueueVec_18_deq_ready & reorderQueueVec_18_deq_valid;
  wire               reorderQueueAllocate_release_18 = _write1HPipe_18_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_18 = readIssueStageEnq ? accessCountEnq_18 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_18 = reorderQueueAllocate_counter_18 + {1'h0, reorderQueueAllocate_allocate_18} - {6'h0, reorderQueueAllocate_release_18};
  reg  [6:0]         reorderQueueAllocate_counter_19;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_19;
  wire               _write1HPipe_19_T = reorderQueueVec_19_deq_ready & reorderQueueVec_19_deq_valid;
  wire               reorderQueueAllocate_release_19 = _write1HPipe_19_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_19 = readIssueStageEnq ? accessCountEnq_19 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_19 = reorderQueueAllocate_counter_19 + {1'h0, reorderQueueAllocate_allocate_19} - {6'h0, reorderQueueAllocate_release_19};
  reg  [6:0]         reorderQueueAllocate_counter_20;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_20;
  wire               _write1HPipe_20_T = reorderQueueVec_20_deq_ready & reorderQueueVec_20_deq_valid;
  wire               reorderQueueAllocate_release_20 = _write1HPipe_20_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_20 = readIssueStageEnq ? accessCountEnq_20 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_20 = reorderQueueAllocate_counter_20 + {1'h0, reorderQueueAllocate_allocate_20} - {6'h0, reorderQueueAllocate_release_20};
  reg  [6:0]         reorderQueueAllocate_counter_21;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_21;
  wire               _write1HPipe_21_T = reorderQueueVec_21_deq_ready & reorderQueueVec_21_deq_valid;
  wire               reorderQueueAllocate_release_21 = _write1HPipe_21_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_21 = readIssueStageEnq ? accessCountEnq_21 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_21 = reorderQueueAllocate_counter_21 + {1'h0, reorderQueueAllocate_allocate_21} - {6'h0, reorderQueueAllocate_release_21};
  reg  [6:0]         reorderQueueAllocate_counter_22;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_22;
  wire               _write1HPipe_22_T = reorderQueueVec_22_deq_ready & reorderQueueVec_22_deq_valid;
  wire               reorderQueueAllocate_release_22 = _write1HPipe_22_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_22 = readIssueStageEnq ? accessCountEnq_22 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_22 = reorderQueueAllocate_counter_22 + {1'h0, reorderQueueAllocate_allocate_22} - {6'h0, reorderQueueAllocate_release_22};
  reg  [6:0]         reorderQueueAllocate_counter_23;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_23;
  wire               _write1HPipe_23_T = reorderQueueVec_23_deq_ready & reorderQueueVec_23_deq_valid;
  wire               reorderQueueAllocate_release_23 = _write1HPipe_23_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_23 = readIssueStageEnq ? accessCountEnq_23 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_23 = reorderQueueAllocate_counter_23 + {1'h0, reorderQueueAllocate_allocate_23} - {6'h0, reorderQueueAllocate_release_23};
  reg  [6:0]         reorderQueueAllocate_counter_24;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_24;
  wire               _write1HPipe_24_T = reorderQueueVec_24_deq_ready & reorderQueueVec_24_deq_valid;
  wire               reorderQueueAllocate_release_24 = _write1HPipe_24_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_24 = readIssueStageEnq ? accessCountEnq_24 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_24 = reorderQueueAllocate_counter_24 + {1'h0, reorderQueueAllocate_allocate_24} - {6'h0, reorderQueueAllocate_release_24};
  reg  [6:0]         reorderQueueAllocate_counter_25;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_25;
  wire               _write1HPipe_25_T = reorderQueueVec_25_deq_ready & reorderQueueVec_25_deq_valid;
  wire               reorderQueueAllocate_release_25 = _write1HPipe_25_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_25 = readIssueStageEnq ? accessCountEnq_25 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_25 = reorderQueueAllocate_counter_25 + {1'h0, reorderQueueAllocate_allocate_25} - {6'h0, reorderQueueAllocate_release_25};
  reg  [6:0]         reorderQueueAllocate_counter_26;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_26;
  wire               _write1HPipe_26_T = reorderQueueVec_26_deq_ready & reorderQueueVec_26_deq_valid;
  wire               reorderQueueAllocate_release_26 = _write1HPipe_26_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_26 = readIssueStageEnq ? accessCountEnq_26 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_26 = reorderQueueAllocate_counter_26 + {1'h0, reorderQueueAllocate_allocate_26} - {6'h0, reorderQueueAllocate_release_26};
  reg  [6:0]         reorderQueueAllocate_counter_27;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_27;
  wire               _write1HPipe_27_T = reorderQueueVec_27_deq_ready & reorderQueueVec_27_deq_valid;
  wire               reorderQueueAllocate_release_27 = _write1HPipe_27_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_27 = readIssueStageEnq ? accessCountEnq_27 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_27 = reorderQueueAllocate_counter_27 + {1'h0, reorderQueueAllocate_allocate_27} - {6'h0, reorderQueueAllocate_release_27};
  reg  [6:0]         reorderQueueAllocate_counter_28;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_28;
  wire               _write1HPipe_28_T = reorderQueueVec_28_deq_ready & reorderQueueVec_28_deq_valid;
  wire               reorderQueueAllocate_release_28 = _write1HPipe_28_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_28 = readIssueStageEnq ? accessCountEnq_28 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_28 = reorderQueueAllocate_counter_28 + {1'h0, reorderQueueAllocate_allocate_28} - {6'h0, reorderQueueAllocate_release_28};
  reg  [6:0]         reorderQueueAllocate_counter_29;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_29;
  wire               _write1HPipe_29_T = reorderQueueVec_29_deq_ready & reorderQueueVec_29_deq_valid;
  wire               reorderQueueAllocate_release_29 = _write1HPipe_29_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_29 = readIssueStageEnq ? accessCountEnq_29 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_29 = reorderQueueAllocate_counter_29 + {1'h0, reorderQueueAllocate_allocate_29} - {6'h0, reorderQueueAllocate_release_29};
  reg  [6:0]         reorderQueueAllocate_counter_30;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_30;
  wire               _write1HPipe_30_T = reorderQueueVec_30_deq_ready & reorderQueueVec_30_deq_valid;
  wire               reorderQueueAllocate_release_30 = _write1HPipe_30_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_30 = readIssueStageEnq ? accessCountEnq_30 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_30 = reorderQueueAllocate_counter_30 + {1'h0, reorderQueueAllocate_allocate_30} - {6'h0, reorderQueueAllocate_release_30};
  reg  [6:0]         reorderQueueAllocate_counter_31;
  reg  [6:0]         reorderQueueAllocate_counterWillUpdate_31;
  wire               _write1HPipe_31_T = reorderQueueVec_31_deq_ready & reorderQueueVec_31_deq_valid;
  wire               reorderQueueAllocate_release_31 = _write1HPipe_31_T & readValid;
  wire [5:0]         reorderQueueAllocate_allocate_31 = readIssueStageEnq ? accessCountEnq_31 : 6'h0;
  wire [6:0]         reorderQueueAllocate_counterUpdate_31 = reorderQueueAllocate_counter_31 + {1'h0, reorderQueueAllocate_allocate_31} - {6'h0, reorderQueueAllocate_release_31};
  assign reorderQueueAllocate =
    ~(reorderQueueAllocate_counterWillUpdate[6]) & ~(reorderQueueAllocate_counterWillUpdate_1[6]) & ~(reorderQueueAllocate_counterWillUpdate_2[6]) & ~(reorderQueueAllocate_counterWillUpdate_3[6])
    & ~(reorderQueueAllocate_counterWillUpdate_4[6]) & ~(reorderQueueAllocate_counterWillUpdate_5[6]) & ~(reorderQueueAllocate_counterWillUpdate_6[6]) & ~(reorderQueueAllocate_counterWillUpdate_7[6])
    & ~(reorderQueueAllocate_counterWillUpdate_8[6]) & ~(reorderQueueAllocate_counterWillUpdate_9[6]) & ~(reorderQueueAllocate_counterWillUpdate_10[6]) & ~(reorderQueueAllocate_counterWillUpdate_11[6])
    & ~(reorderQueueAllocate_counterWillUpdate_12[6]) & ~(reorderQueueAllocate_counterWillUpdate_13[6]) & ~(reorderQueueAllocate_counterWillUpdate_14[6]) & ~(reorderQueueAllocate_counterWillUpdate_15[6])
    & ~(reorderQueueAllocate_counterWillUpdate_16[6]) & ~(reorderQueueAllocate_counterWillUpdate_17[6]) & ~(reorderQueueAllocate_counterWillUpdate_18[6]) & ~(reorderQueueAllocate_counterWillUpdate_19[6])
    & ~(reorderQueueAllocate_counterWillUpdate_20[6]) & ~(reorderQueueAllocate_counterWillUpdate_21[6]) & ~(reorderQueueAllocate_counterWillUpdate_22[6]) & ~(reorderQueueAllocate_counterWillUpdate_23[6])
    & ~(reorderQueueAllocate_counterWillUpdate_24[6]) & ~(reorderQueueAllocate_counterWillUpdate_25[6]) & ~(reorderQueueAllocate_counterWillUpdate_26[6]) & ~(reorderQueueAllocate_counterWillUpdate_27[6])
    & ~(reorderQueueAllocate_counterWillUpdate_28[6]) & ~(reorderQueueAllocate_counterWillUpdate_29[6]) & ~(reorderQueueAllocate_counterWillUpdate_30[6]) & ~(reorderQueueAllocate_counterWillUpdate_31[6]);
  reg                reorderStageValid;
  reg  [5:0]         reorderStageState_0;
  reg  [5:0]         reorderStageState_1;
  reg  [5:0]         reorderStageState_2;
  reg  [5:0]         reorderStageState_3;
  reg  [5:0]         reorderStageState_4;
  reg  [5:0]         reorderStageState_5;
  reg  [5:0]         reorderStageState_6;
  reg  [5:0]         reorderStageState_7;
  reg  [5:0]         reorderStageState_8;
  reg  [5:0]         reorderStageState_9;
  reg  [5:0]         reorderStageState_10;
  reg  [5:0]         reorderStageState_11;
  reg  [5:0]         reorderStageState_12;
  reg  [5:0]         reorderStageState_13;
  reg  [5:0]         reorderStageState_14;
  reg  [5:0]         reorderStageState_15;
  reg  [5:0]         reorderStageState_16;
  reg  [5:0]         reorderStageState_17;
  reg  [5:0]         reorderStageState_18;
  reg  [5:0]         reorderStageState_19;
  reg  [5:0]         reorderStageState_20;
  reg  [5:0]         reorderStageState_21;
  reg  [5:0]         reorderStageState_22;
  reg  [5:0]         reorderStageState_23;
  reg  [5:0]         reorderStageState_24;
  reg  [5:0]         reorderStageState_25;
  reg  [5:0]         reorderStageState_26;
  reg  [5:0]         reorderStageState_27;
  reg  [5:0]         reorderStageState_28;
  reg  [5:0]         reorderStageState_29;
  reg  [5:0]         reorderStageState_30;
  reg  [5:0]         reorderStageState_31;
  reg  [5:0]         reorderStageNeed_0;
  reg  [5:0]         reorderStageNeed_1;
  reg  [5:0]         reorderStageNeed_2;
  reg  [5:0]         reorderStageNeed_3;
  reg  [5:0]         reorderStageNeed_4;
  reg  [5:0]         reorderStageNeed_5;
  reg  [5:0]         reorderStageNeed_6;
  reg  [5:0]         reorderStageNeed_7;
  reg  [5:0]         reorderStageNeed_8;
  reg  [5:0]         reorderStageNeed_9;
  reg  [5:0]         reorderStageNeed_10;
  reg  [5:0]         reorderStageNeed_11;
  reg  [5:0]         reorderStageNeed_12;
  reg  [5:0]         reorderStageNeed_13;
  reg  [5:0]         reorderStageNeed_14;
  reg  [5:0]         reorderStageNeed_15;
  reg  [5:0]         reorderStageNeed_16;
  reg  [5:0]         reorderStageNeed_17;
  reg  [5:0]         reorderStageNeed_18;
  reg  [5:0]         reorderStageNeed_19;
  reg  [5:0]         reorderStageNeed_20;
  reg  [5:0]         reorderStageNeed_21;
  reg  [5:0]         reorderStageNeed_22;
  reg  [5:0]         reorderStageNeed_23;
  reg  [5:0]         reorderStageNeed_24;
  reg  [5:0]         reorderStageNeed_25;
  reg  [5:0]         reorderStageNeed_26;
  reg  [5:0]         reorderStageNeed_27;
  reg  [5:0]         reorderStageNeed_28;
  reg  [5:0]         reorderStageNeed_29;
  reg  [5:0]         reorderStageNeed_30;
  reg  [5:0]         reorderStageNeed_31;
  wire               stateCheck =
    reorderStageState_0 == reorderStageNeed_0 & reorderStageState_1 == reorderStageNeed_1 & reorderStageState_2 == reorderStageNeed_2 & reorderStageState_3 == reorderStageNeed_3 & reorderStageState_4 == reorderStageNeed_4
    & reorderStageState_5 == reorderStageNeed_5 & reorderStageState_6 == reorderStageNeed_6 & reorderStageState_7 == reorderStageNeed_7 & reorderStageState_8 == reorderStageNeed_8 & reorderStageState_9 == reorderStageNeed_9
    & reorderStageState_10 == reorderStageNeed_10 & reorderStageState_11 == reorderStageNeed_11 & reorderStageState_12 == reorderStageNeed_12 & reorderStageState_13 == reorderStageNeed_13 & reorderStageState_14 == reorderStageNeed_14
    & reorderStageState_15 == reorderStageNeed_15 & reorderStageState_16 == reorderStageNeed_16 & reorderStageState_17 == reorderStageNeed_17 & reorderStageState_18 == reorderStageNeed_18 & reorderStageState_19 == reorderStageNeed_19
    & reorderStageState_20 == reorderStageNeed_20 & reorderStageState_21 == reorderStageNeed_21 & reorderStageState_22 == reorderStageNeed_22 & reorderStageState_23 == reorderStageNeed_23 & reorderStageState_24 == reorderStageNeed_24
    & reorderStageState_25 == reorderStageNeed_25 & reorderStageState_26 == reorderStageNeed_26 & reorderStageState_27 == reorderStageNeed_27 & reorderStageState_28 == reorderStageNeed_28 & reorderStageState_29 == reorderStageNeed_29
    & reorderStageState_30 == reorderStageNeed_30 & reorderStageState_31 == reorderStageNeed_31;
  assign accessCountQueue_deq_ready = ~reorderStageValid | stateCheck;
  wire               reorderStageEnqFire = accessCountQueue_deq_ready & accessCountQueue_deq_valid;
  wire               reorderStageDeqFire = stateCheck & reorderStageValid;
  wire [31:0]        sourceLane;
  wire               readMessageQueue_deq_valid;
  assign readMessageQueue_deq_valid = ~_readMessageQueue_fifo_empty;
  wire [31:0]        readMessageQueue_dataOut_readSource;
  assign reorderQueueVec_0_enq_bits_write1H = readMessageQueue_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_dataOffset;
  wire [31:0]        readMessageQueue_enq_bits_readSource;
  wire [1:0]         readMessageQueue_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn = {readMessageQueue_enq_bits_readSource, readMessageQueue_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_dataOffset = _readMessageQueue_fifo_data_out[1:0];
  assign readMessageQueue_dataOut_readSource = _readMessageQueue_fifo_data_out[33:2];
  assign readMessageQueue_deq_bits_readSource = readMessageQueue_dataOut_readSource;
  wire [1:0]         readMessageQueue_deq_bits_dataOffset = readMessageQueue_dataOut_dataOffset;
  wire               readMessageQueue_enq_ready = ~_readMessageQueue_fifo_full;
  wire               readMessageQueue_enq_valid;
  assign deqAllocate = ~readValid | reorderStageValid & reorderStageState_0 != reorderStageNeed_0;
  assign reorderQueueVec_0_deq_ready = deqAllocate;
  assign sourceLane = 32'h1 << _readCrossBar_output_0_bits_writeIndex;
  assign readMessageQueue_enq_bits_readSource = sourceLane;
  wire               readChannel_0_valid_0 = maskDestinationType ? _maskedWrite_readChannel_0_valid : _readCrossBar_output_0_valid & readMessageQueue_enq_ready;
  wire [4:0]         readChannel_0_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_0_bits_vs : _readCrossBar_output_0_bits_vs;
  wire               readChannel_0_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_0_bits_offset : _readCrossBar_output_0_bits_offset;
  assign readMessageQueue_enq_valid = readChannel_0_ready_0 & readChannel_0_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_0_enq_bits_data = readResult_0_bits >> {27'h0, readMessageQueue_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_0 = _write1HPipe_0_T & ~maskDestinationType ? reorderQueueVec_0_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_1;
  wire               readMessageQueue_1_deq_valid;
  assign readMessageQueue_1_deq_valid = ~_readMessageQueue_fifo_1_empty;
  wire [31:0]        readMessageQueue_dataOut_1_readSource;
  assign reorderQueueVec_1_enq_bits_write1H = readMessageQueue_1_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_1_dataOffset;
  wire [31:0]        readMessageQueue_1_enq_bits_readSource;
  wire [1:0]         readMessageQueue_1_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_1 = {readMessageQueue_1_enq_bits_readSource, readMessageQueue_1_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_1_dataOffset = _readMessageQueue_fifo_1_data_out[1:0];
  assign readMessageQueue_dataOut_1_readSource = _readMessageQueue_fifo_1_data_out[33:2];
  assign readMessageQueue_1_deq_bits_readSource = readMessageQueue_dataOut_1_readSource;
  wire [1:0]         readMessageQueue_1_deq_bits_dataOffset = readMessageQueue_dataOut_1_dataOffset;
  wire               readMessageQueue_1_enq_ready = ~_readMessageQueue_fifo_1_full;
  wire               readMessageQueue_1_enq_valid;
  assign deqAllocate_1 = ~readValid | reorderStageValid & reorderStageState_1 != reorderStageNeed_1;
  assign reorderQueueVec_1_deq_ready = deqAllocate_1;
  assign sourceLane_1 = 32'h1 << _readCrossBar_output_1_bits_writeIndex;
  assign readMessageQueue_1_enq_bits_readSource = sourceLane_1;
  wire               readChannel_1_valid_0 = maskDestinationType ? _maskedWrite_readChannel_1_valid : _readCrossBar_output_1_valid & readMessageQueue_1_enq_ready;
  wire [4:0]         readChannel_1_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_1_bits_vs : _readCrossBar_output_1_bits_vs;
  wire               readChannel_1_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_1_bits_offset : _readCrossBar_output_1_bits_offset;
  assign readMessageQueue_1_enq_valid = readChannel_1_ready_0 & readChannel_1_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_1_enq_bits_data = readResult_1_bits >> {27'h0, readMessageQueue_1_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_1 = _write1HPipe_1_T & ~maskDestinationType ? reorderQueueVec_1_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_2;
  wire               readMessageQueue_2_deq_valid;
  assign readMessageQueue_2_deq_valid = ~_readMessageQueue_fifo_2_empty;
  wire [31:0]        readMessageQueue_dataOut_2_readSource;
  assign reorderQueueVec_2_enq_bits_write1H = readMessageQueue_2_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_2_dataOffset;
  wire [31:0]        readMessageQueue_2_enq_bits_readSource;
  wire [1:0]         readMessageQueue_2_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_2 = {readMessageQueue_2_enq_bits_readSource, readMessageQueue_2_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_2_dataOffset = _readMessageQueue_fifo_2_data_out[1:0];
  assign readMessageQueue_dataOut_2_readSource = _readMessageQueue_fifo_2_data_out[33:2];
  assign readMessageQueue_2_deq_bits_readSource = readMessageQueue_dataOut_2_readSource;
  wire [1:0]         readMessageQueue_2_deq_bits_dataOffset = readMessageQueue_dataOut_2_dataOffset;
  wire               readMessageQueue_2_enq_ready = ~_readMessageQueue_fifo_2_full;
  wire               readMessageQueue_2_enq_valid;
  assign deqAllocate_2 = ~readValid | reorderStageValid & reorderStageState_2 != reorderStageNeed_2;
  assign reorderQueueVec_2_deq_ready = deqAllocate_2;
  assign sourceLane_2 = 32'h1 << _readCrossBar_output_2_bits_writeIndex;
  assign readMessageQueue_2_enq_bits_readSource = sourceLane_2;
  wire               readChannel_2_valid_0 = maskDestinationType ? _maskedWrite_readChannel_2_valid : _readCrossBar_output_2_valid & readMessageQueue_2_enq_ready;
  wire [4:0]         readChannel_2_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_2_bits_vs : _readCrossBar_output_2_bits_vs;
  wire               readChannel_2_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_2_bits_offset : _readCrossBar_output_2_bits_offset;
  assign readMessageQueue_2_enq_valid = readChannel_2_ready_0 & readChannel_2_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_2_enq_bits_data = readResult_2_bits >> {27'h0, readMessageQueue_2_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_2 = _write1HPipe_2_T & ~maskDestinationType ? reorderQueueVec_2_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_3;
  wire               readMessageQueue_3_deq_valid;
  assign readMessageQueue_3_deq_valid = ~_readMessageQueue_fifo_3_empty;
  wire [31:0]        readMessageQueue_dataOut_3_readSource;
  assign reorderQueueVec_3_enq_bits_write1H = readMessageQueue_3_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_3_dataOffset;
  wire [31:0]        readMessageQueue_3_enq_bits_readSource;
  wire [1:0]         readMessageQueue_3_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_3 = {readMessageQueue_3_enq_bits_readSource, readMessageQueue_3_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_3_dataOffset = _readMessageQueue_fifo_3_data_out[1:0];
  assign readMessageQueue_dataOut_3_readSource = _readMessageQueue_fifo_3_data_out[33:2];
  assign readMessageQueue_3_deq_bits_readSource = readMessageQueue_dataOut_3_readSource;
  wire [1:0]         readMessageQueue_3_deq_bits_dataOffset = readMessageQueue_dataOut_3_dataOffset;
  wire               readMessageQueue_3_enq_ready = ~_readMessageQueue_fifo_3_full;
  wire               readMessageQueue_3_enq_valid;
  assign deqAllocate_3 = ~readValid | reorderStageValid & reorderStageState_3 != reorderStageNeed_3;
  assign reorderQueueVec_3_deq_ready = deqAllocate_3;
  assign sourceLane_3 = 32'h1 << _readCrossBar_output_3_bits_writeIndex;
  assign readMessageQueue_3_enq_bits_readSource = sourceLane_3;
  wire               readChannel_3_valid_0 = maskDestinationType ? _maskedWrite_readChannel_3_valid : _readCrossBar_output_3_valid & readMessageQueue_3_enq_ready;
  wire [4:0]         readChannel_3_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_3_bits_vs : _readCrossBar_output_3_bits_vs;
  wire               readChannel_3_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_3_bits_offset : _readCrossBar_output_3_bits_offset;
  assign readMessageQueue_3_enq_valid = readChannel_3_ready_0 & readChannel_3_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_3_enq_bits_data = readResult_3_bits >> {27'h0, readMessageQueue_3_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_3 = _write1HPipe_3_T & ~maskDestinationType ? reorderQueueVec_3_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_4;
  wire               readMessageQueue_4_deq_valid;
  assign readMessageQueue_4_deq_valid = ~_readMessageQueue_fifo_4_empty;
  wire [31:0]        readMessageQueue_dataOut_4_readSource;
  assign reorderQueueVec_4_enq_bits_write1H = readMessageQueue_4_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_4_dataOffset;
  wire [31:0]        readMessageQueue_4_enq_bits_readSource;
  wire [1:0]         readMessageQueue_4_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_4 = {readMessageQueue_4_enq_bits_readSource, readMessageQueue_4_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_4_dataOffset = _readMessageQueue_fifo_4_data_out[1:0];
  assign readMessageQueue_dataOut_4_readSource = _readMessageQueue_fifo_4_data_out[33:2];
  assign readMessageQueue_4_deq_bits_readSource = readMessageQueue_dataOut_4_readSource;
  wire [1:0]         readMessageQueue_4_deq_bits_dataOffset = readMessageQueue_dataOut_4_dataOffset;
  wire               readMessageQueue_4_enq_ready = ~_readMessageQueue_fifo_4_full;
  wire               readMessageQueue_4_enq_valid;
  assign deqAllocate_4 = ~readValid | reorderStageValid & reorderStageState_4 != reorderStageNeed_4;
  assign reorderQueueVec_4_deq_ready = deqAllocate_4;
  assign sourceLane_4 = 32'h1 << _readCrossBar_output_4_bits_writeIndex;
  assign readMessageQueue_4_enq_bits_readSource = sourceLane_4;
  wire               readChannel_4_valid_0 = maskDestinationType ? _maskedWrite_readChannel_4_valid : _readCrossBar_output_4_valid & readMessageQueue_4_enq_ready;
  wire [4:0]         readChannel_4_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_4_bits_vs : _readCrossBar_output_4_bits_vs;
  wire               readChannel_4_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_4_bits_offset : _readCrossBar_output_4_bits_offset;
  assign readMessageQueue_4_enq_valid = readChannel_4_ready_0 & readChannel_4_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_4_enq_bits_data = readResult_4_bits >> {27'h0, readMessageQueue_4_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_4 = _write1HPipe_4_T & ~maskDestinationType ? reorderQueueVec_4_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_5;
  wire               readMessageQueue_5_deq_valid;
  assign readMessageQueue_5_deq_valid = ~_readMessageQueue_fifo_5_empty;
  wire [31:0]        readMessageQueue_dataOut_5_readSource;
  assign reorderQueueVec_5_enq_bits_write1H = readMessageQueue_5_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_5_dataOffset;
  wire [31:0]        readMessageQueue_5_enq_bits_readSource;
  wire [1:0]         readMessageQueue_5_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_5 = {readMessageQueue_5_enq_bits_readSource, readMessageQueue_5_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_5_dataOffset = _readMessageQueue_fifo_5_data_out[1:0];
  assign readMessageQueue_dataOut_5_readSource = _readMessageQueue_fifo_5_data_out[33:2];
  assign readMessageQueue_5_deq_bits_readSource = readMessageQueue_dataOut_5_readSource;
  wire [1:0]         readMessageQueue_5_deq_bits_dataOffset = readMessageQueue_dataOut_5_dataOffset;
  wire               readMessageQueue_5_enq_ready = ~_readMessageQueue_fifo_5_full;
  wire               readMessageQueue_5_enq_valid;
  assign deqAllocate_5 = ~readValid | reorderStageValid & reorderStageState_5 != reorderStageNeed_5;
  assign reorderQueueVec_5_deq_ready = deqAllocate_5;
  assign sourceLane_5 = 32'h1 << _readCrossBar_output_5_bits_writeIndex;
  assign readMessageQueue_5_enq_bits_readSource = sourceLane_5;
  wire               readChannel_5_valid_0 = maskDestinationType ? _maskedWrite_readChannel_5_valid : _readCrossBar_output_5_valid & readMessageQueue_5_enq_ready;
  wire [4:0]         readChannel_5_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_5_bits_vs : _readCrossBar_output_5_bits_vs;
  wire               readChannel_5_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_5_bits_offset : _readCrossBar_output_5_bits_offset;
  assign readMessageQueue_5_enq_valid = readChannel_5_ready_0 & readChannel_5_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_5_enq_bits_data = readResult_5_bits >> {27'h0, readMessageQueue_5_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_5 = _write1HPipe_5_T & ~maskDestinationType ? reorderQueueVec_5_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_6;
  wire               readMessageQueue_6_deq_valid;
  assign readMessageQueue_6_deq_valid = ~_readMessageQueue_fifo_6_empty;
  wire [31:0]        readMessageQueue_dataOut_6_readSource;
  assign reorderQueueVec_6_enq_bits_write1H = readMessageQueue_6_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_6_dataOffset;
  wire [31:0]        readMessageQueue_6_enq_bits_readSource;
  wire [1:0]         readMessageQueue_6_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_6 = {readMessageQueue_6_enq_bits_readSource, readMessageQueue_6_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_6_dataOffset = _readMessageQueue_fifo_6_data_out[1:0];
  assign readMessageQueue_dataOut_6_readSource = _readMessageQueue_fifo_6_data_out[33:2];
  assign readMessageQueue_6_deq_bits_readSource = readMessageQueue_dataOut_6_readSource;
  wire [1:0]         readMessageQueue_6_deq_bits_dataOffset = readMessageQueue_dataOut_6_dataOffset;
  wire               readMessageQueue_6_enq_ready = ~_readMessageQueue_fifo_6_full;
  wire               readMessageQueue_6_enq_valid;
  assign deqAllocate_6 = ~readValid | reorderStageValid & reorderStageState_6 != reorderStageNeed_6;
  assign reorderQueueVec_6_deq_ready = deqAllocate_6;
  assign sourceLane_6 = 32'h1 << _readCrossBar_output_6_bits_writeIndex;
  assign readMessageQueue_6_enq_bits_readSource = sourceLane_6;
  wire               readChannel_6_valid_0 = maskDestinationType ? _maskedWrite_readChannel_6_valid : _readCrossBar_output_6_valid & readMessageQueue_6_enq_ready;
  wire [4:0]         readChannel_6_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_6_bits_vs : _readCrossBar_output_6_bits_vs;
  wire               readChannel_6_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_6_bits_offset : _readCrossBar_output_6_bits_offset;
  assign readMessageQueue_6_enq_valid = readChannel_6_ready_0 & readChannel_6_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_6_enq_bits_data = readResult_6_bits >> {27'h0, readMessageQueue_6_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_6 = _write1HPipe_6_T & ~maskDestinationType ? reorderQueueVec_6_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_7;
  wire               readMessageQueue_7_deq_valid;
  assign readMessageQueue_7_deq_valid = ~_readMessageQueue_fifo_7_empty;
  wire [31:0]        readMessageQueue_dataOut_7_readSource;
  assign reorderQueueVec_7_enq_bits_write1H = readMessageQueue_7_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_7_dataOffset;
  wire [31:0]        readMessageQueue_7_enq_bits_readSource;
  wire [1:0]         readMessageQueue_7_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_7 = {readMessageQueue_7_enq_bits_readSource, readMessageQueue_7_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_7_dataOffset = _readMessageQueue_fifo_7_data_out[1:0];
  assign readMessageQueue_dataOut_7_readSource = _readMessageQueue_fifo_7_data_out[33:2];
  assign readMessageQueue_7_deq_bits_readSource = readMessageQueue_dataOut_7_readSource;
  wire [1:0]         readMessageQueue_7_deq_bits_dataOffset = readMessageQueue_dataOut_7_dataOffset;
  wire               readMessageQueue_7_enq_ready = ~_readMessageQueue_fifo_7_full;
  wire               readMessageQueue_7_enq_valid;
  assign deqAllocate_7 = ~readValid | reorderStageValid & reorderStageState_7 != reorderStageNeed_7;
  assign reorderQueueVec_7_deq_ready = deqAllocate_7;
  assign sourceLane_7 = 32'h1 << _readCrossBar_output_7_bits_writeIndex;
  assign readMessageQueue_7_enq_bits_readSource = sourceLane_7;
  wire               readChannel_7_valid_0 = maskDestinationType ? _maskedWrite_readChannel_7_valid : _readCrossBar_output_7_valid & readMessageQueue_7_enq_ready;
  wire [4:0]         readChannel_7_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_7_bits_vs : _readCrossBar_output_7_bits_vs;
  wire               readChannel_7_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_7_bits_offset : _readCrossBar_output_7_bits_offset;
  assign readMessageQueue_7_enq_valid = readChannel_7_ready_0 & readChannel_7_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_7_enq_bits_data = readResult_7_bits >> {27'h0, readMessageQueue_7_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_7 = _write1HPipe_7_T & ~maskDestinationType ? reorderQueueVec_7_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_8;
  wire               readMessageQueue_8_deq_valid;
  assign readMessageQueue_8_deq_valid = ~_readMessageQueue_fifo_8_empty;
  wire [31:0]        readMessageQueue_dataOut_8_readSource;
  assign reorderQueueVec_8_enq_bits_write1H = readMessageQueue_8_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_8_dataOffset;
  wire [31:0]        readMessageQueue_8_enq_bits_readSource;
  wire [1:0]         readMessageQueue_8_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_8 = {readMessageQueue_8_enq_bits_readSource, readMessageQueue_8_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_8_dataOffset = _readMessageQueue_fifo_8_data_out[1:0];
  assign readMessageQueue_dataOut_8_readSource = _readMessageQueue_fifo_8_data_out[33:2];
  assign readMessageQueue_8_deq_bits_readSource = readMessageQueue_dataOut_8_readSource;
  wire [1:0]         readMessageQueue_8_deq_bits_dataOffset = readMessageQueue_dataOut_8_dataOffset;
  wire               readMessageQueue_8_enq_ready = ~_readMessageQueue_fifo_8_full;
  wire               readMessageQueue_8_enq_valid;
  assign deqAllocate_8 = ~readValid | reorderStageValid & reorderStageState_8 != reorderStageNeed_8;
  assign reorderQueueVec_8_deq_ready = deqAllocate_8;
  assign sourceLane_8 = 32'h1 << _readCrossBar_output_8_bits_writeIndex;
  assign readMessageQueue_8_enq_bits_readSource = sourceLane_8;
  wire               readChannel_8_valid_0 = maskDestinationType ? _maskedWrite_readChannel_8_valid : _readCrossBar_output_8_valid & readMessageQueue_8_enq_ready;
  wire [4:0]         readChannel_8_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_8_bits_vs : _readCrossBar_output_8_bits_vs;
  wire               readChannel_8_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_8_bits_offset : _readCrossBar_output_8_bits_offset;
  assign readMessageQueue_8_enq_valid = readChannel_8_ready_0 & readChannel_8_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_8_enq_bits_data = readResult_8_bits >> {27'h0, readMessageQueue_8_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_8 = _write1HPipe_8_T & ~maskDestinationType ? reorderQueueVec_8_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_9;
  wire               readMessageQueue_9_deq_valid;
  assign readMessageQueue_9_deq_valid = ~_readMessageQueue_fifo_9_empty;
  wire [31:0]        readMessageQueue_dataOut_9_readSource;
  assign reorderQueueVec_9_enq_bits_write1H = readMessageQueue_9_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_9_dataOffset;
  wire [31:0]        readMessageQueue_9_enq_bits_readSource;
  wire [1:0]         readMessageQueue_9_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_9 = {readMessageQueue_9_enq_bits_readSource, readMessageQueue_9_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_9_dataOffset = _readMessageQueue_fifo_9_data_out[1:0];
  assign readMessageQueue_dataOut_9_readSource = _readMessageQueue_fifo_9_data_out[33:2];
  assign readMessageQueue_9_deq_bits_readSource = readMessageQueue_dataOut_9_readSource;
  wire [1:0]         readMessageQueue_9_deq_bits_dataOffset = readMessageQueue_dataOut_9_dataOffset;
  wire               readMessageQueue_9_enq_ready = ~_readMessageQueue_fifo_9_full;
  wire               readMessageQueue_9_enq_valid;
  assign deqAllocate_9 = ~readValid | reorderStageValid & reorderStageState_9 != reorderStageNeed_9;
  assign reorderQueueVec_9_deq_ready = deqAllocate_9;
  assign sourceLane_9 = 32'h1 << _readCrossBar_output_9_bits_writeIndex;
  assign readMessageQueue_9_enq_bits_readSource = sourceLane_9;
  wire               readChannel_9_valid_0 = maskDestinationType ? _maskedWrite_readChannel_9_valid : _readCrossBar_output_9_valid & readMessageQueue_9_enq_ready;
  wire [4:0]         readChannel_9_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_9_bits_vs : _readCrossBar_output_9_bits_vs;
  wire               readChannel_9_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_9_bits_offset : _readCrossBar_output_9_bits_offset;
  assign readMessageQueue_9_enq_valid = readChannel_9_ready_0 & readChannel_9_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_9_enq_bits_data = readResult_9_bits >> {27'h0, readMessageQueue_9_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_9 = _write1HPipe_9_T & ~maskDestinationType ? reorderQueueVec_9_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_10;
  wire               readMessageQueue_10_deq_valid;
  assign readMessageQueue_10_deq_valid = ~_readMessageQueue_fifo_10_empty;
  wire [31:0]        readMessageQueue_dataOut_10_readSource;
  assign reorderQueueVec_10_enq_bits_write1H = readMessageQueue_10_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_10_dataOffset;
  wire [31:0]        readMessageQueue_10_enq_bits_readSource;
  wire [1:0]         readMessageQueue_10_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_10 = {readMessageQueue_10_enq_bits_readSource, readMessageQueue_10_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_10_dataOffset = _readMessageQueue_fifo_10_data_out[1:0];
  assign readMessageQueue_dataOut_10_readSource = _readMessageQueue_fifo_10_data_out[33:2];
  assign readMessageQueue_10_deq_bits_readSource = readMessageQueue_dataOut_10_readSource;
  wire [1:0]         readMessageQueue_10_deq_bits_dataOffset = readMessageQueue_dataOut_10_dataOffset;
  wire               readMessageQueue_10_enq_ready = ~_readMessageQueue_fifo_10_full;
  wire               readMessageQueue_10_enq_valid;
  assign deqAllocate_10 = ~readValid | reorderStageValid & reorderStageState_10 != reorderStageNeed_10;
  assign reorderQueueVec_10_deq_ready = deqAllocate_10;
  assign sourceLane_10 = 32'h1 << _readCrossBar_output_10_bits_writeIndex;
  assign readMessageQueue_10_enq_bits_readSource = sourceLane_10;
  wire               readChannel_10_valid_0 = maskDestinationType ? _maskedWrite_readChannel_10_valid : _readCrossBar_output_10_valid & readMessageQueue_10_enq_ready;
  wire [4:0]         readChannel_10_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_10_bits_vs : _readCrossBar_output_10_bits_vs;
  wire               readChannel_10_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_10_bits_offset : _readCrossBar_output_10_bits_offset;
  assign readMessageQueue_10_enq_valid = readChannel_10_ready_0 & readChannel_10_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_10_enq_bits_data = readResult_10_bits >> {27'h0, readMessageQueue_10_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_10 = _write1HPipe_10_T & ~maskDestinationType ? reorderQueueVec_10_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_11;
  wire               readMessageQueue_11_deq_valid;
  assign readMessageQueue_11_deq_valid = ~_readMessageQueue_fifo_11_empty;
  wire [31:0]        readMessageQueue_dataOut_11_readSource;
  assign reorderQueueVec_11_enq_bits_write1H = readMessageQueue_11_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_11_dataOffset;
  wire [31:0]        readMessageQueue_11_enq_bits_readSource;
  wire [1:0]         readMessageQueue_11_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_11 = {readMessageQueue_11_enq_bits_readSource, readMessageQueue_11_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_11_dataOffset = _readMessageQueue_fifo_11_data_out[1:0];
  assign readMessageQueue_dataOut_11_readSource = _readMessageQueue_fifo_11_data_out[33:2];
  assign readMessageQueue_11_deq_bits_readSource = readMessageQueue_dataOut_11_readSource;
  wire [1:0]         readMessageQueue_11_deq_bits_dataOffset = readMessageQueue_dataOut_11_dataOffset;
  wire               readMessageQueue_11_enq_ready = ~_readMessageQueue_fifo_11_full;
  wire               readMessageQueue_11_enq_valid;
  assign deqAllocate_11 = ~readValid | reorderStageValid & reorderStageState_11 != reorderStageNeed_11;
  assign reorderQueueVec_11_deq_ready = deqAllocate_11;
  assign sourceLane_11 = 32'h1 << _readCrossBar_output_11_bits_writeIndex;
  assign readMessageQueue_11_enq_bits_readSource = sourceLane_11;
  wire               readChannel_11_valid_0 = maskDestinationType ? _maskedWrite_readChannel_11_valid : _readCrossBar_output_11_valid & readMessageQueue_11_enq_ready;
  wire [4:0]         readChannel_11_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_11_bits_vs : _readCrossBar_output_11_bits_vs;
  wire               readChannel_11_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_11_bits_offset : _readCrossBar_output_11_bits_offset;
  assign readMessageQueue_11_enq_valid = readChannel_11_ready_0 & readChannel_11_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_11_enq_bits_data = readResult_11_bits >> {27'h0, readMessageQueue_11_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_11 = _write1HPipe_11_T & ~maskDestinationType ? reorderQueueVec_11_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_12;
  wire               readMessageQueue_12_deq_valid;
  assign readMessageQueue_12_deq_valid = ~_readMessageQueue_fifo_12_empty;
  wire [31:0]        readMessageQueue_dataOut_12_readSource;
  assign reorderQueueVec_12_enq_bits_write1H = readMessageQueue_12_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_12_dataOffset;
  wire [31:0]        readMessageQueue_12_enq_bits_readSource;
  wire [1:0]         readMessageQueue_12_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_12 = {readMessageQueue_12_enq_bits_readSource, readMessageQueue_12_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_12_dataOffset = _readMessageQueue_fifo_12_data_out[1:0];
  assign readMessageQueue_dataOut_12_readSource = _readMessageQueue_fifo_12_data_out[33:2];
  assign readMessageQueue_12_deq_bits_readSource = readMessageQueue_dataOut_12_readSource;
  wire [1:0]         readMessageQueue_12_deq_bits_dataOffset = readMessageQueue_dataOut_12_dataOffset;
  wire               readMessageQueue_12_enq_ready = ~_readMessageQueue_fifo_12_full;
  wire               readMessageQueue_12_enq_valid;
  assign deqAllocate_12 = ~readValid | reorderStageValid & reorderStageState_12 != reorderStageNeed_12;
  assign reorderQueueVec_12_deq_ready = deqAllocate_12;
  assign sourceLane_12 = 32'h1 << _readCrossBar_output_12_bits_writeIndex;
  assign readMessageQueue_12_enq_bits_readSource = sourceLane_12;
  wire               readChannel_12_valid_0 = maskDestinationType ? _maskedWrite_readChannel_12_valid : _readCrossBar_output_12_valid & readMessageQueue_12_enq_ready;
  wire [4:0]         readChannel_12_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_12_bits_vs : _readCrossBar_output_12_bits_vs;
  wire               readChannel_12_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_12_bits_offset : _readCrossBar_output_12_bits_offset;
  assign readMessageQueue_12_enq_valid = readChannel_12_ready_0 & readChannel_12_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_12_enq_bits_data = readResult_12_bits >> {27'h0, readMessageQueue_12_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_12 = _write1HPipe_12_T & ~maskDestinationType ? reorderQueueVec_12_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_13;
  wire               readMessageQueue_13_deq_valid;
  assign readMessageQueue_13_deq_valid = ~_readMessageQueue_fifo_13_empty;
  wire [31:0]        readMessageQueue_dataOut_13_readSource;
  assign reorderQueueVec_13_enq_bits_write1H = readMessageQueue_13_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_13_dataOffset;
  wire [31:0]        readMessageQueue_13_enq_bits_readSource;
  wire [1:0]         readMessageQueue_13_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_13 = {readMessageQueue_13_enq_bits_readSource, readMessageQueue_13_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_13_dataOffset = _readMessageQueue_fifo_13_data_out[1:0];
  assign readMessageQueue_dataOut_13_readSource = _readMessageQueue_fifo_13_data_out[33:2];
  assign readMessageQueue_13_deq_bits_readSource = readMessageQueue_dataOut_13_readSource;
  wire [1:0]         readMessageQueue_13_deq_bits_dataOffset = readMessageQueue_dataOut_13_dataOffset;
  wire               readMessageQueue_13_enq_ready = ~_readMessageQueue_fifo_13_full;
  wire               readMessageQueue_13_enq_valid;
  assign deqAllocate_13 = ~readValid | reorderStageValid & reorderStageState_13 != reorderStageNeed_13;
  assign reorderQueueVec_13_deq_ready = deqAllocate_13;
  assign sourceLane_13 = 32'h1 << _readCrossBar_output_13_bits_writeIndex;
  assign readMessageQueue_13_enq_bits_readSource = sourceLane_13;
  wire               readChannel_13_valid_0 = maskDestinationType ? _maskedWrite_readChannel_13_valid : _readCrossBar_output_13_valid & readMessageQueue_13_enq_ready;
  wire [4:0]         readChannel_13_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_13_bits_vs : _readCrossBar_output_13_bits_vs;
  wire               readChannel_13_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_13_bits_offset : _readCrossBar_output_13_bits_offset;
  assign readMessageQueue_13_enq_valid = readChannel_13_ready_0 & readChannel_13_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_13_enq_bits_data = readResult_13_bits >> {27'h0, readMessageQueue_13_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_13 = _write1HPipe_13_T & ~maskDestinationType ? reorderQueueVec_13_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_14;
  wire               readMessageQueue_14_deq_valid;
  assign readMessageQueue_14_deq_valid = ~_readMessageQueue_fifo_14_empty;
  wire [31:0]        readMessageQueue_dataOut_14_readSource;
  assign reorderQueueVec_14_enq_bits_write1H = readMessageQueue_14_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_14_dataOffset;
  wire [31:0]        readMessageQueue_14_enq_bits_readSource;
  wire [1:0]         readMessageQueue_14_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_14 = {readMessageQueue_14_enq_bits_readSource, readMessageQueue_14_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_14_dataOffset = _readMessageQueue_fifo_14_data_out[1:0];
  assign readMessageQueue_dataOut_14_readSource = _readMessageQueue_fifo_14_data_out[33:2];
  assign readMessageQueue_14_deq_bits_readSource = readMessageQueue_dataOut_14_readSource;
  wire [1:0]         readMessageQueue_14_deq_bits_dataOffset = readMessageQueue_dataOut_14_dataOffset;
  wire               readMessageQueue_14_enq_ready = ~_readMessageQueue_fifo_14_full;
  wire               readMessageQueue_14_enq_valid;
  assign deqAllocate_14 = ~readValid | reorderStageValid & reorderStageState_14 != reorderStageNeed_14;
  assign reorderQueueVec_14_deq_ready = deqAllocate_14;
  assign sourceLane_14 = 32'h1 << _readCrossBar_output_14_bits_writeIndex;
  assign readMessageQueue_14_enq_bits_readSource = sourceLane_14;
  wire               readChannel_14_valid_0 = maskDestinationType ? _maskedWrite_readChannel_14_valid : _readCrossBar_output_14_valid & readMessageQueue_14_enq_ready;
  wire [4:0]         readChannel_14_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_14_bits_vs : _readCrossBar_output_14_bits_vs;
  wire               readChannel_14_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_14_bits_offset : _readCrossBar_output_14_bits_offset;
  assign readMessageQueue_14_enq_valid = readChannel_14_ready_0 & readChannel_14_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_14_enq_bits_data = readResult_14_bits >> {27'h0, readMessageQueue_14_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_14 = _write1HPipe_14_T & ~maskDestinationType ? reorderQueueVec_14_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_15;
  wire               readMessageQueue_15_deq_valid;
  assign readMessageQueue_15_deq_valid = ~_readMessageQueue_fifo_15_empty;
  wire [31:0]        readMessageQueue_dataOut_15_readSource;
  assign reorderQueueVec_15_enq_bits_write1H = readMessageQueue_15_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_15_dataOffset;
  wire [31:0]        readMessageQueue_15_enq_bits_readSource;
  wire [1:0]         readMessageQueue_15_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_15 = {readMessageQueue_15_enq_bits_readSource, readMessageQueue_15_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_15_dataOffset = _readMessageQueue_fifo_15_data_out[1:0];
  assign readMessageQueue_dataOut_15_readSource = _readMessageQueue_fifo_15_data_out[33:2];
  assign readMessageQueue_15_deq_bits_readSource = readMessageQueue_dataOut_15_readSource;
  wire [1:0]         readMessageQueue_15_deq_bits_dataOffset = readMessageQueue_dataOut_15_dataOffset;
  wire               readMessageQueue_15_enq_ready = ~_readMessageQueue_fifo_15_full;
  wire               readMessageQueue_15_enq_valid;
  assign deqAllocate_15 = ~readValid | reorderStageValid & reorderStageState_15 != reorderStageNeed_15;
  assign reorderQueueVec_15_deq_ready = deqAllocate_15;
  assign sourceLane_15 = 32'h1 << _readCrossBar_output_15_bits_writeIndex;
  assign readMessageQueue_15_enq_bits_readSource = sourceLane_15;
  wire               readChannel_15_valid_0 = maskDestinationType ? _maskedWrite_readChannel_15_valid : _readCrossBar_output_15_valid & readMessageQueue_15_enq_ready;
  wire [4:0]         readChannel_15_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_15_bits_vs : _readCrossBar_output_15_bits_vs;
  wire               readChannel_15_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_15_bits_offset : _readCrossBar_output_15_bits_offset;
  assign readMessageQueue_15_enq_valid = readChannel_15_ready_0 & readChannel_15_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_15_enq_bits_data = readResult_15_bits >> {27'h0, readMessageQueue_15_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_15 = _write1HPipe_15_T & ~maskDestinationType ? reorderQueueVec_15_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_16;
  wire               readMessageQueue_16_deq_valid;
  assign readMessageQueue_16_deq_valid = ~_readMessageQueue_fifo_16_empty;
  wire [31:0]        readMessageQueue_dataOut_16_readSource;
  assign reorderQueueVec_16_enq_bits_write1H = readMessageQueue_16_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_16_dataOffset;
  wire [31:0]        readMessageQueue_16_enq_bits_readSource;
  wire [1:0]         readMessageQueue_16_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_16 = {readMessageQueue_16_enq_bits_readSource, readMessageQueue_16_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_16_dataOffset = _readMessageQueue_fifo_16_data_out[1:0];
  assign readMessageQueue_dataOut_16_readSource = _readMessageQueue_fifo_16_data_out[33:2];
  assign readMessageQueue_16_deq_bits_readSource = readMessageQueue_dataOut_16_readSource;
  wire [1:0]         readMessageQueue_16_deq_bits_dataOffset = readMessageQueue_dataOut_16_dataOffset;
  wire               readMessageQueue_16_enq_ready = ~_readMessageQueue_fifo_16_full;
  wire               readMessageQueue_16_enq_valid;
  assign deqAllocate_16 = ~readValid | reorderStageValid & reorderStageState_16 != reorderStageNeed_16;
  assign reorderQueueVec_16_deq_ready = deqAllocate_16;
  assign sourceLane_16 = 32'h1 << _readCrossBar_output_16_bits_writeIndex;
  assign readMessageQueue_16_enq_bits_readSource = sourceLane_16;
  wire               readChannel_16_valid_0 = maskDestinationType ? _maskedWrite_readChannel_16_valid : _readCrossBar_output_16_valid & readMessageQueue_16_enq_ready;
  wire [4:0]         readChannel_16_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_16_bits_vs : _readCrossBar_output_16_bits_vs;
  wire               readChannel_16_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_16_bits_offset : _readCrossBar_output_16_bits_offset;
  assign readMessageQueue_16_enq_valid = readChannel_16_ready_0 & readChannel_16_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_16_enq_bits_data = readResult_16_bits >> {27'h0, readMessageQueue_16_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_16 = _write1HPipe_16_T & ~maskDestinationType ? reorderQueueVec_16_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_17;
  wire               readMessageQueue_17_deq_valid;
  assign readMessageQueue_17_deq_valid = ~_readMessageQueue_fifo_17_empty;
  wire [31:0]        readMessageQueue_dataOut_17_readSource;
  assign reorderQueueVec_17_enq_bits_write1H = readMessageQueue_17_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_17_dataOffset;
  wire [31:0]        readMessageQueue_17_enq_bits_readSource;
  wire [1:0]         readMessageQueue_17_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_17 = {readMessageQueue_17_enq_bits_readSource, readMessageQueue_17_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_17_dataOffset = _readMessageQueue_fifo_17_data_out[1:0];
  assign readMessageQueue_dataOut_17_readSource = _readMessageQueue_fifo_17_data_out[33:2];
  assign readMessageQueue_17_deq_bits_readSource = readMessageQueue_dataOut_17_readSource;
  wire [1:0]         readMessageQueue_17_deq_bits_dataOffset = readMessageQueue_dataOut_17_dataOffset;
  wire               readMessageQueue_17_enq_ready = ~_readMessageQueue_fifo_17_full;
  wire               readMessageQueue_17_enq_valid;
  assign deqAllocate_17 = ~readValid | reorderStageValid & reorderStageState_17 != reorderStageNeed_17;
  assign reorderQueueVec_17_deq_ready = deqAllocate_17;
  assign sourceLane_17 = 32'h1 << _readCrossBar_output_17_bits_writeIndex;
  assign readMessageQueue_17_enq_bits_readSource = sourceLane_17;
  wire               readChannel_17_valid_0 = maskDestinationType ? _maskedWrite_readChannel_17_valid : _readCrossBar_output_17_valid & readMessageQueue_17_enq_ready;
  wire [4:0]         readChannel_17_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_17_bits_vs : _readCrossBar_output_17_bits_vs;
  wire               readChannel_17_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_17_bits_offset : _readCrossBar_output_17_bits_offset;
  assign readMessageQueue_17_enq_valid = readChannel_17_ready_0 & readChannel_17_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_17_enq_bits_data = readResult_17_bits >> {27'h0, readMessageQueue_17_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_17 = _write1HPipe_17_T & ~maskDestinationType ? reorderQueueVec_17_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_18;
  wire               readMessageQueue_18_deq_valid;
  assign readMessageQueue_18_deq_valid = ~_readMessageQueue_fifo_18_empty;
  wire [31:0]        readMessageQueue_dataOut_18_readSource;
  assign reorderQueueVec_18_enq_bits_write1H = readMessageQueue_18_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_18_dataOffset;
  wire [31:0]        readMessageQueue_18_enq_bits_readSource;
  wire [1:0]         readMessageQueue_18_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_18 = {readMessageQueue_18_enq_bits_readSource, readMessageQueue_18_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_18_dataOffset = _readMessageQueue_fifo_18_data_out[1:0];
  assign readMessageQueue_dataOut_18_readSource = _readMessageQueue_fifo_18_data_out[33:2];
  assign readMessageQueue_18_deq_bits_readSource = readMessageQueue_dataOut_18_readSource;
  wire [1:0]         readMessageQueue_18_deq_bits_dataOffset = readMessageQueue_dataOut_18_dataOffset;
  wire               readMessageQueue_18_enq_ready = ~_readMessageQueue_fifo_18_full;
  wire               readMessageQueue_18_enq_valid;
  assign deqAllocate_18 = ~readValid | reorderStageValid & reorderStageState_18 != reorderStageNeed_18;
  assign reorderQueueVec_18_deq_ready = deqAllocate_18;
  assign sourceLane_18 = 32'h1 << _readCrossBar_output_18_bits_writeIndex;
  assign readMessageQueue_18_enq_bits_readSource = sourceLane_18;
  wire               readChannel_18_valid_0 = maskDestinationType ? _maskedWrite_readChannel_18_valid : _readCrossBar_output_18_valid & readMessageQueue_18_enq_ready;
  wire [4:0]         readChannel_18_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_18_bits_vs : _readCrossBar_output_18_bits_vs;
  wire               readChannel_18_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_18_bits_offset : _readCrossBar_output_18_bits_offset;
  assign readMessageQueue_18_enq_valid = readChannel_18_ready_0 & readChannel_18_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_18_enq_bits_data = readResult_18_bits >> {27'h0, readMessageQueue_18_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_18 = _write1HPipe_18_T & ~maskDestinationType ? reorderQueueVec_18_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_19;
  wire               readMessageQueue_19_deq_valid;
  assign readMessageQueue_19_deq_valid = ~_readMessageQueue_fifo_19_empty;
  wire [31:0]        readMessageQueue_dataOut_19_readSource;
  assign reorderQueueVec_19_enq_bits_write1H = readMessageQueue_19_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_19_dataOffset;
  wire [31:0]        readMessageQueue_19_enq_bits_readSource;
  wire [1:0]         readMessageQueue_19_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_19 = {readMessageQueue_19_enq_bits_readSource, readMessageQueue_19_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_19_dataOffset = _readMessageQueue_fifo_19_data_out[1:0];
  assign readMessageQueue_dataOut_19_readSource = _readMessageQueue_fifo_19_data_out[33:2];
  assign readMessageQueue_19_deq_bits_readSource = readMessageQueue_dataOut_19_readSource;
  wire [1:0]         readMessageQueue_19_deq_bits_dataOffset = readMessageQueue_dataOut_19_dataOffset;
  wire               readMessageQueue_19_enq_ready = ~_readMessageQueue_fifo_19_full;
  wire               readMessageQueue_19_enq_valid;
  assign deqAllocate_19 = ~readValid | reorderStageValid & reorderStageState_19 != reorderStageNeed_19;
  assign reorderQueueVec_19_deq_ready = deqAllocate_19;
  assign sourceLane_19 = 32'h1 << _readCrossBar_output_19_bits_writeIndex;
  assign readMessageQueue_19_enq_bits_readSource = sourceLane_19;
  wire               readChannel_19_valid_0 = maskDestinationType ? _maskedWrite_readChannel_19_valid : _readCrossBar_output_19_valid & readMessageQueue_19_enq_ready;
  wire [4:0]         readChannel_19_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_19_bits_vs : _readCrossBar_output_19_bits_vs;
  wire               readChannel_19_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_19_bits_offset : _readCrossBar_output_19_bits_offset;
  assign readMessageQueue_19_enq_valid = readChannel_19_ready_0 & readChannel_19_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_19_enq_bits_data = readResult_19_bits >> {27'h0, readMessageQueue_19_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_19 = _write1HPipe_19_T & ~maskDestinationType ? reorderQueueVec_19_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_20;
  wire               readMessageQueue_20_deq_valid;
  assign readMessageQueue_20_deq_valid = ~_readMessageQueue_fifo_20_empty;
  wire [31:0]        readMessageQueue_dataOut_20_readSource;
  assign reorderQueueVec_20_enq_bits_write1H = readMessageQueue_20_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_20_dataOffset;
  wire [31:0]        readMessageQueue_20_enq_bits_readSource;
  wire [1:0]         readMessageQueue_20_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_20 = {readMessageQueue_20_enq_bits_readSource, readMessageQueue_20_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_20_dataOffset = _readMessageQueue_fifo_20_data_out[1:0];
  assign readMessageQueue_dataOut_20_readSource = _readMessageQueue_fifo_20_data_out[33:2];
  assign readMessageQueue_20_deq_bits_readSource = readMessageQueue_dataOut_20_readSource;
  wire [1:0]         readMessageQueue_20_deq_bits_dataOffset = readMessageQueue_dataOut_20_dataOffset;
  wire               readMessageQueue_20_enq_ready = ~_readMessageQueue_fifo_20_full;
  wire               readMessageQueue_20_enq_valid;
  assign deqAllocate_20 = ~readValid | reorderStageValid & reorderStageState_20 != reorderStageNeed_20;
  assign reorderQueueVec_20_deq_ready = deqAllocate_20;
  assign sourceLane_20 = 32'h1 << _readCrossBar_output_20_bits_writeIndex;
  assign readMessageQueue_20_enq_bits_readSource = sourceLane_20;
  wire               readChannel_20_valid_0 = maskDestinationType ? _maskedWrite_readChannel_20_valid : _readCrossBar_output_20_valid & readMessageQueue_20_enq_ready;
  wire [4:0]         readChannel_20_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_20_bits_vs : _readCrossBar_output_20_bits_vs;
  wire               readChannel_20_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_20_bits_offset : _readCrossBar_output_20_bits_offset;
  assign readMessageQueue_20_enq_valid = readChannel_20_ready_0 & readChannel_20_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_20_enq_bits_data = readResult_20_bits >> {27'h0, readMessageQueue_20_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_20 = _write1HPipe_20_T & ~maskDestinationType ? reorderQueueVec_20_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_21;
  wire               readMessageQueue_21_deq_valid;
  assign readMessageQueue_21_deq_valid = ~_readMessageQueue_fifo_21_empty;
  wire [31:0]        readMessageQueue_dataOut_21_readSource;
  assign reorderQueueVec_21_enq_bits_write1H = readMessageQueue_21_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_21_dataOffset;
  wire [31:0]        readMessageQueue_21_enq_bits_readSource;
  wire [1:0]         readMessageQueue_21_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_21 = {readMessageQueue_21_enq_bits_readSource, readMessageQueue_21_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_21_dataOffset = _readMessageQueue_fifo_21_data_out[1:0];
  assign readMessageQueue_dataOut_21_readSource = _readMessageQueue_fifo_21_data_out[33:2];
  assign readMessageQueue_21_deq_bits_readSource = readMessageQueue_dataOut_21_readSource;
  wire [1:0]         readMessageQueue_21_deq_bits_dataOffset = readMessageQueue_dataOut_21_dataOffset;
  wire               readMessageQueue_21_enq_ready = ~_readMessageQueue_fifo_21_full;
  wire               readMessageQueue_21_enq_valid;
  assign deqAllocate_21 = ~readValid | reorderStageValid & reorderStageState_21 != reorderStageNeed_21;
  assign reorderQueueVec_21_deq_ready = deqAllocate_21;
  assign sourceLane_21 = 32'h1 << _readCrossBar_output_21_bits_writeIndex;
  assign readMessageQueue_21_enq_bits_readSource = sourceLane_21;
  wire               readChannel_21_valid_0 = maskDestinationType ? _maskedWrite_readChannel_21_valid : _readCrossBar_output_21_valid & readMessageQueue_21_enq_ready;
  wire [4:0]         readChannel_21_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_21_bits_vs : _readCrossBar_output_21_bits_vs;
  wire               readChannel_21_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_21_bits_offset : _readCrossBar_output_21_bits_offset;
  assign readMessageQueue_21_enq_valid = readChannel_21_ready_0 & readChannel_21_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_21_enq_bits_data = readResult_21_bits >> {27'h0, readMessageQueue_21_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_21 = _write1HPipe_21_T & ~maskDestinationType ? reorderQueueVec_21_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_22;
  wire               readMessageQueue_22_deq_valid;
  assign readMessageQueue_22_deq_valid = ~_readMessageQueue_fifo_22_empty;
  wire [31:0]        readMessageQueue_dataOut_22_readSource;
  assign reorderQueueVec_22_enq_bits_write1H = readMessageQueue_22_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_22_dataOffset;
  wire [31:0]        readMessageQueue_22_enq_bits_readSource;
  wire [1:0]         readMessageQueue_22_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_22 = {readMessageQueue_22_enq_bits_readSource, readMessageQueue_22_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_22_dataOffset = _readMessageQueue_fifo_22_data_out[1:0];
  assign readMessageQueue_dataOut_22_readSource = _readMessageQueue_fifo_22_data_out[33:2];
  assign readMessageQueue_22_deq_bits_readSource = readMessageQueue_dataOut_22_readSource;
  wire [1:0]         readMessageQueue_22_deq_bits_dataOffset = readMessageQueue_dataOut_22_dataOffset;
  wire               readMessageQueue_22_enq_ready = ~_readMessageQueue_fifo_22_full;
  wire               readMessageQueue_22_enq_valid;
  assign deqAllocate_22 = ~readValid | reorderStageValid & reorderStageState_22 != reorderStageNeed_22;
  assign reorderQueueVec_22_deq_ready = deqAllocate_22;
  assign sourceLane_22 = 32'h1 << _readCrossBar_output_22_bits_writeIndex;
  assign readMessageQueue_22_enq_bits_readSource = sourceLane_22;
  wire               readChannel_22_valid_0 = maskDestinationType ? _maskedWrite_readChannel_22_valid : _readCrossBar_output_22_valid & readMessageQueue_22_enq_ready;
  wire [4:0]         readChannel_22_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_22_bits_vs : _readCrossBar_output_22_bits_vs;
  wire               readChannel_22_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_22_bits_offset : _readCrossBar_output_22_bits_offset;
  assign readMessageQueue_22_enq_valid = readChannel_22_ready_0 & readChannel_22_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_22_enq_bits_data = readResult_22_bits >> {27'h0, readMessageQueue_22_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_22 = _write1HPipe_22_T & ~maskDestinationType ? reorderQueueVec_22_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_23;
  wire               readMessageQueue_23_deq_valid;
  assign readMessageQueue_23_deq_valid = ~_readMessageQueue_fifo_23_empty;
  wire [31:0]        readMessageQueue_dataOut_23_readSource;
  assign reorderQueueVec_23_enq_bits_write1H = readMessageQueue_23_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_23_dataOffset;
  wire [31:0]        readMessageQueue_23_enq_bits_readSource;
  wire [1:0]         readMessageQueue_23_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_23 = {readMessageQueue_23_enq_bits_readSource, readMessageQueue_23_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_23_dataOffset = _readMessageQueue_fifo_23_data_out[1:0];
  assign readMessageQueue_dataOut_23_readSource = _readMessageQueue_fifo_23_data_out[33:2];
  assign readMessageQueue_23_deq_bits_readSource = readMessageQueue_dataOut_23_readSource;
  wire [1:0]         readMessageQueue_23_deq_bits_dataOffset = readMessageQueue_dataOut_23_dataOffset;
  wire               readMessageQueue_23_enq_ready = ~_readMessageQueue_fifo_23_full;
  wire               readMessageQueue_23_enq_valid;
  assign deqAllocate_23 = ~readValid | reorderStageValid & reorderStageState_23 != reorderStageNeed_23;
  assign reorderQueueVec_23_deq_ready = deqAllocate_23;
  assign sourceLane_23 = 32'h1 << _readCrossBar_output_23_bits_writeIndex;
  assign readMessageQueue_23_enq_bits_readSource = sourceLane_23;
  wire               readChannel_23_valid_0 = maskDestinationType ? _maskedWrite_readChannel_23_valid : _readCrossBar_output_23_valid & readMessageQueue_23_enq_ready;
  wire [4:0]         readChannel_23_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_23_bits_vs : _readCrossBar_output_23_bits_vs;
  wire               readChannel_23_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_23_bits_offset : _readCrossBar_output_23_bits_offset;
  assign readMessageQueue_23_enq_valid = readChannel_23_ready_0 & readChannel_23_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_23_enq_bits_data = readResult_23_bits >> {27'h0, readMessageQueue_23_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_23 = _write1HPipe_23_T & ~maskDestinationType ? reorderQueueVec_23_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_24;
  wire               readMessageQueue_24_deq_valid;
  assign readMessageQueue_24_deq_valid = ~_readMessageQueue_fifo_24_empty;
  wire [31:0]        readMessageQueue_dataOut_24_readSource;
  assign reorderQueueVec_24_enq_bits_write1H = readMessageQueue_24_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_24_dataOffset;
  wire [31:0]        readMessageQueue_24_enq_bits_readSource;
  wire [1:0]         readMessageQueue_24_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_24 = {readMessageQueue_24_enq_bits_readSource, readMessageQueue_24_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_24_dataOffset = _readMessageQueue_fifo_24_data_out[1:0];
  assign readMessageQueue_dataOut_24_readSource = _readMessageQueue_fifo_24_data_out[33:2];
  assign readMessageQueue_24_deq_bits_readSource = readMessageQueue_dataOut_24_readSource;
  wire [1:0]         readMessageQueue_24_deq_bits_dataOffset = readMessageQueue_dataOut_24_dataOffset;
  wire               readMessageQueue_24_enq_ready = ~_readMessageQueue_fifo_24_full;
  wire               readMessageQueue_24_enq_valid;
  assign deqAllocate_24 = ~readValid | reorderStageValid & reorderStageState_24 != reorderStageNeed_24;
  assign reorderQueueVec_24_deq_ready = deqAllocate_24;
  assign sourceLane_24 = 32'h1 << _readCrossBar_output_24_bits_writeIndex;
  assign readMessageQueue_24_enq_bits_readSource = sourceLane_24;
  wire               readChannel_24_valid_0 = maskDestinationType ? _maskedWrite_readChannel_24_valid : _readCrossBar_output_24_valid & readMessageQueue_24_enq_ready;
  wire [4:0]         readChannel_24_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_24_bits_vs : _readCrossBar_output_24_bits_vs;
  wire               readChannel_24_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_24_bits_offset : _readCrossBar_output_24_bits_offset;
  assign readMessageQueue_24_enq_valid = readChannel_24_ready_0 & readChannel_24_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_24_enq_bits_data = readResult_24_bits >> {27'h0, readMessageQueue_24_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_24 = _write1HPipe_24_T & ~maskDestinationType ? reorderQueueVec_24_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_25;
  wire               readMessageQueue_25_deq_valid;
  assign readMessageQueue_25_deq_valid = ~_readMessageQueue_fifo_25_empty;
  wire [31:0]        readMessageQueue_dataOut_25_readSource;
  assign reorderQueueVec_25_enq_bits_write1H = readMessageQueue_25_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_25_dataOffset;
  wire [31:0]        readMessageQueue_25_enq_bits_readSource;
  wire [1:0]         readMessageQueue_25_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_25 = {readMessageQueue_25_enq_bits_readSource, readMessageQueue_25_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_25_dataOffset = _readMessageQueue_fifo_25_data_out[1:0];
  assign readMessageQueue_dataOut_25_readSource = _readMessageQueue_fifo_25_data_out[33:2];
  assign readMessageQueue_25_deq_bits_readSource = readMessageQueue_dataOut_25_readSource;
  wire [1:0]         readMessageQueue_25_deq_bits_dataOffset = readMessageQueue_dataOut_25_dataOffset;
  wire               readMessageQueue_25_enq_ready = ~_readMessageQueue_fifo_25_full;
  wire               readMessageQueue_25_enq_valid;
  assign deqAllocate_25 = ~readValid | reorderStageValid & reorderStageState_25 != reorderStageNeed_25;
  assign reorderQueueVec_25_deq_ready = deqAllocate_25;
  assign sourceLane_25 = 32'h1 << _readCrossBar_output_25_bits_writeIndex;
  assign readMessageQueue_25_enq_bits_readSource = sourceLane_25;
  wire               readChannel_25_valid_0 = maskDestinationType ? _maskedWrite_readChannel_25_valid : _readCrossBar_output_25_valid & readMessageQueue_25_enq_ready;
  wire [4:0]         readChannel_25_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_25_bits_vs : _readCrossBar_output_25_bits_vs;
  wire               readChannel_25_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_25_bits_offset : _readCrossBar_output_25_bits_offset;
  assign readMessageQueue_25_enq_valid = readChannel_25_ready_0 & readChannel_25_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_25_enq_bits_data = readResult_25_bits >> {27'h0, readMessageQueue_25_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_25 = _write1HPipe_25_T & ~maskDestinationType ? reorderQueueVec_25_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_26;
  wire               readMessageQueue_26_deq_valid;
  assign readMessageQueue_26_deq_valid = ~_readMessageQueue_fifo_26_empty;
  wire [31:0]        readMessageQueue_dataOut_26_readSource;
  assign reorderQueueVec_26_enq_bits_write1H = readMessageQueue_26_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_26_dataOffset;
  wire [31:0]        readMessageQueue_26_enq_bits_readSource;
  wire [1:0]         readMessageQueue_26_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_26 = {readMessageQueue_26_enq_bits_readSource, readMessageQueue_26_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_26_dataOffset = _readMessageQueue_fifo_26_data_out[1:0];
  assign readMessageQueue_dataOut_26_readSource = _readMessageQueue_fifo_26_data_out[33:2];
  assign readMessageQueue_26_deq_bits_readSource = readMessageQueue_dataOut_26_readSource;
  wire [1:0]         readMessageQueue_26_deq_bits_dataOffset = readMessageQueue_dataOut_26_dataOffset;
  wire               readMessageQueue_26_enq_ready = ~_readMessageQueue_fifo_26_full;
  wire               readMessageQueue_26_enq_valid;
  assign deqAllocate_26 = ~readValid | reorderStageValid & reorderStageState_26 != reorderStageNeed_26;
  assign reorderQueueVec_26_deq_ready = deqAllocate_26;
  assign sourceLane_26 = 32'h1 << _readCrossBar_output_26_bits_writeIndex;
  assign readMessageQueue_26_enq_bits_readSource = sourceLane_26;
  wire               readChannel_26_valid_0 = maskDestinationType ? _maskedWrite_readChannel_26_valid : _readCrossBar_output_26_valid & readMessageQueue_26_enq_ready;
  wire [4:0]         readChannel_26_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_26_bits_vs : _readCrossBar_output_26_bits_vs;
  wire               readChannel_26_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_26_bits_offset : _readCrossBar_output_26_bits_offset;
  assign readMessageQueue_26_enq_valid = readChannel_26_ready_0 & readChannel_26_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_26_enq_bits_data = readResult_26_bits >> {27'h0, readMessageQueue_26_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_26 = _write1HPipe_26_T & ~maskDestinationType ? reorderQueueVec_26_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_27;
  wire               readMessageQueue_27_deq_valid;
  assign readMessageQueue_27_deq_valid = ~_readMessageQueue_fifo_27_empty;
  wire [31:0]        readMessageQueue_dataOut_27_readSource;
  assign reorderQueueVec_27_enq_bits_write1H = readMessageQueue_27_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_27_dataOffset;
  wire [31:0]        readMessageQueue_27_enq_bits_readSource;
  wire [1:0]         readMessageQueue_27_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_27 = {readMessageQueue_27_enq_bits_readSource, readMessageQueue_27_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_27_dataOffset = _readMessageQueue_fifo_27_data_out[1:0];
  assign readMessageQueue_dataOut_27_readSource = _readMessageQueue_fifo_27_data_out[33:2];
  assign readMessageQueue_27_deq_bits_readSource = readMessageQueue_dataOut_27_readSource;
  wire [1:0]         readMessageQueue_27_deq_bits_dataOffset = readMessageQueue_dataOut_27_dataOffset;
  wire               readMessageQueue_27_enq_ready = ~_readMessageQueue_fifo_27_full;
  wire               readMessageQueue_27_enq_valid;
  assign deqAllocate_27 = ~readValid | reorderStageValid & reorderStageState_27 != reorderStageNeed_27;
  assign reorderQueueVec_27_deq_ready = deqAllocate_27;
  assign sourceLane_27 = 32'h1 << _readCrossBar_output_27_bits_writeIndex;
  assign readMessageQueue_27_enq_bits_readSource = sourceLane_27;
  wire               readChannel_27_valid_0 = maskDestinationType ? _maskedWrite_readChannel_27_valid : _readCrossBar_output_27_valid & readMessageQueue_27_enq_ready;
  wire [4:0]         readChannel_27_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_27_bits_vs : _readCrossBar_output_27_bits_vs;
  wire               readChannel_27_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_27_bits_offset : _readCrossBar_output_27_bits_offset;
  assign readMessageQueue_27_enq_valid = readChannel_27_ready_0 & readChannel_27_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_27_enq_bits_data = readResult_27_bits >> {27'h0, readMessageQueue_27_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_27 = _write1HPipe_27_T & ~maskDestinationType ? reorderQueueVec_27_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_28;
  wire               readMessageQueue_28_deq_valid;
  assign readMessageQueue_28_deq_valid = ~_readMessageQueue_fifo_28_empty;
  wire [31:0]        readMessageQueue_dataOut_28_readSource;
  assign reorderQueueVec_28_enq_bits_write1H = readMessageQueue_28_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_28_dataOffset;
  wire [31:0]        readMessageQueue_28_enq_bits_readSource;
  wire [1:0]         readMessageQueue_28_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_28 = {readMessageQueue_28_enq_bits_readSource, readMessageQueue_28_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_28_dataOffset = _readMessageQueue_fifo_28_data_out[1:0];
  assign readMessageQueue_dataOut_28_readSource = _readMessageQueue_fifo_28_data_out[33:2];
  assign readMessageQueue_28_deq_bits_readSource = readMessageQueue_dataOut_28_readSource;
  wire [1:0]         readMessageQueue_28_deq_bits_dataOffset = readMessageQueue_dataOut_28_dataOffset;
  wire               readMessageQueue_28_enq_ready = ~_readMessageQueue_fifo_28_full;
  wire               readMessageQueue_28_enq_valid;
  assign deqAllocate_28 = ~readValid | reorderStageValid & reorderStageState_28 != reorderStageNeed_28;
  assign reorderQueueVec_28_deq_ready = deqAllocate_28;
  assign sourceLane_28 = 32'h1 << _readCrossBar_output_28_bits_writeIndex;
  assign readMessageQueue_28_enq_bits_readSource = sourceLane_28;
  wire               readChannel_28_valid_0 = maskDestinationType ? _maskedWrite_readChannel_28_valid : _readCrossBar_output_28_valid & readMessageQueue_28_enq_ready;
  wire [4:0]         readChannel_28_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_28_bits_vs : _readCrossBar_output_28_bits_vs;
  wire               readChannel_28_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_28_bits_offset : _readCrossBar_output_28_bits_offset;
  assign readMessageQueue_28_enq_valid = readChannel_28_ready_0 & readChannel_28_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_28_enq_bits_data = readResult_28_bits >> {27'h0, readMessageQueue_28_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_28 = _write1HPipe_28_T & ~maskDestinationType ? reorderQueueVec_28_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_29;
  wire               readMessageQueue_29_deq_valid;
  assign readMessageQueue_29_deq_valid = ~_readMessageQueue_fifo_29_empty;
  wire [31:0]        readMessageQueue_dataOut_29_readSource;
  assign reorderQueueVec_29_enq_bits_write1H = readMessageQueue_29_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_29_dataOffset;
  wire [31:0]        readMessageQueue_29_enq_bits_readSource;
  wire [1:0]         readMessageQueue_29_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_29 = {readMessageQueue_29_enq_bits_readSource, readMessageQueue_29_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_29_dataOffset = _readMessageQueue_fifo_29_data_out[1:0];
  assign readMessageQueue_dataOut_29_readSource = _readMessageQueue_fifo_29_data_out[33:2];
  assign readMessageQueue_29_deq_bits_readSource = readMessageQueue_dataOut_29_readSource;
  wire [1:0]         readMessageQueue_29_deq_bits_dataOffset = readMessageQueue_dataOut_29_dataOffset;
  wire               readMessageQueue_29_enq_ready = ~_readMessageQueue_fifo_29_full;
  wire               readMessageQueue_29_enq_valid;
  assign deqAllocate_29 = ~readValid | reorderStageValid & reorderStageState_29 != reorderStageNeed_29;
  assign reorderQueueVec_29_deq_ready = deqAllocate_29;
  assign sourceLane_29 = 32'h1 << _readCrossBar_output_29_bits_writeIndex;
  assign readMessageQueue_29_enq_bits_readSource = sourceLane_29;
  wire               readChannel_29_valid_0 = maskDestinationType ? _maskedWrite_readChannel_29_valid : _readCrossBar_output_29_valid & readMessageQueue_29_enq_ready;
  wire [4:0]         readChannel_29_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_29_bits_vs : _readCrossBar_output_29_bits_vs;
  wire               readChannel_29_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_29_bits_offset : _readCrossBar_output_29_bits_offset;
  assign readMessageQueue_29_enq_valid = readChannel_29_ready_0 & readChannel_29_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_29_enq_bits_data = readResult_29_bits >> {27'h0, readMessageQueue_29_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_29 = _write1HPipe_29_T & ~maskDestinationType ? reorderQueueVec_29_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_30;
  wire               readMessageQueue_30_deq_valid;
  assign readMessageQueue_30_deq_valid = ~_readMessageQueue_fifo_30_empty;
  wire [31:0]        readMessageQueue_dataOut_30_readSource;
  assign reorderQueueVec_30_enq_bits_write1H = readMessageQueue_30_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_30_dataOffset;
  wire [31:0]        readMessageQueue_30_enq_bits_readSource;
  wire [1:0]         readMessageQueue_30_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_30 = {readMessageQueue_30_enq_bits_readSource, readMessageQueue_30_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_30_dataOffset = _readMessageQueue_fifo_30_data_out[1:0];
  assign readMessageQueue_dataOut_30_readSource = _readMessageQueue_fifo_30_data_out[33:2];
  assign readMessageQueue_30_deq_bits_readSource = readMessageQueue_dataOut_30_readSource;
  wire [1:0]         readMessageQueue_30_deq_bits_dataOffset = readMessageQueue_dataOut_30_dataOffset;
  wire               readMessageQueue_30_enq_ready = ~_readMessageQueue_fifo_30_full;
  wire               readMessageQueue_30_enq_valid;
  assign deqAllocate_30 = ~readValid | reorderStageValid & reorderStageState_30 != reorderStageNeed_30;
  assign reorderQueueVec_30_deq_ready = deqAllocate_30;
  assign sourceLane_30 = 32'h1 << _readCrossBar_output_30_bits_writeIndex;
  assign readMessageQueue_30_enq_bits_readSource = sourceLane_30;
  wire               readChannel_30_valid_0 = maskDestinationType ? _maskedWrite_readChannel_30_valid : _readCrossBar_output_30_valid & readMessageQueue_30_enq_ready;
  wire [4:0]         readChannel_30_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_30_bits_vs : _readCrossBar_output_30_bits_vs;
  wire               readChannel_30_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_30_bits_offset : _readCrossBar_output_30_bits_offset;
  assign readMessageQueue_30_enq_valid = readChannel_30_ready_0 & readChannel_30_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_30_enq_bits_data = readResult_30_bits >> {27'h0, readMessageQueue_30_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_30 = _write1HPipe_30_T & ~maskDestinationType ? reorderQueueVec_30_deq_bits_write1H : 32'h0;
  wire [31:0]        sourceLane_31;
  wire               readMessageQueue_31_deq_valid;
  assign readMessageQueue_31_deq_valid = ~_readMessageQueue_fifo_31_empty;
  wire [31:0]        readMessageQueue_dataOut_31_readSource;
  assign reorderQueueVec_31_enq_bits_write1H = readMessageQueue_31_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_31_dataOffset;
  wire [31:0]        readMessageQueue_31_enq_bits_readSource;
  wire [1:0]         readMessageQueue_31_enq_bits_dataOffset;
  wire [33:0]        readMessageQueue_dataIn_31 = {readMessageQueue_31_enq_bits_readSource, readMessageQueue_31_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_31_dataOffset = _readMessageQueue_fifo_31_data_out[1:0];
  assign readMessageQueue_dataOut_31_readSource = _readMessageQueue_fifo_31_data_out[33:2];
  assign readMessageQueue_31_deq_bits_readSource = readMessageQueue_dataOut_31_readSource;
  wire [1:0]         readMessageQueue_31_deq_bits_dataOffset = readMessageQueue_dataOut_31_dataOffset;
  wire               readMessageQueue_31_enq_ready = ~_readMessageQueue_fifo_31_full;
  wire               readMessageQueue_31_enq_valid;
  assign deqAllocate_31 = ~readValid | reorderStageValid & reorderStageState_31 != reorderStageNeed_31;
  assign reorderQueueVec_31_deq_ready = deqAllocate_31;
  assign sourceLane_31 = 32'h1 << _readCrossBar_output_31_bits_writeIndex;
  assign readMessageQueue_31_enq_bits_readSource = sourceLane_31;
  wire               readChannel_31_valid_0 = maskDestinationType ? _maskedWrite_readChannel_31_valid : _readCrossBar_output_31_valid & readMessageQueue_31_enq_ready;
  wire [4:0]         readChannel_31_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_31_bits_vs : _readCrossBar_output_31_bits_vs;
  wire               readChannel_31_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_31_bits_offset : _readCrossBar_output_31_bits_offset;
  assign readMessageQueue_31_enq_valid = readChannel_31_ready_0 & readChannel_31_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_31_enq_bits_data = readResult_31_bits >> {27'h0, readMessageQueue_31_deq_bits_dataOffset, 3'h0};
  wire [31:0]        write1HPipe_31 = _write1HPipe_31_T & ~maskDestinationType ? reorderQueueVec_31_deq_bits_write1H : 32'h0;
  wire [31:0]        readData_data;
  wire               readData_readDataQueue_enq_ready = ~_readData_readDataQueue_fifo_full;
  wire               readData_readDataQueue_deq_ready;
  wire               readData_readDataQueue_enq_valid;
  wire               readData_readDataQueue_deq_valid = ~_readData_readDataQueue_fifo_empty | readData_readDataQueue_enq_valid;
  wire [31:0]        readData_readDataQueue_enq_bits;
  wire [31:0]        readData_readDataQueue_deq_bits = _readData_readDataQueue_fifo_empty ? readData_readDataQueue_enq_bits : _readData_readDataQueue_fifo_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo = {write1HPipe_1[0], write1HPipe_0[0]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi = {write1HPipe_3[0], write1HPipe_2[0]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo = {readData_readResultSelect_lo_lo_lo_hi, readData_readResultSelect_lo_lo_lo_lo};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo = {write1HPipe_5[0], write1HPipe_4[0]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi = {write1HPipe_7[0], write1HPipe_6[0]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi = {readData_readResultSelect_lo_lo_hi_hi, readData_readResultSelect_lo_lo_hi_lo};
  wire [7:0]         readData_readResultSelect_lo_lo = {readData_readResultSelect_lo_lo_hi, readData_readResultSelect_lo_lo_lo};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo = {write1HPipe_9[0], write1HPipe_8[0]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi = {write1HPipe_11[0], write1HPipe_10[0]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo = {readData_readResultSelect_lo_hi_lo_hi, readData_readResultSelect_lo_hi_lo_lo};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo = {write1HPipe_13[0], write1HPipe_12[0]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi = {write1HPipe_15[0], write1HPipe_14[0]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi = {readData_readResultSelect_lo_hi_hi_hi, readData_readResultSelect_lo_hi_hi_lo};
  wire [7:0]         readData_readResultSelect_lo_hi = {readData_readResultSelect_lo_hi_hi, readData_readResultSelect_lo_hi_lo};
  wire [15:0]        readData_readResultSelect_lo = {readData_readResultSelect_lo_hi, readData_readResultSelect_lo_lo};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo = {write1HPipe_17[0], write1HPipe_16[0]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi = {write1HPipe_19[0], write1HPipe_18[0]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo = {readData_readResultSelect_hi_lo_lo_hi, readData_readResultSelect_hi_lo_lo_lo};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo = {write1HPipe_21[0], write1HPipe_20[0]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi = {write1HPipe_23[0], write1HPipe_22[0]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi = {readData_readResultSelect_hi_lo_hi_hi, readData_readResultSelect_hi_lo_hi_lo};
  wire [7:0]         readData_readResultSelect_hi_lo = {readData_readResultSelect_hi_lo_hi, readData_readResultSelect_hi_lo_lo};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo = {write1HPipe_25[0], write1HPipe_24[0]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi = {write1HPipe_27[0], write1HPipe_26[0]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo = {readData_readResultSelect_hi_hi_lo_hi, readData_readResultSelect_hi_hi_lo_lo};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo = {write1HPipe_29[0], write1HPipe_28[0]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi = {write1HPipe_31[0], write1HPipe_30[0]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi = {readData_readResultSelect_hi_hi_hi_hi, readData_readResultSelect_hi_hi_hi_lo};
  wire [7:0]         readData_readResultSelect_hi_hi = {readData_readResultSelect_hi_hi_hi, readData_readResultSelect_hi_hi_lo};
  wire [15:0]        readData_readResultSelect_hi = {readData_readResultSelect_hi_hi, readData_readResultSelect_hi_lo};
  wire [31:0]        readData_readResultSelect = {readData_readResultSelect_hi, readData_readResultSelect_lo};
  assign readData_data =
    (readData_readResultSelect[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_enq_bits = readData_data;
  wire               readTokenRelease_0 = readData_readDataQueue_deq_ready & readData_readDataQueue_deq_valid;
  assign readData_readDataQueue_enq_valid = |readData_readResultSelect;
  wire [31:0]        readData_data_1;
  wire               isWaiteForThisData_1;
  wire               readData_readDataQueue_1_enq_ready = ~_readData_readDataQueue_fifo_1_full;
  wire               readData_readDataQueue_1_deq_ready;
  wire               readData_readDataQueue_1_enq_valid;
  wire               readData_readDataQueue_1_deq_valid = ~_readData_readDataQueue_fifo_1_empty | readData_readDataQueue_1_enq_valid;
  wire [31:0]        readData_readDataQueue_1_enq_bits;
  wire [31:0]        readData_readDataQueue_1_deq_bits = _readData_readDataQueue_fifo_1_empty ? readData_readDataQueue_1_enq_bits : _readData_readDataQueue_fifo_1_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_1 = {write1HPipe_1[1], write1HPipe_0[1]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_1 = {write1HPipe_3[1], write1HPipe_2[1]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_1 = {readData_readResultSelect_lo_lo_lo_hi_1, readData_readResultSelect_lo_lo_lo_lo_1};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_1 = {write1HPipe_5[1], write1HPipe_4[1]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_1 = {write1HPipe_7[1], write1HPipe_6[1]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_1 = {readData_readResultSelect_lo_lo_hi_hi_1, readData_readResultSelect_lo_lo_hi_lo_1};
  wire [7:0]         readData_readResultSelect_lo_lo_1 = {readData_readResultSelect_lo_lo_hi_1, readData_readResultSelect_lo_lo_lo_1};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_1 = {write1HPipe_9[1], write1HPipe_8[1]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_1 = {write1HPipe_11[1], write1HPipe_10[1]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_1 = {readData_readResultSelect_lo_hi_lo_hi_1, readData_readResultSelect_lo_hi_lo_lo_1};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_1 = {write1HPipe_13[1], write1HPipe_12[1]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_1 = {write1HPipe_15[1], write1HPipe_14[1]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_1 = {readData_readResultSelect_lo_hi_hi_hi_1, readData_readResultSelect_lo_hi_hi_lo_1};
  wire [7:0]         readData_readResultSelect_lo_hi_1 = {readData_readResultSelect_lo_hi_hi_1, readData_readResultSelect_lo_hi_lo_1};
  wire [15:0]        readData_readResultSelect_lo_1 = {readData_readResultSelect_lo_hi_1, readData_readResultSelect_lo_lo_1};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_1 = {write1HPipe_17[1], write1HPipe_16[1]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_1 = {write1HPipe_19[1], write1HPipe_18[1]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_1 = {readData_readResultSelect_hi_lo_lo_hi_1, readData_readResultSelect_hi_lo_lo_lo_1};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_1 = {write1HPipe_21[1], write1HPipe_20[1]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_1 = {write1HPipe_23[1], write1HPipe_22[1]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_1 = {readData_readResultSelect_hi_lo_hi_hi_1, readData_readResultSelect_hi_lo_hi_lo_1};
  wire [7:0]         readData_readResultSelect_hi_lo_1 = {readData_readResultSelect_hi_lo_hi_1, readData_readResultSelect_hi_lo_lo_1};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_1 = {write1HPipe_25[1], write1HPipe_24[1]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_1 = {write1HPipe_27[1], write1HPipe_26[1]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_1 = {readData_readResultSelect_hi_hi_lo_hi_1, readData_readResultSelect_hi_hi_lo_lo_1};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_1 = {write1HPipe_29[1], write1HPipe_28[1]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_1 = {write1HPipe_31[1], write1HPipe_30[1]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_1 = {readData_readResultSelect_hi_hi_hi_hi_1, readData_readResultSelect_hi_hi_hi_lo_1};
  wire [7:0]         readData_readResultSelect_hi_hi_1 = {readData_readResultSelect_hi_hi_hi_1, readData_readResultSelect_hi_hi_lo_1};
  wire [15:0]        readData_readResultSelect_hi_1 = {readData_readResultSelect_hi_hi_1, readData_readResultSelect_hi_lo_1};
  wire [31:0]        readData_readResultSelect_1 = {readData_readResultSelect_hi_1, readData_readResultSelect_lo_1};
  assign readData_data_1 =
    (readData_readResultSelect_1[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_1[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_1[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_1[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_1[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_1[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_1[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_1[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_1[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_1[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_1[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_1[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_1[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_1[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_1[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_1[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_1[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_1[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_1[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_1[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_1[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_1[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_1[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_1[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_1[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_1[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_1[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_1[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_1[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_1[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_1[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_1[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_1_enq_bits = readData_data_1;
  wire               readTokenRelease_1 = readData_readDataQueue_1_deq_ready & readData_readDataQueue_1_deq_valid;
  assign readData_readDataQueue_1_enq_valid = |readData_readResultSelect_1;
  wire [31:0]        readData_data_2;
  wire               isWaiteForThisData_2;
  wire               readData_readDataQueue_2_enq_ready = ~_readData_readDataQueue_fifo_2_full;
  wire               readData_readDataQueue_2_deq_ready;
  wire               readData_readDataQueue_2_enq_valid;
  wire               readData_readDataQueue_2_deq_valid = ~_readData_readDataQueue_fifo_2_empty | readData_readDataQueue_2_enq_valid;
  wire [31:0]        readData_readDataQueue_2_enq_bits;
  wire [31:0]        readData_readDataQueue_2_deq_bits = _readData_readDataQueue_fifo_2_empty ? readData_readDataQueue_2_enq_bits : _readData_readDataQueue_fifo_2_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_2 = {write1HPipe_1[2], write1HPipe_0[2]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_2 = {write1HPipe_3[2], write1HPipe_2[2]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_2 = {readData_readResultSelect_lo_lo_lo_hi_2, readData_readResultSelect_lo_lo_lo_lo_2};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_2 = {write1HPipe_5[2], write1HPipe_4[2]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_2 = {write1HPipe_7[2], write1HPipe_6[2]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_2 = {readData_readResultSelect_lo_lo_hi_hi_2, readData_readResultSelect_lo_lo_hi_lo_2};
  wire [7:0]         readData_readResultSelect_lo_lo_2 = {readData_readResultSelect_lo_lo_hi_2, readData_readResultSelect_lo_lo_lo_2};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_2 = {write1HPipe_9[2], write1HPipe_8[2]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_2 = {write1HPipe_11[2], write1HPipe_10[2]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_2 = {readData_readResultSelect_lo_hi_lo_hi_2, readData_readResultSelect_lo_hi_lo_lo_2};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_2 = {write1HPipe_13[2], write1HPipe_12[2]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_2 = {write1HPipe_15[2], write1HPipe_14[2]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_2 = {readData_readResultSelect_lo_hi_hi_hi_2, readData_readResultSelect_lo_hi_hi_lo_2};
  wire [7:0]         readData_readResultSelect_lo_hi_2 = {readData_readResultSelect_lo_hi_hi_2, readData_readResultSelect_lo_hi_lo_2};
  wire [15:0]        readData_readResultSelect_lo_2 = {readData_readResultSelect_lo_hi_2, readData_readResultSelect_lo_lo_2};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_2 = {write1HPipe_17[2], write1HPipe_16[2]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_2 = {write1HPipe_19[2], write1HPipe_18[2]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_2 = {readData_readResultSelect_hi_lo_lo_hi_2, readData_readResultSelect_hi_lo_lo_lo_2};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_2 = {write1HPipe_21[2], write1HPipe_20[2]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_2 = {write1HPipe_23[2], write1HPipe_22[2]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_2 = {readData_readResultSelect_hi_lo_hi_hi_2, readData_readResultSelect_hi_lo_hi_lo_2};
  wire [7:0]         readData_readResultSelect_hi_lo_2 = {readData_readResultSelect_hi_lo_hi_2, readData_readResultSelect_hi_lo_lo_2};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_2 = {write1HPipe_25[2], write1HPipe_24[2]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_2 = {write1HPipe_27[2], write1HPipe_26[2]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_2 = {readData_readResultSelect_hi_hi_lo_hi_2, readData_readResultSelect_hi_hi_lo_lo_2};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_2 = {write1HPipe_29[2], write1HPipe_28[2]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_2 = {write1HPipe_31[2], write1HPipe_30[2]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_2 = {readData_readResultSelect_hi_hi_hi_hi_2, readData_readResultSelect_hi_hi_hi_lo_2};
  wire [7:0]         readData_readResultSelect_hi_hi_2 = {readData_readResultSelect_hi_hi_hi_2, readData_readResultSelect_hi_hi_lo_2};
  wire [15:0]        readData_readResultSelect_hi_2 = {readData_readResultSelect_hi_hi_2, readData_readResultSelect_hi_lo_2};
  wire [31:0]        readData_readResultSelect_2 = {readData_readResultSelect_hi_2, readData_readResultSelect_lo_2};
  assign readData_data_2 =
    (readData_readResultSelect_2[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_2[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_2[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_2[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_2[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_2[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_2[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_2[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_2[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_2[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_2[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_2[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_2[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_2[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_2[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_2[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_2[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_2[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_2[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_2[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_2[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_2[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_2[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_2[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_2[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_2[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_2[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_2[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_2[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_2[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_2[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_2[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_2_enq_bits = readData_data_2;
  wire               readTokenRelease_2 = readData_readDataQueue_2_deq_ready & readData_readDataQueue_2_deq_valid;
  assign readData_readDataQueue_2_enq_valid = |readData_readResultSelect_2;
  wire [31:0]        readData_data_3;
  wire               isWaiteForThisData_3;
  wire               readData_readDataQueue_3_enq_ready = ~_readData_readDataQueue_fifo_3_full;
  wire               readData_readDataQueue_3_deq_ready;
  wire               readData_readDataQueue_3_enq_valid;
  wire               readData_readDataQueue_3_deq_valid = ~_readData_readDataQueue_fifo_3_empty | readData_readDataQueue_3_enq_valid;
  wire [31:0]        readData_readDataQueue_3_enq_bits;
  wire [31:0]        readData_readDataQueue_3_deq_bits = _readData_readDataQueue_fifo_3_empty ? readData_readDataQueue_3_enq_bits : _readData_readDataQueue_fifo_3_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_3 = {write1HPipe_1[3], write1HPipe_0[3]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_3 = {write1HPipe_3[3], write1HPipe_2[3]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_3 = {readData_readResultSelect_lo_lo_lo_hi_3, readData_readResultSelect_lo_lo_lo_lo_3};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_3 = {write1HPipe_5[3], write1HPipe_4[3]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_3 = {write1HPipe_7[3], write1HPipe_6[3]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_3 = {readData_readResultSelect_lo_lo_hi_hi_3, readData_readResultSelect_lo_lo_hi_lo_3};
  wire [7:0]         readData_readResultSelect_lo_lo_3 = {readData_readResultSelect_lo_lo_hi_3, readData_readResultSelect_lo_lo_lo_3};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_3 = {write1HPipe_9[3], write1HPipe_8[3]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_3 = {write1HPipe_11[3], write1HPipe_10[3]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_3 = {readData_readResultSelect_lo_hi_lo_hi_3, readData_readResultSelect_lo_hi_lo_lo_3};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_3 = {write1HPipe_13[3], write1HPipe_12[3]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_3 = {write1HPipe_15[3], write1HPipe_14[3]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_3 = {readData_readResultSelect_lo_hi_hi_hi_3, readData_readResultSelect_lo_hi_hi_lo_3};
  wire [7:0]         readData_readResultSelect_lo_hi_3 = {readData_readResultSelect_lo_hi_hi_3, readData_readResultSelect_lo_hi_lo_3};
  wire [15:0]        readData_readResultSelect_lo_3 = {readData_readResultSelect_lo_hi_3, readData_readResultSelect_lo_lo_3};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_3 = {write1HPipe_17[3], write1HPipe_16[3]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_3 = {write1HPipe_19[3], write1HPipe_18[3]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_3 = {readData_readResultSelect_hi_lo_lo_hi_3, readData_readResultSelect_hi_lo_lo_lo_3};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_3 = {write1HPipe_21[3], write1HPipe_20[3]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_3 = {write1HPipe_23[3], write1HPipe_22[3]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_3 = {readData_readResultSelect_hi_lo_hi_hi_3, readData_readResultSelect_hi_lo_hi_lo_3};
  wire [7:0]         readData_readResultSelect_hi_lo_3 = {readData_readResultSelect_hi_lo_hi_3, readData_readResultSelect_hi_lo_lo_3};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_3 = {write1HPipe_25[3], write1HPipe_24[3]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_3 = {write1HPipe_27[3], write1HPipe_26[3]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_3 = {readData_readResultSelect_hi_hi_lo_hi_3, readData_readResultSelect_hi_hi_lo_lo_3};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_3 = {write1HPipe_29[3], write1HPipe_28[3]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_3 = {write1HPipe_31[3], write1HPipe_30[3]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_3 = {readData_readResultSelect_hi_hi_hi_hi_3, readData_readResultSelect_hi_hi_hi_lo_3};
  wire [7:0]         readData_readResultSelect_hi_hi_3 = {readData_readResultSelect_hi_hi_hi_3, readData_readResultSelect_hi_hi_lo_3};
  wire [15:0]        readData_readResultSelect_hi_3 = {readData_readResultSelect_hi_hi_3, readData_readResultSelect_hi_lo_3};
  wire [31:0]        readData_readResultSelect_3 = {readData_readResultSelect_hi_3, readData_readResultSelect_lo_3};
  assign readData_data_3 =
    (readData_readResultSelect_3[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_3[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_3[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_3[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_3[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_3[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_3[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_3[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_3[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_3[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_3[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_3[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_3[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_3[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_3[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_3[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_3[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_3[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_3[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_3[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_3[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_3[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_3[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_3[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_3[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_3[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_3[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_3[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_3[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_3[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_3[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_3[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_3_enq_bits = readData_data_3;
  wire               readTokenRelease_3 = readData_readDataQueue_3_deq_ready & readData_readDataQueue_3_deq_valid;
  assign readData_readDataQueue_3_enq_valid = |readData_readResultSelect_3;
  wire [31:0]        readData_data_4;
  wire               isWaiteForThisData_4;
  wire               readData_readDataQueue_4_enq_ready = ~_readData_readDataQueue_fifo_4_full;
  wire               readData_readDataQueue_4_deq_ready;
  wire               readData_readDataQueue_4_enq_valid;
  wire               readData_readDataQueue_4_deq_valid = ~_readData_readDataQueue_fifo_4_empty | readData_readDataQueue_4_enq_valid;
  wire [31:0]        readData_readDataQueue_4_enq_bits;
  wire [31:0]        readData_readDataQueue_4_deq_bits = _readData_readDataQueue_fifo_4_empty ? readData_readDataQueue_4_enq_bits : _readData_readDataQueue_fifo_4_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_4 = {write1HPipe_1[4], write1HPipe_0[4]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_4 = {write1HPipe_3[4], write1HPipe_2[4]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_4 = {readData_readResultSelect_lo_lo_lo_hi_4, readData_readResultSelect_lo_lo_lo_lo_4};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_4 = {write1HPipe_5[4], write1HPipe_4[4]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_4 = {write1HPipe_7[4], write1HPipe_6[4]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_4 = {readData_readResultSelect_lo_lo_hi_hi_4, readData_readResultSelect_lo_lo_hi_lo_4};
  wire [7:0]         readData_readResultSelect_lo_lo_4 = {readData_readResultSelect_lo_lo_hi_4, readData_readResultSelect_lo_lo_lo_4};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_4 = {write1HPipe_9[4], write1HPipe_8[4]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_4 = {write1HPipe_11[4], write1HPipe_10[4]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_4 = {readData_readResultSelect_lo_hi_lo_hi_4, readData_readResultSelect_lo_hi_lo_lo_4};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_4 = {write1HPipe_13[4], write1HPipe_12[4]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_4 = {write1HPipe_15[4], write1HPipe_14[4]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_4 = {readData_readResultSelect_lo_hi_hi_hi_4, readData_readResultSelect_lo_hi_hi_lo_4};
  wire [7:0]         readData_readResultSelect_lo_hi_4 = {readData_readResultSelect_lo_hi_hi_4, readData_readResultSelect_lo_hi_lo_4};
  wire [15:0]        readData_readResultSelect_lo_4 = {readData_readResultSelect_lo_hi_4, readData_readResultSelect_lo_lo_4};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_4 = {write1HPipe_17[4], write1HPipe_16[4]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_4 = {write1HPipe_19[4], write1HPipe_18[4]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_4 = {readData_readResultSelect_hi_lo_lo_hi_4, readData_readResultSelect_hi_lo_lo_lo_4};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_4 = {write1HPipe_21[4], write1HPipe_20[4]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_4 = {write1HPipe_23[4], write1HPipe_22[4]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_4 = {readData_readResultSelect_hi_lo_hi_hi_4, readData_readResultSelect_hi_lo_hi_lo_4};
  wire [7:0]         readData_readResultSelect_hi_lo_4 = {readData_readResultSelect_hi_lo_hi_4, readData_readResultSelect_hi_lo_lo_4};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_4 = {write1HPipe_25[4], write1HPipe_24[4]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_4 = {write1HPipe_27[4], write1HPipe_26[4]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_4 = {readData_readResultSelect_hi_hi_lo_hi_4, readData_readResultSelect_hi_hi_lo_lo_4};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_4 = {write1HPipe_29[4], write1HPipe_28[4]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_4 = {write1HPipe_31[4], write1HPipe_30[4]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_4 = {readData_readResultSelect_hi_hi_hi_hi_4, readData_readResultSelect_hi_hi_hi_lo_4};
  wire [7:0]         readData_readResultSelect_hi_hi_4 = {readData_readResultSelect_hi_hi_hi_4, readData_readResultSelect_hi_hi_lo_4};
  wire [15:0]        readData_readResultSelect_hi_4 = {readData_readResultSelect_hi_hi_4, readData_readResultSelect_hi_lo_4};
  wire [31:0]        readData_readResultSelect_4 = {readData_readResultSelect_hi_4, readData_readResultSelect_lo_4};
  assign readData_data_4 =
    (readData_readResultSelect_4[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_4[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_4[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_4[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_4[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_4[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_4[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_4[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_4[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_4[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_4[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_4[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_4[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_4[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_4[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_4[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_4[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_4[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_4[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_4[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_4[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_4[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_4[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_4[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_4[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_4[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_4[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_4[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_4[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_4[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_4[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_4[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_4_enq_bits = readData_data_4;
  wire               readTokenRelease_4 = readData_readDataQueue_4_deq_ready & readData_readDataQueue_4_deq_valid;
  assign readData_readDataQueue_4_enq_valid = |readData_readResultSelect_4;
  wire [31:0]        readData_data_5;
  wire               isWaiteForThisData_5;
  wire               readData_readDataQueue_5_enq_ready = ~_readData_readDataQueue_fifo_5_full;
  wire               readData_readDataQueue_5_deq_ready;
  wire               readData_readDataQueue_5_enq_valid;
  wire               readData_readDataQueue_5_deq_valid = ~_readData_readDataQueue_fifo_5_empty | readData_readDataQueue_5_enq_valid;
  wire [31:0]        readData_readDataQueue_5_enq_bits;
  wire [31:0]        readData_readDataQueue_5_deq_bits = _readData_readDataQueue_fifo_5_empty ? readData_readDataQueue_5_enq_bits : _readData_readDataQueue_fifo_5_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_5 = {write1HPipe_1[5], write1HPipe_0[5]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_5 = {write1HPipe_3[5], write1HPipe_2[5]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_5 = {readData_readResultSelect_lo_lo_lo_hi_5, readData_readResultSelect_lo_lo_lo_lo_5};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_5 = {write1HPipe_5[5], write1HPipe_4[5]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_5 = {write1HPipe_7[5], write1HPipe_6[5]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_5 = {readData_readResultSelect_lo_lo_hi_hi_5, readData_readResultSelect_lo_lo_hi_lo_5};
  wire [7:0]         readData_readResultSelect_lo_lo_5 = {readData_readResultSelect_lo_lo_hi_5, readData_readResultSelect_lo_lo_lo_5};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_5 = {write1HPipe_9[5], write1HPipe_8[5]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_5 = {write1HPipe_11[5], write1HPipe_10[5]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_5 = {readData_readResultSelect_lo_hi_lo_hi_5, readData_readResultSelect_lo_hi_lo_lo_5};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_5 = {write1HPipe_13[5], write1HPipe_12[5]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_5 = {write1HPipe_15[5], write1HPipe_14[5]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_5 = {readData_readResultSelect_lo_hi_hi_hi_5, readData_readResultSelect_lo_hi_hi_lo_5};
  wire [7:0]         readData_readResultSelect_lo_hi_5 = {readData_readResultSelect_lo_hi_hi_5, readData_readResultSelect_lo_hi_lo_5};
  wire [15:0]        readData_readResultSelect_lo_5 = {readData_readResultSelect_lo_hi_5, readData_readResultSelect_lo_lo_5};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_5 = {write1HPipe_17[5], write1HPipe_16[5]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_5 = {write1HPipe_19[5], write1HPipe_18[5]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_5 = {readData_readResultSelect_hi_lo_lo_hi_5, readData_readResultSelect_hi_lo_lo_lo_5};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_5 = {write1HPipe_21[5], write1HPipe_20[5]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_5 = {write1HPipe_23[5], write1HPipe_22[5]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_5 = {readData_readResultSelect_hi_lo_hi_hi_5, readData_readResultSelect_hi_lo_hi_lo_5};
  wire [7:0]         readData_readResultSelect_hi_lo_5 = {readData_readResultSelect_hi_lo_hi_5, readData_readResultSelect_hi_lo_lo_5};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_5 = {write1HPipe_25[5], write1HPipe_24[5]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_5 = {write1HPipe_27[5], write1HPipe_26[5]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_5 = {readData_readResultSelect_hi_hi_lo_hi_5, readData_readResultSelect_hi_hi_lo_lo_5};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_5 = {write1HPipe_29[5], write1HPipe_28[5]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_5 = {write1HPipe_31[5], write1HPipe_30[5]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_5 = {readData_readResultSelect_hi_hi_hi_hi_5, readData_readResultSelect_hi_hi_hi_lo_5};
  wire [7:0]         readData_readResultSelect_hi_hi_5 = {readData_readResultSelect_hi_hi_hi_5, readData_readResultSelect_hi_hi_lo_5};
  wire [15:0]        readData_readResultSelect_hi_5 = {readData_readResultSelect_hi_hi_5, readData_readResultSelect_hi_lo_5};
  wire [31:0]        readData_readResultSelect_5 = {readData_readResultSelect_hi_5, readData_readResultSelect_lo_5};
  assign readData_data_5 =
    (readData_readResultSelect_5[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_5[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_5[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_5[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_5[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_5[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_5[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_5[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_5[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_5[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_5[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_5[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_5[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_5[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_5[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_5[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_5[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_5[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_5[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_5[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_5[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_5[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_5[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_5[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_5[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_5[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_5[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_5[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_5[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_5[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_5[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_5[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_5_enq_bits = readData_data_5;
  wire               readTokenRelease_5 = readData_readDataQueue_5_deq_ready & readData_readDataQueue_5_deq_valid;
  assign readData_readDataQueue_5_enq_valid = |readData_readResultSelect_5;
  wire [31:0]        readData_data_6;
  wire               isWaiteForThisData_6;
  wire               readData_readDataQueue_6_enq_ready = ~_readData_readDataQueue_fifo_6_full;
  wire               readData_readDataQueue_6_deq_ready;
  wire               readData_readDataQueue_6_enq_valid;
  wire               readData_readDataQueue_6_deq_valid = ~_readData_readDataQueue_fifo_6_empty | readData_readDataQueue_6_enq_valid;
  wire [31:0]        readData_readDataQueue_6_enq_bits;
  wire [31:0]        readData_readDataQueue_6_deq_bits = _readData_readDataQueue_fifo_6_empty ? readData_readDataQueue_6_enq_bits : _readData_readDataQueue_fifo_6_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_6 = {write1HPipe_1[6], write1HPipe_0[6]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_6 = {write1HPipe_3[6], write1HPipe_2[6]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_6 = {readData_readResultSelect_lo_lo_lo_hi_6, readData_readResultSelect_lo_lo_lo_lo_6};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_6 = {write1HPipe_5[6], write1HPipe_4[6]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_6 = {write1HPipe_7[6], write1HPipe_6[6]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_6 = {readData_readResultSelect_lo_lo_hi_hi_6, readData_readResultSelect_lo_lo_hi_lo_6};
  wire [7:0]         readData_readResultSelect_lo_lo_6 = {readData_readResultSelect_lo_lo_hi_6, readData_readResultSelect_lo_lo_lo_6};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_6 = {write1HPipe_9[6], write1HPipe_8[6]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_6 = {write1HPipe_11[6], write1HPipe_10[6]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_6 = {readData_readResultSelect_lo_hi_lo_hi_6, readData_readResultSelect_lo_hi_lo_lo_6};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_6 = {write1HPipe_13[6], write1HPipe_12[6]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_6 = {write1HPipe_15[6], write1HPipe_14[6]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_6 = {readData_readResultSelect_lo_hi_hi_hi_6, readData_readResultSelect_lo_hi_hi_lo_6};
  wire [7:0]         readData_readResultSelect_lo_hi_6 = {readData_readResultSelect_lo_hi_hi_6, readData_readResultSelect_lo_hi_lo_6};
  wire [15:0]        readData_readResultSelect_lo_6 = {readData_readResultSelect_lo_hi_6, readData_readResultSelect_lo_lo_6};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_6 = {write1HPipe_17[6], write1HPipe_16[6]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_6 = {write1HPipe_19[6], write1HPipe_18[6]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_6 = {readData_readResultSelect_hi_lo_lo_hi_6, readData_readResultSelect_hi_lo_lo_lo_6};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_6 = {write1HPipe_21[6], write1HPipe_20[6]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_6 = {write1HPipe_23[6], write1HPipe_22[6]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_6 = {readData_readResultSelect_hi_lo_hi_hi_6, readData_readResultSelect_hi_lo_hi_lo_6};
  wire [7:0]         readData_readResultSelect_hi_lo_6 = {readData_readResultSelect_hi_lo_hi_6, readData_readResultSelect_hi_lo_lo_6};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_6 = {write1HPipe_25[6], write1HPipe_24[6]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_6 = {write1HPipe_27[6], write1HPipe_26[6]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_6 = {readData_readResultSelect_hi_hi_lo_hi_6, readData_readResultSelect_hi_hi_lo_lo_6};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_6 = {write1HPipe_29[6], write1HPipe_28[6]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_6 = {write1HPipe_31[6], write1HPipe_30[6]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_6 = {readData_readResultSelect_hi_hi_hi_hi_6, readData_readResultSelect_hi_hi_hi_lo_6};
  wire [7:0]         readData_readResultSelect_hi_hi_6 = {readData_readResultSelect_hi_hi_hi_6, readData_readResultSelect_hi_hi_lo_6};
  wire [15:0]        readData_readResultSelect_hi_6 = {readData_readResultSelect_hi_hi_6, readData_readResultSelect_hi_lo_6};
  wire [31:0]        readData_readResultSelect_6 = {readData_readResultSelect_hi_6, readData_readResultSelect_lo_6};
  assign readData_data_6 =
    (readData_readResultSelect_6[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_6[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_6[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_6[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_6[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_6[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_6[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_6[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_6[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_6[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_6[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_6[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_6[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_6[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_6[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_6[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_6[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_6[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_6[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_6[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_6[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_6[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_6[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_6[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_6[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_6[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_6[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_6[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_6[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_6[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_6[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_6[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_6_enq_bits = readData_data_6;
  wire               readTokenRelease_6 = readData_readDataQueue_6_deq_ready & readData_readDataQueue_6_deq_valid;
  assign readData_readDataQueue_6_enq_valid = |readData_readResultSelect_6;
  wire [31:0]        readData_data_7;
  wire               isWaiteForThisData_7;
  wire               readData_readDataQueue_7_enq_ready = ~_readData_readDataQueue_fifo_7_full;
  wire               readData_readDataQueue_7_deq_ready;
  wire               readData_readDataQueue_7_enq_valid;
  wire               readData_readDataQueue_7_deq_valid = ~_readData_readDataQueue_fifo_7_empty | readData_readDataQueue_7_enq_valid;
  wire [31:0]        readData_readDataQueue_7_enq_bits;
  wire [31:0]        readData_readDataQueue_7_deq_bits = _readData_readDataQueue_fifo_7_empty ? readData_readDataQueue_7_enq_bits : _readData_readDataQueue_fifo_7_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_7 = {write1HPipe_1[7], write1HPipe_0[7]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_7 = {write1HPipe_3[7], write1HPipe_2[7]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_7 = {readData_readResultSelect_lo_lo_lo_hi_7, readData_readResultSelect_lo_lo_lo_lo_7};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_7 = {write1HPipe_5[7], write1HPipe_4[7]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_7 = {write1HPipe_7[7], write1HPipe_6[7]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_7 = {readData_readResultSelect_lo_lo_hi_hi_7, readData_readResultSelect_lo_lo_hi_lo_7};
  wire [7:0]         readData_readResultSelect_lo_lo_7 = {readData_readResultSelect_lo_lo_hi_7, readData_readResultSelect_lo_lo_lo_7};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_7 = {write1HPipe_9[7], write1HPipe_8[7]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_7 = {write1HPipe_11[7], write1HPipe_10[7]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_7 = {readData_readResultSelect_lo_hi_lo_hi_7, readData_readResultSelect_lo_hi_lo_lo_7};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_7 = {write1HPipe_13[7], write1HPipe_12[7]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_7 = {write1HPipe_15[7], write1HPipe_14[7]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_7 = {readData_readResultSelect_lo_hi_hi_hi_7, readData_readResultSelect_lo_hi_hi_lo_7};
  wire [7:0]         readData_readResultSelect_lo_hi_7 = {readData_readResultSelect_lo_hi_hi_7, readData_readResultSelect_lo_hi_lo_7};
  wire [15:0]        readData_readResultSelect_lo_7 = {readData_readResultSelect_lo_hi_7, readData_readResultSelect_lo_lo_7};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_7 = {write1HPipe_17[7], write1HPipe_16[7]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_7 = {write1HPipe_19[7], write1HPipe_18[7]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_7 = {readData_readResultSelect_hi_lo_lo_hi_7, readData_readResultSelect_hi_lo_lo_lo_7};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_7 = {write1HPipe_21[7], write1HPipe_20[7]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_7 = {write1HPipe_23[7], write1HPipe_22[7]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_7 = {readData_readResultSelect_hi_lo_hi_hi_7, readData_readResultSelect_hi_lo_hi_lo_7};
  wire [7:0]         readData_readResultSelect_hi_lo_7 = {readData_readResultSelect_hi_lo_hi_7, readData_readResultSelect_hi_lo_lo_7};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_7 = {write1HPipe_25[7], write1HPipe_24[7]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_7 = {write1HPipe_27[7], write1HPipe_26[7]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_7 = {readData_readResultSelect_hi_hi_lo_hi_7, readData_readResultSelect_hi_hi_lo_lo_7};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_7 = {write1HPipe_29[7], write1HPipe_28[7]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_7 = {write1HPipe_31[7], write1HPipe_30[7]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_7 = {readData_readResultSelect_hi_hi_hi_hi_7, readData_readResultSelect_hi_hi_hi_lo_7};
  wire [7:0]         readData_readResultSelect_hi_hi_7 = {readData_readResultSelect_hi_hi_hi_7, readData_readResultSelect_hi_hi_lo_7};
  wire [15:0]        readData_readResultSelect_hi_7 = {readData_readResultSelect_hi_hi_7, readData_readResultSelect_hi_lo_7};
  wire [31:0]        readData_readResultSelect_7 = {readData_readResultSelect_hi_7, readData_readResultSelect_lo_7};
  assign readData_data_7 =
    (readData_readResultSelect_7[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_7[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_7[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_7[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_7[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_7[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_7[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_7[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_7[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_7[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_7[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_7[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_7[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_7[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_7[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_7[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_7[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_7[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_7[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_7[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_7[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_7[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_7[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_7[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_7[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_7[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_7[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_7[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_7[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_7[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_7[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_7[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_7_enq_bits = readData_data_7;
  wire               readTokenRelease_7 = readData_readDataQueue_7_deq_ready & readData_readDataQueue_7_deq_valid;
  assign readData_readDataQueue_7_enq_valid = |readData_readResultSelect_7;
  wire [31:0]        readData_data_8;
  wire               isWaiteForThisData_8;
  wire               readData_readDataQueue_8_enq_ready = ~_readData_readDataQueue_fifo_8_full;
  wire               readData_readDataQueue_8_deq_ready;
  wire               readData_readDataQueue_8_enq_valid;
  wire               readData_readDataQueue_8_deq_valid = ~_readData_readDataQueue_fifo_8_empty | readData_readDataQueue_8_enq_valid;
  wire [31:0]        readData_readDataQueue_8_enq_bits;
  wire [31:0]        readData_readDataQueue_8_deq_bits = _readData_readDataQueue_fifo_8_empty ? readData_readDataQueue_8_enq_bits : _readData_readDataQueue_fifo_8_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_8 = {write1HPipe_1[8], write1HPipe_0[8]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_8 = {write1HPipe_3[8], write1HPipe_2[8]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_8 = {readData_readResultSelect_lo_lo_lo_hi_8, readData_readResultSelect_lo_lo_lo_lo_8};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_8 = {write1HPipe_5[8], write1HPipe_4[8]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_8 = {write1HPipe_7[8], write1HPipe_6[8]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_8 = {readData_readResultSelect_lo_lo_hi_hi_8, readData_readResultSelect_lo_lo_hi_lo_8};
  wire [7:0]         readData_readResultSelect_lo_lo_8 = {readData_readResultSelect_lo_lo_hi_8, readData_readResultSelect_lo_lo_lo_8};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_8 = {write1HPipe_9[8], write1HPipe_8[8]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_8 = {write1HPipe_11[8], write1HPipe_10[8]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_8 = {readData_readResultSelect_lo_hi_lo_hi_8, readData_readResultSelect_lo_hi_lo_lo_8};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_8 = {write1HPipe_13[8], write1HPipe_12[8]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_8 = {write1HPipe_15[8], write1HPipe_14[8]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_8 = {readData_readResultSelect_lo_hi_hi_hi_8, readData_readResultSelect_lo_hi_hi_lo_8};
  wire [7:0]         readData_readResultSelect_lo_hi_8 = {readData_readResultSelect_lo_hi_hi_8, readData_readResultSelect_lo_hi_lo_8};
  wire [15:0]        readData_readResultSelect_lo_8 = {readData_readResultSelect_lo_hi_8, readData_readResultSelect_lo_lo_8};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_8 = {write1HPipe_17[8], write1HPipe_16[8]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_8 = {write1HPipe_19[8], write1HPipe_18[8]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_8 = {readData_readResultSelect_hi_lo_lo_hi_8, readData_readResultSelect_hi_lo_lo_lo_8};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_8 = {write1HPipe_21[8], write1HPipe_20[8]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_8 = {write1HPipe_23[8], write1HPipe_22[8]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_8 = {readData_readResultSelect_hi_lo_hi_hi_8, readData_readResultSelect_hi_lo_hi_lo_8};
  wire [7:0]         readData_readResultSelect_hi_lo_8 = {readData_readResultSelect_hi_lo_hi_8, readData_readResultSelect_hi_lo_lo_8};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_8 = {write1HPipe_25[8], write1HPipe_24[8]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_8 = {write1HPipe_27[8], write1HPipe_26[8]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_8 = {readData_readResultSelect_hi_hi_lo_hi_8, readData_readResultSelect_hi_hi_lo_lo_8};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_8 = {write1HPipe_29[8], write1HPipe_28[8]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_8 = {write1HPipe_31[8], write1HPipe_30[8]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_8 = {readData_readResultSelect_hi_hi_hi_hi_8, readData_readResultSelect_hi_hi_hi_lo_8};
  wire [7:0]         readData_readResultSelect_hi_hi_8 = {readData_readResultSelect_hi_hi_hi_8, readData_readResultSelect_hi_hi_lo_8};
  wire [15:0]        readData_readResultSelect_hi_8 = {readData_readResultSelect_hi_hi_8, readData_readResultSelect_hi_lo_8};
  wire [31:0]        readData_readResultSelect_8 = {readData_readResultSelect_hi_8, readData_readResultSelect_lo_8};
  assign readData_data_8 =
    (readData_readResultSelect_8[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_8[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_8[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_8[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_8[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_8[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_8[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_8[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_8[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_8[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_8[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_8[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_8[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_8[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_8[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_8[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_8[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_8[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_8[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_8[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_8[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_8[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_8[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_8[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_8[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_8[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_8[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_8[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_8[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_8[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_8[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_8[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_8_enq_bits = readData_data_8;
  wire               readTokenRelease_8 = readData_readDataQueue_8_deq_ready & readData_readDataQueue_8_deq_valid;
  assign readData_readDataQueue_8_enq_valid = |readData_readResultSelect_8;
  wire [31:0]        readData_data_9;
  wire               isWaiteForThisData_9;
  wire               readData_readDataQueue_9_enq_ready = ~_readData_readDataQueue_fifo_9_full;
  wire               readData_readDataQueue_9_deq_ready;
  wire               readData_readDataQueue_9_enq_valid;
  wire               readData_readDataQueue_9_deq_valid = ~_readData_readDataQueue_fifo_9_empty | readData_readDataQueue_9_enq_valid;
  wire [31:0]        readData_readDataQueue_9_enq_bits;
  wire [31:0]        readData_readDataQueue_9_deq_bits = _readData_readDataQueue_fifo_9_empty ? readData_readDataQueue_9_enq_bits : _readData_readDataQueue_fifo_9_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_9 = {write1HPipe_1[9], write1HPipe_0[9]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_9 = {write1HPipe_3[9], write1HPipe_2[9]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_9 = {readData_readResultSelect_lo_lo_lo_hi_9, readData_readResultSelect_lo_lo_lo_lo_9};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_9 = {write1HPipe_5[9], write1HPipe_4[9]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_9 = {write1HPipe_7[9], write1HPipe_6[9]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_9 = {readData_readResultSelect_lo_lo_hi_hi_9, readData_readResultSelect_lo_lo_hi_lo_9};
  wire [7:0]         readData_readResultSelect_lo_lo_9 = {readData_readResultSelect_lo_lo_hi_9, readData_readResultSelect_lo_lo_lo_9};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_9 = {write1HPipe_9[9], write1HPipe_8[9]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_9 = {write1HPipe_11[9], write1HPipe_10[9]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_9 = {readData_readResultSelect_lo_hi_lo_hi_9, readData_readResultSelect_lo_hi_lo_lo_9};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_9 = {write1HPipe_13[9], write1HPipe_12[9]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_9 = {write1HPipe_15[9], write1HPipe_14[9]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_9 = {readData_readResultSelect_lo_hi_hi_hi_9, readData_readResultSelect_lo_hi_hi_lo_9};
  wire [7:0]         readData_readResultSelect_lo_hi_9 = {readData_readResultSelect_lo_hi_hi_9, readData_readResultSelect_lo_hi_lo_9};
  wire [15:0]        readData_readResultSelect_lo_9 = {readData_readResultSelect_lo_hi_9, readData_readResultSelect_lo_lo_9};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_9 = {write1HPipe_17[9], write1HPipe_16[9]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_9 = {write1HPipe_19[9], write1HPipe_18[9]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_9 = {readData_readResultSelect_hi_lo_lo_hi_9, readData_readResultSelect_hi_lo_lo_lo_9};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_9 = {write1HPipe_21[9], write1HPipe_20[9]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_9 = {write1HPipe_23[9], write1HPipe_22[9]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_9 = {readData_readResultSelect_hi_lo_hi_hi_9, readData_readResultSelect_hi_lo_hi_lo_9};
  wire [7:0]         readData_readResultSelect_hi_lo_9 = {readData_readResultSelect_hi_lo_hi_9, readData_readResultSelect_hi_lo_lo_9};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_9 = {write1HPipe_25[9], write1HPipe_24[9]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_9 = {write1HPipe_27[9], write1HPipe_26[9]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_9 = {readData_readResultSelect_hi_hi_lo_hi_9, readData_readResultSelect_hi_hi_lo_lo_9};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_9 = {write1HPipe_29[9], write1HPipe_28[9]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_9 = {write1HPipe_31[9], write1HPipe_30[9]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_9 = {readData_readResultSelect_hi_hi_hi_hi_9, readData_readResultSelect_hi_hi_hi_lo_9};
  wire [7:0]         readData_readResultSelect_hi_hi_9 = {readData_readResultSelect_hi_hi_hi_9, readData_readResultSelect_hi_hi_lo_9};
  wire [15:0]        readData_readResultSelect_hi_9 = {readData_readResultSelect_hi_hi_9, readData_readResultSelect_hi_lo_9};
  wire [31:0]        readData_readResultSelect_9 = {readData_readResultSelect_hi_9, readData_readResultSelect_lo_9};
  assign readData_data_9 =
    (readData_readResultSelect_9[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_9[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_9[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_9[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_9[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_9[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_9[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_9[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_9[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_9[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_9[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_9[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_9[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_9[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_9[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_9[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_9[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_9[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_9[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_9[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_9[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_9[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_9[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_9[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_9[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_9[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_9[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_9[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_9[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_9[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_9[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_9[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_9_enq_bits = readData_data_9;
  wire               readTokenRelease_9 = readData_readDataQueue_9_deq_ready & readData_readDataQueue_9_deq_valid;
  assign readData_readDataQueue_9_enq_valid = |readData_readResultSelect_9;
  wire [31:0]        readData_data_10;
  wire               isWaiteForThisData_10;
  wire               readData_readDataQueue_10_enq_ready = ~_readData_readDataQueue_fifo_10_full;
  wire               readData_readDataQueue_10_deq_ready;
  wire               readData_readDataQueue_10_enq_valid;
  wire               readData_readDataQueue_10_deq_valid = ~_readData_readDataQueue_fifo_10_empty | readData_readDataQueue_10_enq_valid;
  wire [31:0]        readData_readDataQueue_10_enq_bits;
  wire [31:0]        readData_readDataQueue_10_deq_bits = _readData_readDataQueue_fifo_10_empty ? readData_readDataQueue_10_enq_bits : _readData_readDataQueue_fifo_10_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_10 = {write1HPipe_1[10], write1HPipe_0[10]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_10 = {write1HPipe_3[10], write1HPipe_2[10]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_10 = {readData_readResultSelect_lo_lo_lo_hi_10, readData_readResultSelect_lo_lo_lo_lo_10};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_10 = {write1HPipe_5[10], write1HPipe_4[10]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_10 = {write1HPipe_7[10], write1HPipe_6[10]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_10 = {readData_readResultSelect_lo_lo_hi_hi_10, readData_readResultSelect_lo_lo_hi_lo_10};
  wire [7:0]         readData_readResultSelect_lo_lo_10 = {readData_readResultSelect_lo_lo_hi_10, readData_readResultSelect_lo_lo_lo_10};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_10 = {write1HPipe_9[10], write1HPipe_8[10]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_10 = {write1HPipe_11[10], write1HPipe_10[10]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_10 = {readData_readResultSelect_lo_hi_lo_hi_10, readData_readResultSelect_lo_hi_lo_lo_10};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_10 = {write1HPipe_13[10], write1HPipe_12[10]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_10 = {write1HPipe_15[10], write1HPipe_14[10]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_10 = {readData_readResultSelect_lo_hi_hi_hi_10, readData_readResultSelect_lo_hi_hi_lo_10};
  wire [7:0]         readData_readResultSelect_lo_hi_10 = {readData_readResultSelect_lo_hi_hi_10, readData_readResultSelect_lo_hi_lo_10};
  wire [15:0]        readData_readResultSelect_lo_10 = {readData_readResultSelect_lo_hi_10, readData_readResultSelect_lo_lo_10};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_10 = {write1HPipe_17[10], write1HPipe_16[10]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_10 = {write1HPipe_19[10], write1HPipe_18[10]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_10 = {readData_readResultSelect_hi_lo_lo_hi_10, readData_readResultSelect_hi_lo_lo_lo_10};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_10 = {write1HPipe_21[10], write1HPipe_20[10]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_10 = {write1HPipe_23[10], write1HPipe_22[10]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_10 = {readData_readResultSelect_hi_lo_hi_hi_10, readData_readResultSelect_hi_lo_hi_lo_10};
  wire [7:0]         readData_readResultSelect_hi_lo_10 = {readData_readResultSelect_hi_lo_hi_10, readData_readResultSelect_hi_lo_lo_10};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_10 = {write1HPipe_25[10], write1HPipe_24[10]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_10 = {write1HPipe_27[10], write1HPipe_26[10]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_10 = {readData_readResultSelect_hi_hi_lo_hi_10, readData_readResultSelect_hi_hi_lo_lo_10};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_10 = {write1HPipe_29[10], write1HPipe_28[10]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_10 = {write1HPipe_31[10], write1HPipe_30[10]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_10 = {readData_readResultSelect_hi_hi_hi_hi_10, readData_readResultSelect_hi_hi_hi_lo_10};
  wire [7:0]         readData_readResultSelect_hi_hi_10 = {readData_readResultSelect_hi_hi_hi_10, readData_readResultSelect_hi_hi_lo_10};
  wire [15:0]        readData_readResultSelect_hi_10 = {readData_readResultSelect_hi_hi_10, readData_readResultSelect_hi_lo_10};
  wire [31:0]        readData_readResultSelect_10 = {readData_readResultSelect_hi_10, readData_readResultSelect_lo_10};
  assign readData_data_10 =
    (readData_readResultSelect_10[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_10[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_10[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_10[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_10[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_10[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_10[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_10[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_10[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_10[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_10[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_10[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_10[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_10[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_10[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_10[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_10[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_10[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_10[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_10[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_10[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_10[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_10[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_10[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_10[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_10[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_10[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_10[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_10[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_10[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_10[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_10[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_10_enq_bits = readData_data_10;
  wire               readTokenRelease_10 = readData_readDataQueue_10_deq_ready & readData_readDataQueue_10_deq_valid;
  assign readData_readDataQueue_10_enq_valid = |readData_readResultSelect_10;
  wire [31:0]        readData_data_11;
  wire               isWaiteForThisData_11;
  wire               readData_readDataQueue_11_enq_ready = ~_readData_readDataQueue_fifo_11_full;
  wire               readData_readDataQueue_11_deq_ready;
  wire               readData_readDataQueue_11_enq_valid;
  wire               readData_readDataQueue_11_deq_valid = ~_readData_readDataQueue_fifo_11_empty | readData_readDataQueue_11_enq_valid;
  wire [31:0]        readData_readDataQueue_11_enq_bits;
  wire [31:0]        readData_readDataQueue_11_deq_bits = _readData_readDataQueue_fifo_11_empty ? readData_readDataQueue_11_enq_bits : _readData_readDataQueue_fifo_11_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_11 = {write1HPipe_1[11], write1HPipe_0[11]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_11 = {write1HPipe_3[11], write1HPipe_2[11]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_11 = {readData_readResultSelect_lo_lo_lo_hi_11, readData_readResultSelect_lo_lo_lo_lo_11};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_11 = {write1HPipe_5[11], write1HPipe_4[11]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_11 = {write1HPipe_7[11], write1HPipe_6[11]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_11 = {readData_readResultSelect_lo_lo_hi_hi_11, readData_readResultSelect_lo_lo_hi_lo_11};
  wire [7:0]         readData_readResultSelect_lo_lo_11 = {readData_readResultSelect_lo_lo_hi_11, readData_readResultSelect_lo_lo_lo_11};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_11 = {write1HPipe_9[11], write1HPipe_8[11]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_11 = {write1HPipe_11[11], write1HPipe_10[11]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_11 = {readData_readResultSelect_lo_hi_lo_hi_11, readData_readResultSelect_lo_hi_lo_lo_11};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_11 = {write1HPipe_13[11], write1HPipe_12[11]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_11 = {write1HPipe_15[11], write1HPipe_14[11]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_11 = {readData_readResultSelect_lo_hi_hi_hi_11, readData_readResultSelect_lo_hi_hi_lo_11};
  wire [7:0]         readData_readResultSelect_lo_hi_11 = {readData_readResultSelect_lo_hi_hi_11, readData_readResultSelect_lo_hi_lo_11};
  wire [15:0]        readData_readResultSelect_lo_11 = {readData_readResultSelect_lo_hi_11, readData_readResultSelect_lo_lo_11};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_11 = {write1HPipe_17[11], write1HPipe_16[11]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_11 = {write1HPipe_19[11], write1HPipe_18[11]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_11 = {readData_readResultSelect_hi_lo_lo_hi_11, readData_readResultSelect_hi_lo_lo_lo_11};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_11 = {write1HPipe_21[11], write1HPipe_20[11]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_11 = {write1HPipe_23[11], write1HPipe_22[11]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_11 = {readData_readResultSelect_hi_lo_hi_hi_11, readData_readResultSelect_hi_lo_hi_lo_11};
  wire [7:0]         readData_readResultSelect_hi_lo_11 = {readData_readResultSelect_hi_lo_hi_11, readData_readResultSelect_hi_lo_lo_11};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_11 = {write1HPipe_25[11], write1HPipe_24[11]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_11 = {write1HPipe_27[11], write1HPipe_26[11]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_11 = {readData_readResultSelect_hi_hi_lo_hi_11, readData_readResultSelect_hi_hi_lo_lo_11};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_11 = {write1HPipe_29[11], write1HPipe_28[11]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_11 = {write1HPipe_31[11], write1HPipe_30[11]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_11 = {readData_readResultSelect_hi_hi_hi_hi_11, readData_readResultSelect_hi_hi_hi_lo_11};
  wire [7:0]         readData_readResultSelect_hi_hi_11 = {readData_readResultSelect_hi_hi_hi_11, readData_readResultSelect_hi_hi_lo_11};
  wire [15:0]        readData_readResultSelect_hi_11 = {readData_readResultSelect_hi_hi_11, readData_readResultSelect_hi_lo_11};
  wire [31:0]        readData_readResultSelect_11 = {readData_readResultSelect_hi_11, readData_readResultSelect_lo_11};
  assign readData_data_11 =
    (readData_readResultSelect_11[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_11[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_11[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_11[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_11[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_11[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_11[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_11[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_11[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_11[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_11[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_11[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_11[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_11[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_11[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_11[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_11[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_11[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_11[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_11[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_11[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_11[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_11[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_11[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_11[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_11[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_11[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_11[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_11[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_11[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_11[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_11[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_11_enq_bits = readData_data_11;
  wire               readTokenRelease_11 = readData_readDataQueue_11_deq_ready & readData_readDataQueue_11_deq_valid;
  assign readData_readDataQueue_11_enq_valid = |readData_readResultSelect_11;
  wire [31:0]        readData_data_12;
  wire               isWaiteForThisData_12;
  wire               readData_readDataQueue_12_enq_ready = ~_readData_readDataQueue_fifo_12_full;
  wire               readData_readDataQueue_12_deq_ready;
  wire               readData_readDataQueue_12_enq_valid;
  wire               readData_readDataQueue_12_deq_valid = ~_readData_readDataQueue_fifo_12_empty | readData_readDataQueue_12_enq_valid;
  wire [31:0]        readData_readDataQueue_12_enq_bits;
  wire [31:0]        readData_readDataQueue_12_deq_bits = _readData_readDataQueue_fifo_12_empty ? readData_readDataQueue_12_enq_bits : _readData_readDataQueue_fifo_12_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_12 = {write1HPipe_1[12], write1HPipe_0[12]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_12 = {write1HPipe_3[12], write1HPipe_2[12]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_12 = {readData_readResultSelect_lo_lo_lo_hi_12, readData_readResultSelect_lo_lo_lo_lo_12};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_12 = {write1HPipe_5[12], write1HPipe_4[12]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_12 = {write1HPipe_7[12], write1HPipe_6[12]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_12 = {readData_readResultSelect_lo_lo_hi_hi_12, readData_readResultSelect_lo_lo_hi_lo_12};
  wire [7:0]         readData_readResultSelect_lo_lo_12 = {readData_readResultSelect_lo_lo_hi_12, readData_readResultSelect_lo_lo_lo_12};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_12 = {write1HPipe_9[12], write1HPipe_8[12]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_12 = {write1HPipe_11[12], write1HPipe_10[12]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_12 = {readData_readResultSelect_lo_hi_lo_hi_12, readData_readResultSelect_lo_hi_lo_lo_12};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_12 = {write1HPipe_13[12], write1HPipe_12[12]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_12 = {write1HPipe_15[12], write1HPipe_14[12]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_12 = {readData_readResultSelect_lo_hi_hi_hi_12, readData_readResultSelect_lo_hi_hi_lo_12};
  wire [7:0]         readData_readResultSelect_lo_hi_12 = {readData_readResultSelect_lo_hi_hi_12, readData_readResultSelect_lo_hi_lo_12};
  wire [15:0]        readData_readResultSelect_lo_12 = {readData_readResultSelect_lo_hi_12, readData_readResultSelect_lo_lo_12};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_12 = {write1HPipe_17[12], write1HPipe_16[12]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_12 = {write1HPipe_19[12], write1HPipe_18[12]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_12 = {readData_readResultSelect_hi_lo_lo_hi_12, readData_readResultSelect_hi_lo_lo_lo_12};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_12 = {write1HPipe_21[12], write1HPipe_20[12]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_12 = {write1HPipe_23[12], write1HPipe_22[12]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_12 = {readData_readResultSelect_hi_lo_hi_hi_12, readData_readResultSelect_hi_lo_hi_lo_12};
  wire [7:0]         readData_readResultSelect_hi_lo_12 = {readData_readResultSelect_hi_lo_hi_12, readData_readResultSelect_hi_lo_lo_12};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_12 = {write1HPipe_25[12], write1HPipe_24[12]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_12 = {write1HPipe_27[12], write1HPipe_26[12]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_12 = {readData_readResultSelect_hi_hi_lo_hi_12, readData_readResultSelect_hi_hi_lo_lo_12};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_12 = {write1HPipe_29[12], write1HPipe_28[12]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_12 = {write1HPipe_31[12], write1HPipe_30[12]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_12 = {readData_readResultSelect_hi_hi_hi_hi_12, readData_readResultSelect_hi_hi_hi_lo_12};
  wire [7:0]         readData_readResultSelect_hi_hi_12 = {readData_readResultSelect_hi_hi_hi_12, readData_readResultSelect_hi_hi_lo_12};
  wire [15:0]        readData_readResultSelect_hi_12 = {readData_readResultSelect_hi_hi_12, readData_readResultSelect_hi_lo_12};
  wire [31:0]        readData_readResultSelect_12 = {readData_readResultSelect_hi_12, readData_readResultSelect_lo_12};
  assign readData_data_12 =
    (readData_readResultSelect_12[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_12[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_12[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_12[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_12[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_12[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_12[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_12[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_12[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_12[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_12[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_12[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_12[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_12[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_12[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_12[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_12[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_12[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_12[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_12[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_12[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_12[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_12[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_12[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_12[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_12[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_12[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_12[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_12[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_12[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_12[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_12[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_12_enq_bits = readData_data_12;
  wire               readTokenRelease_12 = readData_readDataQueue_12_deq_ready & readData_readDataQueue_12_deq_valid;
  assign readData_readDataQueue_12_enq_valid = |readData_readResultSelect_12;
  wire [31:0]        readData_data_13;
  wire               isWaiteForThisData_13;
  wire               readData_readDataQueue_13_enq_ready = ~_readData_readDataQueue_fifo_13_full;
  wire               readData_readDataQueue_13_deq_ready;
  wire               readData_readDataQueue_13_enq_valid;
  wire               readData_readDataQueue_13_deq_valid = ~_readData_readDataQueue_fifo_13_empty | readData_readDataQueue_13_enq_valid;
  wire [31:0]        readData_readDataQueue_13_enq_bits;
  wire [31:0]        readData_readDataQueue_13_deq_bits = _readData_readDataQueue_fifo_13_empty ? readData_readDataQueue_13_enq_bits : _readData_readDataQueue_fifo_13_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_13 = {write1HPipe_1[13], write1HPipe_0[13]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_13 = {write1HPipe_3[13], write1HPipe_2[13]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_13 = {readData_readResultSelect_lo_lo_lo_hi_13, readData_readResultSelect_lo_lo_lo_lo_13};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_13 = {write1HPipe_5[13], write1HPipe_4[13]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_13 = {write1HPipe_7[13], write1HPipe_6[13]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_13 = {readData_readResultSelect_lo_lo_hi_hi_13, readData_readResultSelect_lo_lo_hi_lo_13};
  wire [7:0]         readData_readResultSelect_lo_lo_13 = {readData_readResultSelect_lo_lo_hi_13, readData_readResultSelect_lo_lo_lo_13};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_13 = {write1HPipe_9[13], write1HPipe_8[13]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_13 = {write1HPipe_11[13], write1HPipe_10[13]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_13 = {readData_readResultSelect_lo_hi_lo_hi_13, readData_readResultSelect_lo_hi_lo_lo_13};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_13 = {write1HPipe_13[13], write1HPipe_12[13]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_13 = {write1HPipe_15[13], write1HPipe_14[13]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_13 = {readData_readResultSelect_lo_hi_hi_hi_13, readData_readResultSelect_lo_hi_hi_lo_13};
  wire [7:0]         readData_readResultSelect_lo_hi_13 = {readData_readResultSelect_lo_hi_hi_13, readData_readResultSelect_lo_hi_lo_13};
  wire [15:0]        readData_readResultSelect_lo_13 = {readData_readResultSelect_lo_hi_13, readData_readResultSelect_lo_lo_13};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_13 = {write1HPipe_17[13], write1HPipe_16[13]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_13 = {write1HPipe_19[13], write1HPipe_18[13]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_13 = {readData_readResultSelect_hi_lo_lo_hi_13, readData_readResultSelect_hi_lo_lo_lo_13};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_13 = {write1HPipe_21[13], write1HPipe_20[13]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_13 = {write1HPipe_23[13], write1HPipe_22[13]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_13 = {readData_readResultSelect_hi_lo_hi_hi_13, readData_readResultSelect_hi_lo_hi_lo_13};
  wire [7:0]         readData_readResultSelect_hi_lo_13 = {readData_readResultSelect_hi_lo_hi_13, readData_readResultSelect_hi_lo_lo_13};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_13 = {write1HPipe_25[13], write1HPipe_24[13]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_13 = {write1HPipe_27[13], write1HPipe_26[13]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_13 = {readData_readResultSelect_hi_hi_lo_hi_13, readData_readResultSelect_hi_hi_lo_lo_13};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_13 = {write1HPipe_29[13], write1HPipe_28[13]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_13 = {write1HPipe_31[13], write1HPipe_30[13]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_13 = {readData_readResultSelect_hi_hi_hi_hi_13, readData_readResultSelect_hi_hi_hi_lo_13};
  wire [7:0]         readData_readResultSelect_hi_hi_13 = {readData_readResultSelect_hi_hi_hi_13, readData_readResultSelect_hi_hi_lo_13};
  wire [15:0]        readData_readResultSelect_hi_13 = {readData_readResultSelect_hi_hi_13, readData_readResultSelect_hi_lo_13};
  wire [31:0]        readData_readResultSelect_13 = {readData_readResultSelect_hi_13, readData_readResultSelect_lo_13};
  assign readData_data_13 =
    (readData_readResultSelect_13[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_13[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_13[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_13[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_13[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_13[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_13[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_13[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_13[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_13[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_13[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_13[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_13[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_13[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_13[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_13[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_13[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_13[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_13[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_13[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_13[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_13[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_13[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_13[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_13[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_13[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_13[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_13[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_13[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_13[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_13[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_13[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_13_enq_bits = readData_data_13;
  wire               readTokenRelease_13 = readData_readDataQueue_13_deq_ready & readData_readDataQueue_13_deq_valid;
  assign readData_readDataQueue_13_enq_valid = |readData_readResultSelect_13;
  wire [31:0]        readData_data_14;
  wire               isWaiteForThisData_14;
  wire               readData_readDataQueue_14_enq_ready = ~_readData_readDataQueue_fifo_14_full;
  wire               readData_readDataQueue_14_deq_ready;
  wire               readData_readDataQueue_14_enq_valid;
  wire               readData_readDataQueue_14_deq_valid = ~_readData_readDataQueue_fifo_14_empty | readData_readDataQueue_14_enq_valid;
  wire [31:0]        readData_readDataQueue_14_enq_bits;
  wire [31:0]        readData_readDataQueue_14_deq_bits = _readData_readDataQueue_fifo_14_empty ? readData_readDataQueue_14_enq_bits : _readData_readDataQueue_fifo_14_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_14 = {write1HPipe_1[14], write1HPipe_0[14]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_14 = {write1HPipe_3[14], write1HPipe_2[14]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_14 = {readData_readResultSelect_lo_lo_lo_hi_14, readData_readResultSelect_lo_lo_lo_lo_14};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_14 = {write1HPipe_5[14], write1HPipe_4[14]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_14 = {write1HPipe_7[14], write1HPipe_6[14]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_14 = {readData_readResultSelect_lo_lo_hi_hi_14, readData_readResultSelect_lo_lo_hi_lo_14};
  wire [7:0]         readData_readResultSelect_lo_lo_14 = {readData_readResultSelect_lo_lo_hi_14, readData_readResultSelect_lo_lo_lo_14};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_14 = {write1HPipe_9[14], write1HPipe_8[14]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_14 = {write1HPipe_11[14], write1HPipe_10[14]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_14 = {readData_readResultSelect_lo_hi_lo_hi_14, readData_readResultSelect_lo_hi_lo_lo_14};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_14 = {write1HPipe_13[14], write1HPipe_12[14]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_14 = {write1HPipe_15[14], write1HPipe_14[14]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_14 = {readData_readResultSelect_lo_hi_hi_hi_14, readData_readResultSelect_lo_hi_hi_lo_14};
  wire [7:0]         readData_readResultSelect_lo_hi_14 = {readData_readResultSelect_lo_hi_hi_14, readData_readResultSelect_lo_hi_lo_14};
  wire [15:0]        readData_readResultSelect_lo_14 = {readData_readResultSelect_lo_hi_14, readData_readResultSelect_lo_lo_14};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_14 = {write1HPipe_17[14], write1HPipe_16[14]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_14 = {write1HPipe_19[14], write1HPipe_18[14]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_14 = {readData_readResultSelect_hi_lo_lo_hi_14, readData_readResultSelect_hi_lo_lo_lo_14};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_14 = {write1HPipe_21[14], write1HPipe_20[14]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_14 = {write1HPipe_23[14], write1HPipe_22[14]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_14 = {readData_readResultSelect_hi_lo_hi_hi_14, readData_readResultSelect_hi_lo_hi_lo_14};
  wire [7:0]         readData_readResultSelect_hi_lo_14 = {readData_readResultSelect_hi_lo_hi_14, readData_readResultSelect_hi_lo_lo_14};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_14 = {write1HPipe_25[14], write1HPipe_24[14]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_14 = {write1HPipe_27[14], write1HPipe_26[14]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_14 = {readData_readResultSelect_hi_hi_lo_hi_14, readData_readResultSelect_hi_hi_lo_lo_14};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_14 = {write1HPipe_29[14], write1HPipe_28[14]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_14 = {write1HPipe_31[14], write1HPipe_30[14]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_14 = {readData_readResultSelect_hi_hi_hi_hi_14, readData_readResultSelect_hi_hi_hi_lo_14};
  wire [7:0]         readData_readResultSelect_hi_hi_14 = {readData_readResultSelect_hi_hi_hi_14, readData_readResultSelect_hi_hi_lo_14};
  wire [15:0]        readData_readResultSelect_hi_14 = {readData_readResultSelect_hi_hi_14, readData_readResultSelect_hi_lo_14};
  wire [31:0]        readData_readResultSelect_14 = {readData_readResultSelect_hi_14, readData_readResultSelect_lo_14};
  assign readData_data_14 =
    (readData_readResultSelect_14[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_14[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_14[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_14[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_14[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_14[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_14[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_14[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_14[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_14[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_14[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_14[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_14[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_14[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_14[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_14[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_14[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_14[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_14[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_14[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_14[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_14[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_14[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_14[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_14[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_14[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_14[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_14[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_14[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_14[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_14[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_14[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_14_enq_bits = readData_data_14;
  wire               readTokenRelease_14 = readData_readDataQueue_14_deq_ready & readData_readDataQueue_14_deq_valid;
  assign readData_readDataQueue_14_enq_valid = |readData_readResultSelect_14;
  wire [31:0]        readData_data_15;
  wire               isWaiteForThisData_15;
  wire               readData_readDataQueue_15_enq_ready = ~_readData_readDataQueue_fifo_15_full;
  wire               readData_readDataQueue_15_deq_ready;
  wire               readData_readDataQueue_15_enq_valid;
  wire               readData_readDataQueue_15_deq_valid = ~_readData_readDataQueue_fifo_15_empty | readData_readDataQueue_15_enq_valid;
  wire [31:0]        readData_readDataQueue_15_enq_bits;
  wire [31:0]        readData_readDataQueue_15_deq_bits = _readData_readDataQueue_fifo_15_empty ? readData_readDataQueue_15_enq_bits : _readData_readDataQueue_fifo_15_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_15 = {write1HPipe_1[15], write1HPipe_0[15]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_15 = {write1HPipe_3[15], write1HPipe_2[15]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_15 = {readData_readResultSelect_lo_lo_lo_hi_15, readData_readResultSelect_lo_lo_lo_lo_15};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_15 = {write1HPipe_5[15], write1HPipe_4[15]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_15 = {write1HPipe_7[15], write1HPipe_6[15]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_15 = {readData_readResultSelect_lo_lo_hi_hi_15, readData_readResultSelect_lo_lo_hi_lo_15};
  wire [7:0]         readData_readResultSelect_lo_lo_15 = {readData_readResultSelect_lo_lo_hi_15, readData_readResultSelect_lo_lo_lo_15};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_15 = {write1HPipe_9[15], write1HPipe_8[15]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_15 = {write1HPipe_11[15], write1HPipe_10[15]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_15 = {readData_readResultSelect_lo_hi_lo_hi_15, readData_readResultSelect_lo_hi_lo_lo_15};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_15 = {write1HPipe_13[15], write1HPipe_12[15]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_15 = {write1HPipe_15[15], write1HPipe_14[15]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_15 = {readData_readResultSelect_lo_hi_hi_hi_15, readData_readResultSelect_lo_hi_hi_lo_15};
  wire [7:0]         readData_readResultSelect_lo_hi_15 = {readData_readResultSelect_lo_hi_hi_15, readData_readResultSelect_lo_hi_lo_15};
  wire [15:0]        readData_readResultSelect_lo_15 = {readData_readResultSelect_lo_hi_15, readData_readResultSelect_lo_lo_15};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_15 = {write1HPipe_17[15], write1HPipe_16[15]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_15 = {write1HPipe_19[15], write1HPipe_18[15]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_15 = {readData_readResultSelect_hi_lo_lo_hi_15, readData_readResultSelect_hi_lo_lo_lo_15};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_15 = {write1HPipe_21[15], write1HPipe_20[15]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_15 = {write1HPipe_23[15], write1HPipe_22[15]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_15 = {readData_readResultSelect_hi_lo_hi_hi_15, readData_readResultSelect_hi_lo_hi_lo_15};
  wire [7:0]         readData_readResultSelect_hi_lo_15 = {readData_readResultSelect_hi_lo_hi_15, readData_readResultSelect_hi_lo_lo_15};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_15 = {write1HPipe_25[15], write1HPipe_24[15]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_15 = {write1HPipe_27[15], write1HPipe_26[15]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_15 = {readData_readResultSelect_hi_hi_lo_hi_15, readData_readResultSelect_hi_hi_lo_lo_15};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_15 = {write1HPipe_29[15], write1HPipe_28[15]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_15 = {write1HPipe_31[15], write1HPipe_30[15]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_15 = {readData_readResultSelect_hi_hi_hi_hi_15, readData_readResultSelect_hi_hi_hi_lo_15};
  wire [7:0]         readData_readResultSelect_hi_hi_15 = {readData_readResultSelect_hi_hi_hi_15, readData_readResultSelect_hi_hi_lo_15};
  wire [15:0]        readData_readResultSelect_hi_15 = {readData_readResultSelect_hi_hi_15, readData_readResultSelect_hi_lo_15};
  wire [31:0]        readData_readResultSelect_15 = {readData_readResultSelect_hi_15, readData_readResultSelect_lo_15};
  assign readData_data_15 =
    (readData_readResultSelect_15[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_15[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_15[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_15[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_15[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_15[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_15[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_15[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_15[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_15[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_15[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_15[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_15[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_15[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_15[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_15[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_15[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_15[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_15[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_15[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_15[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_15[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_15[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_15[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_15[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_15[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_15[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_15[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_15[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_15[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_15[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_15[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_15_enq_bits = readData_data_15;
  wire               readTokenRelease_15 = readData_readDataQueue_15_deq_ready & readData_readDataQueue_15_deq_valid;
  assign readData_readDataQueue_15_enq_valid = |readData_readResultSelect_15;
  wire [31:0]        readData_data_16;
  wire               isWaiteForThisData_16;
  wire               readData_readDataQueue_16_enq_ready = ~_readData_readDataQueue_fifo_16_full;
  wire               readData_readDataQueue_16_deq_ready;
  wire               readData_readDataQueue_16_enq_valid;
  wire               readData_readDataQueue_16_deq_valid = ~_readData_readDataQueue_fifo_16_empty | readData_readDataQueue_16_enq_valid;
  wire [31:0]        readData_readDataQueue_16_enq_bits;
  wire [31:0]        readData_readDataQueue_16_deq_bits = _readData_readDataQueue_fifo_16_empty ? readData_readDataQueue_16_enq_bits : _readData_readDataQueue_fifo_16_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_16 = {write1HPipe_1[16], write1HPipe_0[16]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_16 = {write1HPipe_3[16], write1HPipe_2[16]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_16 = {readData_readResultSelect_lo_lo_lo_hi_16, readData_readResultSelect_lo_lo_lo_lo_16};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_16 = {write1HPipe_5[16], write1HPipe_4[16]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_16 = {write1HPipe_7[16], write1HPipe_6[16]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_16 = {readData_readResultSelect_lo_lo_hi_hi_16, readData_readResultSelect_lo_lo_hi_lo_16};
  wire [7:0]         readData_readResultSelect_lo_lo_16 = {readData_readResultSelect_lo_lo_hi_16, readData_readResultSelect_lo_lo_lo_16};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_16 = {write1HPipe_9[16], write1HPipe_8[16]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_16 = {write1HPipe_11[16], write1HPipe_10[16]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_16 = {readData_readResultSelect_lo_hi_lo_hi_16, readData_readResultSelect_lo_hi_lo_lo_16};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_16 = {write1HPipe_13[16], write1HPipe_12[16]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_16 = {write1HPipe_15[16], write1HPipe_14[16]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_16 = {readData_readResultSelect_lo_hi_hi_hi_16, readData_readResultSelect_lo_hi_hi_lo_16};
  wire [7:0]         readData_readResultSelect_lo_hi_16 = {readData_readResultSelect_lo_hi_hi_16, readData_readResultSelect_lo_hi_lo_16};
  wire [15:0]        readData_readResultSelect_lo_16 = {readData_readResultSelect_lo_hi_16, readData_readResultSelect_lo_lo_16};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_16 = {write1HPipe_17[16], write1HPipe_16[16]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_16 = {write1HPipe_19[16], write1HPipe_18[16]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_16 = {readData_readResultSelect_hi_lo_lo_hi_16, readData_readResultSelect_hi_lo_lo_lo_16};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_16 = {write1HPipe_21[16], write1HPipe_20[16]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_16 = {write1HPipe_23[16], write1HPipe_22[16]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_16 = {readData_readResultSelect_hi_lo_hi_hi_16, readData_readResultSelect_hi_lo_hi_lo_16};
  wire [7:0]         readData_readResultSelect_hi_lo_16 = {readData_readResultSelect_hi_lo_hi_16, readData_readResultSelect_hi_lo_lo_16};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_16 = {write1HPipe_25[16], write1HPipe_24[16]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_16 = {write1HPipe_27[16], write1HPipe_26[16]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_16 = {readData_readResultSelect_hi_hi_lo_hi_16, readData_readResultSelect_hi_hi_lo_lo_16};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_16 = {write1HPipe_29[16], write1HPipe_28[16]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_16 = {write1HPipe_31[16], write1HPipe_30[16]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_16 = {readData_readResultSelect_hi_hi_hi_hi_16, readData_readResultSelect_hi_hi_hi_lo_16};
  wire [7:0]         readData_readResultSelect_hi_hi_16 = {readData_readResultSelect_hi_hi_hi_16, readData_readResultSelect_hi_hi_lo_16};
  wire [15:0]        readData_readResultSelect_hi_16 = {readData_readResultSelect_hi_hi_16, readData_readResultSelect_hi_lo_16};
  wire [31:0]        readData_readResultSelect_16 = {readData_readResultSelect_hi_16, readData_readResultSelect_lo_16};
  assign readData_data_16 =
    (readData_readResultSelect_16[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_16[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_16[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_16[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_16[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_16[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_16[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_16[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_16[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_16[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_16[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_16[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_16[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_16[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_16[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_16[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_16[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_16[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_16[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_16[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_16[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_16[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_16[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_16[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_16[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_16[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_16[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_16[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_16[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_16[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_16[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_16[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_16_enq_bits = readData_data_16;
  wire               readTokenRelease_16 = readData_readDataQueue_16_deq_ready & readData_readDataQueue_16_deq_valid;
  assign readData_readDataQueue_16_enq_valid = |readData_readResultSelect_16;
  wire [31:0]        readData_data_17;
  wire               isWaiteForThisData_17;
  wire               readData_readDataQueue_17_enq_ready = ~_readData_readDataQueue_fifo_17_full;
  wire               readData_readDataQueue_17_deq_ready;
  wire               readData_readDataQueue_17_enq_valid;
  wire               readData_readDataQueue_17_deq_valid = ~_readData_readDataQueue_fifo_17_empty | readData_readDataQueue_17_enq_valid;
  wire [31:0]        readData_readDataQueue_17_enq_bits;
  wire [31:0]        readData_readDataQueue_17_deq_bits = _readData_readDataQueue_fifo_17_empty ? readData_readDataQueue_17_enq_bits : _readData_readDataQueue_fifo_17_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_17 = {write1HPipe_1[17], write1HPipe_0[17]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_17 = {write1HPipe_3[17], write1HPipe_2[17]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_17 = {readData_readResultSelect_lo_lo_lo_hi_17, readData_readResultSelect_lo_lo_lo_lo_17};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_17 = {write1HPipe_5[17], write1HPipe_4[17]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_17 = {write1HPipe_7[17], write1HPipe_6[17]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_17 = {readData_readResultSelect_lo_lo_hi_hi_17, readData_readResultSelect_lo_lo_hi_lo_17};
  wire [7:0]         readData_readResultSelect_lo_lo_17 = {readData_readResultSelect_lo_lo_hi_17, readData_readResultSelect_lo_lo_lo_17};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_17 = {write1HPipe_9[17], write1HPipe_8[17]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_17 = {write1HPipe_11[17], write1HPipe_10[17]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_17 = {readData_readResultSelect_lo_hi_lo_hi_17, readData_readResultSelect_lo_hi_lo_lo_17};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_17 = {write1HPipe_13[17], write1HPipe_12[17]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_17 = {write1HPipe_15[17], write1HPipe_14[17]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_17 = {readData_readResultSelect_lo_hi_hi_hi_17, readData_readResultSelect_lo_hi_hi_lo_17};
  wire [7:0]         readData_readResultSelect_lo_hi_17 = {readData_readResultSelect_lo_hi_hi_17, readData_readResultSelect_lo_hi_lo_17};
  wire [15:0]        readData_readResultSelect_lo_17 = {readData_readResultSelect_lo_hi_17, readData_readResultSelect_lo_lo_17};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_17 = {write1HPipe_17[17], write1HPipe_16[17]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_17 = {write1HPipe_19[17], write1HPipe_18[17]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_17 = {readData_readResultSelect_hi_lo_lo_hi_17, readData_readResultSelect_hi_lo_lo_lo_17};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_17 = {write1HPipe_21[17], write1HPipe_20[17]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_17 = {write1HPipe_23[17], write1HPipe_22[17]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_17 = {readData_readResultSelect_hi_lo_hi_hi_17, readData_readResultSelect_hi_lo_hi_lo_17};
  wire [7:0]         readData_readResultSelect_hi_lo_17 = {readData_readResultSelect_hi_lo_hi_17, readData_readResultSelect_hi_lo_lo_17};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_17 = {write1HPipe_25[17], write1HPipe_24[17]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_17 = {write1HPipe_27[17], write1HPipe_26[17]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_17 = {readData_readResultSelect_hi_hi_lo_hi_17, readData_readResultSelect_hi_hi_lo_lo_17};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_17 = {write1HPipe_29[17], write1HPipe_28[17]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_17 = {write1HPipe_31[17], write1HPipe_30[17]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_17 = {readData_readResultSelect_hi_hi_hi_hi_17, readData_readResultSelect_hi_hi_hi_lo_17};
  wire [7:0]         readData_readResultSelect_hi_hi_17 = {readData_readResultSelect_hi_hi_hi_17, readData_readResultSelect_hi_hi_lo_17};
  wire [15:0]        readData_readResultSelect_hi_17 = {readData_readResultSelect_hi_hi_17, readData_readResultSelect_hi_lo_17};
  wire [31:0]        readData_readResultSelect_17 = {readData_readResultSelect_hi_17, readData_readResultSelect_lo_17};
  assign readData_data_17 =
    (readData_readResultSelect_17[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_17[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_17[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_17[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_17[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_17[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_17[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_17[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_17[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_17[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_17[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_17[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_17[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_17[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_17[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_17[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_17[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_17[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_17[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_17[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_17[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_17[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_17[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_17[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_17[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_17[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_17[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_17[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_17[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_17[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_17[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_17[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_17_enq_bits = readData_data_17;
  wire               readTokenRelease_17 = readData_readDataQueue_17_deq_ready & readData_readDataQueue_17_deq_valid;
  assign readData_readDataQueue_17_enq_valid = |readData_readResultSelect_17;
  wire [31:0]        readData_data_18;
  wire               isWaiteForThisData_18;
  wire               readData_readDataQueue_18_enq_ready = ~_readData_readDataQueue_fifo_18_full;
  wire               readData_readDataQueue_18_deq_ready;
  wire               readData_readDataQueue_18_enq_valid;
  wire               readData_readDataQueue_18_deq_valid = ~_readData_readDataQueue_fifo_18_empty | readData_readDataQueue_18_enq_valid;
  wire [31:0]        readData_readDataQueue_18_enq_bits;
  wire [31:0]        readData_readDataQueue_18_deq_bits = _readData_readDataQueue_fifo_18_empty ? readData_readDataQueue_18_enq_bits : _readData_readDataQueue_fifo_18_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_18 = {write1HPipe_1[18], write1HPipe_0[18]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_18 = {write1HPipe_3[18], write1HPipe_2[18]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_18 = {readData_readResultSelect_lo_lo_lo_hi_18, readData_readResultSelect_lo_lo_lo_lo_18};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_18 = {write1HPipe_5[18], write1HPipe_4[18]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_18 = {write1HPipe_7[18], write1HPipe_6[18]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_18 = {readData_readResultSelect_lo_lo_hi_hi_18, readData_readResultSelect_lo_lo_hi_lo_18};
  wire [7:0]         readData_readResultSelect_lo_lo_18 = {readData_readResultSelect_lo_lo_hi_18, readData_readResultSelect_lo_lo_lo_18};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_18 = {write1HPipe_9[18], write1HPipe_8[18]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_18 = {write1HPipe_11[18], write1HPipe_10[18]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_18 = {readData_readResultSelect_lo_hi_lo_hi_18, readData_readResultSelect_lo_hi_lo_lo_18};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_18 = {write1HPipe_13[18], write1HPipe_12[18]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_18 = {write1HPipe_15[18], write1HPipe_14[18]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_18 = {readData_readResultSelect_lo_hi_hi_hi_18, readData_readResultSelect_lo_hi_hi_lo_18};
  wire [7:0]         readData_readResultSelect_lo_hi_18 = {readData_readResultSelect_lo_hi_hi_18, readData_readResultSelect_lo_hi_lo_18};
  wire [15:0]        readData_readResultSelect_lo_18 = {readData_readResultSelect_lo_hi_18, readData_readResultSelect_lo_lo_18};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_18 = {write1HPipe_17[18], write1HPipe_16[18]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_18 = {write1HPipe_19[18], write1HPipe_18[18]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_18 = {readData_readResultSelect_hi_lo_lo_hi_18, readData_readResultSelect_hi_lo_lo_lo_18};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_18 = {write1HPipe_21[18], write1HPipe_20[18]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_18 = {write1HPipe_23[18], write1HPipe_22[18]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_18 = {readData_readResultSelect_hi_lo_hi_hi_18, readData_readResultSelect_hi_lo_hi_lo_18};
  wire [7:0]         readData_readResultSelect_hi_lo_18 = {readData_readResultSelect_hi_lo_hi_18, readData_readResultSelect_hi_lo_lo_18};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_18 = {write1HPipe_25[18], write1HPipe_24[18]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_18 = {write1HPipe_27[18], write1HPipe_26[18]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_18 = {readData_readResultSelect_hi_hi_lo_hi_18, readData_readResultSelect_hi_hi_lo_lo_18};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_18 = {write1HPipe_29[18], write1HPipe_28[18]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_18 = {write1HPipe_31[18], write1HPipe_30[18]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_18 = {readData_readResultSelect_hi_hi_hi_hi_18, readData_readResultSelect_hi_hi_hi_lo_18};
  wire [7:0]         readData_readResultSelect_hi_hi_18 = {readData_readResultSelect_hi_hi_hi_18, readData_readResultSelect_hi_hi_lo_18};
  wire [15:0]        readData_readResultSelect_hi_18 = {readData_readResultSelect_hi_hi_18, readData_readResultSelect_hi_lo_18};
  wire [31:0]        readData_readResultSelect_18 = {readData_readResultSelect_hi_18, readData_readResultSelect_lo_18};
  assign readData_data_18 =
    (readData_readResultSelect_18[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_18[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_18[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_18[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_18[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_18[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_18[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_18[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_18[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_18[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_18[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_18[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_18[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_18[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_18[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_18[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_18[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_18[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_18[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_18[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_18[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_18[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_18[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_18[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_18[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_18[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_18[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_18[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_18[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_18[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_18[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_18[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_18_enq_bits = readData_data_18;
  wire               readTokenRelease_18 = readData_readDataQueue_18_deq_ready & readData_readDataQueue_18_deq_valid;
  assign readData_readDataQueue_18_enq_valid = |readData_readResultSelect_18;
  wire [31:0]        readData_data_19;
  wire               isWaiteForThisData_19;
  wire               readData_readDataQueue_19_enq_ready = ~_readData_readDataQueue_fifo_19_full;
  wire               readData_readDataQueue_19_deq_ready;
  wire               readData_readDataQueue_19_enq_valid;
  wire               readData_readDataQueue_19_deq_valid = ~_readData_readDataQueue_fifo_19_empty | readData_readDataQueue_19_enq_valid;
  wire [31:0]        readData_readDataQueue_19_enq_bits;
  wire [31:0]        readData_readDataQueue_19_deq_bits = _readData_readDataQueue_fifo_19_empty ? readData_readDataQueue_19_enq_bits : _readData_readDataQueue_fifo_19_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_19 = {write1HPipe_1[19], write1HPipe_0[19]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_19 = {write1HPipe_3[19], write1HPipe_2[19]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_19 = {readData_readResultSelect_lo_lo_lo_hi_19, readData_readResultSelect_lo_lo_lo_lo_19};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_19 = {write1HPipe_5[19], write1HPipe_4[19]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_19 = {write1HPipe_7[19], write1HPipe_6[19]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_19 = {readData_readResultSelect_lo_lo_hi_hi_19, readData_readResultSelect_lo_lo_hi_lo_19};
  wire [7:0]         readData_readResultSelect_lo_lo_19 = {readData_readResultSelect_lo_lo_hi_19, readData_readResultSelect_lo_lo_lo_19};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_19 = {write1HPipe_9[19], write1HPipe_8[19]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_19 = {write1HPipe_11[19], write1HPipe_10[19]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_19 = {readData_readResultSelect_lo_hi_lo_hi_19, readData_readResultSelect_lo_hi_lo_lo_19};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_19 = {write1HPipe_13[19], write1HPipe_12[19]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_19 = {write1HPipe_15[19], write1HPipe_14[19]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_19 = {readData_readResultSelect_lo_hi_hi_hi_19, readData_readResultSelect_lo_hi_hi_lo_19};
  wire [7:0]         readData_readResultSelect_lo_hi_19 = {readData_readResultSelect_lo_hi_hi_19, readData_readResultSelect_lo_hi_lo_19};
  wire [15:0]        readData_readResultSelect_lo_19 = {readData_readResultSelect_lo_hi_19, readData_readResultSelect_lo_lo_19};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_19 = {write1HPipe_17[19], write1HPipe_16[19]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_19 = {write1HPipe_19[19], write1HPipe_18[19]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_19 = {readData_readResultSelect_hi_lo_lo_hi_19, readData_readResultSelect_hi_lo_lo_lo_19};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_19 = {write1HPipe_21[19], write1HPipe_20[19]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_19 = {write1HPipe_23[19], write1HPipe_22[19]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_19 = {readData_readResultSelect_hi_lo_hi_hi_19, readData_readResultSelect_hi_lo_hi_lo_19};
  wire [7:0]         readData_readResultSelect_hi_lo_19 = {readData_readResultSelect_hi_lo_hi_19, readData_readResultSelect_hi_lo_lo_19};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_19 = {write1HPipe_25[19], write1HPipe_24[19]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_19 = {write1HPipe_27[19], write1HPipe_26[19]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_19 = {readData_readResultSelect_hi_hi_lo_hi_19, readData_readResultSelect_hi_hi_lo_lo_19};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_19 = {write1HPipe_29[19], write1HPipe_28[19]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_19 = {write1HPipe_31[19], write1HPipe_30[19]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_19 = {readData_readResultSelect_hi_hi_hi_hi_19, readData_readResultSelect_hi_hi_hi_lo_19};
  wire [7:0]         readData_readResultSelect_hi_hi_19 = {readData_readResultSelect_hi_hi_hi_19, readData_readResultSelect_hi_hi_lo_19};
  wire [15:0]        readData_readResultSelect_hi_19 = {readData_readResultSelect_hi_hi_19, readData_readResultSelect_hi_lo_19};
  wire [31:0]        readData_readResultSelect_19 = {readData_readResultSelect_hi_19, readData_readResultSelect_lo_19};
  assign readData_data_19 =
    (readData_readResultSelect_19[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_19[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_19[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_19[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_19[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_19[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_19[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_19[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_19[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_19[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_19[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_19[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_19[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_19[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_19[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_19[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_19[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_19[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_19[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_19[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_19[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_19[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_19[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_19[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_19[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_19[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_19[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_19[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_19[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_19[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_19[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_19[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_19_enq_bits = readData_data_19;
  wire               readTokenRelease_19 = readData_readDataQueue_19_deq_ready & readData_readDataQueue_19_deq_valid;
  assign readData_readDataQueue_19_enq_valid = |readData_readResultSelect_19;
  wire [31:0]        readData_data_20;
  wire               isWaiteForThisData_20;
  wire               readData_readDataQueue_20_enq_ready = ~_readData_readDataQueue_fifo_20_full;
  wire               readData_readDataQueue_20_deq_ready;
  wire               readData_readDataQueue_20_enq_valid;
  wire               readData_readDataQueue_20_deq_valid = ~_readData_readDataQueue_fifo_20_empty | readData_readDataQueue_20_enq_valid;
  wire [31:0]        readData_readDataQueue_20_enq_bits;
  wire [31:0]        readData_readDataQueue_20_deq_bits = _readData_readDataQueue_fifo_20_empty ? readData_readDataQueue_20_enq_bits : _readData_readDataQueue_fifo_20_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_20 = {write1HPipe_1[20], write1HPipe_0[20]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_20 = {write1HPipe_3[20], write1HPipe_2[20]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_20 = {readData_readResultSelect_lo_lo_lo_hi_20, readData_readResultSelect_lo_lo_lo_lo_20};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_20 = {write1HPipe_5[20], write1HPipe_4[20]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_20 = {write1HPipe_7[20], write1HPipe_6[20]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_20 = {readData_readResultSelect_lo_lo_hi_hi_20, readData_readResultSelect_lo_lo_hi_lo_20};
  wire [7:0]         readData_readResultSelect_lo_lo_20 = {readData_readResultSelect_lo_lo_hi_20, readData_readResultSelect_lo_lo_lo_20};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_20 = {write1HPipe_9[20], write1HPipe_8[20]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_20 = {write1HPipe_11[20], write1HPipe_10[20]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_20 = {readData_readResultSelect_lo_hi_lo_hi_20, readData_readResultSelect_lo_hi_lo_lo_20};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_20 = {write1HPipe_13[20], write1HPipe_12[20]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_20 = {write1HPipe_15[20], write1HPipe_14[20]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_20 = {readData_readResultSelect_lo_hi_hi_hi_20, readData_readResultSelect_lo_hi_hi_lo_20};
  wire [7:0]         readData_readResultSelect_lo_hi_20 = {readData_readResultSelect_lo_hi_hi_20, readData_readResultSelect_lo_hi_lo_20};
  wire [15:0]        readData_readResultSelect_lo_20 = {readData_readResultSelect_lo_hi_20, readData_readResultSelect_lo_lo_20};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_20 = {write1HPipe_17[20], write1HPipe_16[20]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_20 = {write1HPipe_19[20], write1HPipe_18[20]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_20 = {readData_readResultSelect_hi_lo_lo_hi_20, readData_readResultSelect_hi_lo_lo_lo_20};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_20 = {write1HPipe_21[20], write1HPipe_20[20]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_20 = {write1HPipe_23[20], write1HPipe_22[20]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_20 = {readData_readResultSelect_hi_lo_hi_hi_20, readData_readResultSelect_hi_lo_hi_lo_20};
  wire [7:0]         readData_readResultSelect_hi_lo_20 = {readData_readResultSelect_hi_lo_hi_20, readData_readResultSelect_hi_lo_lo_20};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_20 = {write1HPipe_25[20], write1HPipe_24[20]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_20 = {write1HPipe_27[20], write1HPipe_26[20]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_20 = {readData_readResultSelect_hi_hi_lo_hi_20, readData_readResultSelect_hi_hi_lo_lo_20};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_20 = {write1HPipe_29[20], write1HPipe_28[20]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_20 = {write1HPipe_31[20], write1HPipe_30[20]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_20 = {readData_readResultSelect_hi_hi_hi_hi_20, readData_readResultSelect_hi_hi_hi_lo_20};
  wire [7:0]         readData_readResultSelect_hi_hi_20 = {readData_readResultSelect_hi_hi_hi_20, readData_readResultSelect_hi_hi_lo_20};
  wire [15:0]        readData_readResultSelect_hi_20 = {readData_readResultSelect_hi_hi_20, readData_readResultSelect_hi_lo_20};
  wire [31:0]        readData_readResultSelect_20 = {readData_readResultSelect_hi_20, readData_readResultSelect_lo_20};
  assign readData_data_20 =
    (readData_readResultSelect_20[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_20[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_20[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_20[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_20[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_20[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_20[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_20[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_20[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_20[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_20[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_20[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_20[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_20[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_20[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_20[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_20[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_20[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_20[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_20[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_20[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_20[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_20[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_20[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_20[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_20[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_20[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_20[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_20[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_20[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_20[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_20[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_20_enq_bits = readData_data_20;
  wire               readTokenRelease_20 = readData_readDataQueue_20_deq_ready & readData_readDataQueue_20_deq_valid;
  assign readData_readDataQueue_20_enq_valid = |readData_readResultSelect_20;
  wire [31:0]        readData_data_21;
  wire               isWaiteForThisData_21;
  wire               readData_readDataQueue_21_enq_ready = ~_readData_readDataQueue_fifo_21_full;
  wire               readData_readDataQueue_21_deq_ready;
  wire               readData_readDataQueue_21_enq_valid;
  wire               readData_readDataQueue_21_deq_valid = ~_readData_readDataQueue_fifo_21_empty | readData_readDataQueue_21_enq_valid;
  wire [31:0]        readData_readDataQueue_21_enq_bits;
  wire [31:0]        readData_readDataQueue_21_deq_bits = _readData_readDataQueue_fifo_21_empty ? readData_readDataQueue_21_enq_bits : _readData_readDataQueue_fifo_21_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_21 = {write1HPipe_1[21], write1HPipe_0[21]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_21 = {write1HPipe_3[21], write1HPipe_2[21]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_21 = {readData_readResultSelect_lo_lo_lo_hi_21, readData_readResultSelect_lo_lo_lo_lo_21};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_21 = {write1HPipe_5[21], write1HPipe_4[21]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_21 = {write1HPipe_7[21], write1HPipe_6[21]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_21 = {readData_readResultSelect_lo_lo_hi_hi_21, readData_readResultSelect_lo_lo_hi_lo_21};
  wire [7:0]         readData_readResultSelect_lo_lo_21 = {readData_readResultSelect_lo_lo_hi_21, readData_readResultSelect_lo_lo_lo_21};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_21 = {write1HPipe_9[21], write1HPipe_8[21]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_21 = {write1HPipe_11[21], write1HPipe_10[21]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_21 = {readData_readResultSelect_lo_hi_lo_hi_21, readData_readResultSelect_lo_hi_lo_lo_21};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_21 = {write1HPipe_13[21], write1HPipe_12[21]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_21 = {write1HPipe_15[21], write1HPipe_14[21]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_21 = {readData_readResultSelect_lo_hi_hi_hi_21, readData_readResultSelect_lo_hi_hi_lo_21};
  wire [7:0]         readData_readResultSelect_lo_hi_21 = {readData_readResultSelect_lo_hi_hi_21, readData_readResultSelect_lo_hi_lo_21};
  wire [15:0]        readData_readResultSelect_lo_21 = {readData_readResultSelect_lo_hi_21, readData_readResultSelect_lo_lo_21};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_21 = {write1HPipe_17[21], write1HPipe_16[21]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_21 = {write1HPipe_19[21], write1HPipe_18[21]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_21 = {readData_readResultSelect_hi_lo_lo_hi_21, readData_readResultSelect_hi_lo_lo_lo_21};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_21 = {write1HPipe_21[21], write1HPipe_20[21]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_21 = {write1HPipe_23[21], write1HPipe_22[21]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_21 = {readData_readResultSelect_hi_lo_hi_hi_21, readData_readResultSelect_hi_lo_hi_lo_21};
  wire [7:0]         readData_readResultSelect_hi_lo_21 = {readData_readResultSelect_hi_lo_hi_21, readData_readResultSelect_hi_lo_lo_21};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_21 = {write1HPipe_25[21], write1HPipe_24[21]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_21 = {write1HPipe_27[21], write1HPipe_26[21]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_21 = {readData_readResultSelect_hi_hi_lo_hi_21, readData_readResultSelect_hi_hi_lo_lo_21};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_21 = {write1HPipe_29[21], write1HPipe_28[21]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_21 = {write1HPipe_31[21], write1HPipe_30[21]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_21 = {readData_readResultSelect_hi_hi_hi_hi_21, readData_readResultSelect_hi_hi_hi_lo_21};
  wire [7:0]         readData_readResultSelect_hi_hi_21 = {readData_readResultSelect_hi_hi_hi_21, readData_readResultSelect_hi_hi_lo_21};
  wire [15:0]        readData_readResultSelect_hi_21 = {readData_readResultSelect_hi_hi_21, readData_readResultSelect_hi_lo_21};
  wire [31:0]        readData_readResultSelect_21 = {readData_readResultSelect_hi_21, readData_readResultSelect_lo_21};
  assign readData_data_21 =
    (readData_readResultSelect_21[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_21[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_21[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_21[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_21[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_21[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_21[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_21[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_21[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_21[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_21[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_21[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_21[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_21[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_21[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_21[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_21[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_21[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_21[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_21[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_21[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_21[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_21[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_21[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_21[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_21[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_21[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_21[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_21[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_21[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_21[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_21[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_21_enq_bits = readData_data_21;
  wire               readTokenRelease_21 = readData_readDataQueue_21_deq_ready & readData_readDataQueue_21_deq_valid;
  assign readData_readDataQueue_21_enq_valid = |readData_readResultSelect_21;
  wire [31:0]        readData_data_22;
  wire               isWaiteForThisData_22;
  wire               readData_readDataQueue_22_enq_ready = ~_readData_readDataQueue_fifo_22_full;
  wire               readData_readDataQueue_22_deq_ready;
  wire               readData_readDataQueue_22_enq_valid;
  wire               readData_readDataQueue_22_deq_valid = ~_readData_readDataQueue_fifo_22_empty | readData_readDataQueue_22_enq_valid;
  wire [31:0]        readData_readDataQueue_22_enq_bits;
  wire [31:0]        readData_readDataQueue_22_deq_bits = _readData_readDataQueue_fifo_22_empty ? readData_readDataQueue_22_enq_bits : _readData_readDataQueue_fifo_22_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_22 = {write1HPipe_1[22], write1HPipe_0[22]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_22 = {write1HPipe_3[22], write1HPipe_2[22]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_22 = {readData_readResultSelect_lo_lo_lo_hi_22, readData_readResultSelect_lo_lo_lo_lo_22};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_22 = {write1HPipe_5[22], write1HPipe_4[22]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_22 = {write1HPipe_7[22], write1HPipe_6[22]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_22 = {readData_readResultSelect_lo_lo_hi_hi_22, readData_readResultSelect_lo_lo_hi_lo_22};
  wire [7:0]         readData_readResultSelect_lo_lo_22 = {readData_readResultSelect_lo_lo_hi_22, readData_readResultSelect_lo_lo_lo_22};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_22 = {write1HPipe_9[22], write1HPipe_8[22]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_22 = {write1HPipe_11[22], write1HPipe_10[22]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_22 = {readData_readResultSelect_lo_hi_lo_hi_22, readData_readResultSelect_lo_hi_lo_lo_22};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_22 = {write1HPipe_13[22], write1HPipe_12[22]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_22 = {write1HPipe_15[22], write1HPipe_14[22]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_22 = {readData_readResultSelect_lo_hi_hi_hi_22, readData_readResultSelect_lo_hi_hi_lo_22};
  wire [7:0]         readData_readResultSelect_lo_hi_22 = {readData_readResultSelect_lo_hi_hi_22, readData_readResultSelect_lo_hi_lo_22};
  wire [15:0]        readData_readResultSelect_lo_22 = {readData_readResultSelect_lo_hi_22, readData_readResultSelect_lo_lo_22};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_22 = {write1HPipe_17[22], write1HPipe_16[22]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_22 = {write1HPipe_19[22], write1HPipe_18[22]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_22 = {readData_readResultSelect_hi_lo_lo_hi_22, readData_readResultSelect_hi_lo_lo_lo_22};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_22 = {write1HPipe_21[22], write1HPipe_20[22]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_22 = {write1HPipe_23[22], write1HPipe_22[22]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_22 = {readData_readResultSelect_hi_lo_hi_hi_22, readData_readResultSelect_hi_lo_hi_lo_22};
  wire [7:0]         readData_readResultSelect_hi_lo_22 = {readData_readResultSelect_hi_lo_hi_22, readData_readResultSelect_hi_lo_lo_22};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_22 = {write1HPipe_25[22], write1HPipe_24[22]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_22 = {write1HPipe_27[22], write1HPipe_26[22]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_22 = {readData_readResultSelect_hi_hi_lo_hi_22, readData_readResultSelect_hi_hi_lo_lo_22};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_22 = {write1HPipe_29[22], write1HPipe_28[22]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_22 = {write1HPipe_31[22], write1HPipe_30[22]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_22 = {readData_readResultSelect_hi_hi_hi_hi_22, readData_readResultSelect_hi_hi_hi_lo_22};
  wire [7:0]         readData_readResultSelect_hi_hi_22 = {readData_readResultSelect_hi_hi_hi_22, readData_readResultSelect_hi_hi_lo_22};
  wire [15:0]        readData_readResultSelect_hi_22 = {readData_readResultSelect_hi_hi_22, readData_readResultSelect_hi_lo_22};
  wire [31:0]        readData_readResultSelect_22 = {readData_readResultSelect_hi_22, readData_readResultSelect_lo_22};
  assign readData_data_22 =
    (readData_readResultSelect_22[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_22[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_22[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_22[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_22[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_22[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_22[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_22[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_22[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_22[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_22[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_22[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_22[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_22[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_22[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_22[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_22[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_22[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_22[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_22[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_22[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_22[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_22[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_22[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_22[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_22[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_22[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_22[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_22[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_22[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_22[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_22[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_22_enq_bits = readData_data_22;
  wire               readTokenRelease_22 = readData_readDataQueue_22_deq_ready & readData_readDataQueue_22_deq_valid;
  assign readData_readDataQueue_22_enq_valid = |readData_readResultSelect_22;
  wire [31:0]        readData_data_23;
  wire               isWaiteForThisData_23;
  wire               readData_readDataQueue_23_enq_ready = ~_readData_readDataQueue_fifo_23_full;
  wire               readData_readDataQueue_23_deq_ready;
  wire               readData_readDataQueue_23_enq_valid;
  wire               readData_readDataQueue_23_deq_valid = ~_readData_readDataQueue_fifo_23_empty | readData_readDataQueue_23_enq_valid;
  wire [31:0]        readData_readDataQueue_23_enq_bits;
  wire [31:0]        readData_readDataQueue_23_deq_bits = _readData_readDataQueue_fifo_23_empty ? readData_readDataQueue_23_enq_bits : _readData_readDataQueue_fifo_23_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_23 = {write1HPipe_1[23], write1HPipe_0[23]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_23 = {write1HPipe_3[23], write1HPipe_2[23]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_23 = {readData_readResultSelect_lo_lo_lo_hi_23, readData_readResultSelect_lo_lo_lo_lo_23};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_23 = {write1HPipe_5[23], write1HPipe_4[23]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_23 = {write1HPipe_7[23], write1HPipe_6[23]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_23 = {readData_readResultSelect_lo_lo_hi_hi_23, readData_readResultSelect_lo_lo_hi_lo_23};
  wire [7:0]         readData_readResultSelect_lo_lo_23 = {readData_readResultSelect_lo_lo_hi_23, readData_readResultSelect_lo_lo_lo_23};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_23 = {write1HPipe_9[23], write1HPipe_8[23]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_23 = {write1HPipe_11[23], write1HPipe_10[23]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_23 = {readData_readResultSelect_lo_hi_lo_hi_23, readData_readResultSelect_lo_hi_lo_lo_23};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_23 = {write1HPipe_13[23], write1HPipe_12[23]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_23 = {write1HPipe_15[23], write1HPipe_14[23]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_23 = {readData_readResultSelect_lo_hi_hi_hi_23, readData_readResultSelect_lo_hi_hi_lo_23};
  wire [7:0]         readData_readResultSelect_lo_hi_23 = {readData_readResultSelect_lo_hi_hi_23, readData_readResultSelect_lo_hi_lo_23};
  wire [15:0]        readData_readResultSelect_lo_23 = {readData_readResultSelect_lo_hi_23, readData_readResultSelect_lo_lo_23};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_23 = {write1HPipe_17[23], write1HPipe_16[23]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_23 = {write1HPipe_19[23], write1HPipe_18[23]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_23 = {readData_readResultSelect_hi_lo_lo_hi_23, readData_readResultSelect_hi_lo_lo_lo_23};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_23 = {write1HPipe_21[23], write1HPipe_20[23]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_23 = {write1HPipe_23[23], write1HPipe_22[23]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_23 = {readData_readResultSelect_hi_lo_hi_hi_23, readData_readResultSelect_hi_lo_hi_lo_23};
  wire [7:0]         readData_readResultSelect_hi_lo_23 = {readData_readResultSelect_hi_lo_hi_23, readData_readResultSelect_hi_lo_lo_23};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_23 = {write1HPipe_25[23], write1HPipe_24[23]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_23 = {write1HPipe_27[23], write1HPipe_26[23]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_23 = {readData_readResultSelect_hi_hi_lo_hi_23, readData_readResultSelect_hi_hi_lo_lo_23};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_23 = {write1HPipe_29[23], write1HPipe_28[23]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_23 = {write1HPipe_31[23], write1HPipe_30[23]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_23 = {readData_readResultSelect_hi_hi_hi_hi_23, readData_readResultSelect_hi_hi_hi_lo_23};
  wire [7:0]         readData_readResultSelect_hi_hi_23 = {readData_readResultSelect_hi_hi_hi_23, readData_readResultSelect_hi_hi_lo_23};
  wire [15:0]        readData_readResultSelect_hi_23 = {readData_readResultSelect_hi_hi_23, readData_readResultSelect_hi_lo_23};
  wire [31:0]        readData_readResultSelect_23 = {readData_readResultSelect_hi_23, readData_readResultSelect_lo_23};
  assign readData_data_23 =
    (readData_readResultSelect_23[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_23[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_23[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_23[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_23[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_23[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_23[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_23[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_23[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_23[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_23[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_23[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_23[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_23[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_23[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_23[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_23[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_23[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_23[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_23[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_23[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_23[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_23[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_23[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_23[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_23[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_23[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_23[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_23[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_23[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_23[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_23[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_23_enq_bits = readData_data_23;
  wire               readTokenRelease_23 = readData_readDataQueue_23_deq_ready & readData_readDataQueue_23_deq_valid;
  assign readData_readDataQueue_23_enq_valid = |readData_readResultSelect_23;
  wire [31:0]        readData_data_24;
  wire               isWaiteForThisData_24;
  wire               readData_readDataQueue_24_enq_ready = ~_readData_readDataQueue_fifo_24_full;
  wire               readData_readDataQueue_24_deq_ready;
  wire               readData_readDataQueue_24_enq_valid;
  wire               readData_readDataQueue_24_deq_valid = ~_readData_readDataQueue_fifo_24_empty | readData_readDataQueue_24_enq_valid;
  wire [31:0]        readData_readDataQueue_24_enq_bits;
  wire [31:0]        readData_readDataQueue_24_deq_bits = _readData_readDataQueue_fifo_24_empty ? readData_readDataQueue_24_enq_bits : _readData_readDataQueue_fifo_24_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_24 = {write1HPipe_1[24], write1HPipe_0[24]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_24 = {write1HPipe_3[24], write1HPipe_2[24]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_24 = {readData_readResultSelect_lo_lo_lo_hi_24, readData_readResultSelect_lo_lo_lo_lo_24};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_24 = {write1HPipe_5[24], write1HPipe_4[24]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_24 = {write1HPipe_7[24], write1HPipe_6[24]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_24 = {readData_readResultSelect_lo_lo_hi_hi_24, readData_readResultSelect_lo_lo_hi_lo_24};
  wire [7:0]         readData_readResultSelect_lo_lo_24 = {readData_readResultSelect_lo_lo_hi_24, readData_readResultSelect_lo_lo_lo_24};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_24 = {write1HPipe_9[24], write1HPipe_8[24]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_24 = {write1HPipe_11[24], write1HPipe_10[24]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_24 = {readData_readResultSelect_lo_hi_lo_hi_24, readData_readResultSelect_lo_hi_lo_lo_24};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_24 = {write1HPipe_13[24], write1HPipe_12[24]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_24 = {write1HPipe_15[24], write1HPipe_14[24]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_24 = {readData_readResultSelect_lo_hi_hi_hi_24, readData_readResultSelect_lo_hi_hi_lo_24};
  wire [7:0]         readData_readResultSelect_lo_hi_24 = {readData_readResultSelect_lo_hi_hi_24, readData_readResultSelect_lo_hi_lo_24};
  wire [15:0]        readData_readResultSelect_lo_24 = {readData_readResultSelect_lo_hi_24, readData_readResultSelect_lo_lo_24};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_24 = {write1HPipe_17[24], write1HPipe_16[24]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_24 = {write1HPipe_19[24], write1HPipe_18[24]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_24 = {readData_readResultSelect_hi_lo_lo_hi_24, readData_readResultSelect_hi_lo_lo_lo_24};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_24 = {write1HPipe_21[24], write1HPipe_20[24]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_24 = {write1HPipe_23[24], write1HPipe_22[24]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_24 = {readData_readResultSelect_hi_lo_hi_hi_24, readData_readResultSelect_hi_lo_hi_lo_24};
  wire [7:0]         readData_readResultSelect_hi_lo_24 = {readData_readResultSelect_hi_lo_hi_24, readData_readResultSelect_hi_lo_lo_24};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_24 = {write1HPipe_25[24], write1HPipe_24[24]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_24 = {write1HPipe_27[24], write1HPipe_26[24]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_24 = {readData_readResultSelect_hi_hi_lo_hi_24, readData_readResultSelect_hi_hi_lo_lo_24};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_24 = {write1HPipe_29[24], write1HPipe_28[24]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_24 = {write1HPipe_31[24], write1HPipe_30[24]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_24 = {readData_readResultSelect_hi_hi_hi_hi_24, readData_readResultSelect_hi_hi_hi_lo_24};
  wire [7:0]         readData_readResultSelect_hi_hi_24 = {readData_readResultSelect_hi_hi_hi_24, readData_readResultSelect_hi_hi_lo_24};
  wire [15:0]        readData_readResultSelect_hi_24 = {readData_readResultSelect_hi_hi_24, readData_readResultSelect_hi_lo_24};
  wire [31:0]        readData_readResultSelect_24 = {readData_readResultSelect_hi_24, readData_readResultSelect_lo_24};
  assign readData_data_24 =
    (readData_readResultSelect_24[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_24[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_24[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_24[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_24[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_24[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_24[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_24[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_24[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_24[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_24[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_24[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_24[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_24[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_24[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_24[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_24[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_24[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_24[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_24[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_24[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_24[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_24[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_24[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_24[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_24[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_24[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_24[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_24[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_24[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_24[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_24[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_24_enq_bits = readData_data_24;
  wire               readTokenRelease_24 = readData_readDataQueue_24_deq_ready & readData_readDataQueue_24_deq_valid;
  assign readData_readDataQueue_24_enq_valid = |readData_readResultSelect_24;
  wire [31:0]        readData_data_25;
  wire               isWaiteForThisData_25;
  wire               readData_readDataQueue_25_enq_ready = ~_readData_readDataQueue_fifo_25_full;
  wire               readData_readDataQueue_25_deq_ready;
  wire               readData_readDataQueue_25_enq_valid;
  wire               readData_readDataQueue_25_deq_valid = ~_readData_readDataQueue_fifo_25_empty | readData_readDataQueue_25_enq_valid;
  wire [31:0]        readData_readDataQueue_25_enq_bits;
  wire [31:0]        readData_readDataQueue_25_deq_bits = _readData_readDataQueue_fifo_25_empty ? readData_readDataQueue_25_enq_bits : _readData_readDataQueue_fifo_25_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_25 = {write1HPipe_1[25], write1HPipe_0[25]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_25 = {write1HPipe_3[25], write1HPipe_2[25]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_25 = {readData_readResultSelect_lo_lo_lo_hi_25, readData_readResultSelect_lo_lo_lo_lo_25};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_25 = {write1HPipe_5[25], write1HPipe_4[25]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_25 = {write1HPipe_7[25], write1HPipe_6[25]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_25 = {readData_readResultSelect_lo_lo_hi_hi_25, readData_readResultSelect_lo_lo_hi_lo_25};
  wire [7:0]         readData_readResultSelect_lo_lo_25 = {readData_readResultSelect_lo_lo_hi_25, readData_readResultSelect_lo_lo_lo_25};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_25 = {write1HPipe_9[25], write1HPipe_8[25]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_25 = {write1HPipe_11[25], write1HPipe_10[25]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_25 = {readData_readResultSelect_lo_hi_lo_hi_25, readData_readResultSelect_lo_hi_lo_lo_25};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_25 = {write1HPipe_13[25], write1HPipe_12[25]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_25 = {write1HPipe_15[25], write1HPipe_14[25]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_25 = {readData_readResultSelect_lo_hi_hi_hi_25, readData_readResultSelect_lo_hi_hi_lo_25};
  wire [7:0]         readData_readResultSelect_lo_hi_25 = {readData_readResultSelect_lo_hi_hi_25, readData_readResultSelect_lo_hi_lo_25};
  wire [15:0]        readData_readResultSelect_lo_25 = {readData_readResultSelect_lo_hi_25, readData_readResultSelect_lo_lo_25};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_25 = {write1HPipe_17[25], write1HPipe_16[25]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_25 = {write1HPipe_19[25], write1HPipe_18[25]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_25 = {readData_readResultSelect_hi_lo_lo_hi_25, readData_readResultSelect_hi_lo_lo_lo_25};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_25 = {write1HPipe_21[25], write1HPipe_20[25]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_25 = {write1HPipe_23[25], write1HPipe_22[25]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_25 = {readData_readResultSelect_hi_lo_hi_hi_25, readData_readResultSelect_hi_lo_hi_lo_25};
  wire [7:0]         readData_readResultSelect_hi_lo_25 = {readData_readResultSelect_hi_lo_hi_25, readData_readResultSelect_hi_lo_lo_25};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_25 = {write1HPipe_25[25], write1HPipe_24[25]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_25 = {write1HPipe_27[25], write1HPipe_26[25]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_25 = {readData_readResultSelect_hi_hi_lo_hi_25, readData_readResultSelect_hi_hi_lo_lo_25};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_25 = {write1HPipe_29[25], write1HPipe_28[25]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_25 = {write1HPipe_31[25], write1HPipe_30[25]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_25 = {readData_readResultSelect_hi_hi_hi_hi_25, readData_readResultSelect_hi_hi_hi_lo_25};
  wire [7:0]         readData_readResultSelect_hi_hi_25 = {readData_readResultSelect_hi_hi_hi_25, readData_readResultSelect_hi_hi_lo_25};
  wire [15:0]        readData_readResultSelect_hi_25 = {readData_readResultSelect_hi_hi_25, readData_readResultSelect_hi_lo_25};
  wire [31:0]        readData_readResultSelect_25 = {readData_readResultSelect_hi_25, readData_readResultSelect_lo_25};
  assign readData_data_25 =
    (readData_readResultSelect_25[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_25[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_25[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_25[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_25[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_25[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_25[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_25[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_25[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_25[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_25[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_25[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_25[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_25[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_25[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_25[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_25[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_25[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_25[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_25[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_25[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_25[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_25[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_25[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_25[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_25[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_25[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_25[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_25[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_25[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_25[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_25[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_25_enq_bits = readData_data_25;
  wire               readTokenRelease_25 = readData_readDataQueue_25_deq_ready & readData_readDataQueue_25_deq_valid;
  assign readData_readDataQueue_25_enq_valid = |readData_readResultSelect_25;
  wire [31:0]        readData_data_26;
  wire               isWaiteForThisData_26;
  wire               readData_readDataQueue_26_enq_ready = ~_readData_readDataQueue_fifo_26_full;
  wire               readData_readDataQueue_26_deq_ready;
  wire               readData_readDataQueue_26_enq_valid;
  wire               readData_readDataQueue_26_deq_valid = ~_readData_readDataQueue_fifo_26_empty | readData_readDataQueue_26_enq_valid;
  wire [31:0]        readData_readDataQueue_26_enq_bits;
  wire [31:0]        readData_readDataQueue_26_deq_bits = _readData_readDataQueue_fifo_26_empty ? readData_readDataQueue_26_enq_bits : _readData_readDataQueue_fifo_26_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_26 = {write1HPipe_1[26], write1HPipe_0[26]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_26 = {write1HPipe_3[26], write1HPipe_2[26]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_26 = {readData_readResultSelect_lo_lo_lo_hi_26, readData_readResultSelect_lo_lo_lo_lo_26};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_26 = {write1HPipe_5[26], write1HPipe_4[26]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_26 = {write1HPipe_7[26], write1HPipe_6[26]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_26 = {readData_readResultSelect_lo_lo_hi_hi_26, readData_readResultSelect_lo_lo_hi_lo_26};
  wire [7:0]         readData_readResultSelect_lo_lo_26 = {readData_readResultSelect_lo_lo_hi_26, readData_readResultSelect_lo_lo_lo_26};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_26 = {write1HPipe_9[26], write1HPipe_8[26]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_26 = {write1HPipe_11[26], write1HPipe_10[26]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_26 = {readData_readResultSelect_lo_hi_lo_hi_26, readData_readResultSelect_lo_hi_lo_lo_26};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_26 = {write1HPipe_13[26], write1HPipe_12[26]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_26 = {write1HPipe_15[26], write1HPipe_14[26]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_26 = {readData_readResultSelect_lo_hi_hi_hi_26, readData_readResultSelect_lo_hi_hi_lo_26};
  wire [7:0]         readData_readResultSelect_lo_hi_26 = {readData_readResultSelect_lo_hi_hi_26, readData_readResultSelect_lo_hi_lo_26};
  wire [15:0]        readData_readResultSelect_lo_26 = {readData_readResultSelect_lo_hi_26, readData_readResultSelect_lo_lo_26};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_26 = {write1HPipe_17[26], write1HPipe_16[26]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_26 = {write1HPipe_19[26], write1HPipe_18[26]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_26 = {readData_readResultSelect_hi_lo_lo_hi_26, readData_readResultSelect_hi_lo_lo_lo_26};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_26 = {write1HPipe_21[26], write1HPipe_20[26]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_26 = {write1HPipe_23[26], write1HPipe_22[26]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_26 = {readData_readResultSelect_hi_lo_hi_hi_26, readData_readResultSelect_hi_lo_hi_lo_26};
  wire [7:0]         readData_readResultSelect_hi_lo_26 = {readData_readResultSelect_hi_lo_hi_26, readData_readResultSelect_hi_lo_lo_26};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_26 = {write1HPipe_25[26], write1HPipe_24[26]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_26 = {write1HPipe_27[26], write1HPipe_26[26]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_26 = {readData_readResultSelect_hi_hi_lo_hi_26, readData_readResultSelect_hi_hi_lo_lo_26};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_26 = {write1HPipe_29[26], write1HPipe_28[26]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_26 = {write1HPipe_31[26], write1HPipe_30[26]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_26 = {readData_readResultSelect_hi_hi_hi_hi_26, readData_readResultSelect_hi_hi_hi_lo_26};
  wire [7:0]         readData_readResultSelect_hi_hi_26 = {readData_readResultSelect_hi_hi_hi_26, readData_readResultSelect_hi_hi_lo_26};
  wire [15:0]        readData_readResultSelect_hi_26 = {readData_readResultSelect_hi_hi_26, readData_readResultSelect_hi_lo_26};
  wire [31:0]        readData_readResultSelect_26 = {readData_readResultSelect_hi_26, readData_readResultSelect_lo_26};
  assign readData_data_26 =
    (readData_readResultSelect_26[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_26[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_26[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_26[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_26[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_26[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_26[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_26[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_26[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_26[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_26[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_26[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_26[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_26[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_26[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_26[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_26[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_26[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_26[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_26[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_26[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_26[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_26[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_26[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_26[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_26[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_26[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_26[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_26[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_26[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_26[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_26[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_26_enq_bits = readData_data_26;
  wire               readTokenRelease_26 = readData_readDataQueue_26_deq_ready & readData_readDataQueue_26_deq_valid;
  assign readData_readDataQueue_26_enq_valid = |readData_readResultSelect_26;
  wire [31:0]        readData_data_27;
  wire               isWaiteForThisData_27;
  wire               readData_readDataQueue_27_enq_ready = ~_readData_readDataQueue_fifo_27_full;
  wire               readData_readDataQueue_27_deq_ready;
  wire               readData_readDataQueue_27_enq_valid;
  wire               readData_readDataQueue_27_deq_valid = ~_readData_readDataQueue_fifo_27_empty | readData_readDataQueue_27_enq_valid;
  wire [31:0]        readData_readDataQueue_27_enq_bits;
  wire [31:0]        readData_readDataQueue_27_deq_bits = _readData_readDataQueue_fifo_27_empty ? readData_readDataQueue_27_enq_bits : _readData_readDataQueue_fifo_27_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_27 = {write1HPipe_1[27], write1HPipe_0[27]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_27 = {write1HPipe_3[27], write1HPipe_2[27]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_27 = {readData_readResultSelect_lo_lo_lo_hi_27, readData_readResultSelect_lo_lo_lo_lo_27};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_27 = {write1HPipe_5[27], write1HPipe_4[27]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_27 = {write1HPipe_7[27], write1HPipe_6[27]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_27 = {readData_readResultSelect_lo_lo_hi_hi_27, readData_readResultSelect_lo_lo_hi_lo_27};
  wire [7:0]         readData_readResultSelect_lo_lo_27 = {readData_readResultSelect_lo_lo_hi_27, readData_readResultSelect_lo_lo_lo_27};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_27 = {write1HPipe_9[27], write1HPipe_8[27]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_27 = {write1HPipe_11[27], write1HPipe_10[27]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_27 = {readData_readResultSelect_lo_hi_lo_hi_27, readData_readResultSelect_lo_hi_lo_lo_27};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_27 = {write1HPipe_13[27], write1HPipe_12[27]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_27 = {write1HPipe_15[27], write1HPipe_14[27]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_27 = {readData_readResultSelect_lo_hi_hi_hi_27, readData_readResultSelect_lo_hi_hi_lo_27};
  wire [7:0]         readData_readResultSelect_lo_hi_27 = {readData_readResultSelect_lo_hi_hi_27, readData_readResultSelect_lo_hi_lo_27};
  wire [15:0]        readData_readResultSelect_lo_27 = {readData_readResultSelect_lo_hi_27, readData_readResultSelect_lo_lo_27};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_27 = {write1HPipe_17[27], write1HPipe_16[27]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_27 = {write1HPipe_19[27], write1HPipe_18[27]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_27 = {readData_readResultSelect_hi_lo_lo_hi_27, readData_readResultSelect_hi_lo_lo_lo_27};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_27 = {write1HPipe_21[27], write1HPipe_20[27]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_27 = {write1HPipe_23[27], write1HPipe_22[27]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_27 = {readData_readResultSelect_hi_lo_hi_hi_27, readData_readResultSelect_hi_lo_hi_lo_27};
  wire [7:0]         readData_readResultSelect_hi_lo_27 = {readData_readResultSelect_hi_lo_hi_27, readData_readResultSelect_hi_lo_lo_27};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_27 = {write1HPipe_25[27], write1HPipe_24[27]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_27 = {write1HPipe_27[27], write1HPipe_26[27]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_27 = {readData_readResultSelect_hi_hi_lo_hi_27, readData_readResultSelect_hi_hi_lo_lo_27};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_27 = {write1HPipe_29[27], write1HPipe_28[27]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_27 = {write1HPipe_31[27], write1HPipe_30[27]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_27 = {readData_readResultSelect_hi_hi_hi_hi_27, readData_readResultSelect_hi_hi_hi_lo_27};
  wire [7:0]         readData_readResultSelect_hi_hi_27 = {readData_readResultSelect_hi_hi_hi_27, readData_readResultSelect_hi_hi_lo_27};
  wire [15:0]        readData_readResultSelect_hi_27 = {readData_readResultSelect_hi_hi_27, readData_readResultSelect_hi_lo_27};
  wire [31:0]        readData_readResultSelect_27 = {readData_readResultSelect_hi_27, readData_readResultSelect_lo_27};
  assign readData_data_27 =
    (readData_readResultSelect_27[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_27[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_27[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_27[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_27[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_27[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_27[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_27[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_27[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_27[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_27[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_27[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_27[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_27[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_27[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_27[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_27[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_27[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_27[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_27[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_27[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_27[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_27[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_27[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_27[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_27[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_27[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_27[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_27[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_27[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_27[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_27[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_27_enq_bits = readData_data_27;
  wire               readTokenRelease_27 = readData_readDataQueue_27_deq_ready & readData_readDataQueue_27_deq_valid;
  assign readData_readDataQueue_27_enq_valid = |readData_readResultSelect_27;
  wire [31:0]        readData_data_28;
  wire               isWaiteForThisData_28;
  wire               readData_readDataQueue_28_enq_ready = ~_readData_readDataQueue_fifo_28_full;
  wire               readData_readDataQueue_28_deq_ready;
  wire               readData_readDataQueue_28_enq_valid;
  wire               readData_readDataQueue_28_deq_valid = ~_readData_readDataQueue_fifo_28_empty | readData_readDataQueue_28_enq_valid;
  wire [31:0]        readData_readDataQueue_28_enq_bits;
  wire [31:0]        readData_readDataQueue_28_deq_bits = _readData_readDataQueue_fifo_28_empty ? readData_readDataQueue_28_enq_bits : _readData_readDataQueue_fifo_28_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_28 = {write1HPipe_1[28], write1HPipe_0[28]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_28 = {write1HPipe_3[28], write1HPipe_2[28]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_28 = {readData_readResultSelect_lo_lo_lo_hi_28, readData_readResultSelect_lo_lo_lo_lo_28};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_28 = {write1HPipe_5[28], write1HPipe_4[28]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_28 = {write1HPipe_7[28], write1HPipe_6[28]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_28 = {readData_readResultSelect_lo_lo_hi_hi_28, readData_readResultSelect_lo_lo_hi_lo_28};
  wire [7:0]         readData_readResultSelect_lo_lo_28 = {readData_readResultSelect_lo_lo_hi_28, readData_readResultSelect_lo_lo_lo_28};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_28 = {write1HPipe_9[28], write1HPipe_8[28]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_28 = {write1HPipe_11[28], write1HPipe_10[28]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_28 = {readData_readResultSelect_lo_hi_lo_hi_28, readData_readResultSelect_lo_hi_lo_lo_28};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_28 = {write1HPipe_13[28], write1HPipe_12[28]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_28 = {write1HPipe_15[28], write1HPipe_14[28]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_28 = {readData_readResultSelect_lo_hi_hi_hi_28, readData_readResultSelect_lo_hi_hi_lo_28};
  wire [7:0]         readData_readResultSelect_lo_hi_28 = {readData_readResultSelect_lo_hi_hi_28, readData_readResultSelect_lo_hi_lo_28};
  wire [15:0]        readData_readResultSelect_lo_28 = {readData_readResultSelect_lo_hi_28, readData_readResultSelect_lo_lo_28};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_28 = {write1HPipe_17[28], write1HPipe_16[28]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_28 = {write1HPipe_19[28], write1HPipe_18[28]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_28 = {readData_readResultSelect_hi_lo_lo_hi_28, readData_readResultSelect_hi_lo_lo_lo_28};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_28 = {write1HPipe_21[28], write1HPipe_20[28]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_28 = {write1HPipe_23[28], write1HPipe_22[28]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_28 = {readData_readResultSelect_hi_lo_hi_hi_28, readData_readResultSelect_hi_lo_hi_lo_28};
  wire [7:0]         readData_readResultSelect_hi_lo_28 = {readData_readResultSelect_hi_lo_hi_28, readData_readResultSelect_hi_lo_lo_28};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_28 = {write1HPipe_25[28], write1HPipe_24[28]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_28 = {write1HPipe_27[28], write1HPipe_26[28]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_28 = {readData_readResultSelect_hi_hi_lo_hi_28, readData_readResultSelect_hi_hi_lo_lo_28};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_28 = {write1HPipe_29[28], write1HPipe_28[28]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_28 = {write1HPipe_31[28], write1HPipe_30[28]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_28 = {readData_readResultSelect_hi_hi_hi_hi_28, readData_readResultSelect_hi_hi_hi_lo_28};
  wire [7:0]         readData_readResultSelect_hi_hi_28 = {readData_readResultSelect_hi_hi_hi_28, readData_readResultSelect_hi_hi_lo_28};
  wire [15:0]        readData_readResultSelect_hi_28 = {readData_readResultSelect_hi_hi_28, readData_readResultSelect_hi_lo_28};
  wire [31:0]        readData_readResultSelect_28 = {readData_readResultSelect_hi_28, readData_readResultSelect_lo_28};
  assign readData_data_28 =
    (readData_readResultSelect_28[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_28[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_28[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_28[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_28[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_28[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_28[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_28[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_28[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_28[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_28[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_28[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_28[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_28[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_28[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_28[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_28[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_28[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_28[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_28[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_28[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_28[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_28[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_28[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_28[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_28[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_28[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_28[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_28[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_28[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_28[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_28[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_28_enq_bits = readData_data_28;
  wire               readTokenRelease_28 = readData_readDataQueue_28_deq_ready & readData_readDataQueue_28_deq_valid;
  assign readData_readDataQueue_28_enq_valid = |readData_readResultSelect_28;
  wire [31:0]        readData_data_29;
  wire               isWaiteForThisData_29;
  wire               readData_readDataQueue_29_enq_ready = ~_readData_readDataQueue_fifo_29_full;
  wire               readData_readDataQueue_29_deq_ready;
  wire               readData_readDataQueue_29_enq_valid;
  wire               readData_readDataQueue_29_deq_valid = ~_readData_readDataQueue_fifo_29_empty | readData_readDataQueue_29_enq_valid;
  wire [31:0]        readData_readDataQueue_29_enq_bits;
  wire [31:0]        readData_readDataQueue_29_deq_bits = _readData_readDataQueue_fifo_29_empty ? readData_readDataQueue_29_enq_bits : _readData_readDataQueue_fifo_29_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_29 = {write1HPipe_1[29], write1HPipe_0[29]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_29 = {write1HPipe_3[29], write1HPipe_2[29]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_29 = {readData_readResultSelect_lo_lo_lo_hi_29, readData_readResultSelect_lo_lo_lo_lo_29};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_29 = {write1HPipe_5[29], write1HPipe_4[29]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_29 = {write1HPipe_7[29], write1HPipe_6[29]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_29 = {readData_readResultSelect_lo_lo_hi_hi_29, readData_readResultSelect_lo_lo_hi_lo_29};
  wire [7:0]         readData_readResultSelect_lo_lo_29 = {readData_readResultSelect_lo_lo_hi_29, readData_readResultSelect_lo_lo_lo_29};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_29 = {write1HPipe_9[29], write1HPipe_8[29]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_29 = {write1HPipe_11[29], write1HPipe_10[29]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_29 = {readData_readResultSelect_lo_hi_lo_hi_29, readData_readResultSelect_lo_hi_lo_lo_29};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_29 = {write1HPipe_13[29], write1HPipe_12[29]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_29 = {write1HPipe_15[29], write1HPipe_14[29]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_29 = {readData_readResultSelect_lo_hi_hi_hi_29, readData_readResultSelect_lo_hi_hi_lo_29};
  wire [7:0]         readData_readResultSelect_lo_hi_29 = {readData_readResultSelect_lo_hi_hi_29, readData_readResultSelect_lo_hi_lo_29};
  wire [15:0]        readData_readResultSelect_lo_29 = {readData_readResultSelect_lo_hi_29, readData_readResultSelect_lo_lo_29};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_29 = {write1HPipe_17[29], write1HPipe_16[29]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_29 = {write1HPipe_19[29], write1HPipe_18[29]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_29 = {readData_readResultSelect_hi_lo_lo_hi_29, readData_readResultSelect_hi_lo_lo_lo_29};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_29 = {write1HPipe_21[29], write1HPipe_20[29]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_29 = {write1HPipe_23[29], write1HPipe_22[29]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_29 = {readData_readResultSelect_hi_lo_hi_hi_29, readData_readResultSelect_hi_lo_hi_lo_29};
  wire [7:0]         readData_readResultSelect_hi_lo_29 = {readData_readResultSelect_hi_lo_hi_29, readData_readResultSelect_hi_lo_lo_29};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_29 = {write1HPipe_25[29], write1HPipe_24[29]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_29 = {write1HPipe_27[29], write1HPipe_26[29]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_29 = {readData_readResultSelect_hi_hi_lo_hi_29, readData_readResultSelect_hi_hi_lo_lo_29};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_29 = {write1HPipe_29[29], write1HPipe_28[29]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_29 = {write1HPipe_31[29], write1HPipe_30[29]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_29 = {readData_readResultSelect_hi_hi_hi_hi_29, readData_readResultSelect_hi_hi_hi_lo_29};
  wire [7:0]         readData_readResultSelect_hi_hi_29 = {readData_readResultSelect_hi_hi_hi_29, readData_readResultSelect_hi_hi_lo_29};
  wire [15:0]        readData_readResultSelect_hi_29 = {readData_readResultSelect_hi_hi_29, readData_readResultSelect_hi_lo_29};
  wire [31:0]        readData_readResultSelect_29 = {readData_readResultSelect_hi_29, readData_readResultSelect_lo_29};
  assign readData_data_29 =
    (readData_readResultSelect_29[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_29[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_29[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_29[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_29[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_29[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_29[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_29[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_29[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_29[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_29[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_29[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_29[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_29[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_29[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_29[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_29[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_29[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_29[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_29[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_29[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_29[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_29[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_29[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_29[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_29[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_29[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_29[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_29[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_29[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_29[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_29[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_29_enq_bits = readData_data_29;
  wire               readTokenRelease_29 = readData_readDataQueue_29_deq_ready & readData_readDataQueue_29_deq_valid;
  assign readData_readDataQueue_29_enq_valid = |readData_readResultSelect_29;
  wire [31:0]        readData_data_30;
  wire               isWaiteForThisData_30;
  wire               readData_readDataQueue_30_enq_ready = ~_readData_readDataQueue_fifo_30_full;
  wire               readData_readDataQueue_30_deq_ready;
  wire               readData_readDataQueue_30_enq_valid;
  wire               readData_readDataQueue_30_deq_valid = ~_readData_readDataQueue_fifo_30_empty | readData_readDataQueue_30_enq_valid;
  wire [31:0]        readData_readDataQueue_30_enq_bits;
  wire [31:0]        readData_readDataQueue_30_deq_bits = _readData_readDataQueue_fifo_30_empty ? readData_readDataQueue_30_enq_bits : _readData_readDataQueue_fifo_30_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_30 = {write1HPipe_1[30], write1HPipe_0[30]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_30 = {write1HPipe_3[30], write1HPipe_2[30]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_30 = {readData_readResultSelect_lo_lo_lo_hi_30, readData_readResultSelect_lo_lo_lo_lo_30};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_30 = {write1HPipe_5[30], write1HPipe_4[30]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_30 = {write1HPipe_7[30], write1HPipe_6[30]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_30 = {readData_readResultSelect_lo_lo_hi_hi_30, readData_readResultSelect_lo_lo_hi_lo_30};
  wire [7:0]         readData_readResultSelect_lo_lo_30 = {readData_readResultSelect_lo_lo_hi_30, readData_readResultSelect_lo_lo_lo_30};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_30 = {write1HPipe_9[30], write1HPipe_8[30]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_30 = {write1HPipe_11[30], write1HPipe_10[30]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_30 = {readData_readResultSelect_lo_hi_lo_hi_30, readData_readResultSelect_lo_hi_lo_lo_30};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_30 = {write1HPipe_13[30], write1HPipe_12[30]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_30 = {write1HPipe_15[30], write1HPipe_14[30]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_30 = {readData_readResultSelect_lo_hi_hi_hi_30, readData_readResultSelect_lo_hi_hi_lo_30};
  wire [7:0]         readData_readResultSelect_lo_hi_30 = {readData_readResultSelect_lo_hi_hi_30, readData_readResultSelect_lo_hi_lo_30};
  wire [15:0]        readData_readResultSelect_lo_30 = {readData_readResultSelect_lo_hi_30, readData_readResultSelect_lo_lo_30};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_30 = {write1HPipe_17[30], write1HPipe_16[30]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_30 = {write1HPipe_19[30], write1HPipe_18[30]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_30 = {readData_readResultSelect_hi_lo_lo_hi_30, readData_readResultSelect_hi_lo_lo_lo_30};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_30 = {write1HPipe_21[30], write1HPipe_20[30]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_30 = {write1HPipe_23[30], write1HPipe_22[30]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_30 = {readData_readResultSelect_hi_lo_hi_hi_30, readData_readResultSelect_hi_lo_hi_lo_30};
  wire [7:0]         readData_readResultSelect_hi_lo_30 = {readData_readResultSelect_hi_lo_hi_30, readData_readResultSelect_hi_lo_lo_30};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_30 = {write1HPipe_25[30], write1HPipe_24[30]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_30 = {write1HPipe_27[30], write1HPipe_26[30]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_30 = {readData_readResultSelect_hi_hi_lo_hi_30, readData_readResultSelect_hi_hi_lo_lo_30};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_30 = {write1HPipe_29[30], write1HPipe_28[30]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_30 = {write1HPipe_31[30], write1HPipe_30[30]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_30 = {readData_readResultSelect_hi_hi_hi_hi_30, readData_readResultSelect_hi_hi_hi_lo_30};
  wire [7:0]         readData_readResultSelect_hi_hi_30 = {readData_readResultSelect_hi_hi_hi_30, readData_readResultSelect_hi_hi_lo_30};
  wire [15:0]        readData_readResultSelect_hi_30 = {readData_readResultSelect_hi_hi_30, readData_readResultSelect_hi_lo_30};
  wire [31:0]        readData_readResultSelect_30 = {readData_readResultSelect_hi_30, readData_readResultSelect_lo_30};
  assign readData_data_30 =
    (readData_readResultSelect_30[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_30[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_30[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_30[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_30[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_30[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_30[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_30[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_30[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_30[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_30[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_30[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_30[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_30[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_30[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_30[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_30[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_30[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_30[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_30[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_30[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_30[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_30[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_30[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_30[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_30[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_30[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_30[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_30[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_30[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_30[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_30[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_30_enq_bits = readData_data_30;
  wire               readTokenRelease_30 = readData_readDataQueue_30_deq_ready & readData_readDataQueue_30_deq_valid;
  assign readData_readDataQueue_30_enq_valid = |readData_readResultSelect_30;
  wire [31:0]        readData_data_31;
  wire               isWaiteForThisData_31;
  wire               readData_readDataQueue_31_enq_ready = ~_readData_readDataQueue_fifo_31_full;
  wire               readData_readDataQueue_31_deq_ready;
  wire               readData_readDataQueue_31_enq_valid;
  wire               readData_readDataQueue_31_deq_valid = ~_readData_readDataQueue_fifo_31_empty | readData_readDataQueue_31_enq_valid;
  wire [31:0]        readData_readDataQueue_31_enq_bits;
  wire [31:0]        readData_readDataQueue_31_deq_bits = _readData_readDataQueue_fifo_31_empty ? readData_readDataQueue_31_enq_bits : _readData_readDataQueue_fifo_31_data_out;
  wire [1:0]         readData_readResultSelect_lo_lo_lo_lo_31 = {write1HPipe_1[31], write1HPipe_0[31]};
  wire [1:0]         readData_readResultSelect_lo_lo_lo_hi_31 = {write1HPipe_3[31], write1HPipe_2[31]};
  wire [3:0]         readData_readResultSelect_lo_lo_lo_31 = {readData_readResultSelect_lo_lo_lo_hi_31, readData_readResultSelect_lo_lo_lo_lo_31};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_lo_31 = {write1HPipe_5[31], write1HPipe_4[31]};
  wire [1:0]         readData_readResultSelect_lo_lo_hi_hi_31 = {write1HPipe_7[31], write1HPipe_6[31]};
  wire [3:0]         readData_readResultSelect_lo_lo_hi_31 = {readData_readResultSelect_lo_lo_hi_hi_31, readData_readResultSelect_lo_lo_hi_lo_31};
  wire [7:0]         readData_readResultSelect_lo_lo_31 = {readData_readResultSelect_lo_lo_hi_31, readData_readResultSelect_lo_lo_lo_31};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_lo_31 = {write1HPipe_9[31], write1HPipe_8[31]};
  wire [1:0]         readData_readResultSelect_lo_hi_lo_hi_31 = {write1HPipe_11[31], write1HPipe_10[31]};
  wire [3:0]         readData_readResultSelect_lo_hi_lo_31 = {readData_readResultSelect_lo_hi_lo_hi_31, readData_readResultSelect_lo_hi_lo_lo_31};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_lo_31 = {write1HPipe_13[31], write1HPipe_12[31]};
  wire [1:0]         readData_readResultSelect_lo_hi_hi_hi_31 = {write1HPipe_15[31], write1HPipe_14[31]};
  wire [3:0]         readData_readResultSelect_lo_hi_hi_31 = {readData_readResultSelect_lo_hi_hi_hi_31, readData_readResultSelect_lo_hi_hi_lo_31};
  wire [7:0]         readData_readResultSelect_lo_hi_31 = {readData_readResultSelect_lo_hi_hi_31, readData_readResultSelect_lo_hi_lo_31};
  wire [15:0]        readData_readResultSelect_lo_31 = {readData_readResultSelect_lo_hi_31, readData_readResultSelect_lo_lo_31};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_lo_31 = {write1HPipe_17[31], write1HPipe_16[31]};
  wire [1:0]         readData_readResultSelect_hi_lo_lo_hi_31 = {write1HPipe_19[31], write1HPipe_18[31]};
  wire [3:0]         readData_readResultSelect_hi_lo_lo_31 = {readData_readResultSelect_hi_lo_lo_hi_31, readData_readResultSelect_hi_lo_lo_lo_31};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_lo_31 = {write1HPipe_21[31], write1HPipe_20[31]};
  wire [1:0]         readData_readResultSelect_hi_lo_hi_hi_31 = {write1HPipe_23[31], write1HPipe_22[31]};
  wire [3:0]         readData_readResultSelect_hi_lo_hi_31 = {readData_readResultSelect_hi_lo_hi_hi_31, readData_readResultSelect_hi_lo_hi_lo_31};
  wire [7:0]         readData_readResultSelect_hi_lo_31 = {readData_readResultSelect_hi_lo_hi_31, readData_readResultSelect_hi_lo_lo_31};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_lo_31 = {write1HPipe_25[31], write1HPipe_24[31]};
  wire [1:0]         readData_readResultSelect_hi_hi_lo_hi_31 = {write1HPipe_27[31], write1HPipe_26[31]};
  wire [3:0]         readData_readResultSelect_hi_hi_lo_31 = {readData_readResultSelect_hi_hi_lo_hi_31, readData_readResultSelect_hi_hi_lo_lo_31};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_lo_31 = {write1HPipe_29[31], write1HPipe_28[31]};
  wire [1:0]         readData_readResultSelect_hi_hi_hi_hi_31 = {write1HPipe_31[31], write1HPipe_30[31]};
  wire [3:0]         readData_readResultSelect_hi_hi_hi_31 = {readData_readResultSelect_hi_hi_hi_hi_31, readData_readResultSelect_hi_hi_hi_lo_31};
  wire [7:0]         readData_readResultSelect_hi_hi_31 = {readData_readResultSelect_hi_hi_hi_31, readData_readResultSelect_hi_hi_lo_31};
  wire [15:0]        readData_readResultSelect_hi_31 = {readData_readResultSelect_hi_hi_31, readData_readResultSelect_hi_lo_31};
  wire [31:0]        readData_readResultSelect_31 = {readData_readResultSelect_hi_31, readData_readResultSelect_lo_31};
  assign readData_data_31 =
    (readData_readResultSelect_31[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_31[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_31[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_31[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_31[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_31[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_31[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_31[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_31[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_31[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_31[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_31[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_31[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_31[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_31[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_31[15] ? dataAfterReorderCheck_15 : 32'h0) | (readData_readResultSelect_31[16] ? dataAfterReorderCheck_16 : 32'h0) | (readData_readResultSelect_31[17] ? dataAfterReorderCheck_17 : 32'h0)
    | (readData_readResultSelect_31[18] ? dataAfterReorderCheck_18 : 32'h0) | (readData_readResultSelect_31[19] ? dataAfterReorderCheck_19 : 32'h0) | (readData_readResultSelect_31[20] ? dataAfterReorderCheck_20 : 32'h0)
    | (readData_readResultSelect_31[21] ? dataAfterReorderCheck_21 : 32'h0) | (readData_readResultSelect_31[22] ? dataAfterReorderCheck_22 : 32'h0) | (readData_readResultSelect_31[23] ? dataAfterReorderCheck_23 : 32'h0)
    | (readData_readResultSelect_31[24] ? dataAfterReorderCheck_24 : 32'h0) | (readData_readResultSelect_31[25] ? dataAfterReorderCheck_25 : 32'h0) | (readData_readResultSelect_31[26] ? dataAfterReorderCheck_26 : 32'h0)
    | (readData_readResultSelect_31[27] ? dataAfterReorderCheck_27 : 32'h0) | (readData_readResultSelect_31[28] ? dataAfterReorderCheck_28 : 32'h0) | (readData_readResultSelect_31[29] ? dataAfterReorderCheck_29 : 32'h0)
    | (readData_readResultSelect_31[30] ? dataAfterReorderCheck_30 : 32'h0) | (readData_readResultSelect_31[31] ? dataAfterReorderCheck_31 : 32'h0);
  assign readData_readDataQueue_31_enq_bits = readData_data_31;
  wire               readTokenRelease_31 = readData_readDataQueue_31_deq_ready & readData_readDataQueue_31_deq_valid;
  assign readData_readDataQueue_31_enq_valid = |readData_readResultSelect_31;
  reg  [6:0]         waiteReadDataPipeReg_executeGroup;
  reg  [31:0]        waiteReadDataPipeReg_sourceValid;
  reg  [31:0]        waiteReadDataPipeReg_replaceVs1;
  reg  [31:0]        waiteReadDataPipeReg_needRead;
  reg                waiteReadDataPipeReg_last;
  reg  [31:0]        waiteReadData_0;
  reg  [31:0]        waiteReadData_1;
  reg  [31:0]        waiteReadData_2;
  reg  [31:0]        waiteReadData_3;
  reg  [31:0]        waiteReadData_4;
  reg  [31:0]        waiteReadData_5;
  reg  [31:0]        waiteReadData_6;
  reg  [31:0]        waiteReadData_7;
  reg  [31:0]        waiteReadData_8;
  reg  [31:0]        waiteReadData_9;
  reg  [31:0]        waiteReadData_10;
  reg  [31:0]        waiteReadData_11;
  reg  [31:0]        waiteReadData_12;
  reg  [31:0]        waiteReadData_13;
  reg  [31:0]        waiteReadData_14;
  reg  [31:0]        waiteReadData_15;
  reg  [31:0]        waiteReadData_16;
  reg  [31:0]        waiteReadData_17;
  reg  [31:0]        waiteReadData_18;
  reg  [31:0]        waiteReadData_19;
  reg  [31:0]        waiteReadData_20;
  reg  [31:0]        waiteReadData_21;
  reg  [31:0]        waiteReadData_22;
  reg  [31:0]        waiteReadData_23;
  reg  [31:0]        waiteReadData_24;
  reg  [31:0]        waiteReadData_25;
  reg  [31:0]        waiteReadData_26;
  reg  [31:0]        waiteReadData_27;
  reg  [31:0]        waiteReadData_28;
  reg  [31:0]        waiteReadData_29;
  reg  [31:0]        waiteReadData_30;
  reg  [31:0]        waiteReadData_31;
  reg  [31:0]        waiteReadSate;
  reg                waiteReadStageValid;
  wire [1:0]         executeIndexVec_0 = waiteReadDataPipeReg_executeGroup[1:0];
  wire [1:0]         executeIndexVec_1 = {waiteReadDataPipeReg_executeGroup[0], 1'h0};
  wire               writeDataVec_data_dataIsRead = waiteReadDataPipeReg_needRead[0];
  wire               writeDataVec_data_dataIsRead_32 = waiteReadDataPipeReg_needRead[0];
  wire               writeDataVec_data_dataIsRead_64 = waiteReadDataPipeReg_needRead[0];
  wire [31:0]        _GEN_141 = waiteReadDataPipeReg_replaceVs1[0] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData;
  assign writeDataVec_data_unreadData = _GEN_141;
  wire [31:0]        writeDataVec_data_unreadData_32;
  assign writeDataVec_data_unreadData_32 = _GEN_141;
  wire [31:0]        writeDataVec_data_unreadData_64;
  assign writeDataVec_data_unreadData_64 = _GEN_141;
  wire [7:0]         writeDataVec_data_dataElement = writeDataVec_data_dataIsRead ? waiteReadData_0[7:0] : writeDataVec_data_unreadData[7:0];
  wire               writeDataVec_data_dataIsRead_1 = waiteReadDataPipeReg_needRead[1];
  wire               writeDataVec_data_dataIsRead_33 = waiteReadDataPipeReg_needRead[1];
  wire               writeDataVec_data_dataIsRead_65 = waiteReadDataPipeReg_needRead[1];
  wire [31:0]        _GEN_142 = waiteReadDataPipeReg_replaceVs1[1] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_1;
  assign writeDataVec_data_unreadData_1 = _GEN_142;
  wire [31:0]        writeDataVec_data_unreadData_33;
  assign writeDataVec_data_unreadData_33 = _GEN_142;
  wire [31:0]        writeDataVec_data_unreadData_65;
  assign writeDataVec_data_unreadData_65 = _GEN_142;
  wire [7:0]         writeDataVec_data_dataElement_1 = writeDataVec_data_dataIsRead_1 ? waiteReadData_1[7:0] : writeDataVec_data_unreadData_1[7:0];
  wire               writeDataVec_data_dataIsRead_2 = waiteReadDataPipeReg_needRead[2];
  wire               writeDataVec_data_dataIsRead_34 = waiteReadDataPipeReg_needRead[2];
  wire               writeDataVec_data_dataIsRead_66 = waiteReadDataPipeReg_needRead[2];
  wire [31:0]        _GEN_143 = waiteReadDataPipeReg_replaceVs1[2] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_2;
  assign writeDataVec_data_unreadData_2 = _GEN_143;
  wire [31:0]        writeDataVec_data_unreadData_34;
  assign writeDataVec_data_unreadData_34 = _GEN_143;
  wire [31:0]        writeDataVec_data_unreadData_66;
  assign writeDataVec_data_unreadData_66 = _GEN_143;
  wire [7:0]         writeDataVec_data_dataElement_2 = writeDataVec_data_dataIsRead_2 ? waiteReadData_2[7:0] : writeDataVec_data_unreadData_2[7:0];
  wire               writeDataVec_data_dataIsRead_3 = waiteReadDataPipeReg_needRead[3];
  wire               writeDataVec_data_dataIsRead_35 = waiteReadDataPipeReg_needRead[3];
  wire               writeDataVec_data_dataIsRead_67 = waiteReadDataPipeReg_needRead[3];
  wire [31:0]        _GEN_144 = waiteReadDataPipeReg_replaceVs1[3] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_3;
  assign writeDataVec_data_unreadData_3 = _GEN_144;
  wire [31:0]        writeDataVec_data_unreadData_35;
  assign writeDataVec_data_unreadData_35 = _GEN_144;
  wire [31:0]        writeDataVec_data_unreadData_67;
  assign writeDataVec_data_unreadData_67 = _GEN_144;
  wire [7:0]         writeDataVec_data_dataElement_3 = writeDataVec_data_dataIsRead_3 ? waiteReadData_3[7:0] : writeDataVec_data_unreadData_3[7:0];
  wire               writeDataVec_data_dataIsRead_4 = waiteReadDataPipeReg_needRead[4];
  wire               writeDataVec_data_dataIsRead_36 = waiteReadDataPipeReg_needRead[4];
  wire               writeDataVec_data_dataIsRead_68 = waiteReadDataPipeReg_needRead[4];
  wire [31:0]        _GEN_145 = waiteReadDataPipeReg_replaceVs1[4] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_4;
  assign writeDataVec_data_unreadData_4 = _GEN_145;
  wire [31:0]        writeDataVec_data_unreadData_36;
  assign writeDataVec_data_unreadData_36 = _GEN_145;
  wire [31:0]        writeDataVec_data_unreadData_68;
  assign writeDataVec_data_unreadData_68 = _GEN_145;
  wire [7:0]         writeDataVec_data_dataElement_4 = writeDataVec_data_dataIsRead_4 ? waiteReadData_4[7:0] : writeDataVec_data_unreadData_4[7:0];
  wire               writeDataVec_data_dataIsRead_5 = waiteReadDataPipeReg_needRead[5];
  wire               writeDataVec_data_dataIsRead_37 = waiteReadDataPipeReg_needRead[5];
  wire               writeDataVec_data_dataIsRead_69 = waiteReadDataPipeReg_needRead[5];
  wire [31:0]        _GEN_146 = waiteReadDataPipeReg_replaceVs1[5] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_5;
  assign writeDataVec_data_unreadData_5 = _GEN_146;
  wire [31:0]        writeDataVec_data_unreadData_37;
  assign writeDataVec_data_unreadData_37 = _GEN_146;
  wire [31:0]        writeDataVec_data_unreadData_69;
  assign writeDataVec_data_unreadData_69 = _GEN_146;
  wire [7:0]         writeDataVec_data_dataElement_5 = writeDataVec_data_dataIsRead_5 ? waiteReadData_5[7:0] : writeDataVec_data_unreadData_5[7:0];
  wire               writeDataVec_data_dataIsRead_6 = waiteReadDataPipeReg_needRead[6];
  wire               writeDataVec_data_dataIsRead_38 = waiteReadDataPipeReg_needRead[6];
  wire               writeDataVec_data_dataIsRead_70 = waiteReadDataPipeReg_needRead[6];
  wire [31:0]        _GEN_147 = waiteReadDataPipeReg_replaceVs1[6] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_6;
  assign writeDataVec_data_unreadData_6 = _GEN_147;
  wire [31:0]        writeDataVec_data_unreadData_38;
  assign writeDataVec_data_unreadData_38 = _GEN_147;
  wire [31:0]        writeDataVec_data_unreadData_70;
  assign writeDataVec_data_unreadData_70 = _GEN_147;
  wire [7:0]         writeDataVec_data_dataElement_6 = writeDataVec_data_dataIsRead_6 ? waiteReadData_6[7:0] : writeDataVec_data_unreadData_6[7:0];
  wire               writeDataVec_data_dataIsRead_7 = waiteReadDataPipeReg_needRead[7];
  wire               writeDataVec_data_dataIsRead_39 = waiteReadDataPipeReg_needRead[7];
  wire               writeDataVec_data_dataIsRead_71 = waiteReadDataPipeReg_needRead[7];
  wire [31:0]        _GEN_148 = waiteReadDataPipeReg_replaceVs1[7] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_7;
  assign writeDataVec_data_unreadData_7 = _GEN_148;
  wire [31:0]        writeDataVec_data_unreadData_39;
  assign writeDataVec_data_unreadData_39 = _GEN_148;
  wire [31:0]        writeDataVec_data_unreadData_71;
  assign writeDataVec_data_unreadData_71 = _GEN_148;
  wire [7:0]         writeDataVec_data_dataElement_7 = writeDataVec_data_dataIsRead_7 ? waiteReadData_7[7:0] : writeDataVec_data_unreadData_7[7:0];
  wire               writeDataVec_data_dataIsRead_8 = waiteReadDataPipeReg_needRead[8];
  wire               writeDataVec_data_dataIsRead_40 = waiteReadDataPipeReg_needRead[8];
  wire               writeDataVec_data_dataIsRead_72 = waiteReadDataPipeReg_needRead[8];
  wire [31:0]        _GEN_149 = waiteReadDataPipeReg_replaceVs1[8] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_8;
  assign writeDataVec_data_unreadData_8 = _GEN_149;
  wire [31:0]        writeDataVec_data_unreadData_40;
  assign writeDataVec_data_unreadData_40 = _GEN_149;
  wire [31:0]        writeDataVec_data_unreadData_72;
  assign writeDataVec_data_unreadData_72 = _GEN_149;
  wire [7:0]         writeDataVec_data_dataElement_8 = writeDataVec_data_dataIsRead_8 ? waiteReadData_8[7:0] : writeDataVec_data_unreadData_8[7:0];
  wire               writeDataVec_data_dataIsRead_9 = waiteReadDataPipeReg_needRead[9];
  wire               writeDataVec_data_dataIsRead_41 = waiteReadDataPipeReg_needRead[9];
  wire               writeDataVec_data_dataIsRead_73 = waiteReadDataPipeReg_needRead[9];
  wire [31:0]        _GEN_150 = waiteReadDataPipeReg_replaceVs1[9] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_9;
  assign writeDataVec_data_unreadData_9 = _GEN_150;
  wire [31:0]        writeDataVec_data_unreadData_41;
  assign writeDataVec_data_unreadData_41 = _GEN_150;
  wire [31:0]        writeDataVec_data_unreadData_73;
  assign writeDataVec_data_unreadData_73 = _GEN_150;
  wire [7:0]         writeDataVec_data_dataElement_9 = writeDataVec_data_dataIsRead_9 ? waiteReadData_9[7:0] : writeDataVec_data_unreadData_9[7:0];
  wire               writeDataVec_data_dataIsRead_10 = waiteReadDataPipeReg_needRead[10];
  wire               writeDataVec_data_dataIsRead_42 = waiteReadDataPipeReg_needRead[10];
  wire               writeDataVec_data_dataIsRead_74 = waiteReadDataPipeReg_needRead[10];
  wire [31:0]        _GEN_151 = waiteReadDataPipeReg_replaceVs1[10] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_10;
  assign writeDataVec_data_unreadData_10 = _GEN_151;
  wire [31:0]        writeDataVec_data_unreadData_42;
  assign writeDataVec_data_unreadData_42 = _GEN_151;
  wire [31:0]        writeDataVec_data_unreadData_74;
  assign writeDataVec_data_unreadData_74 = _GEN_151;
  wire [7:0]         writeDataVec_data_dataElement_10 = writeDataVec_data_dataIsRead_10 ? waiteReadData_10[7:0] : writeDataVec_data_unreadData_10[7:0];
  wire               writeDataVec_data_dataIsRead_11 = waiteReadDataPipeReg_needRead[11];
  wire               writeDataVec_data_dataIsRead_43 = waiteReadDataPipeReg_needRead[11];
  wire               writeDataVec_data_dataIsRead_75 = waiteReadDataPipeReg_needRead[11];
  wire [31:0]        _GEN_152 = waiteReadDataPipeReg_replaceVs1[11] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_11;
  assign writeDataVec_data_unreadData_11 = _GEN_152;
  wire [31:0]        writeDataVec_data_unreadData_43;
  assign writeDataVec_data_unreadData_43 = _GEN_152;
  wire [31:0]        writeDataVec_data_unreadData_75;
  assign writeDataVec_data_unreadData_75 = _GEN_152;
  wire [7:0]         writeDataVec_data_dataElement_11 = writeDataVec_data_dataIsRead_11 ? waiteReadData_11[7:0] : writeDataVec_data_unreadData_11[7:0];
  wire               writeDataVec_data_dataIsRead_12 = waiteReadDataPipeReg_needRead[12];
  wire               writeDataVec_data_dataIsRead_44 = waiteReadDataPipeReg_needRead[12];
  wire               writeDataVec_data_dataIsRead_76 = waiteReadDataPipeReg_needRead[12];
  wire [31:0]        _GEN_153 = waiteReadDataPipeReg_replaceVs1[12] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_12;
  assign writeDataVec_data_unreadData_12 = _GEN_153;
  wire [31:0]        writeDataVec_data_unreadData_44;
  assign writeDataVec_data_unreadData_44 = _GEN_153;
  wire [31:0]        writeDataVec_data_unreadData_76;
  assign writeDataVec_data_unreadData_76 = _GEN_153;
  wire [7:0]         writeDataVec_data_dataElement_12 = writeDataVec_data_dataIsRead_12 ? waiteReadData_12[7:0] : writeDataVec_data_unreadData_12[7:0];
  wire               writeDataVec_data_dataIsRead_13 = waiteReadDataPipeReg_needRead[13];
  wire               writeDataVec_data_dataIsRead_45 = waiteReadDataPipeReg_needRead[13];
  wire               writeDataVec_data_dataIsRead_77 = waiteReadDataPipeReg_needRead[13];
  wire [31:0]        _GEN_154 = waiteReadDataPipeReg_replaceVs1[13] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_13;
  assign writeDataVec_data_unreadData_13 = _GEN_154;
  wire [31:0]        writeDataVec_data_unreadData_45;
  assign writeDataVec_data_unreadData_45 = _GEN_154;
  wire [31:0]        writeDataVec_data_unreadData_77;
  assign writeDataVec_data_unreadData_77 = _GEN_154;
  wire [7:0]         writeDataVec_data_dataElement_13 = writeDataVec_data_dataIsRead_13 ? waiteReadData_13[7:0] : writeDataVec_data_unreadData_13[7:0];
  wire               writeDataVec_data_dataIsRead_14 = waiteReadDataPipeReg_needRead[14];
  wire               writeDataVec_data_dataIsRead_46 = waiteReadDataPipeReg_needRead[14];
  wire               writeDataVec_data_dataIsRead_78 = waiteReadDataPipeReg_needRead[14];
  wire [31:0]        _GEN_155 = waiteReadDataPipeReg_replaceVs1[14] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_14;
  assign writeDataVec_data_unreadData_14 = _GEN_155;
  wire [31:0]        writeDataVec_data_unreadData_46;
  assign writeDataVec_data_unreadData_46 = _GEN_155;
  wire [31:0]        writeDataVec_data_unreadData_78;
  assign writeDataVec_data_unreadData_78 = _GEN_155;
  wire [7:0]         writeDataVec_data_dataElement_14 = writeDataVec_data_dataIsRead_14 ? waiteReadData_14[7:0] : writeDataVec_data_unreadData_14[7:0];
  wire               writeDataVec_data_dataIsRead_15 = waiteReadDataPipeReg_needRead[15];
  wire               writeDataVec_data_dataIsRead_47 = waiteReadDataPipeReg_needRead[15];
  wire               writeDataVec_data_dataIsRead_79 = waiteReadDataPipeReg_needRead[15];
  wire [31:0]        _GEN_156 = waiteReadDataPipeReg_replaceVs1[15] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_15;
  assign writeDataVec_data_unreadData_15 = _GEN_156;
  wire [31:0]        writeDataVec_data_unreadData_47;
  assign writeDataVec_data_unreadData_47 = _GEN_156;
  wire [31:0]        writeDataVec_data_unreadData_79;
  assign writeDataVec_data_unreadData_79 = _GEN_156;
  wire [7:0]         writeDataVec_data_dataElement_15 = writeDataVec_data_dataIsRead_15 ? waiteReadData_15[7:0] : writeDataVec_data_unreadData_15[7:0];
  wire               writeDataVec_data_dataIsRead_16 = waiteReadDataPipeReg_needRead[16];
  wire               writeDataVec_data_dataIsRead_48 = waiteReadDataPipeReg_needRead[16];
  wire               writeDataVec_data_dataIsRead_80 = waiteReadDataPipeReg_needRead[16];
  wire [31:0]        _GEN_157 = waiteReadDataPipeReg_replaceVs1[16] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_16;
  assign writeDataVec_data_unreadData_16 = _GEN_157;
  wire [31:0]        writeDataVec_data_unreadData_48;
  assign writeDataVec_data_unreadData_48 = _GEN_157;
  wire [31:0]        writeDataVec_data_unreadData_80;
  assign writeDataVec_data_unreadData_80 = _GEN_157;
  wire [7:0]         writeDataVec_data_dataElement_16 = writeDataVec_data_dataIsRead_16 ? waiteReadData_16[7:0] : writeDataVec_data_unreadData_16[7:0];
  wire               writeDataVec_data_dataIsRead_17 = waiteReadDataPipeReg_needRead[17];
  wire               writeDataVec_data_dataIsRead_49 = waiteReadDataPipeReg_needRead[17];
  wire               writeDataVec_data_dataIsRead_81 = waiteReadDataPipeReg_needRead[17];
  wire [31:0]        _GEN_158 = waiteReadDataPipeReg_replaceVs1[17] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_17;
  assign writeDataVec_data_unreadData_17 = _GEN_158;
  wire [31:0]        writeDataVec_data_unreadData_49;
  assign writeDataVec_data_unreadData_49 = _GEN_158;
  wire [31:0]        writeDataVec_data_unreadData_81;
  assign writeDataVec_data_unreadData_81 = _GEN_158;
  wire [7:0]         writeDataVec_data_dataElement_17 = writeDataVec_data_dataIsRead_17 ? waiteReadData_17[7:0] : writeDataVec_data_unreadData_17[7:0];
  wire               writeDataVec_data_dataIsRead_18 = waiteReadDataPipeReg_needRead[18];
  wire               writeDataVec_data_dataIsRead_50 = waiteReadDataPipeReg_needRead[18];
  wire               writeDataVec_data_dataIsRead_82 = waiteReadDataPipeReg_needRead[18];
  wire [31:0]        _GEN_159 = waiteReadDataPipeReg_replaceVs1[18] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_18;
  assign writeDataVec_data_unreadData_18 = _GEN_159;
  wire [31:0]        writeDataVec_data_unreadData_50;
  assign writeDataVec_data_unreadData_50 = _GEN_159;
  wire [31:0]        writeDataVec_data_unreadData_82;
  assign writeDataVec_data_unreadData_82 = _GEN_159;
  wire [7:0]         writeDataVec_data_dataElement_18 = writeDataVec_data_dataIsRead_18 ? waiteReadData_18[7:0] : writeDataVec_data_unreadData_18[7:0];
  wire               writeDataVec_data_dataIsRead_19 = waiteReadDataPipeReg_needRead[19];
  wire               writeDataVec_data_dataIsRead_51 = waiteReadDataPipeReg_needRead[19];
  wire               writeDataVec_data_dataIsRead_83 = waiteReadDataPipeReg_needRead[19];
  wire [31:0]        _GEN_160 = waiteReadDataPipeReg_replaceVs1[19] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_19;
  assign writeDataVec_data_unreadData_19 = _GEN_160;
  wire [31:0]        writeDataVec_data_unreadData_51;
  assign writeDataVec_data_unreadData_51 = _GEN_160;
  wire [31:0]        writeDataVec_data_unreadData_83;
  assign writeDataVec_data_unreadData_83 = _GEN_160;
  wire [7:0]         writeDataVec_data_dataElement_19 = writeDataVec_data_dataIsRead_19 ? waiteReadData_19[7:0] : writeDataVec_data_unreadData_19[7:0];
  wire               writeDataVec_data_dataIsRead_20 = waiteReadDataPipeReg_needRead[20];
  wire               writeDataVec_data_dataIsRead_52 = waiteReadDataPipeReg_needRead[20];
  wire               writeDataVec_data_dataIsRead_84 = waiteReadDataPipeReg_needRead[20];
  wire [31:0]        _GEN_161 = waiteReadDataPipeReg_replaceVs1[20] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_20;
  assign writeDataVec_data_unreadData_20 = _GEN_161;
  wire [31:0]        writeDataVec_data_unreadData_52;
  assign writeDataVec_data_unreadData_52 = _GEN_161;
  wire [31:0]        writeDataVec_data_unreadData_84;
  assign writeDataVec_data_unreadData_84 = _GEN_161;
  wire [7:0]         writeDataVec_data_dataElement_20 = writeDataVec_data_dataIsRead_20 ? waiteReadData_20[7:0] : writeDataVec_data_unreadData_20[7:0];
  wire               writeDataVec_data_dataIsRead_21 = waiteReadDataPipeReg_needRead[21];
  wire               writeDataVec_data_dataIsRead_53 = waiteReadDataPipeReg_needRead[21];
  wire               writeDataVec_data_dataIsRead_85 = waiteReadDataPipeReg_needRead[21];
  wire [31:0]        _GEN_162 = waiteReadDataPipeReg_replaceVs1[21] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_21;
  assign writeDataVec_data_unreadData_21 = _GEN_162;
  wire [31:0]        writeDataVec_data_unreadData_53;
  assign writeDataVec_data_unreadData_53 = _GEN_162;
  wire [31:0]        writeDataVec_data_unreadData_85;
  assign writeDataVec_data_unreadData_85 = _GEN_162;
  wire [7:0]         writeDataVec_data_dataElement_21 = writeDataVec_data_dataIsRead_21 ? waiteReadData_21[7:0] : writeDataVec_data_unreadData_21[7:0];
  wire               writeDataVec_data_dataIsRead_22 = waiteReadDataPipeReg_needRead[22];
  wire               writeDataVec_data_dataIsRead_54 = waiteReadDataPipeReg_needRead[22];
  wire               writeDataVec_data_dataIsRead_86 = waiteReadDataPipeReg_needRead[22];
  wire [31:0]        _GEN_163 = waiteReadDataPipeReg_replaceVs1[22] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_22;
  assign writeDataVec_data_unreadData_22 = _GEN_163;
  wire [31:0]        writeDataVec_data_unreadData_54;
  assign writeDataVec_data_unreadData_54 = _GEN_163;
  wire [31:0]        writeDataVec_data_unreadData_86;
  assign writeDataVec_data_unreadData_86 = _GEN_163;
  wire [7:0]         writeDataVec_data_dataElement_22 = writeDataVec_data_dataIsRead_22 ? waiteReadData_22[7:0] : writeDataVec_data_unreadData_22[7:0];
  wire               writeDataVec_data_dataIsRead_23 = waiteReadDataPipeReg_needRead[23];
  wire               writeDataVec_data_dataIsRead_55 = waiteReadDataPipeReg_needRead[23];
  wire               writeDataVec_data_dataIsRead_87 = waiteReadDataPipeReg_needRead[23];
  wire [31:0]        _GEN_164 = waiteReadDataPipeReg_replaceVs1[23] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_23;
  assign writeDataVec_data_unreadData_23 = _GEN_164;
  wire [31:0]        writeDataVec_data_unreadData_55;
  assign writeDataVec_data_unreadData_55 = _GEN_164;
  wire [31:0]        writeDataVec_data_unreadData_87;
  assign writeDataVec_data_unreadData_87 = _GEN_164;
  wire [7:0]         writeDataVec_data_dataElement_23 = writeDataVec_data_dataIsRead_23 ? waiteReadData_23[7:0] : writeDataVec_data_unreadData_23[7:0];
  wire               writeDataVec_data_dataIsRead_24 = waiteReadDataPipeReg_needRead[24];
  wire               writeDataVec_data_dataIsRead_56 = waiteReadDataPipeReg_needRead[24];
  wire               writeDataVec_data_dataIsRead_88 = waiteReadDataPipeReg_needRead[24];
  wire [31:0]        _GEN_165 = waiteReadDataPipeReg_replaceVs1[24] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_24;
  assign writeDataVec_data_unreadData_24 = _GEN_165;
  wire [31:0]        writeDataVec_data_unreadData_56;
  assign writeDataVec_data_unreadData_56 = _GEN_165;
  wire [31:0]        writeDataVec_data_unreadData_88;
  assign writeDataVec_data_unreadData_88 = _GEN_165;
  wire [7:0]         writeDataVec_data_dataElement_24 = writeDataVec_data_dataIsRead_24 ? waiteReadData_24[7:0] : writeDataVec_data_unreadData_24[7:0];
  wire               writeDataVec_data_dataIsRead_25 = waiteReadDataPipeReg_needRead[25];
  wire               writeDataVec_data_dataIsRead_57 = waiteReadDataPipeReg_needRead[25];
  wire               writeDataVec_data_dataIsRead_89 = waiteReadDataPipeReg_needRead[25];
  wire [31:0]        _GEN_166 = waiteReadDataPipeReg_replaceVs1[25] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_25;
  assign writeDataVec_data_unreadData_25 = _GEN_166;
  wire [31:0]        writeDataVec_data_unreadData_57;
  assign writeDataVec_data_unreadData_57 = _GEN_166;
  wire [31:0]        writeDataVec_data_unreadData_89;
  assign writeDataVec_data_unreadData_89 = _GEN_166;
  wire [7:0]         writeDataVec_data_dataElement_25 = writeDataVec_data_dataIsRead_25 ? waiteReadData_25[7:0] : writeDataVec_data_unreadData_25[7:0];
  wire               writeDataVec_data_dataIsRead_26 = waiteReadDataPipeReg_needRead[26];
  wire               writeDataVec_data_dataIsRead_58 = waiteReadDataPipeReg_needRead[26];
  wire               writeDataVec_data_dataIsRead_90 = waiteReadDataPipeReg_needRead[26];
  wire [31:0]        _GEN_167 = waiteReadDataPipeReg_replaceVs1[26] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_26;
  assign writeDataVec_data_unreadData_26 = _GEN_167;
  wire [31:0]        writeDataVec_data_unreadData_58;
  assign writeDataVec_data_unreadData_58 = _GEN_167;
  wire [31:0]        writeDataVec_data_unreadData_90;
  assign writeDataVec_data_unreadData_90 = _GEN_167;
  wire [7:0]         writeDataVec_data_dataElement_26 = writeDataVec_data_dataIsRead_26 ? waiteReadData_26[7:0] : writeDataVec_data_unreadData_26[7:0];
  wire               writeDataVec_data_dataIsRead_27 = waiteReadDataPipeReg_needRead[27];
  wire               writeDataVec_data_dataIsRead_59 = waiteReadDataPipeReg_needRead[27];
  wire               writeDataVec_data_dataIsRead_91 = waiteReadDataPipeReg_needRead[27];
  wire [31:0]        _GEN_168 = waiteReadDataPipeReg_replaceVs1[27] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_27;
  assign writeDataVec_data_unreadData_27 = _GEN_168;
  wire [31:0]        writeDataVec_data_unreadData_59;
  assign writeDataVec_data_unreadData_59 = _GEN_168;
  wire [31:0]        writeDataVec_data_unreadData_91;
  assign writeDataVec_data_unreadData_91 = _GEN_168;
  wire [7:0]         writeDataVec_data_dataElement_27 = writeDataVec_data_dataIsRead_27 ? waiteReadData_27[7:0] : writeDataVec_data_unreadData_27[7:0];
  wire               writeDataVec_data_dataIsRead_28 = waiteReadDataPipeReg_needRead[28];
  wire               writeDataVec_data_dataIsRead_60 = waiteReadDataPipeReg_needRead[28];
  wire               writeDataVec_data_dataIsRead_92 = waiteReadDataPipeReg_needRead[28];
  wire [31:0]        _GEN_169 = waiteReadDataPipeReg_replaceVs1[28] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_28;
  assign writeDataVec_data_unreadData_28 = _GEN_169;
  wire [31:0]        writeDataVec_data_unreadData_60;
  assign writeDataVec_data_unreadData_60 = _GEN_169;
  wire [31:0]        writeDataVec_data_unreadData_92;
  assign writeDataVec_data_unreadData_92 = _GEN_169;
  wire [7:0]         writeDataVec_data_dataElement_28 = writeDataVec_data_dataIsRead_28 ? waiteReadData_28[7:0] : writeDataVec_data_unreadData_28[7:0];
  wire               writeDataVec_data_dataIsRead_29 = waiteReadDataPipeReg_needRead[29];
  wire               writeDataVec_data_dataIsRead_61 = waiteReadDataPipeReg_needRead[29];
  wire               writeDataVec_data_dataIsRead_93 = waiteReadDataPipeReg_needRead[29];
  wire [31:0]        _GEN_170 = waiteReadDataPipeReg_replaceVs1[29] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_29;
  assign writeDataVec_data_unreadData_29 = _GEN_170;
  wire [31:0]        writeDataVec_data_unreadData_61;
  assign writeDataVec_data_unreadData_61 = _GEN_170;
  wire [31:0]        writeDataVec_data_unreadData_93;
  assign writeDataVec_data_unreadData_93 = _GEN_170;
  wire [7:0]         writeDataVec_data_dataElement_29 = writeDataVec_data_dataIsRead_29 ? waiteReadData_29[7:0] : writeDataVec_data_unreadData_29[7:0];
  wire               writeDataVec_data_dataIsRead_30 = waiteReadDataPipeReg_needRead[30];
  wire               writeDataVec_data_dataIsRead_62 = waiteReadDataPipeReg_needRead[30];
  wire               writeDataVec_data_dataIsRead_94 = waiteReadDataPipeReg_needRead[30];
  wire [31:0]        _GEN_174 = waiteReadDataPipeReg_replaceVs1[30] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_30;
  assign writeDataVec_data_unreadData_30 = _GEN_174;
  wire [31:0]        writeDataVec_data_unreadData_62;
  assign writeDataVec_data_unreadData_62 = _GEN_174;
  wire [31:0]        writeDataVec_data_unreadData_94;
  assign writeDataVec_data_unreadData_94 = _GEN_174;
  wire [7:0]         writeDataVec_data_dataElement_30 = writeDataVec_data_dataIsRead_30 ? waiteReadData_30[7:0] : writeDataVec_data_unreadData_30[7:0];
  wire               writeDataVec_data_dataIsRead_31 = waiteReadDataPipeReg_needRead[31];
  wire               writeDataVec_data_dataIsRead_63 = waiteReadDataPipeReg_needRead[31];
  wire               writeDataVec_data_dataIsRead_95 = waiteReadDataPipeReg_needRead[31];
  wire [31:0]        _GEN_175 = waiteReadDataPipeReg_replaceVs1[31] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_31;
  assign writeDataVec_data_unreadData_31 = _GEN_175;
  wire [31:0]        writeDataVec_data_unreadData_63;
  assign writeDataVec_data_unreadData_63 = _GEN_175;
  wire [31:0]        writeDataVec_data_unreadData_95;
  assign writeDataVec_data_unreadData_95 = _GEN_175;
  wire [7:0]         writeDataVec_data_dataElement_31 = writeDataVec_data_dataIsRead_31 ? waiteReadData_31[7:0] : writeDataVec_data_unreadData_31[7:0];
  wire [15:0]        writeDataVec_data_lo_lo_lo_lo = {writeDataVec_data_dataElement_1, writeDataVec_data_dataElement};
  wire [15:0]        writeDataVec_data_lo_lo_lo_hi = {writeDataVec_data_dataElement_3, writeDataVec_data_dataElement_2};
  wire [31:0]        writeDataVec_data_lo_lo_lo = {writeDataVec_data_lo_lo_lo_hi, writeDataVec_data_lo_lo_lo_lo};
  wire [15:0]        writeDataVec_data_lo_lo_hi_lo = {writeDataVec_data_dataElement_5, writeDataVec_data_dataElement_4};
  wire [15:0]        writeDataVec_data_lo_lo_hi_hi = {writeDataVec_data_dataElement_7, writeDataVec_data_dataElement_6};
  wire [31:0]        writeDataVec_data_lo_lo_hi = {writeDataVec_data_lo_lo_hi_hi, writeDataVec_data_lo_lo_hi_lo};
  wire [63:0]        writeDataVec_data_lo_lo = {writeDataVec_data_lo_lo_hi, writeDataVec_data_lo_lo_lo};
  wire [15:0]        writeDataVec_data_lo_hi_lo_lo = {writeDataVec_data_dataElement_9, writeDataVec_data_dataElement_8};
  wire [15:0]        writeDataVec_data_lo_hi_lo_hi = {writeDataVec_data_dataElement_11, writeDataVec_data_dataElement_10};
  wire [31:0]        writeDataVec_data_lo_hi_lo = {writeDataVec_data_lo_hi_lo_hi, writeDataVec_data_lo_hi_lo_lo};
  wire [15:0]        writeDataVec_data_lo_hi_hi_lo = {writeDataVec_data_dataElement_13, writeDataVec_data_dataElement_12};
  wire [15:0]        writeDataVec_data_lo_hi_hi_hi = {writeDataVec_data_dataElement_15, writeDataVec_data_dataElement_14};
  wire [31:0]        writeDataVec_data_lo_hi_hi = {writeDataVec_data_lo_hi_hi_hi, writeDataVec_data_lo_hi_hi_lo};
  wire [63:0]        writeDataVec_data_lo_hi = {writeDataVec_data_lo_hi_hi, writeDataVec_data_lo_hi_lo};
  wire [127:0]       writeDataVec_data_lo = {writeDataVec_data_lo_hi, writeDataVec_data_lo_lo};
  wire [15:0]        writeDataVec_data_hi_lo_lo_lo = {writeDataVec_data_dataElement_17, writeDataVec_data_dataElement_16};
  wire [15:0]        writeDataVec_data_hi_lo_lo_hi = {writeDataVec_data_dataElement_19, writeDataVec_data_dataElement_18};
  wire [31:0]        writeDataVec_data_hi_lo_lo = {writeDataVec_data_hi_lo_lo_hi, writeDataVec_data_hi_lo_lo_lo};
  wire [15:0]        writeDataVec_data_hi_lo_hi_lo = {writeDataVec_data_dataElement_21, writeDataVec_data_dataElement_20};
  wire [15:0]        writeDataVec_data_hi_lo_hi_hi = {writeDataVec_data_dataElement_23, writeDataVec_data_dataElement_22};
  wire [31:0]        writeDataVec_data_hi_lo_hi = {writeDataVec_data_hi_lo_hi_hi, writeDataVec_data_hi_lo_hi_lo};
  wire [63:0]        writeDataVec_data_hi_lo = {writeDataVec_data_hi_lo_hi, writeDataVec_data_hi_lo_lo};
  wire [15:0]        writeDataVec_data_hi_hi_lo_lo = {writeDataVec_data_dataElement_25, writeDataVec_data_dataElement_24};
  wire [15:0]        writeDataVec_data_hi_hi_lo_hi = {writeDataVec_data_dataElement_27, writeDataVec_data_dataElement_26};
  wire [31:0]        writeDataVec_data_hi_hi_lo = {writeDataVec_data_hi_hi_lo_hi, writeDataVec_data_hi_hi_lo_lo};
  wire [15:0]        writeDataVec_data_hi_hi_hi_lo = {writeDataVec_data_dataElement_29, writeDataVec_data_dataElement_28};
  wire [15:0]        writeDataVec_data_hi_hi_hi_hi = {writeDataVec_data_dataElement_31, writeDataVec_data_dataElement_30};
  wire [31:0]        writeDataVec_data_hi_hi_hi = {writeDataVec_data_hi_hi_hi_hi, writeDataVec_data_hi_hi_hi_lo};
  wire [63:0]        writeDataVec_data_hi_hi = {writeDataVec_data_hi_hi_hi, writeDataVec_data_hi_hi_lo};
  wire [127:0]       writeDataVec_data_hi = {writeDataVec_data_hi_hi, writeDataVec_data_hi_lo};
  wire [255:0]       writeDataVec_data = {writeDataVec_data_hi, writeDataVec_data_lo};
  wire [1278:0]      writeDataVec_shifterData = {1023'h0, writeDataVec_data} << {1269'h0, executeIndexVec_0, 8'h0};
  wire [1023:0]      writeDataVec_0 = writeDataVec_shifterData[1023:0];
  wire [15:0]        writeDataVec_data_dataElement_32 = writeDataVec_data_dataIsRead_32 ? waiteReadData_0[15:0] : writeDataVec_data_unreadData_32[15:0];
  wire [15:0]        writeDataVec_data_dataElement_33 = writeDataVec_data_dataIsRead_33 ? waiteReadData_1[15:0] : writeDataVec_data_unreadData_33[15:0];
  wire [15:0]        writeDataVec_data_dataElement_34 = writeDataVec_data_dataIsRead_34 ? waiteReadData_2[15:0] : writeDataVec_data_unreadData_34[15:0];
  wire [15:0]        writeDataVec_data_dataElement_35 = writeDataVec_data_dataIsRead_35 ? waiteReadData_3[15:0] : writeDataVec_data_unreadData_35[15:0];
  wire [15:0]        writeDataVec_data_dataElement_36 = writeDataVec_data_dataIsRead_36 ? waiteReadData_4[15:0] : writeDataVec_data_unreadData_36[15:0];
  wire [15:0]        writeDataVec_data_dataElement_37 = writeDataVec_data_dataIsRead_37 ? waiteReadData_5[15:0] : writeDataVec_data_unreadData_37[15:0];
  wire [15:0]        writeDataVec_data_dataElement_38 = writeDataVec_data_dataIsRead_38 ? waiteReadData_6[15:0] : writeDataVec_data_unreadData_38[15:0];
  wire [15:0]        writeDataVec_data_dataElement_39 = writeDataVec_data_dataIsRead_39 ? waiteReadData_7[15:0] : writeDataVec_data_unreadData_39[15:0];
  wire [15:0]        writeDataVec_data_dataElement_40 = writeDataVec_data_dataIsRead_40 ? waiteReadData_8[15:0] : writeDataVec_data_unreadData_40[15:0];
  wire [15:0]        writeDataVec_data_dataElement_41 = writeDataVec_data_dataIsRead_41 ? waiteReadData_9[15:0] : writeDataVec_data_unreadData_41[15:0];
  wire [15:0]        writeDataVec_data_dataElement_42 = writeDataVec_data_dataIsRead_42 ? waiteReadData_10[15:0] : writeDataVec_data_unreadData_42[15:0];
  wire [15:0]        writeDataVec_data_dataElement_43 = writeDataVec_data_dataIsRead_43 ? waiteReadData_11[15:0] : writeDataVec_data_unreadData_43[15:0];
  wire [15:0]        writeDataVec_data_dataElement_44 = writeDataVec_data_dataIsRead_44 ? waiteReadData_12[15:0] : writeDataVec_data_unreadData_44[15:0];
  wire [15:0]        writeDataVec_data_dataElement_45 = writeDataVec_data_dataIsRead_45 ? waiteReadData_13[15:0] : writeDataVec_data_unreadData_45[15:0];
  wire [15:0]        writeDataVec_data_dataElement_46 = writeDataVec_data_dataIsRead_46 ? waiteReadData_14[15:0] : writeDataVec_data_unreadData_46[15:0];
  wire [15:0]        writeDataVec_data_dataElement_47 = writeDataVec_data_dataIsRead_47 ? waiteReadData_15[15:0] : writeDataVec_data_unreadData_47[15:0];
  wire [15:0]        writeDataVec_data_dataElement_48 = writeDataVec_data_dataIsRead_48 ? waiteReadData_16[15:0] : writeDataVec_data_unreadData_48[15:0];
  wire [15:0]        writeDataVec_data_dataElement_49 = writeDataVec_data_dataIsRead_49 ? waiteReadData_17[15:0] : writeDataVec_data_unreadData_49[15:0];
  wire [15:0]        writeDataVec_data_dataElement_50 = writeDataVec_data_dataIsRead_50 ? waiteReadData_18[15:0] : writeDataVec_data_unreadData_50[15:0];
  wire [15:0]        writeDataVec_data_dataElement_51 = writeDataVec_data_dataIsRead_51 ? waiteReadData_19[15:0] : writeDataVec_data_unreadData_51[15:0];
  wire [15:0]        writeDataVec_data_dataElement_52 = writeDataVec_data_dataIsRead_52 ? waiteReadData_20[15:0] : writeDataVec_data_unreadData_52[15:0];
  wire [15:0]        writeDataVec_data_dataElement_53 = writeDataVec_data_dataIsRead_53 ? waiteReadData_21[15:0] : writeDataVec_data_unreadData_53[15:0];
  wire [15:0]        writeDataVec_data_dataElement_54 = writeDataVec_data_dataIsRead_54 ? waiteReadData_22[15:0] : writeDataVec_data_unreadData_54[15:0];
  wire [15:0]        writeDataVec_data_dataElement_55 = writeDataVec_data_dataIsRead_55 ? waiteReadData_23[15:0] : writeDataVec_data_unreadData_55[15:0];
  wire [15:0]        writeDataVec_data_dataElement_56 = writeDataVec_data_dataIsRead_56 ? waiteReadData_24[15:0] : writeDataVec_data_unreadData_56[15:0];
  wire [15:0]        writeDataVec_data_dataElement_57 = writeDataVec_data_dataIsRead_57 ? waiteReadData_25[15:0] : writeDataVec_data_unreadData_57[15:0];
  wire [15:0]        writeDataVec_data_dataElement_58 = writeDataVec_data_dataIsRead_58 ? waiteReadData_26[15:0] : writeDataVec_data_unreadData_58[15:0];
  wire [15:0]        writeDataVec_data_dataElement_59 = writeDataVec_data_dataIsRead_59 ? waiteReadData_27[15:0] : writeDataVec_data_unreadData_59[15:0];
  wire [15:0]        writeDataVec_data_dataElement_60 = writeDataVec_data_dataIsRead_60 ? waiteReadData_28[15:0] : writeDataVec_data_unreadData_60[15:0];
  wire [15:0]        writeDataVec_data_dataElement_61 = writeDataVec_data_dataIsRead_61 ? waiteReadData_29[15:0] : writeDataVec_data_unreadData_61[15:0];
  wire [15:0]        writeDataVec_data_dataElement_62 = writeDataVec_data_dataIsRead_62 ? waiteReadData_30[15:0] : writeDataVec_data_unreadData_62[15:0];
  wire [15:0]        writeDataVec_data_dataElement_63 = writeDataVec_data_dataIsRead_63 ? waiteReadData_31[15:0] : writeDataVec_data_unreadData_63[15:0];
  wire [31:0]        writeDataVec_data_lo_lo_lo_lo_1 = {writeDataVec_data_dataElement_33, writeDataVec_data_dataElement_32};
  wire [31:0]        writeDataVec_data_lo_lo_lo_hi_1 = {writeDataVec_data_dataElement_35, writeDataVec_data_dataElement_34};
  wire [63:0]        writeDataVec_data_lo_lo_lo_1 = {writeDataVec_data_lo_lo_lo_hi_1, writeDataVec_data_lo_lo_lo_lo_1};
  wire [31:0]        writeDataVec_data_lo_lo_hi_lo_1 = {writeDataVec_data_dataElement_37, writeDataVec_data_dataElement_36};
  wire [31:0]        writeDataVec_data_lo_lo_hi_hi_1 = {writeDataVec_data_dataElement_39, writeDataVec_data_dataElement_38};
  wire [63:0]        writeDataVec_data_lo_lo_hi_1 = {writeDataVec_data_lo_lo_hi_hi_1, writeDataVec_data_lo_lo_hi_lo_1};
  wire [127:0]       writeDataVec_data_lo_lo_1 = {writeDataVec_data_lo_lo_hi_1, writeDataVec_data_lo_lo_lo_1};
  wire [31:0]        writeDataVec_data_lo_hi_lo_lo_1 = {writeDataVec_data_dataElement_41, writeDataVec_data_dataElement_40};
  wire [31:0]        writeDataVec_data_lo_hi_lo_hi_1 = {writeDataVec_data_dataElement_43, writeDataVec_data_dataElement_42};
  wire [63:0]        writeDataVec_data_lo_hi_lo_1 = {writeDataVec_data_lo_hi_lo_hi_1, writeDataVec_data_lo_hi_lo_lo_1};
  wire [31:0]        writeDataVec_data_lo_hi_hi_lo_1 = {writeDataVec_data_dataElement_45, writeDataVec_data_dataElement_44};
  wire [31:0]        writeDataVec_data_lo_hi_hi_hi_1 = {writeDataVec_data_dataElement_47, writeDataVec_data_dataElement_46};
  wire [63:0]        writeDataVec_data_lo_hi_hi_1 = {writeDataVec_data_lo_hi_hi_hi_1, writeDataVec_data_lo_hi_hi_lo_1};
  wire [127:0]       writeDataVec_data_lo_hi_1 = {writeDataVec_data_lo_hi_hi_1, writeDataVec_data_lo_hi_lo_1};
  wire [255:0]       writeDataVec_data_lo_1 = {writeDataVec_data_lo_hi_1, writeDataVec_data_lo_lo_1};
  wire [31:0]        writeDataVec_data_hi_lo_lo_lo_1 = {writeDataVec_data_dataElement_49, writeDataVec_data_dataElement_48};
  wire [31:0]        writeDataVec_data_hi_lo_lo_hi_1 = {writeDataVec_data_dataElement_51, writeDataVec_data_dataElement_50};
  wire [63:0]        writeDataVec_data_hi_lo_lo_1 = {writeDataVec_data_hi_lo_lo_hi_1, writeDataVec_data_hi_lo_lo_lo_1};
  wire [31:0]        writeDataVec_data_hi_lo_hi_lo_1 = {writeDataVec_data_dataElement_53, writeDataVec_data_dataElement_52};
  wire [31:0]        writeDataVec_data_hi_lo_hi_hi_1 = {writeDataVec_data_dataElement_55, writeDataVec_data_dataElement_54};
  wire [63:0]        writeDataVec_data_hi_lo_hi_1 = {writeDataVec_data_hi_lo_hi_hi_1, writeDataVec_data_hi_lo_hi_lo_1};
  wire [127:0]       writeDataVec_data_hi_lo_1 = {writeDataVec_data_hi_lo_hi_1, writeDataVec_data_hi_lo_lo_1};
  wire [31:0]        writeDataVec_data_hi_hi_lo_lo_1 = {writeDataVec_data_dataElement_57, writeDataVec_data_dataElement_56};
  wire [31:0]        writeDataVec_data_hi_hi_lo_hi_1 = {writeDataVec_data_dataElement_59, writeDataVec_data_dataElement_58};
  wire [63:0]        writeDataVec_data_hi_hi_lo_1 = {writeDataVec_data_hi_hi_lo_hi_1, writeDataVec_data_hi_hi_lo_lo_1};
  wire [31:0]        writeDataVec_data_hi_hi_hi_lo_1 = {writeDataVec_data_dataElement_61, writeDataVec_data_dataElement_60};
  wire [31:0]        writeDataVec_data_hi_hi_hi_hi_1 = {writeDataVec_data_dataElement_63, writeDataVec_data_dataElement_62};
  wire [63:0]        writeDataVec_data_hi_hi_hi_1 = {writeDataVec_data_hi_hi_hi_hi_1, writeDataVec_data_hi_hi_hi_lo_1};
  wire [127:0]       writeDataVec_data_hi_hi_1 = {writeDataVec_data_hi_hi_hi_1, writeDataVec_data_hi_hi_lo_1};
  wire [255:0]       writeDataVec_data_hi_1 = {writeDataVec_data_hi_hi_1, writeDataVec_data_hi_lo_1};
  wire [511:0]       writeDataVec_data_1 = {writeDataVec_data_hi_1, writeDataVec_data_lo_1};
  wire [1534:0]      writeDataVec_shifterData_1 = {1023'h0, writeDataVec_data_1} << {1525'h0, executeIndexVec_1, 8'h0};
  wire [1023:0]      writeDataVec_1 = writeDataVec_shifterData_1[1023:0];
  wire [31:0]        writeDataVec_data_dataElement_64 = writeDataVec_data_dataIsRead_64 ? waiteReadData_0 : writeDataVec_data_unreadData_64;
  wire [31:0]        writeDataVec_data_dataElement_65 = writeDataVec_data_dataIsRead_65 ? waiteReadData_1 : writeDataVec_data_unreadData_65;
  wire [31:0]        writeDataVec_data_dataElement_66 = writeDataVec_data_dataIsRead_66 ? waiteReadData_2 : writeDataVec_data_unreadData_66;
  wire [31:0]        writeDataVec_data_dataElement_67 = writeDataVec_data_dataIsRead_67 ? waiteReadData_3 : writeDataVec_data_unreadData_67;
  wire [31:0]        writeDataVec_data_dataElement_68 = writeDataVec_data_dataIsRead_68 ? waiteReadData_4 : writeDataVec_data_unreadData_68;
  wire [31:0]        writeDataVec_data_dataElement_69 = writeDataVec_data_dataIsRead_69 ? waiteReadData_5 : writeDataVec_data_unreadData_69;
  wire [31:0]        writeDataVec_data_dataElement_70 = writeDataVec_data_dataIsRead_70 ? waiteReadData_6 : writeDataVec_data_unreadData_70;
  wire [31:0]        writeDataVec_data_dataElement_71 = writeDataVec_data_dataIsRead_71 ? waiteReadData_7 : writeDataVec_data_unreadData_71;
  wire [31:0]        writeDataVec_data_dataElement_72 = writeDataVec_data_dataIsRead_72 ? waiteReadData_8 : writeDataVec_data_unreadData_72;
  wire [31:0]        writeDataVec_data_dataElement_73 = writeDataVec_data_dataIsRead_73 ? waiteReadData_9 : writeDataVec_data_unreadData_73;
  wire [31:0]        writeDataVec_data_dataElement_74 = writeDataVec_data_dataIsRead_74 ? waiteReadData_10 : writeDataVec_data_unreadData_74;
  wire [31:0]        writeDataVec_data_dataElement_75 = writeDataVec_data_dataIsRead_75 ? waiteReadData_11 : writeDataVec_data_unreadData_75;
  wire [31:0]        writeDataVec_data_dataElement_76 = writeDataVec_data_dataIsRead_76 ? waiteReadData_12 : writeDataVec_data_unreadData_76;
  wire [31:0]        writeDataVec_data_dataElement_77 = writeDataVec_data_dataIsRead_77 ? waiteReadData_13 : writeDataVec_data_unreadData_77;
  wire [31:0]        writeDataVec_data_dataElement_78 = writeDataVec_data_dataIsRead_78 ? waiteReadData_14 : writeDataVec_data_unreadData_78;
  wire [31:0]        writeDataVec_data_dataElement_79 = writeDataVec_data_dataIsRead_79 ? waiteReadData_15 : writeDataVec_data_unreadData_79;
  wire [31:0]        writeDataVec_data_dataElement_80 = writeDataVec_data_dataIsRead_80 ? waiteReadData_16 : writeDataVec_data_unreadData_80;
  wire [31:0]        writeDataVec_data_dataElement_81 = writeDataVec_data_dataIsRead_81 ? waiteReadData_17 : writeDataVec_data_unreadData_81;
  wire [31:0]        writeDataVec_data_dataElement_82 = writeDataVec_data_dataIsRead_82 ? waiteReadData_18 : writeDataVec_data_unreadData_82;
  wire [31:0]        writeDataVec_data_dataElement_83 = writeDataVec_data_dataIsRead_83 ? waiteReadData_19 : writeDataVec_data_unreadData_83;
  wire [31:0]        writeDataVec_data_dataElement_84 = writeDataVec_data_dataIsRead_84 ? waiteReadData_20 : writeDataVec_data_unreadData_84;
  wire [31:0]        writeDataVec_data_dataElement_85 = writeDataVec_data_dataIsRead_85 ? waiteReadData_21 : writeDataVec_data_unreadData_85;
  wire [31:0]        writeDataVec_data_dataElement_86 = writeDataVec_data_dataIsRead_86 ? waiteReadData_22 : writeDataVec_data_unreadData_86;
  wire [31:0]        writeDataVec_data_dataElement_87 = writeDataVec_data_dataIsRead_87 ? waiteReadData_23 : writeDataVec_data_unreadData_87;
  wire [31:0]        writeDataVec_data_dataElement_88 = writeDataVec_data_dataIsRead_88 ? waiteReadData_24 : writeDataVec_data_unreadData_88;
  wire [31:0]        writeDataVec_data_dataElement_89 = writeDataVec_data_dataIsRead_89 ? waiteReadData_25 : writeDataVec_data_unreadData_89;
  wire [31:0]        writeDataVec_data_dataElement_90 = writeDataVec_data_dataIsRead_90 ? waiteReadData_26 : writeDataVec_data_unreadData_90;
  wire [31:0]        writeDataVec_data_dataElement_91 = writeDataVec_data_dataIsRead_91 ? waiteReadData_27 : writeDataVec_data_unreadData_91;
  wire [31:0]        writeDataVec_data_dataElement_92 = writeDataVec_data_dataIsRead_92 ? waiteReadData_28 : writeDataVec_data_unreadData_92;
  wire [31:0]        writeDataVec_data_dataElement_93 = writeDataVec_data_dataIsRead_93 ? waiteReadData_29 : writeDataVec_data_unreadData_93;
  wire [31:0]        writeDataVec_data_dataElement_94 = writeDataVec_data_dataIsRead_94 ? waiteReadData_30 : writeDataVec_data_unreadData_94;
  wire [31:0]        writeDataVec_data_dataElement_95 = writeDataVec_data_dataIsRead_95 ? waiteReadData_31 : writeDataVec_data_unreadData_95;
  wire [63:0]        writeDataVec_data_lo_lo_lo_lo_2 = {writeDataVec_data_dataElement_65, writeDataVec_data_dataElement_64};
  wire [63:0]        writeDataVec_data_lo_lo_lo_hi_2 = {writeDataVec_data_dataElement_67, writeDataVec_data_dataElement_66};
  wire [127:0]       writeDataVec_data_lo_lo_lo_2 = {writeDataVec_data_lo_lo_lo_hi_2, writeDataVec_data_lo_lo_lo_lo_2};
  wire [63:0]        writeDataVec_data_lo_lo_hi_lo_2 = {writeDataVec_data_dataElement_69, writeDataVec_data_dataElement_68};
  wire [63:0]        writeDataVec_data_lo_lo_hi_hi_2 = {writeDataVec_data_dataElement_71, writeDataVec_data_dataElement_70};
  wire [127:0]       writeDataVec_data_lo_lo_hi_2 = {writeDataVec_data_lo_lo_hi_hi_2, writeDataVec_data_lo_lo_hi_lo_2};
  wire [255:0]       writeDataVec_data_lo_lo_2 = {writeDataVec_data_lo_lo_hi_2, writeDataVec_data_lo_lo_lo_2};
  wire [63:0]        writeDataVec_data_lo_hi_lo_lo_2 = {writeDataVec_data_dataElement_73, writeDataVec_data_dataElement_72};
  wire [63:0]        writeDataVec_data_lo_hi_lo_hi_2 = {writeDataVec_data_dataElement_75, writeDataVec_data_dataElement_74};
  wire [127:0]       writeDataVec_data_lo_hi_lo_2 = {writeDataVec_data_lo_hi_lo_hi_2, writeDataVec_data_lo_hi_lo_lo_2};
  wire [63:0]        writeDataVec_data_lo_hi_hi_lo_2 = {writeDataVec_data_dataElement_77, writeDataVec_data_dataElement_76};
  wire [63:0]        writeDataVec_data_lo_hi_hi_hi_2 = {writeDataVec_data_dataElement_79, writeDataVec_data_dataElement_78};
  wire [127:0]       writeDataVec_data_lo_hi_hi_2 = {writeDataVec_data_lo_hi_hi_hi_2, writeDataVec_data_lo_hi_hi_lo_2};
  wire [255:0]       writeDataVec_data_lo_hi_2 = {writeDataVec_data_lo_hi_hi_2, writeDataVec_data_lo_hi_lo_2};
  wire [511:0]       writeDataVec_data_lo_2 = {writeDataVec_data_lo_hi_2, writeDataVec_data_lo_lo_2};
  wire [63:0]        writeDataVec_data_hi_lo_lo_lo_2 = {writeDataVec_data_dataElement_81, writeDataVec_data_dataElement_80};
  wire [63:0]        writeDataVec_data_hi_lo_lo_hi_2 = {writeDataVec_data_dataElement_83, writeDataVec_data_dataElement_82};
  wire [127:0]       writeDataVec_data_hi_lo_lo_2 = {writeDataVec_data_hi_lo_lo_hi_2, writeDataVec_data_hi_lo_lo_lo_2};
  wire [63:0]        writeDataVec_data_hi_lo_hi_lo_2 = {writeDataVec_data_dataElement_85, writeDataVec_data_dataElement_84};
  wire [63:0]        writeDataVec_data_hi_lo_hi_hi_2 = {writeDataVec_data_dataElement_87, writeDataVec_data_dataElement_86};
  wire [127:0]       writeDataVec_data_hi_lo_hi_2 = {writeDataVec_data_hi_lo_hi_hi_2, writeDataVec_data_hi_lo_hi_lo_2};
  wire [255:0]       writeDataVec_data_hi_lo_2 = {writeDataVec_data_hi_lo_hi_2, writeDataVec_data_hi_lo_lo_2};
  wire [63:0]        writeDataVec_data_hi_hi_lo_lo_2 = {writeDataVec_data_dataElement_89, writeDataVec_data_dataElement_88};
  wire [63:0]        writeDataVec_data_hi_hi_lo_hi_2 = {writeDataVec_data_dataElement_91, writeDataVec_data_dataElement_90};
  wire [127:0]       writeDataVec_data_hi_hi_lo_2 = {writeDataVec_data_hi_hi_lo_hi_2, writeDataVec_data_hi_hi_lo_lo_2};
  wire [63:0]        writeDataVec_data_hi_hi_hi_lo_2 = {writeDataVec_data_dataElement_93, writeDataVec_data_dataElement_92};
  wire [63:0]        writeDataVec_data_hi_hi_hi_hi_2 = {writeDataVec_data_dataElement_95, writeDataVec_data_dataElement_94};
  wire [127:0]       writeDataVec_data_hi_hi_hi_2 = {writeDataVec_data_hi_hi_hi_hi_2, writeDataVec_data_hi_hi_hi_lo_2};
  wire [255:0]       writeDataVec_data_hi_hi_2 = {writeDataVec_data_hi_hi_hi_2, writeDataVec_data_hi_hi_lo_2};
  wire [511:0]       writeDataVec_data_hi_2 = {writeDataVec_data_hi_hi_2, writeDataVec_data_hi_lo_2};
  wire [1023:0]      writeDataVec_data_2 = {writeDataVec_data_hi_2, writeDataVec_data_lo_2};
  wire [1534:0]      writeDataVec_shifterData_2 = {511'h0, writeDataVec_data_2};
  wire [1023:0]      writeDataVec_2 = writeDataVec_shifterData_2[1023:0];
  wire [1023:0]      writeData = (sew1H[0] ? writeDataVec_0 : 1024'h0) | (sew1H[1] ? writeDataVec_1 : 1024'h0) | (sew1H[2] ? writeDataVec_2 : 1024'h0);
  wire [1:0]         writeMaskVec_mask_lo_lo_lo_lo = waiteReadDataPipeReg_sourceValid[1:0];
  wire [1:0]         writeMaskVec_mask_lo_lo_lo_hi = waiteReadDataPipeReg_sourceValid[3:2];
  wire [3:0]         writeMaskVec_mask_lo_lo_lo = {writeMaskVec_mask_lo_lo_lo_hi, writeMaskVec_mask_lo_lo_lo_lo};
  wire [1:0]         writeMaskVec_mask_lo_lo_hi_lo = waiteReadDataPipeReg_sourceValid[5:4];
  wire [1:0]         writeMaskVec_mask_lo_lo_hi_hi = waiteReadDataPipeReg_sourceValid[7:6];
  wire [3:0]         writeMaskVec_mask_lo_lo_hi = {writeMaskVec_mask_lo_lo_hi_hi, writeMaskVec_mask_lo_lo_hi_lo};
  wire [7:0]         writeMaskVec_mask_lo_lo = {writeMaskVec_mask_lo_lo_hi, writeMaskVec_mask_lo_lo_lo};
  wire [1:0]         writeMaskVec_mask_lo_hi_lo_lo = waiteReadDataPipeReg_sourceValid[9:8];
  wire [1:0]         writeMaskVec_mask_lo_hi_lo_hi = waiteReadDataPipeReg_sourceValid[11:10];
  wire [3:0]         writeMaskVec_mask_lo_hi_lo = {writeMaskVec_mask_lo_hi_lo_hi, writeMaskVec_mask_lo_hi_lo_lo};
  wire [1:0]         writeMaskVec_mask_lo_hi_hi_lo = waiteReadDataPipeReg_sourceValid[13:12];
  wire [1:0]         writeMaskVec_mask_lo_hi_hi_hi = waiteReadDataPipeReg_sourceValid[15:14];
  wire [3:0]         writeMaskVec_mask_lo_hi_hi = {writeMaskVec_mask_lo_hi_hi_hi, writeMaskVec_mask_lo_hi_hi_lo};
  wire [7:0]         writeMaskVec_mask_lo_hi = {writeMaskVec_mask_lo_hi_hi, writeMaskVec_mask_lo_hi_lo};
  wire [15:0]        writeMaskVec_mask_lo = {writeMaskVec_mask_lo_hi, writeMaskVec_mask_lo_lo};
  wire [1:0]         writeMaskVec_mask_hi_lo_lo_lo = waiteReadDataPipeReg_sourceValid[17:16];
  wire [1:0]         writeMaskVec_mask_hi_lo_lo_hi = waiteReadDataPipeReg_sourceValid[19:18];
  wire [3:0]         writeMaskVec_mask_hi_lo_lo = {writeMaskVec_mask_hi_lo_lo_hi, writeMaskVec_mask_hi_lo_lo_lo};
  wire [1:0]         writeMaskVec_mask_hi_lo_hi_lo = waiteReadDataPipeReg_sourceValid[21:20];
  wire [1:0]         writeMaskVec_mask_hi_lo_hi_hi = waiteReadDataPipeReg_sourceValid[23:22];
  wire [3:0]         writeMaskVec_mask_hi_lo_hi = {writeMaskVec_mask_hi_lo_hi_hi, writeMaskVec_mask_hi_lo_hi_lo};
  wire [7:0]         writeMaskVec_mask_hi_lo = {writeMaskVec_mask_hi_lo_hi, writeMaskVec_mask_hi_lo_lo};
  wire [1:0]         writeMaskVec_mask_hi_hi_lo_lo = waiteReadDataPipeReg_sourceValid[25:24];
  wire [1:0]         writeMaskVec_mask_hi_hi_lo_hi = waiteReadDataPipeReg_sourceValid[27:26];
  wire [3:0]         writeMaskVec_mask_hi_hi_lo = {writeMaskVec_mask_hi_hi_lo_hi, writeMaskVec_mask_hi_hi_lo_lo};
  wire [1:0]         writeMaskVec_mask_hi_hi_hi_lo = waiteReadDataPipeReg_sourceValid[29:28];
  wire [1:0]         writeMaskVec_mask_hi_hi_hi_hi = waiteReadDataPipeReg_sourceValid[31:30];
  wire [3:0]         writeMaskVec_mask_hi_hi_hi = {writeMaskVec_mask_hi_hi_hi_hi, writeMaskVec_mask_hi_hi_hi_lo};
  wire [7:0]         writeMaskVec_mask_hi_hi = {writeMaskVec_mask_hi_hi_hi, writeMaskVec_mask_hi_hi_lo};
  wire [15:0]        writeMaskVec_mask_hi = {writeMaskVec_mask_hi_hi, writeMaskVec_mask_hi_lo};
  wire [31:0]        writeMaskVec_mask = {writeMaskVec_mask_hi, writeMaskVec_mask_lo};
  wire [158:0]       writeMaskVec_shifterMask = {127'h0, writeMaskVec_mask} << {152'h0, executeIndexVec_0, 5'h0};
  wire [127:0]       writeMaskVec_0 = writeMaskVec_shifterMask[127:0];
  wire [3:0]         writeMaskVec_mask_lo_lo_lo_lo_1 = {{2{waiteReadDataPipeReg_sourceValid[1]}}, {2{waiteReadDataPipeReg_sourceValid[0]}}};
  wire [3:0]         writeMaskVec_mask_lo_lo_lo_hi_1 = {{2{waiteReadDataPipeReg_sourceValid[3]}}, {2{waiteReadDataPipeReg_sourceValid[2]}}};
  wire [7:0]         writeMaskVec_mask_lo_lo_lo_1 = {writeMaskVec_mask_lo_lo_lo_hi_1, writeMaskVec_mask_lo_lo_lo_lo_1};
  wire [3:0]         writeMaskVec_mask_lo_lo_hi_lo_1 = {{2{waiteReadDataPipeReg_sourceValid[5]}}, {2{waiteReadDataPipeReg_sourceValid[4]}}};
  wire [3:0]         writeMaskVec_mask_lo_lo_hi_hi_1 = {{2{waiteReadDataPipeReg_sourceValid[7]}}, {2{waiteReadDataPipeReg_sourceValid[6]}}};
  wire [7:0]         writeMaskVec_mask_lo_lo_hi_1 = {writeMaskVec_mask_lo_lo_hi_hi_1, writeMaskVec_mask_lo_lo_hi_lo_1};
  wire [15:0]        writeMaskVec_mask_lo_lo_1 = {writeMaskVec_mask_lo_lo_hi_1, writeMaskVec_mask_lo_lo_lo_1};
  wire [3:0]         writeMaskVec_mask_lo_hi_lo_lo_1 = {{2{waiteReadDataPipeReg_sourceValid[9]}}, {2{waiteReadDataPipeReg_sourceValid[8]}}};
  wire [3:0]         writeMaskVec_mask_lo_hi_lo_hi_1 = {{2{waiteReadDataPipeReg_sourceValid[11]}}, {2{waiteReadDataPipeReg_sourceValid[10]}}};
  wire [7:0]         writeMaskVec_mask_lo_hi_lo_1 = {writeMaskVec_mask_lo_hi_lo_hi_1, writeMaskVec_mask_lo_hi_lo_lo_1};
  wire [3:0]         writeMaskVec_mask_lo_hi_hi_lo_1 = {{2{waiteReadDataPipeReg_sourceValid[13]}}, {2{waiteReadDataPipeReg_sourceValid[12]}}};
  wire [3:0]         writeMaskVec_mask_lo_hi_hi_hi_1 = {{2{waiteReadDataPipeReg_sourceValid[15]}}, {2{waiteReadDataPipeReg_sourceValid[14]}}};
  wire [7:0]         writeMaskVec_mask_lo_hi_hi_1 = {writeMaskVec_mask_lo_hi_hi_hi_1, writeMaskVec_mask_lo_hi_hi_lo_1};
  wire [15:0]        writeMaskVec_mask_lo_hi_1 = {writeMaskVec_mask_lo_hi_hi_1, writeMaskVec_mask_lo_hi_lo_1};
  wire [31:0]        writeMaskVec_mask_lo_1 = {writeMaskVec_mask_lo_hi_1, writeMaskVec_mask_lo_lo_1};
  wire [3:0]         writeMaskVec_mask_hi_lo_lo_lo_1 = {{2{waiteReadDataPipeReg_sourceValid[17]}}, {2{waiteReadDataPipeReg_sourceValid[16]}}};
  wire [3:0]         writeMaskVec_mask_hi_lo_lo_hi_1 = {{2{waiteReadDataPipeReg_sourceValid[19]}}, {2{waiteReadDataPipeReg_sourceValid[18]}}};
  wire [7:0]         writeMaskVec_mask_hi_lo_lo_1 = {writeMaskVec_mask_hi_lo_lo_hi_1, writeMaskVec_mask_hi_lo_lo_lo_1};
  wire [3:0]         writeMaskVec_mask_hi_lo_hi_lo_1 = {{2{waiteReadDataPipeReg_sourceValid[21]}}, {2{waiteReadDataPipeReg_sourceValid[20]}}};
  wire [3:0]         writeMaskVec_mask_hi_lo_hi_hi_1 = {{2{waiteReadDataPipeReg_sourceValid[23]}}, {2{waiteReadDataPipeReg_sourceValid[22]}}};
  wire [7:0]         writeMaskVec_mask_hi_lo_hi_1 = {writeMaskVec_mask_hi_lo_hi_hi_1, writeMaskVec_mask_hi_lo_hi_lo_1};
  wire [15:0]        writeMaskVec_mask_hi_lo_1 = {writeMaskVec_mask_hi_lo_hi_1, writeMaskVec_mask_hi_lo_lo_1};
  wire [3:0]         writeMaskVec_mask_hi_hi_lo_lo_1 = {{2{waiteReadDataPipeReg_sourceValid[25]}}, {2{waiteReadDataPipeReg_sourceValid[24]}}};
  wire [3:0]         writeMaskVec_mask_hi_hi_lo_hi_1 = {{2{waiteReadDataPipeReg_sourceValid[27]}}, {2{waiteReadDataPipeReg_sourceValid[26]}}};
  wire [7:0]         writeMaskVec_mask_hi_hi_lo_1 = {writeMaskVec_mask_hi_hi_lo_hi_1, writeMaskVec_mask_hi_hi_lo_lo_1};
  wire [3:0]         writeMaskVec_mask_hi_hi_hi_lo_1 = {{2{waiteReadDataPipeReg_sourceValid[29]}}, {2{waiteReadDataPipeReg_sourceValid[28]}}};
  wire [3:0]         writeMaskVec_mask_hi_hi_hi_hi_1 = {{2{waiteReadDataPipeReg_sourceValid[31]}}, {2{waiteReadDataPipeReg_sourceValid[30]}}};
  wire [7:0]         writeMaskVec_mask_hi_hi_hi_1 = {writeMaskVec_mask_hi_hi_hi_hi_1, writeMaskVec_mask_hi_hi_hi_lo_1};
  wire [15:0]        writeMaskVec_mask_hi_hi_1 = {writeMaskVec_mask_hi_hi_hi_1, writeMaskVec_mask_hi_hi_lo_1};
  wire [31:0]        writeMaskVec_mask_hi_1 = {writeMaskVec_mask_hi_hi_1, writeMaskVec_mask_hi_lo_1};
  wire [63:0]        writeMaskVec_mask_1 = {writeMaskVec_mask_hi_1, writeMaskVec_mask_lo_1};
  wire [190:0]       writeMaskVec_shifterMask_1 = {127'h0, writeMaskVec_mask_1} << {184'h0, executeIndexVec_1, 5'h0};
  wire [127:0]       writeMaskVec_1 = writeMaskVec_shifterMask_1[127:0];
  wire [7:0]         writeMaskVec_mask_lo_lo_lo_lo_2 = {{4{waiteReadDataPipeReg_sourceValid[1]}}, {4{waiteReadDataPipeReg_sourceValid[0]}}};
  wire [7:0]         writeMaskVec_mask_lo_lo_lo_hi_2 = {{4{waiteReadDataPipeReg_sourceValid[3]}}, {4{waiteReadDataPipeReg_sourceValid[2]}}};
  wire [15:0]        writeMaskVec_mask_lo_lo_lo_2 = {writeMaskVec_mask_lo_lo_lo_hi_2, writeMaskVec_mask_lo_lo_lo_lo_2};
  wire [7:0]         writeMaskVec_mask_lo_lo_hi_lo_2 = {{4{waiteReadDataPipeReg_sourceValid[5]}}, {4{waiteReadDataPipeReg_sourceValid[4]}}};
  wire [7:0]         writeMaskVec_mask_lo_lo_hi_hi_2 = {{4{waiteReadDataPipeReg_sourceValid[7]}}, {4{waiteReadDataPipeReg_sourceValid[6]}}};
  wire [15:0]        writeMaskVec_mask_lo_lo_hi_2 = {writeMaskVec_mask_lo_lo_hi_hi_2, writeMaskVec_mask_lo_lo_hi_lo_2};
  wire [31:0]        writeMaskVec_mask_lo_lo_2 = {writeMaskVec_mask_lo_lo_hi_2, writeMaskVec_mask_lo_lo_lo_2};
  wire [7:0]         writeMaskVec_mask_lo_hi_lo_lo_2 = {{4{waiteReadDataPipeReg_sourceValid[9]}}, {4{waiteReadDataPipeReg_sourceValid[8]}}};
  wire [7:0]         writeMaskVec_mask_lo_hi_lo_hi_2 = {{4{waiteReadDataPipeReg_sourceValid[11]}}, {4{waiteReadDataPipeReg_sourceValid[10]}}};
  wire [15:0]        writeMaskVec_mask_lo_hi_lo_2 = {writeMaskVec_mask_lo_hi_lo_hi_2, writeMaskVec_mask_lo_hi_lo_lo_2};
  wire [7:0]         writeMaskVec_mask_lo_hi_hi_lo_2 = {{4{waiteReadDataPipeReg_sourceValid[13]}}, {4{waiteReadDataPipeReg_sourceValid[12]}}};
  wire [7:0]         writeMaskVec_mask_lo_hi_hi_hi_2 = {{4{waiteReadDataPipeReg_sourceValid[15]}}, {4{waiteReadDataPipeReg_sourceValid[14]}}};
  wire [15:0]        writeMaskVec_mask_lo_hi_hi_2 = {writeMaskVec_mask_lo_hi_hi_hi_2, writeMaskVec_mask_lo_hi_hi_lo_2};
  wire [31:0]        writeMaskVec_mask_lo_hi_2 = {writeMaskVec_mask_lo_hi_hi_2, writeMaskVec_mask_lo_hi_lo_2};
  wire [63:0]        writeMaskVec_mask_lo_2 = {writeMaskVec_mask_lo_hi_2, writeMaskVec_mask_lo_lo_2};
  wire [7:0]         writeMaskVec_mask_hi_lo_lo_lo_2 = {{4{waiteReadDataPipeReg_sourceValid[17]}}, {4{waiteReadDataPipeReg_sourceValid[16]}}};
  wire [7:0]         writeMaskVec_mask_hi_lo_lo_hi_2 = {{4{waiteReadDataPipeReg_sourceValid[19]}}, {4{waiteReadDataPipeReg_sourceValid[18]}}};
  wire [15:0]        writeMaskVec_mask_hi_lo_lo_2 = {writeMaskVec_mask_hi_lo_lo_hi_2, writeMaskVec_mask_hi_lo_lo_lo_2};
  wire [7:0]         writeMaskVec_mask_hi_lo_hi_lo_2 = {{4{waiteReadDataPipeReg_sourceValid[21]}}, {4{waiteReadDataPipeReg_sourceValid[20]}}};
  wire [7:0]         writeMaskVec_mask_hi_lo_hi_hi_2 = {{4{waiteReadDataPipeReg_sourceValid[23]}}, {4{waiteReadDataPipeReg_sourceValid[22]}}};
  wire [15:0]        writeMaskVec_mask_hi_lo_hi_2 = {writeMaskVec_mask_hi_lo_hi_hi_2, writeMaskVec_mask_hi_lo_hi_lo_2};
  wire [31:0]        writeMaskVec_mask_hi_lo_2 = {writeMaskVec_mask_hi_lo_hi_2, writeMaskVec_mask_hi_lo_lo_2};
  wire [7:0]         writeMaskVec_mask_hi_hi_lo_lo_2 = {{4{waiteReadDataPipeReg_sourceValid[25]}}, {4{waiteReadDataPipeReg_sourceValid[24]}}};
  wire [7:0]         writeMaskVec_mask_hi_hi_lo_hi_2 = {{4{waiteReadDataPipeReg_sourceValid[27]}}, {4{waiteReadDataPipeReg_sourceValid[26]}}};
  wire [15:0]        writeMaskVec_mask_hi_hi_lo_2 = {writeMaskVec_mask_hi_hi_lo_hi_2, writeMaskVec_mask_hi_hi_lo_lo_2};
  wire [7:0]         writeMaskVec_mask_hi_hi_hi_lo_2 = {{4{waiteReadDataPipeReg_sourceValid[29]}}, {4{waiteReadDataPipeReg_sourceValid[28]}}};
  wire [7:0]         writeMaskVec_mask_hi_hi_hi_hi_2 = {{4{waiteReadDataPipeReg_sourceValid[31]}}, {4{waiteReadDataPipeReg_sourceValid[30]}}};
  wire [15:0]        writeMaskVec_mask_hi_hi_hi_2 = {writeMaskVec_mask_hi_hi_hi_hi_2, writeMaskVec_mask_hi_hi_hi_lo_2};
  wire [31:0]        writeMaskVec_mask_hi_hi_2 = {writeMaskVec_mask_hi_hi_hi_2, writeMaskVec_mask_hi_hi_lo_2};
  wire [63:0]        writeMaskVec_mask_hi_2 = {writeMaskVec_mask_hi_hi_2, writeMaskVec_mask_hi_lo_2};
  wire [127:0]       writeMaskVec_mask_2 = {writeMaskVec_mask_hi_2, writeMaskVec_mask_lo_2};
  wire [190:0]       writeMaskVec_shifterMask_2 = {63'h0, writeMaskVec_mask_2};
  wire [127:0]       writeMaskVec_2 = writeMaskVec_shifterMask_2[127:0];
  wire [127:0]       writeMask = (sew1H[0] ? writeMaskVec_0 : 128'h0) | (sew1H[1] ? writeMaskVec_1 : 128'h0) | (sew1H[2] ? writeMaskVec_2 : 128'h0);
  wire [9:0]         _writeRequest_res_writeData_groupCounter_T_62 = {3'h0, waiteReadDataPipeReg_executeGroup} << instReg_sew;
  wire [4:0]         writeRequest_0_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_1_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_2_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_3_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_4_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_5_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_6_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_7_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_8_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_9_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_10_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_11_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_12_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_13_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_14_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_15_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_16_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_17_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_18_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_19_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_20_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_21_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_22_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_23_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_24_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_25_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_26_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_27_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_28_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_29_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_30_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [4:0]         writeRequest_31_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_62[6:2];
  wire [31:0]        writeRequest_0_writeData_data = writeData[31:0];
  wire [31:0]        writeRequest_1_writeData_data = writeData[63:32];
  wire [31:0]        writeRequest_2_writeData_data = writeData[95:64];
  wire [31:0]        writeRequest_3_writeData_data = writeData[127:96];
  wire [31:0]        writeRequest_4_writeData_data = writeData[159:128];
  wire [31:0]        writeRequest_5_writeData_data = writeData[191:160];
  wire [31:0]        writeRequest_6_writeData_data = writeData[223:192];
  wire [31:0]        writeRequest_7_writeData_data = writeData[255:224];
  wire [31:0]        writeRequest_8_writeData_data = writeData[287:256];
  wire [31:0]        writeRequest_9_writeData_data = writeData[319:288];
  wire [31:0]        writeRequest_10_writeData_data = writeData[351:320];
  wire [31:0]        writeRequest_11_writeData_data = writeData[383:352];
  wire [31:0]        writeRequest_12_writeData_data = writeData[415:384];
  wire [31:0]        writeRequest_13_writeData_data = writeData[447:416];
  wire [31:0]        writeRequest_14_writeData_data = writeData[479:448];
  wire [31:0]        writeRequest_15_writeData_data = writeData[511:480];
  wire [31:0]        writeRequest_16_writeData_data = writeData[543:512];
  wire [31:0]        writeRequest_17_writeData_data = writeData[575:544];
  wire [31:0]        writeRequest_18_writeData_data = writeData[607:576];
  wire [31:0]        writeRequest_19_writeData_data = writeData[639:608];
  wire [31:0]        writeRequest_20_writeData_data = writeData[671:640];
  wire [31:0]        writeRequest_21_writeData_data = writeData[703:672];
  wire [31:0]        writeRequest_22_writeData_data = writeData[735:704];
  wire [31:0]        writeRequest_23_writeData_data = writeData[767:736];
  wire [31:0]        writeRequest_24_writeData_data = writeData[799:768];
  wire [31:0]        writeRequest_25_writeData_data = writeData[831:800];
  wire [31:0]        writeRequest_26_writeData_data = writeData[863:832];
  wire [31:0]        writeRequest_27_writeData_data = writeData[895:864];
  wire [31:0]        writeRequest_28_writeData_data = writeData[927:896];
  wire [31:0]        writeRequest_29_writeData_data = writeData[959:928];
  wire [31:0]        writeRequest_30_writeData_data = writeData[991:960];
  wire [31:0]        writeRequest_31_writeData_data = writeData[1023:992];
  wire [3:0]         writeRequest_0_writeData_mask = writeMask[3:0];
  wire [3:0]         writeRequest_1_writeData_mask = writeMask[7:4];
  wire [3:0]         writeRequest_2_writeData_mask = writeMask[11:8];
  wire [3:0]         writeRequest_3_writeData_mask = writeMask[15:12];
  wire [3:0]         writeRequest_4_writeData_mask = writeMask[19:16];
  wire [3:0]         writeRequest_5_writeData_mask = writeMask[23:20];
  wire [3:0]         writeRequest_6_writeData_mask = writeMask[27:24];
  wire [3:0]         writeRequest_7_writeData_mask = writeMask[31:28];
  wire [3:0]         writeRequest_8_writeData_mask = writeMask[35:32];
  wire [3:0]         writeRequest_9_writeData_mask = writeMask[39:36];
  wire [3:0]         writeRequest_10_writeData_mask = writeMask[43:40];
  wire [3:0]         writeRequest_11_writeData_mask = writeMask[47:44];
  wire [3:0]         writeRequest_12_writeData_mask = writeMask[51:48];
  wire [3:0]         writeRequest_13_writeData_mask = writeMask[55:52];
  wire [3:0]         writeRequest_14_writeData_mask = writeMask[59:56];
  wire [3:0]         writeRequest_15_writeData_mask = writeMask[63:60];
  wire [3:0]         writeRequest_16_writeData_mask = writeMask[67:64];
  wire [3:0]         writeRequest_17_writeData_mask = writeMask[71:68];
  wire [3:0]         writeRequest_18_writeData_mask = writeMask[75:72];
  wire [3:0]         writeRequest_19_writeData_mask = writeMask[79:76];
  wire [3:0]         writeRequest_20_writeData_mask = writeMask[83:80];
  wire [3:0]         writeRequest_21_writeData_mask = writeMask[87:84];
  wire [3:0]         writeRequest_22_writeData_mask = writeMask[91:88];
  wire [3:0]         writeRequest_23_writeData_mask = writeMask[95:92];
  wire [3:0]         writeRequest_24_writeData_mask = writeMask[99:96];
  wire [3:0]         writeRequest_25_writeData_mask = writeMask[103:100];
  wire [3:0]         writeRequest_26_writeData_mask = writeMask[107:104];
  wire [3:0]         writeRequest_27_writeData_mask = writeMask[111:108];
  wire [3:0]         writeRequest_28_writeData_mask = writeMask[115:112];
  wire [3:0]         writeRequest_29_writeData_mask = writeMask[119:116];
  wire [3:0]         writeRequest_30_writeData_mask = writeMask[123:120];
  wire [3:0]         writeRequest_31_writeData_mask = writeMask[127:124];
  wire [1:0]         WillWriteLane_lo_lo_lo_lo = {|writeRequest_1_writeData_mask, |writeRequest_0_writeData_mask};
  wire [1:0]         WillWriteLane_lo_lo_lo_hi = {|writeRequest_3_writeData_mask, |writeRequest_2_writeData_mask};
  wire [3:0]         WillWriteLane_lo_lo_lo = {WillWriteLane_lo_lo_lo_hi, WillWriteLane_lo_lo_lo_lo};
  wire [1:0]         WillWriteLane_lo_lo_hi_lo = {|writeRequest_5_writeData_mask, |writeRequest_4_writeData_mask};
  wire [1:0]         WillWriteLane_lo_lo_hi_hi = {|writeRequest_7_writeData_mask, |writeRequest_6_writeData_mask};
  wire [3:0]         WillWriteLane_lo_lo_hi = {WillWriteLane_lo_lo_hi_hi, WillWriteLane_lo_lo_hi_lo};
  wire [7:0]         WillWriteLane_lo_lo = {WillWriteLane_lo_lo_hi, WillWriteLane_lo_lo_lo};
  wire [1:0]         WillWriteLane_lo_hi_lo_lo = {|writeRequest_9_writeData_mask, |writeRequest_8_writeData_mask};
  wire [1:0]         WillWriteLane_lo_hi_lo_hi = {|writeRequest_11_writeData_mask, |writeRequest_10_writeData_mask};
  wire [3:0]         WillWriteLane_lo_hi_lo = {WillWriteLane_lo_hi_lo_hi, WillWriteLane_lo_hi_lo_lo};
  wire [1:0]         WillWriteLane_lo_hi_hi_lo = {|writeRequest_13_writeData_mask, |writeRequest_12_writeData_mask};
  wire [1:0]         WillWriteLane_lo_hi_hi_hi = {|writeRequest_15_writeData_mask, |writeRequest_14_writeData_mask};
  wire [3:0]         WillWriteLane_lo_hi_hi = {WillWriteLane_lo_hi_hi_hi, WillWriteLane_lo_hi_hi_lo};
  wire [7:0]         WillWriteLane_lo_hi = {WillWriteLane_lo_hi_hi, WillWriteLane_lo_hi_lo};
  wire [15:0]        WillWriteLane_lo = {WillWriteLane_lo_hi, WillWriteLane_lo_lo};
  wire [1:0]         WillWriteLane_hi_lo_lo_lo = {|writeRequest_17_writeData_mask, |writeRequest_16_writeData_mask};
  wire [1:0]         WillWriteLane_hi_lo_lo_hi = {|writeRequest_19_writeData_mask, |writeRequest_18_writeData_mask};
  wire [3:0]         WillWriteLane_hi_lo_lo = {WillWriteLane_hi_lo_lo_hi, WillWriteLane_hi_lo_lo_lo};
  wire [1:0]         WillWriteLane_hi_lo_hi_lo = {|writeRequest_21_writeData_mask, |writeRequest_20_writeData_mask};
  wire [1:0]         WillWriteLane_hi_lo_hi_hi = {|writeRequest_23_writeData_mask, |writeRequest_22_writeData_mask};
  wire [3:0]         WillWriteLane_hi_lo_hi = {WillWriteLane_hi_lo_hi_hi, WillWriteLane_hi_lo_hi_lo};
  wire [7:0]         WillWriteLane_hi_lo = {WillWriteLane_hi_lo_hi, WillWriteLane_hi_lo_lo};
  wire [1:0]         WillWriteLane_hi_hi_lo_lo = {|writeRequest_25_writeData_mask, |writeRequest_24_writeData_mask};
  wire [1:0]         WillWriteLane_hi_hi_lo_hi = {|writeRequest_27_writeData_mask, |writeRequest_26_writeData_mask};
  wire [3:0]         WillWriteLane_hi_hi_lo = {WillWriteLane_hi_hi_lo_hi, WillWriteLane_hi_hi_lo_lo};
  wire [1:0]         WillWriteLane_hi_hi_hi_lo = {|writeRequest_29_writeData_mask, |writeRequest_28_writeData_mask};
  wire [1:0]         WillWriteLane_hi_hi_hi_hi = {|writeRequest_31_writeData_mask, |writeRequest_30_writeData_mask};
  wire [3:0]         WillWriteLane_hi_hi_hi = {WillWriteLane_hi_hi_hi_hi, WillWriteLane_hi_hi_hi_lo};
  wire [7:0]         WillWriteLane_hi_hi = {WillWriteLane_hi_hi_hi, WillWriteLane_hi_hi_lo};
  wire [15:0]        WillWriteLane_hi = {WillWriteLane_hi_hi, WillWriteLane_hi_lo};
  wire [31:0]        WillWriteLane = {WillWriteLane_hi, WillWriteLane_lo};
  wire               waiteStageDeqValid = waiteReadStageValid & (waiteReadSate == waiteReadDataPipeReg_needRead | waiteReadDataPipeReg_needRead == 32'h0);
  wire               waiteStageDeqReady;
  wire               waiteStageDeqFire = waiteStageDeqValid & waiteStageDeqReady;
  assign waiteStageEnqReady = ~waiteReadStageValid | waiteStageDeqFire;
  assign readWaitQueue_deq_ready = waiteStageEnqReady;
  wire               waiteStageEnqFire = readWaitQueue_deq_valid & waiteStageEnqReady;
  wire               isWaiteForThisData = waiteReadDataPipeReg_needRead[0] & ~(waiteReadSate[0]) & waiteReadStageValid;
  assign readData_readDataQueue_deq_ready = isWaiteForThisData | unitType[2] | compress | gatherWaiteRead | mvRd;
  assign isWaiteForThisData_1 = waiteReadDataPipeReg_needRead[1] & ~(waiteReadSate[1]) & waiteReadStageValid;
  assign readData_readDataQueue_1_deq_ready = isWaiteForThisData_1;
  assign isWaiteForThisData_2 = waiteReadDataPipeReg_needRead[2] & ~(waiteReadSate[2]) & waiteReadStageValid;
  assign readData_readDataQueue_2_deq_ready = isWaiteForThisData_2;
  assign isWaiteForThisData_3 = waiteReadDataPipeReg_needRead[3] & ~(waiteReadSate[3]) & waiteReadStageValid;
  assign readData_readDataQueue_3_deq_ready = isWaiteForThisData_3;
  assign isWaiteForThisData_4 = waiteReadDataPipeReg_needRead[4] & ~(waiteReadSate[4]) & waiteReadStageValid;
  assign readData_readDataQueue_4_deq_ready = isWaiteForThisData_4;
  assign isWaiteForThisData_5 = waiteReadDataPipeReg_needRead[5] & ~(waiteReadSate[5]) & waiteReadStageValid;
  assign readData_readDataQueue_5_deq_ready = isWaiteForThisData_5;
  assign isWaiteForThisData_6 = waiteReadDataPipeReg_needRead[6] & ~(waiteReadSate[6]) & waiteReadStageValid;
  assign readData_readDataQueue_6_deq_ready = isWaiteForThisData_6;
  assign isWaiteForThisData_7 = waiteReadDataPipeReg_needRead[7] & ~(waiteReadSate[7]) & waiteReadStageValid;
  assign readData_readDataQueue_7_deq_ready = isWaiteForThisData_7;
  assign isWaiteForThisData_8 = waiteReadDataPipeReg_needRead[8] & ~(waiteReadSate[8]) & waiteReadStageValid;
  assign readData_readDataQueue_8_deq_ready = isWaiteForThisData_8;
  assign isWaiteForThisData_9 = waiteReadDataPipeReg_needRead[9] & ~(waiteReadSate[9]) & waiteReadStageValid;
  assign readData_readDataQueue_9_deq_ready = isWaiteForThisData_9;
  assign isWaiteForThisData_10 = waiteReadDataPipeReg_needRead[10] & ~(waiteReadSate[10]) & waiteReadStageValid;
  assign readData_readDataQueue_10_deq_ready = isWaiteForThisData_10;
  assign isWaiteForThisData_11 = waiteReadDataPipeReg_needRead[11] & ~(waiteReadSate[11]) & waiteReadStageValid;
  assign readData_readDataQueue_11_deq_ready = isWaiteForThisData_11;
  assign isWaiteForThisData_12 = waiteReadDataPipeReg_needRead[12] & ~(waiteReadSate[12]) & waiteReadStageValid;
  assign readData_readDataQueue_12_deq_ready = isWaiteForThisData_12;
  assign isWaiteForThisData_13 = waiteReadDataPipeReg_needRead[13] & ~(waiteReadSate[13]) & waiteReadStageValid;
  assign readData_readDataQueue_13_deq_ready = isWaiteForThisData_13;
  assign isWaiteForThisData_14 = waiteReadDataPipeReg_needRead[14] & ~(waiteReadSate[14]) & waiteReadStageValid;
  assign readData_readDataQueue_14_deq_ready = isWaiteForThisData_14;
  assign isWaiteForThisData_15 = waiteReadDataPipeReg_needRead[15] & ~(waiteReadSate[15]) & waiteReadStageValid;
  assign readData_readDataQueue_15_deq_ready = isWaiteForThisData_15;
  assign isWaiteForThisData_16 = waiteReadDataPipeReg_needRead[16] & ~(waiteReadSate[16]) & waiteReadStageValid;
  assign readData_readDataQueue_16_deq_ready = isWaiteForThisData_16;
  assign isWaiteForThisData_17 = waiteReadDataPipeReg_needRead[17] & ~(waiteReadSate[17]) & waiteReadStageValid;
  assign readData_readDataQueue_17_deq_ready = isWaiteForThisData_17;
  assign isWaiteForThisData_18 = waiteReadDataPipeReg_needRead[18] & ~(waiteReadSate[18]) & waiteReadStageValid;
  assign readData_readDataQueue_18_deq_ready = isWaiteForThisData_18;
  assign isWaiteForThisData_19 = waiteReadDataPipeReg_needRead[19] & ~(waiteReadSate[19]) & waiteReadStageValid;
  assign readData_readDataQueue_19_deq_ready = isWaiteForThisData_19;
  assign isWaiteForThisData_20 = waiteReadDataPipeReg_needRead[20] & ~(waiteReadSate[20]) & waiteReadStageValid;
  assign readData_readDataQueue_20_deq_ready = isWaiteForThisData_20;
  assign isWaiteForThisData_21 = waiteReadDataPipeReg_needRead[21] & ~(waiteReadSate[21]) & waiteReadStageValid;
  assign readData_readDataQueue_21_deq_ready = isWaiteForThisData_21;
  assign isWaiteForThisData_22 = waiteReadDataPipeReg_needRead[22] & ~(waiteReadSate[22]) & waiteReadStageValid;
  assign readData_readDataQueue_22_deq_ready = isWaiteForThisData_22;
  assign isWaiteForThisData_23 = waiteReadDataPipeReg_needRead[23] & ~(waiteReadSate[23]) & waiteReadStageValid;
  assign readData_readDataQueue_23_deq_ready = isWaiteForThisData_23;
  assign isWaiteForThisData_24 = waiteReadDataPipeReg_needRead[24] & ~(waiteReadSate[24]) & waiteReadStageValid;
  assign readData_readDataQueue_24_deq_ready = isWaiteForThisData_24;
  assign isWaiteForThisData_25 = waiteReadDataPipeReg_needRead[25] & ~(waiteReadSate[25]) & waiteReadStageValid;
  assign readData_readDataQueue_25_deq_ready = isWaiteForThisData_25;
  assign isWaiteForThisData_26 = waiteReadDataPipeReg_needRead[26] & ~(waiteReadSate[26]) & waiteReadStageValid;
  assign readData_readDataQueue_26_deq_ready = isWaiteForThisData_26;
  assign isWaiteForThisData_27 = waiteReadDataPipeReg_needRead[27] & ~(waiteReadSate[27]) & waiteReadStageValid;
  assign readData_readDataQueue_27_deq_ready = isWaiteForThisData_27;
  assign isWaiteForThisData_28 = waiteReadDataPipeReg_needRead[28] & ~(waiteReadSate[28]) & waiteReadStageValid;
  assign readData_readDataQueue_28_deq_ready = isWaiteForThisData_28;
  assign isWaiteForThisData_29 = waiteReadDataPipeReg_needRead[29] & ~(waiteReadSate[29]) & waiteReadStageValid;
  assign readData_readDataQueue_29_deq_ready = isWaiteForThisData_29;
  assign isWaiteForThisData_30 = waiteReadDataPipeReg_needRead[30] & ~(waiteReadSate[30]) & waiteReadStageValid;
  assign readData_readDataQueue_30_deq_ready = isWaiteForThisData_30;
  assign isWaiteForThisData_31 = waiteReadDataPipeReg_needRead[31] & ~(waiteReadSate[31]) & waiteReadStageValid;
  assign readData_readDataQueue_31_deq_ready = isWaiteForThisData_31;
  wire [1:0]         readResultValid_lo_lo_lo_lo = {readTokenRelease_1, readTokenRelease_0};
  wire [1:0]         readResultValid_lo_lo_lo_hi = {readTokenRelease_3, readTokenRelease_2};
  wire [3:0]         readResultValid_lo_lo_lo = {readResultValid_lo_lo_lo_hi, readResultValid_lo_lo_lo_lo};
  wire [1:0]         readResultValid_lo_lo_hi_lo = {readTokenRelease_5, readTokenRelease_4};
  wire [1:0]         readResultValid_lo_lo_hi_hi = {readTokenRelease_7, readTokenRelease_6};
  wire [3:0]         readResultValid_lo_lo_hi = {readResultValid_lo_lo_hi_hi, readResultValid_lo_lo_hi_lo};
  wire [7:0]         readResultValid_lo_lo = {readResultValid_lo_lo_hi, readResultValid_lo_lo_lo};
  wire [1:0]         readResultValid_lo_hi_lo_lo = {readTokenRelease_9, readTokenRelease_8};
  wire [1:0]         readResultValid_lo_hi_lo_hi = {readTokenRelease_11, readTokenRelease_10};
  wire [3:0]         readResultValid_lo_hi_lo = {readResultValid_lo_hi_lo_hi, readResultValid_lo_hi_lo_lo};
  wire [1:0]         readResultValid_lo_hi_hi_lo = {readTokenRelease_13, readTokenRelease_12};
  wire [1:0]         readResultValid_lo_hi_hi_hi = {readTokenRelease_15, readTokenRelease_14};
  wire [3:0]         readResultValid_lo_hi_hi = {readResultValid_lo_hi_hi_hi, readResultValid_lo_hi_hi_lo};
  wire [7:0]         readResultValid_lo_hi = {readResultValid_lo_hi_hi, readResultValid_lo_hi_lo};
  wire [15:0]        readResultValid_lo = {readResultValid_lo_hi, readResultValid_lo_lo};
  wire [1:0]         readResultValid_hi_lo_lo_lo = {readTokenRelease_17, readTokenRelease_16};
  wire [1:0]         readResultValid_hi_lo_lo_hi = {readTokenRelease_19, readTokenRelease_18};
  wire [3:0]         readResultValid_hi_lo_lo = {readResultValid_hi_lo_lo_hi, readResultValid_hi_lo_lo_lo};
  wire [1:0]         readResultValid_hi_lo_hi_lo = {readTokenRelease_21, readTokenRelease_20};
  wire [1:0]         readResultValid_hi_lo_hi_hi = {readTokenRelease_23, readTokenRelease_22};
  wire [3:0]         readResultValid_hi_lo_hi = {readResultValid_hi_lo_hi_hi, readResultValid_hi_lo_hi_lo};
  wire [7:0]         readResultValid_hi_lo = {readResultValid_hi_lo_hi, readResultValid_hi_lo_lo};
  wire [1:0]         readResultValid_hi_hi_lo_lo = {readTokenRelease_25, readTokenRelease_24};
  wire [1:0]         readResultValid_hi_hi_lo_hi = {readTokenRelease_27, readTokenRelease_26};
  wire [3:0]         readResultValid_hi_hi_lo = {readResultValid_hi_hi_lo_hi, readResultValid_hi_hi_lo_lo};
  wire [1:0]         readResultValid_hi_hi_hi_lo = {readTokenRelease_29, readTokenRelease_28};
  wire [1:0]         readResultValid_hi_hi_hi_hi = {readTokenRelease_31, readTokenRelease_30};
  wire [3:0]         readResultValid_hi_hi_hi = {readResultValid_hi_hi_hi_hi, readResultValid_hi_hi_hi_lo};
  wire [7:0]         readResultValid_hi_hi = {readResultValid_hi_hi_hi, readResultValid_hi_hi_lo};
  wire [15:0]        readResultValid_hi = {readResultValid_hi_hi, readResultValid_hi_lo};
  wire [31:0]        readResultValid = {readResultValid_hi, readResultValid_lo};
  wire               executeEnqValid = otherTypeRequestDeq & ~readType;
  wire [63:0]        source2_lo_lo_lo_lo = {exeReqReg_1_bits_source2, exeReqReg_0_bits_source2};
  wire [63:0]        source2_lo_lo_lo_hi = {exeReqReg_3_bits_source2, exeReqReg_2_bits_source2};
  wire [127:0]       source2_lo_lo_lo = {source2_lo_lo_lo_hi, source2_lo_lo_lo_lo};
  wire [63:0]        source2_lo_lo_hi_lo = {exeReqReg_5_bits_source2, exeReqReg_4_bits_source2};
  wire [63:0]        source2_lo_lo_hi_hi = {exeReqReg_7_bits_source2, exeReqReg_6_bits_source2};
  wire [127:0]       source2_lo_lo_hi = {source2_lo_lo_hi_hi, source2_lo_lo_hi_lo};
  wire [255:0]       source2_lo_lo = {source2_lo_lo_hi, source2_lo_lo_lo};
  wire [63:0]        source2_lo_hi_lo_lo = {exeReqReg_9_bits_source2, exeReqReg_8_bits_source2};
  wire [63:0]        source2_lo_hi_lo_hi = {exeReqReg_11_bits_source2, exeReqReg_10_bits_source2};
  wire [127:0]       source2_lo_hi_lo = {source2_lo_hi_lo_hi, source2_lo_hi_lo_lo};
  wire [63:0]        source2_lo_hi_hi_lo = {exeReqReg_13_bits_source2, exeReqReg_12_bits_source2};
  wire [63:0]        source2_lo_hi_hi_hi = {exeReqReg_15_bits_source2, exeReqReg_14_bits_source2};
  wire [127:0]       source2_lo_hi_hi = {source2_lo_hi_hi_hi, source2_lo_hi_hi_lo};
  wire [255:0]       source2_lo_hi = {source2_lo_hi_hi, source2_lo_hi_lo};
  wire [511:0]       source2_lo = {source2_lo_hi, source2_lo_lo};
  wire [63:0]        source2_hi_lo_lo_lo = {exeReqReg_17_bits_source2, exeReqReg_16_bits_source2};
  wire [63:0]        source2_hi_lo_lo_hi = {exeReqReg_19_bits_source2, exeReqReg_18_bits_source2};
  wire [127:0]       source2_hi_lo_lo = {source2_hi_lo_lo_hi, source2_hi_lo_lo_lo};
  wire [63:0]        source2_hi_lo_hi_lo = {exeReqReg_21_bits_source2, exeReqReg_20_bits_source2};
  wire [63:0]        source2_hi_lo_hi_hi = {exeReqReg_23_bits_source2, exeReqReg_22_bits_source2};
  wire [127:0]       source2_hi_lo_hi = {source2_hi_lo_hi_hi, source2_hi_lo_hi_lo};
  wire [255:0]       source2_hi_lo = {source2_hi_lo_hi, source2_hi_lo_lo};
  wire [63:0]        source2_hi_hi_lo_lo = {exeReqReg_25_bits_source2, exeReqReg_24_bits_source2};
  wire [63:0]        source2_hi_hi_lo_hi = {exeReqReg_27_bits_source2, exeReqReg_26_bits_source2};
  wire [127:0]       source2_hi_hi_lo = {source2_hi_hi_lo_hi, source2_hi_hi_lo_lo};
  wire [63:0]        source2_hi_hi_hi_lo = {exeReqReg_29_bits_source2, exeReqReg_28_bits_source2};
  wire [63:0]        source2_hi_hi_hi_hi = {exeReqReg_31_bits_source2, exeReqReg_30_bits_source2};
  wire [127:0]       source2_hi_hi_hi = {source2_hi_hi_hi_hi, source2_hi_hi_hi_lo};
  wire [255:0]       source2_hi_hi = {source2_hi_hi_hi, source2_hi_hi_lo};
  wire [511:0]       source2_hi = {source2_hi_hi, source2_hi_lo};
  wire [1023:0]      source2 = {source2_hi, source2_lo};
  wire [127:0]       source1_lo_lo_lo = {source1_lo_lo_lo_hi, source1_lo_lo_lo_lo};
  wire [127:0]       source1_lo_lo_hi = {source1_lo_lo_hi_hi, source1_lo_lo_hi_lo};
  wire [255:0]       source1_lo_lo = {source1_lo_lo_hi, source1_lo_lo_lo};
  wire [127:0]       source1_lo_hi_lo = {source1_lo_hi_lo_hi, source1_lo_hi_lo_lo};
  wire [127:0]       source1_lo_hi_hi = {source1_lo_hi_hi_hi, source1_lo_hi_hi_lo};
  wire [255:0]       source1_lo_hi = {source1_lo_hi_hi, source1_lo_hi_lo};
  wire [511:0]       source1_lo = {source1_lo_hi, source1_lo_lo};
  wire [127:0]       source1_hi_lo_lo = {source1_hi_lo_lo_hi, source1_hi_lo_lo_lo};
  wire [127:0]       source1_hi_lo_hi = {source1_hi_lo_hi_hi, source1_hi_lo_hi_lo};
  wire [255:0]       source1_hi_lo = {source1_hi_lo_hi, source1_hi_lo_lo};
  wire [127:0]       source1_hi_hi_lo = {source1_hi_hi_lo_hi, source1_hi_hi_lo_lo};
  wire [127:0]       source1_hi_hi_hi = {source1_hi_hi_hi_hi, source1_hi_hi_hi_lo};
  wire [255:0]       source1_hi_hi = {source1_hi_hi_hi, source1_hi_hi_lo};
  wire [511:0]       source1_hi = {source1_hi_hi, source1_hi_lo};
  wire [1023:0]      source1 = {source1_hi, source1_lo};
  wire [31:0]        compressSource1 = (|sew1H) ? readVS1Reg_data : 32'h0;
  wire [31:0]        source1Select = mv ? readVS1Reg_data : compressSource1;
  wire               source1Change = |sew1H;
  assign viotaCounterAdd = executeEnqValid & unitType[1];
  wire [1:0]         view__in_bits_ffoInput_lo_lo_lo_lo = {exeReqReg_1_bits_ffo, exeReqReg_0_bits_ffo};
  wire [1:0]         view__in_bits_ffoInput_lo_lo_lo_hi = {exeReqReg_3_bits_ffo, exeReqReg_2_bits_ffo};
  wire [3:0]         view__in_bits_ffoInput_lo_lo_lo = {view__in_bits_ffoInput_lo_lo_lo_hi, view__in_bits_ffoInput_lo_lo_lo_lo};
  wire [1:0]         view__in_bits_ffoInput_lo_lo_hi_lo = {exeReqReg_5_bits_ffo, exeReqReg_4_bits_ffo};
  wire [1:0]         view__in_bits_ffoInput_lo_lo_hi_hi = {exeReqReg_7_bits_ffo, exeReqReg_6_bits_ffo};
  wire [3:0]         view__in_bits_ffoInput_lo_lo_hi = {view__in_bits_ffoInput_lo_lo_hi_hi, view__in_bits_ffoInput_lo_lo_hi_lo};
  wire [7:0]         view__in_bits_ffoInput_lo_lo = {view__in_bits_ffoInput_lo_lo_hi, view__in_bits_ffoInput_lo_lo_lo};
  wire [1:0]         view__in_bits_ffoInput_lo_hi_lo_lo = {exeReqReg_9_bits_ffo, exeReqReg_8_bits_ffo};
  wire [1:0]         view__in_bits_ffoInput_lo_hi_lo_hi = {exeReqReg_11_bits_ffo, exeReqReg_10_bits_ffo};
  wire [3:0]         view__in_bits_ffoInput_lo_hi_lo = {view__in_bits_ffoInput_lo_hi_lo_hi, view__in_bits_ffoInput_lo_hi_lo_lo};
  wire [1:0]         view__in_bits_ffoInput_lo_hi_hi_lo = {exeReqReg_13_bits_ffo, exeReqReg_12_bits_ffo};
  wire [1:0]         view__in_bits_ffoInput_lo_hi_hi_hi = {exeReqReg_15_bits_ffo, exeReqReg_14_bits_ffo};
  wire [3:0]         view__in_bits_ffoInput_lo_hi_hi = {view__in_bits_ffoInput_lo_hi_hi_hi, view__in_bits_ffoInput_lo_hi_hi_lo};
  wire [7:0]         view__in_bits_ffoInput_lo_hi = {view__in_bits_ffoInput_lo_hi_hi, view__in_bits_ffoInput_lo_hi_lo};
  wire [15:0]        view__in_bits_ffoInput_lo = {view__in_bits_ffoInput_lo_hi, view__in_bits_ffoInput_lo_lo};
  wire [1:0]         view__in_bits_ffoInput_hi_lo_lo_lo = {exeReqReg_17_bits_ffo, exeReqReg_16_bits_ffo};
  wire [1:0]         view__in_bits_ffoInput_hi_lo_lo_hi = {exeReqReg_19_bits_ffo, exeReqReg_18_bits_ffo};
  wire [3:0]         view__in_bits_ffoInput_hi_lo_lo = {view__in_bits_ffoInput_hi_lo_lo_hi, view__in_bits_ffoInput_hi_lo_lo_lo};
  wire [1:0]         view__in_bits_ffoInput_hi_lo_hi_lo = {exeReqReg_21_bits_ffo, exeReqReg_20_bits_ffo};
  wire [1:0]         view__in_bits_ffoInput_hi_lo_hi_hi = {exeReqReg_23_bits_ffo, exeReqReg_22_bits_ffo};
  wire [3:0]         view__in_bits_ffoInput_hi_lo_hi = {view__in_bits_ffoInput_hi_lo_hi_hi, view__in_bits_ffoInput_hi_lo_hi_lo};
  wire [7:0]         view__in_bits_ffoInput_hi_lo = {view__in_bits_ffoInput_hi_lo_hi, view__in_bits_ffoInput_hi_lo_lo};
  wire [1:0]         view__in_bits_ffoInput_hi_hi_lo_lo = {exeReqReg_25_bits_ffo, exeReqReg_24_bits_ffo};
  wire [1:0]         view__in_bits_ffoInput_hi_hi_lo_hi = {exeReqReg_27_bits_ffo, exeReqReg_26_bits_ffo};
  wire [3:0]         view__in_bits_ffoInput_hi_hi_lo = {view__in_bits_ffoInput_hi_hi_lo_hi, view__in_bits_ffoInput_hi_hi_lo_lo};
  wire [1:0]         view__in_bits_ffoInput_hi_hi_hi_lo = {exeReqReg_29_bits_ffo, exeReqReg_28_bits_ffo};
  wire [1:0]         view__in_bits_ffoInput_hi_hi_hi_hi = {exeReqReg_31_bits_ffo, exeReqReg_30_bits_ffo};
  wire [3:0]         view__in_bits_ffoInput_hi_hi_hi = {view__in_bits_ffoInput_hi_hi_hi_hi, view__in_bits_ffoInput_hi_hi_hi_lo};
  wire [7:0]         view__in_bits_ffoInput_hi_hi = {view__in_bits_ffoInput_hi_hi_hi, view__in_bits_ffoInput_hi_hi_lo};
  wire [15:0]        view__in_bits_ffoInput_hi = {view__in_bits_ffoInput_hi_hi, view__in_bits_ffoInput_hi_lo};
  wire [3:0]         view__in_bits_validInput_lo_lo_lo = {view__in_bits_validInput_lo_lo_lo_hi, view__in_bits_validInput_lo_lo_lo_lo};
  wire [3:0]         view__in_bits_validInput_lo_lo_hi = {view__in_bits_validInput_lo_lo_hi_hi, view__in_bits_validInput_lo_lo_hi_lo};
  wire [7:0]         view__in_bits_validInput_lo_lo = {view__in_bits_validInput_lo_lo_hi, view__in_bits_validInput_lo_lo_lo};
  wire [3:0]         view__in_bits_validInput_lo_hi_lo = {view__in_bits_validInput_lo_hi_lo_hi, view__in_bits_validInput_lo_hi_lo_lo};
  wire [3:0]         view__in_bits_validInput_lo_hi_hi = {view__in_bits_validInput_lo_hi_hi_hi, view__in_bits_validInput_lo_hi_hi_lo};
  wire [7:0]         view__in_bits_validInput_lo_hi = {view__in_bits_validInput_lo_hi_hi, view__in_bits_validInput_lo_hi_lo};
  wire [15:0]        view__in_bits_validInput_lo = {view__in_bits_validInput_lo_hi, view__in_bits_validInput_lo_lo};
  wire [3:0]         view__in_bits_validInput_hi_lo_lo = {view__in_bits_validInput_hi_lo_lo_hi, view__in_bits_validInput_hi_lo_lo_lo};
  wire [3:0]         view__in_bits_validInput_hi_lo_hi = {view__in_bits_validInput_hi_lo_hi_hi, view__in_bits_validInput_hi_lo_hi_lo};
  wire [7:0]         view__in_bits_validInput_hi_lo = {view__in_bits_validInput_hi_lo_hi, view__in_bits_validInput_hi_lo_lo};
  wire [3:0]         view__in_bits_validInput_hi_hi_lo = {view__in_bits_validInput_hi_hi_lo_hi, view__in_bits_validInput_hi_hi_lo_lo};
  wire [3:0]         view__in_bits_validInput_hi_hi_hi = {view__in_bits_validInput_hi_hi_hi_hi, view__in_bits_validInput_hi_hi_hi_lo};
  wire [7:0]         view__in_bits_validInput_hi_hi = {view__in_bits_validInput_hi_hi_hi, view__in_bits_validInput_hi_hi_lo};
  wire [15:0]        view__in_bits_validInput_hi = {view__in_bits_validInput_hi_hi, view__in_bits_validInput_hi_lo};
  wire               reduceUnit_in_valid = executeEnqValid & unitType[2];
  wire [3:0]         view__in_bits_sourceValid_lo_lo_lo = {view__in_bits_sourceValid_lo_lo_lo_hi, view__in_bits_sourceValid_lo_lo_lo_lo};
  wire [3:0]         view__in_bits_sourceValid_lo_lo_hi = {view__in_bits_sourceValid_lo_lo_hi_hi, view__in_bits_sourceValid_lo_lo_hi_lo};
  wire [7:0]         view__in_bits_sourceValid_lo_lo = {view__in_bits_sourceValid_lo_lo_hi, view__in_bits_sourceValid_lo_lo_lo};
  wire [3:0]         view__in_bits_sourceValid_lo_hi_lo = {view__in_bits_sourceValid_lo_hi_lo_hi, view__in_bits_sourceValid_lo_hi_lo_lo};
  wire [3:0]         view__in_bits_sourceValid_lo_hi_hi = {view__in_bits_sourceValid_lo_hi_hi_hi, view__in_bits_sourceValid_lo_hi_hi_lo};
  wire [7:0]         view__in_bits_sourceValid_lo_hi = {view__in_bits_sourceValid_lo_hi_hi, view__in_bits_sourceValid_lo_hi_lo};
  wire [15:0]        view__in_bits_sourceValid_lo = {view__in_bits_sourceValid_lo_hi, view__in_bits_sourceValid_lo_lo};
  wire [3:0]         view__in_bits_sourceValid_hi_lo_lo = {view__in_bits_sourceValid_hi_lo_lo_hi, view__in_bits_sourceValid_hi_lo_lo_lo};
  wire [3:0]         view__in_bits_sourceValid_hi_lo_hi = {view__in_bits_sourceValid_hi_lo_hi_hi, view__in_bits_sourceValid_hi_lo_hi_lo};
  wire [7:0]         view__in_bits_sourceValid_hi_lo = {view__in_bits_sourceValid_hi_lo_hi, view__in_bits_sourceValid_hi_lo_lo};
  wire [3:0]         view__in_bits_sourceValid_hi_hi_lo = {view__in_bits_sourceValid_hi_hi_lo_hi, view__in_bits_sourceValid_hi_hi_lo_lo};
  wire [3:0]         view__in_bits_sourceValid_hi_hi_hi = {view__in_bits_sourceValid_hi_hi_hi_hi, view__in_bits_sourceValid_hi_hi_hi_lo};
  wire [7:0]         view__in_bits_sourceValid_hi_hi = {view__in_bits_sourceValid_hi_hi_hi, view__in_bits_sourceValid_hi_hi_lo};
  wire [15:0]        view__in_bits_sourceValid_hi = {view__in_bits_sourceValid_hi_hi, view__in_bits_sourceValid_hi_lo};
  wire               _view__firstGroup_T_1 = _reduceUnit_in_ready & reduceUnit_in_valid;
  wire [6:0]         extendGroupCount = extendType ? (subType[2] ? _extendGroupCount_T_1 : {1'h0, requestCounter, executeIndex[1]}) : {2'h0, requestCounter};
  wire [1023:0]      _executeResult_T_4 = unitType[1] ? compressUnitResultQueue_deq_bits_data : 1024'h0;
  wire [1023:0]      executeResult = {_executeResult_T_4[1023:32], _executeResult_T_4[31:0] | (unitType[2] ? _reduceUnit_out_bits_data : 32'h0)} | (unitType[3] ? _extendUnit_out : 1024'h0);
  assign executeReady = readType | unitType[1] | unitType[2] & _reduceUnit_in_ready & readVS1Reg_dataValid | unitType[3] & executeEnqValid;
  wire [3:0]         compressUnitResultQueue_deq_ready_lo_lo_lo = {compressUnitResultQueue_deq_ready_lo_lo_lo_hi, compressUnitResultQueue_deq_ready_lo_lo_lo_lo};
  wire [3:0]         compressUnitResultQueue_deq_ready_lo_lo_hi = {compressUnitResultQueue_deq_ready_lo_lo_hi_hi, compressUnitResultQueue_deq_ready_lo_lo_hi_lo};
  wire [7:0]         compressUnitResultQueue_deq_ready_lo_lo = {compressUnitResultQueue_deq_ready_lo_lo_hi, compressUnitResultQueue_deq_ready_lo_lo_lo};
  wire [3:0]         compressUnitResultQueue_deq_ready_lo_hi_lo = {compressUnitResultQueue_deq_ready_lo_hi_lo_hi, compressUnitResultQueue_deq_ready_lo_hi_lo_lo};
  wire [3:0]         compressUnitResultQueue_deq_ready_lo_hi_hi = {compressUnitResultQueue_deq_ready_lo_hi_hi_hi, compressUnitResultQueue_deq_ready_lo_hi_hi_lo};
  wire [7:0]         compressUnitResultQueue_deq_ready_lo_hi = {compressUnitResultQueue_deq_ready_lo_hi_hi, compressUnitResultQueue_deq_ready_lo_hi_lo};
  wire [15:0]        compressUnitResultQueue_deq_ready_lo = {compressUnitResultQueue_deq_ready_lo_hi, compressUnitResultQueue_deq_ready_lo_lo};
  wire [3:0]         compressUnitResultQueue_deq_ready_hi_lo_lo = {compressUnitResultQueue_deq_ready_hi_lo_lo_hi, compressUnitResultQueue_deq_ready_hi_lo_lo_lo};
  wire [3:0]         compressUnitResultQueue_deq_ready_hi_lo_hi = {compressUnitResultQueue_deq_ready_hi_lo_hi_hi, compressUnitResultQueue_deq_ready_hi_lo_hi_lo};
  wire [7:0]         compressUnitResultQueue_deq_ready_hi_lo = {compressUnitResultQueue_deq_ready_hi_lo_hi, compressUnitResultQueue_deq_ready_hi_lo_lo};
  wire [3:0]         compressUnitResultQueue_deq_ready_hi_hi_lo = {compressUnitResultQueue_deq_ready_hi_hi_lo_hi, compressUnitResultQueue_deq_ready_hi_hi_lo_lo};
  wire [3:0]         compressUnitResultQueue_deq_ready_hi_hi_hi = {compressUnitResultQueue_deq_ready_hi_hi_hi_hi, compressUnitResultQueue_deq_ready_hi_hi_hi_lo};
  wire [7:0]         compressUnitResultQueue_deq_ready_hi_hi = {compressUnitResultQueue_deq_ready_hi_hi_hi, compressUnitResultQueue_deq_ready_hi_hi_lo};
  wire [15:0]        compressUnitResultQueue_deq_ready_hi = {compressUnitResultQueue_deq_ready_hi_hi, compressUnitResultQueue_deq_ready_hi_lo};
  assign compressUnitResultQueue_deq_ready = &{compressUnitResultQueue_deq_ready_hi, compressUnitResultQueue_deq_ready_lo};
  wire               compressDeq = compressUnitResultQueue_deq_ready & compressUnitResultQueue_deq_valid;
  wire               executeValid = unitType[1] & compressDeq | unitType[3] & executeEnqValid;
  assign executeGroupCounter = (unitType[1] | unitType[2] ? requestCounter : 5'h0) | (unitType[3] ? extendGroupCount[4:0] : 5'h0);
  wire [6:0]         executeDeqGroupCounter = {2'h0, (unitType[1] ? compressUnitResultQueue_deq_bits_groupCounter : 5'h0) | (unitType[2] ? requestCounter : 5'h0)} | (unitType[3] ? extendGroupCount : 7'h0);
  wire [127:0]       executeWriteByteMask = compress | ffo | mvVd ? compressUnitResultQueue_deq_bits_mask : executeByteMask;
  wire               maskFilter = |{~maskDestinationType, currentMaskGroupForDestination[31:0]};
  wire               maskFilter_1 = |{~maskDestinationType, currentMaskGroupForDestination[63:32]};
  wire               maskFilter_2 = |{~maskDestinationType, currentMaskGroupForDestination[95:64]};
  wire               maskFilter_3 = |{~maskDestinationType, currentMaskGroupForDestination[127:96]};
  wire               maskFilter_4 = |{~maskDestinationType, currentMaskGroupForDestination[159:128]};
  wire               maskFilter_5 = |{~maskDestinationType, currentMaskGroupForDestination[191:160]};
  wire               maskFilter_6 = |{~maskDestinationType, currentMaskGroupForDestination[223:192]};
  wire               maskFilter_7 = |{~maskDestinationType, currentMaskGroupForDestination[255:224]};
  wire               maskFilter_8 = |{~maskDestinationType, currentMaskGroupForDestination[287:256]};
  wire               maskFilter_9 = |{~maskDestinationType, currentMaskGroupForDestination[319:288]};
  wire               maskFilter_10 = |{~maskDestinationType, currentMaskGroupForDestination[351:320]};
  wire               maskFilter_11 = |{~maskDestinationType, currentMaskGroupForDestination[383:352]};
  wire               maskFilter_12 = |{~maskDestinationType, currentMaskGroupForDestination[415:384]};
  wire               maskFilter_13 = |{~maskDestinationType, currentMaskGroupForDestination[447:416]};
  wire               maskFilter_14 = |{~maskDestinationType, currentMaskGroupForDestination[479:448]};
  wire               maskFilter_15 = |{~maskDestinationType, currentMaskGroupForDestination[511:480]};
  wire               maskFilter_16 = |{~maskDestinationType, currentMaskGroupForDestination[543:512]};
  wire               maskFilter_17 = |{~maskDestinationType, currentMaskGroupForDestination[575:544]};
  wire               maskFilter_18 = |{~maskDestinationType, currentMaskGroupForDestination[607:576]};
  wire               maskFilter_19 = |{~maskDestinationType, currentMaskGroupForDestination[639:608]};
  wire               maskFilter_20 = |{~maskDestinationType, currentMaskGroupForDestination[671:640]};
  wire               maskFilter_21 = |{~maskDestinationType, currentMaskGroupForDestination[703:672]};
  wire               maskFilter_22 = |{~maskDestinationType, currentMaskGroupForDestination[735:704]};
  wire               maskFilter_23 = |{~maskDestinationType, currentMaskGroupForDestination[767:736]};
  wire               maskFilter_24 = |{~maskDestinationType, currentMaskGroupForDestination[799:768]};
  wire               maskFilter_25 = |{~maskDestinationType, currentMaskGroupForDestination[831:800]};
  wire               maskFilter_26 = |{~maskDestinationType, currentMaskGroupForDestination[863:832]};
  wire               maskFilter_27 = |{~maskDestinationType, currentMaskGroupForDestination[895:864]};
  wire               maskFilter_28 = |{~maskDestinationType, currentMaskGroupForDestination[927:896]};
  wire               maskFilter_29 = |{~maskDestinationType, currentMaskGroupForDestination[959:928]};
  wire               maskFilter_30 = |{~maskDestinationType, currentMaskGroupForDestination[991:960]};
  wire               maskFilter_31 = |{~maskDestinationType, currentMaskGroupForDestination[1023:992]};
  assign writeQueue_0_deq_valid = ~_writeQueue_fifo_empty;
  wire               exeResp_0_valid_0 = writeQueue_0_deq_valid;
  wire               writeQueue_dataOut_ffoByOther;
  wire [31:0]        writeQueue_dataOut_writeData_data;
  wire [31:0]        exeResp_0_bits_data_0 = writeQueue_0_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_writeData_mask;
  wire [3:0]         exeResp_0_bits_mask_0 = writeQueue_0_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_writeData_vd;
  wire [2:0]         writeQueue_dataOut_index;
  wire [4:0]         writeQueue_0_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_0_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo = {writeQueue_0_enq_bits_writeData_groupCounter, writeQueue_0_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_0_enq_bits_writeData_data;
  wire [3:0]         writeQueue_0_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi = {writeQueue_0_enq_bits_writeData_data, writeQueue_0_enq_bits_writeData_mask};
  wire               writeQueue_0_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_1 = {writeQueue_0_enq_bits_ffoByOther, writeQueue_dataIn_hi, writeQueue_dataIn_lo};
  wire [49:0]        writeQueue_dataIn = {writeQueue_dataIn_hi_1, writeQueue_0_enq_bits_index};
  assign writeQueue_dataOut_index = _writeQueue_fifo_data_out[2:0];
  assign writeQueue_dataOut_writeData_vd = _writeQueue_fifo_data_out[7:3];
  assign writeQueue_dataOut_writeData_groupCounter = _writeQueue_fifo_data_out[12:8];
  assign writeQueue_dataOut_writeData_mask = _writeQueue_fifo_data_out[16:13];
  assign writeQueue_dataOut_writeData_data = _writeQueue_fifo_data_out[48:17];
  assign writeQueue_dataOut_ffoByOther = _writeQueue_fifo_data_out[49];
  wire               writeQueue_0_deq_bits_ffoByOther = writeQueue_dataOut_ffoByOther;
  assign writeQueue_0_deq_bits_writeData_data = writeQueue_dataOut_writeData_data;
  assign writeQueue_0_deq_bits_writeData_mask = writeQueue_dataOut_writeData_mask;
  wire [4:0]         writeQueue_0_deq_bits_writeData_groupCounter = writeQueue_dataOut_writeData_groupCounter;
  wire [4:0]         writeQueue_0_deq_bits_writeData_vd = writeQueue_dataOut_writeData_vd;
  wire [2:0]         writeQueue_0_deq_bits_index = writeQueue_dataOut_index;
  wire               writeQueue_0_enq_ready = ~_writeQueue_fifo_full;
  wire               writeQueue_0_enq_valid;
  assign writeQueue_1_deq_valid = ~_writeQueue_fifo_1_empty;
  wire               exeResp_1_valid_0 = writeQueue_1_deq_valid;
  wire               writeQueue_dataOut_1_ffoByOther;
  wire [31:0]        writeQueue_dataOut_1_writeData_data;
  wire [31:0]        exeResp_1_bits_data_0 = writeQueue_1_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_1_writeData_mask;
  wire [3:0]         exeResp_1_bits_mask_0 = writeQueue_1_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_1_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_1_writeData_vd;
  wire [2:0]         writeQueue_dataOut_1_index;
  wire [4:0]         writeQueue_1_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_1_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_1 = {writeQueue_1_enq_bits_writeData_groupCounter, writeQueue_1_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_1_enq_bits_writeData_data;
  wire [3:0]         writeQueue_1_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_2 = {writeQueue_1_enq_bits_writeData_data, writeQueue_1_enq_bits_writeData_mask};
  wire               writeQueue_1_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_3 = {writeQueue_1_enq_bits_ffoByOther, writeQueue_dataIn_hi_2, writeQueue_dataIn_lo_1};
  wire [49:0]        writeQueue_dataIn_1 = {writeQueue_dataIn_hi_3, writeQueue_1_enq_bits_index};
  assign writeQueue_dataOut_1_index = _writeQueue_fifo_1_data_out[2:0];
  assign writeQueue_dataOut_1_writeData_vd = _writeQueue_fifo_1_data_out[7:3];
  assign writeQueue_dataOut_1_writeData_groupCounter = _writeQueue_fifo_1_data_out[12:8];
  assign writeQueue_dataOut_1_writeData_mask = _writeQueue_fifo_1_data_out[16:13];
  assign writeQueue_dataOut_1_writeData_data = _writeQueue_fifo_1_data_out[48:17];
  assign writeQueue_dataOut_1_ffoByOther = _writeQueue_fifo_1_data_out[49];
  wire               writeQueue_1_deq_bits_ffoByOther = writeQueue_dataOut_1_ffoByOther;
  assign writeQueue_1_deq_bits_writeData_data = writeQueue_dataOut_1_writeData_data;
  assign writeQueue_1_deq_bits_writeData_mask = writeQueue_dataOut_1_writeData_mask;
  wire [4:0]         writeQueue_1_deq_bits_writeData_groupCounter = writeQueue_dataOut_1_writeData_groupCounter;
  wire [4:0]         writeQueue_1_deq_bits_writeData_vd = writeQueue_dataOut_1_writeData_vd;
  wire [2:0]         writeQueue_1_deq_bits_index = writeQueue_dataOut_1_index;
  wire               writeQueue_1_enq_ready = ~_writeQueue_fifo_1_full;
  wire               writeQueue_1_enq_valid;
  assign writeQueue_2_deq_valid = ~_writeQueue_fifo_2_empty;
  wire               exeResp_2_valid_0 = writeQueue_2_deq_valid;
  wire               writeQueue_dataOut_2_ffoByOther;
  wire [31:0]        writeQueue_dataOut_2_writeData_data;
  wire [31:0]        exeResp_2_bits_data_0 = writeQueue_2_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_2_writeData_mask;
  wire [3:0]         exeResp_2_bits_mask_0 = writeQueue_2_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_2_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_2_writeData_vd;
  wire [2:0]         writeQueue_dataOut_2_index;
  wire [4:0]         writeQueue_2_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_2_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_2 = {writeQueue_2_enq_bits_writeData_groupCounter, writeQueue_2_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_2_enq_bits_writeData_data;
  wire [3:0]         writeQueue_2_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_4 = {writeQueue_2_enq_bits_writeData_data, writeQueue_2_enq_bits_writeData_mask};
  wire               writeQueue_2_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_5 = {writeQueue_2_enq_bits_ffoByOther, writeQueue_dataIn_hi_4, writeQueue_dataIn_lo_2};
  wire [49:0]        writeQueue_dataIn_2 = {writeQueue_dataIn_hi_5, writeQueue_2_enq_bits_index};
  assign writeQueue_dataOut_2_index = _writeQueue_fifo_2_data_out[2:0];
  assign writeQueue_dataOut_2_writeData_vd = _writeQueue_fifo_2_data_out[7:3];
  assign writeQueue_dataOut_2_writeData_groupCounter = _writeQueue_fifo_2_data_out[12:8];
  assign writeQueue_dataOut_2_writeData_mask = _writeQueue_fifo_2_data_out[16:13];
  assign writeQueue_dataOut_2_writeData_data = _writeQueue_fifo_2_data_out[48:17];
  assign writeQueue_dataOut_2_ffoByOther = _writeQueue_fifo_2_data_out[49];
  wire               writeQueue_2_deq_bits_ffoByOther = writeQueue_dataOut_2_ffoByOther;
  assign writeQueue_2_deq_bits_writeData_data = writeQueue_dataOut_2_writeData_data;
  assign writeQueue_2_deq_bits_writeData_mask = writeQueue_dataOut_2_writeData_mask;
  wire [4:0]         writeQueue_2_deq_bits_writeData_groupCounter = writeQueue_dataOut_2_writeData_groupCounter;
  wire [4:0]         writeQueue_2_deq_bits_writeData_vd = writeQueue_dataOut_2_writeData_vd;
  wire [2:0]         writeQueue_2_deq_bits_index = writeQueue_dataOut_2_index;
  wire               writeQueue_2_enq_ready = ~_writeQueue_fifo_2_full;
  wire               writeQueue_2_enq_valid;
  assign writeQueue_3_deq_valid = ~_writeQueue_fifo_3_empty;
  wire               exeResp_3_valid_0 = writeQueue_3_deq_valid;
  wire               writeQueue_dataOut_3_ffoByOther;
  wire [31:0]        writeQueue_dataOut_3_writeData_data;
  wire [31:0]        exeResp_3_bits_data_0 = writeQueue_3_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_3_writeData_mask;
  wire [3:0]         exeResp_3_bits_mask_0 = writeQueue_3_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_3_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_3_writeData_vd;
  wire [2:0]         writeQueue_dataOut_3_index;
  wire [4:0]         writeQueue_3_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_3_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_3 = {writeQueue_3_enq_bits_writeData_groupCounter, writeQueue_3_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_3_enq_bits_writeData_data;
  wire [3:0]         writeQueue_3_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_6 = {writeQueue_3_enq_bits_writeData_data, writeQueue_3_enq_bits_writeData_mask};
  wire               writeQueue_3_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_7 = {writeQueue_3_enq_bits_ffoByOther, writeQueue_dataIn_hi_6, writeQueue_dataIn_lo_3};
  wire [49:0]        writeQueue_dataIn_3 = {writeQueue_dataIn_hi_7, writeQueue_3_enq_bits_index};
  assign writeQueue_dataOut_3_index = _writeQueue_fifo_3_data_out[2:0];
  assign writeQueue_dataOut_3_writeData_vd = _writeQueue_fifo_3_data_out[7:3];
  assign writeQueue_dataOut_3_writeData_groupCounter = _writeQueue_fifo_3_data_out[12:8];
  assign writeQueue_dataOut_3_writeData_mask = _writeQueue_fifo_3_data_out[16:13];
  assign writeQueue_dataOut_3_writeData_data = _writeQueue_fifo_3_data_out[48:17];
  assign writeQueue_dataOut_3_ffoByOther = _writeQueue_fifo_3_data_out[49];
  wire               writeQueue_3_deq_bits_ffoByOther = writeQueue_dataOut_3_ffoByOther;
  assign writeQueue_3_deq_bits_writeData_data = writeQueue_dataOut_3_writeData_data;
  assign writeQueue_3_deq_bits_writeData_mask = writeQueue_dataOut_3_writeData_mask;
  wire [4:0]         writeQueue_3_deq_bits_writeData_groupCounter = writeQueue_dataOut_3_writeData_groupCounter;
  wire [4:0]         writeQueue_3_deq_bits_writeData_vd = writeQueue_dataOut_3_writeData_vd;
  wire [2:0]         writeQueue_3_deq_bits_index = writeQueue_dataOut_3_index;
  wire               writeQueue_3_enq_ready = ~_writeQueue_fifo_3_full;
  wire               writeQueue_3_enq_valid;
  assign writeQueue_4_deq_valid = ~_writeQueue_fifo_4_empty;
  wire               exeResp_4_valid_0 = writeQueue_4_deq_valid;
  wire               writeQueue_dataOut_4_ffoByOther;
  wire [31:0]        writeQueue_dataOut_4_writeData_data;
  wire [31:0]        exeResp_4_bits_data_0 = writeQueue_4_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_4_writeData_mask;
  wire [3:0]         exeResp_4_bits_mask_0 = writeQueue_4_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_4_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_4_writeData_vd;
  wire [2:0]         writeQueue_dataOut_4_index;
  wire [4:0]         writeQueue_4_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_4_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_4 = {writeQueue_4_enq_bits_writeData_groupCounter, writeQueue_4_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_4_enq_bits_writeData_data;
  wire [3:0]         writeQueue_4_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_8 = {writeQueue_4_enq_bits_writeData_data, writeQueue_4_enq_bits_writeData_mask};
  wire               writeQueue_4_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_9 = {writeQueue_4_enq_bits_ffoByOther, writeQueue_dataIn_hi_8, writeQueue_dataIn_lo_4};
  wire [49:0]        writeQueue_dataIn_4 = {writeQueue_dataIn_hi_9, writeQueue_4_enq_bits_index};
  assign writeQueue_dataOut_4_index = _writeQueue_fifo_4_data_out[2:0];
  assign writeQueue_dataOut_4_writeData_vd = _writeQueue_fifo_4_data_out[7:3];
  assign writeQueue_dataOut_4_writeData_groupCounter = _writeQueue_fifo_4_data_out[12:8];
  assign writeQueue_dataOut_4_writeData_mask = _writeQueue_fifo_4_data_out[16:13];
  assign writeQueue_dataOut_4_writeData_data = _writeQueue_fifo_4_data_out[48:17];
  assign writeQueue_dataOut_4_ffoByOther = _writeQueue_fifo_4_data_out[49];
  wire               writeQueue_4_deq_bits_ffoByOther = writeQueue_dataOut_4_ffoByOther;
  assign writeQueue_4_deq_bits_writeData_data = writeQueue_dataOut_4_writeData_data;
  assign writeQueue_4_deq_bits_writeData_mask = writeQueue_dataOut_4_writeData_mask;
  wire [4:0]         writeQueue_4_deq_bits_writeData_groupCounter = writeQueue_dataOut_4_writeData_groupCounter;
  wire [4:0]         writeQueue_4_deq_bits_writeData_vd = writeQueue_dataOut_4_writeData_vd;
  wire [2:0]         writeQueue_4_deq_bits_index = writeQueue_dataOut_4_index;
  wire               writeQueue_4_enq_ready = ~_writeQueue_fifo_4_full;
  wire               writeQueue_4_enq_valid;
  assign writeQueue_5_deq_valid = ~_writeQueue_fifo_5_empty;
  wire               exeResp_5_valid_0 = writeQueue_5_deq_valid;
  wire               writeQueue_dataOut_5_ffoByOther;
  wire [31:0]        writeQueue_dataOut_5_writeData_data;
  wire [31:0]        exeResp_5_bits_data_0 = writeQueue_5_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_5_writeData_mask;
  wire [3:0]         exeResp_5_bits_mask_0 = writeQueue_5_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_5_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_5_writeData_vd;
  wire [2:0]         writeQueue_dataOut_5_index;
  wire [4:0]         writeQueue_5_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_5_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_5 = {writeQueue_5_enq_bits_writeData_groupCounter, writeQueue_5_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_5_enq_bits_writeData_data;
  wire [3:0]         writeQueue_5_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_10 = {writeQueue_5_enq_bits_writeData_data, writeQueue_5_enq_bits_writeData_mask};
  wire               writeQueue_5_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_11 = {writeQueue_5_enq_bits_ffoByOther, writeQueue_dataIn_hi_10, writeQueue_dataIn_lo_5};
  wire [49:0]        writeQueue_dataIn_5 = {writeQueue_dataIn_hi_11, writeQueue_5_enq_bits_index};
  assign writeQueue_dataOut_5_index = _writeQueue_fifo_5_data_out[2:0];
  assign writeQueue_dataOut_5_writeData_vd = _writeQueue_fifo_5_data_out[7:3];
  assign writeQueue_dataOut_5_writeData_groupCounter = _writeQueue_fifo_5_data_out[12:8];
  assign writeQueue_dataOut_5_writeData_mask = _writeQueue_fifo_5_data_out[16:13];
  assign writeQueue_dataOut_5_writeData_data = _writeQueue_fifo_5_data_out[48:17];
  assign writeQueue_dataOut_5_ffoByOther = _writeQueue_fifo_5_data_out[49];
  wire               writeQueue_5_deq_bits_ffoByOther = writeQueue_dataOut_5_ffoByOther;
  assign writeQueue_5_deq_bits_writeData_data = writeQueue_dataOut_5_writeData_data;
  assign writeQueue_5_deq_bits_writeData_mask = writeQueue_dataOut_5_writeData_mask;
  wire [4:0]         writeQueue_5_deq_bits_writeData_groupCounter = writeQueue_dataOut_5_writeData_groupCounter;
  wire [4:0]         writeQueue_5_deq_bits_writeData_vd = writeQueue_dataOut_5_writeData_vd;
  wire [2:0]         writeQueue_5_deq_bits_index = writeQueue_dataOut_5_index;
  wire               writeQueue_5_enq_ready = ~_writeQueue_fifo_5_full;
  wire               writeQueue_5_enq_valid;
  assign writeQueue_6_deq_valid = ~_writeQueue_fifo_6_empty;
  wire               exeResp_6_valid_0 = writeQueue_6_deq_valid;
  wire               writeQueue_dataOut_6_ffoByOther;
  wire [31:0]        writeQueue_dataOut_6_writeData_data;
  wire [31:0]        exeResp_6_bits_data_0 = writeQueue_6_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_6_writeData_mask;
  wire [3:0]         exeResp_6_bits_mask_0 = writeQueue_6_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_6_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_6_writeData_vd;
  wire [2:0]         writeQueue_dataOut_6_index;
  wire [4:0]         writeQueue_6_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_6_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_6 = {writeQueue_6_enq_bits_writeData_groupCounter, writeQueue_6_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_6_enq_bits_writeData_data;
  wire [3:0]         writeQueue_6_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_12 = {writeQueue_6_enq_bits_writeData_data, writeQueue_6_enq_bits_writeData_mask};
  wire               writeQueue_6_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_13 = {writeQueue_6_enq_bits_ffoByOther, writeQueue_dataIn_hi_12, writeQueue_dataIn_lo_6};
  wire [49:0]        writeQueue_dataIn_6 = {writeQueue_dataIn_hi_13, writeQueue_6_enq_bits_index};
  assign writeQueue_dataOut_6_index = _writeQueue_fifo_6_data_out[2:0];
  assign writeQueue_dataOut_6_writeData_vd = _writeQueue_fifo_6_data_out[7:3];
  assign writeQueue_dataOut_6_writeData_groupCounter = _writeQueue_fifo_6_data_out[12:8];
  assign writeQueue_dataOut_6_writeData_mask = _writeQueue_fifo_6_data_out[16:13];
  assign writeQueue_dataOut_6_writeData_data = _writeQueue_fifo_6_data_out[48:17];
  assign writeQueue_dataOut_6_ffoByOther = _writeQueue_fifo_6_data_out[49];
  wire               writeQueue_6_deq_bits_ffoByOther = writeQueue_dataOut_6_ffoByOther;
  assign writeQueue_6_deq_bits_writeData_data = writeQueue_dataOut_6_writeData_data;
  assign writeQueue_6_deq_bits_writeData_mask = writeQueue_dataOut_6_writeData_mask;
  wire [4:0]         writeQueue_6_deq_bits_writeData_groupCounter = writeQueue_dataOut_6_writeData_groupCounter;
  wire [4:0]         writeQueue_6_deq_bits_writeData_vd = writeQueue_dataOut_6_writeData_vd;
  wire [2:0]         writeQueue_6_deq_bits_index = writeQueue_dataOut_6_index;
  wire               writeQueue_6_enq_ready = ~_writeQueue_fifo_6_full;
  wire               writeQueue_6_enq_valid;
  assign writeQueue_7_deq_valid = ~_writeQueue_fifo_7_empty;
  wire               exeResp_7_valid_0 = writeQueue_7_deq_valid;
  wire               writeQueue_dataOut_7_ffoByOther;
  wire [31:0]        writeQueue_dataOut_7_writeData_data;
  wire [31:0]        exeResp_7_bits_data_0 = writeQueue_7_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_7_writeData_mask;
  wire [3:0]         exeResp_7_bits_mask_0 = writeQueue_7_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_7_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_7_writeData_vd;
  wire [2:0]         writeQueue_dataOut_7_index;
  wire [4:0]         writeQueue_7_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_7_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_7 = {writeQueue_7_enq_bits_writeData_groupCounter, writeQueue_7_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_7_enq_bits_writeData_data;
  wire [3:0]         writeQueue_7_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_14 = {writeQueue_7_enq_bits_writeData_data, writeQueue_7_enq_bits_writeData_mask};
  wire               writeQueue_7_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_15 = {writeQueue_7_enq_bits_ffoByOther, writeQueue_dataIn_hi_14, writeQueue_dataIn_lo_7};
  wire [49:0]        writeQueue_dataIn_7 = {writeQueue_dataIn_hi_15, writeQueue_7_enq_bits_index};
  assign writeQueue_dataOut_7_index = _writeQueue_fifo_7_data_out[2:0];
  assign writeQueue_dataOut_7_writeData_vd = _writeQueue_fifo_7_data_out[7:3];
  assign writeQueue_dataOut_7_writeData_groupCounter = _writeQueue_fifo_7_data_out[12:8];
  assign writeQueue_dataOut_7_writeData_mask = _writeQueue_fifo_7_data_out[16:13];
  assign writeQueue_dataOut_7_writeData_data = _writeQueue_fifo_7_data_out[48:17];
  assign writeQueue_dataOut_7_ffoByOther = _writeQueue_fifo_7_data_out[49];
  wire               writeQueue_7_deq_bits_ffoByOther = writeQueue_dataOut_7_ffoByOther;
  assign writeQueue_7_deq_bits_writeData_data = writeQueue_dataOut_7_writeData_data;
  assign writeQueue_7_deq_bits_writeData_mask = writeQueue_dataOut_7_writeData_mask;
  wire [4:0]         writeQueue_7_deq_bits_writeData_groupCounter = writeQueue_dataOut_7_writeData_groupCounter;
  wire [4:0]         writeQueue_7_deq_bits_writeData_vd = writeQueue_dataOut_7_writeData_vd;
  wire [2:0]         writeQueue_7_deq_bits_index = writeQueue_dataOut_7_index;
  wire               writeQueue_7_enq_ready = ~_writeQueue_fifo_7_full;
  wire               writeQueue_7_enq_valid;
  assign writeQueue_8_deq_valid = ~_writeQueue_fifo_8_empty;
  wire               exeResp_8_valid_0 = writeQueue_8_deq_valid;
  wire               writeQueue_dataOut_8_ffoByOther;
  wire [31:0]        writeQueue_dataOut_8_writeData_data;
  wire [31:0]        exeResp_8_bits_data_0 = writeQueue_8_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_8_writeData_mask;
  wire [3:0]         exeResp_8_bits_mask_0 = writeQueue_8_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_8_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_8_writeData_vd;
  wire [2:0]         writeQueue_dataOut_8_index;
  wire [4:0]         writeQueue_8_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_8_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_8 = {writeQueue_8_enq_bits_writeData_groupCounter, writeQueue_8_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_8_enq_bits_writeData_data;
  wire [3:0]         writeQueue_8_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_16 = {writeQueue_8_enq_bits_writeData_data, writeQueue_8_enq_bits_writeData_mask};
  wire               writeQueue_8_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_17 = {writeQueue_8_enq_bits_ffoByOther, writeQueue_dataIn_hi_16, writeQueue_dataIn_lo_8};
  wire [49:0]        writeQueue_dataIn_8 = {writeQueue_dataIn_hi_17, writeQueue_8_enq_bits_index};
  assign writeQueue_dataOut_8_index = _writeQueue_fifo_8_data_out[2:0];
  assign writeQueue_dataOut_8_writeData_vd = _writeQueue_fifo_8_data_out[7:3];
  assign writeQueue_dataOut_8_writeData_groupCounter = _writeQueue_fifo_8_data_out[12:8];
  assign writeQueue_dataOut_8_writeData_mask = _writeQueue_fifo_8_data_out[16:13];
  assign writeQueue_dataOut_8_writeData_data = _writeQueue_fifo_8_data_out[48:17];
  assign writeQueue_dataOut_8_ffoByOther = _writeQueue_fifo_8_data_out[49];
  wire               writeQueue_8_deq_bits_ffoByOther = writeQueue_dataOut_8_ffoByOther;
  assign writeQueue_8_deq_bits_writeData_data = writeQueue_dataOut_8_writeData_data;
  assign writeQueue_8_deq_bits_writeData_mask = writeQueue_dataOut_8_writeData_mask;
  wire [4:0]         writeQueue_8_deq_bits_writeData_groupCounter = writeQueue_dataOut_8_writeData_groupCounter;
  wire [4:0]         writeQueue_8_deq_bits_writeData_vd = writeQueue_dataOut_8_writeData_vd;
  wire [2:0]         writeQueue_8_deq_bits_index = writeQueue_dataOut_8_index;
  wire               writeQueue_8_enq_ready = ~_writeQueue_fifo_8_full;
  wire               writeQueue_8_enq_valid;
  assign writeQueue_9_deq_valid = ~_writeQueue_fifo_9_empty;
  wire               exeResp_9_valid_0 = writeQueue_9_deq_valid;
  wire               writeQueue_dataOut_9_ffoByOther;
  wire [31:0]        writeQueue_dataOut_9_writeData_data;
  wire [31:0]        exeResp_9_bits_data_0 = writeQueue_9_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_9_writeData_mask;
  wire [3:0]         exeResp_9_bits_mask_0 = writeQueue_9_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_9_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_9_writeData_vd;
  wire [2:0]         writeQueue_dataOut_9_index;
  wire [4:0]         writeQueue_9_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_9_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_9 = {writeQueue_9_enq_bits_writeData_groupCounter, writeQueue_9_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_9_enq_bits_writeData_data;
  wire [3:0]         writeQueue_9_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_18 = {writeQueue_9_enq_bits_writeData_data, writeQueue_9_enq_bits_writeData_mask};
  wire               writeQueue_9_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_19 = {writeQueue_9_enq_bits_ffoByOther, writeQueue_dataIn_hi_18, writeQueue_dataIn_lo_9};
  wire [49:0]        writeQueue_dataIn_9 = {writeQueue_dataIn_hi_19, writeQueue_9_enq_bits_index};
  assign writeQueue_dataOut_9_index = _writeQueue_fifo_9_data_out[2:0];
  assign writeQueue_dataOut_9_writeData_vd = _writeQueue_fifo_9_data_out[7:3];
  assign writeQueue_dataOut_9_writeData_groupCounter = _writeQueue_fifo_9_data_out[12:8];
  assign writeQueue_dataOut_9_writeData_mask = _writeQueue_fifo_9_data_out[16:13];
  assign writeQueue_dataOut_9_writeData_data = _writeQueue_fifo_9_data_out[48:17];
  assign writeQueue_dataOut_9_ffoByOther = _writeQueue_fifo_9_data_out[49];
  wire               writeQueue_9_deq_bits_ffoByOther = writeQueue_dataOut_9_ffoByOther;
  assign writeQueue_9_deq_bits_writeData_data = writeQueue_dataOut_9_writeData_data;
  assign writeQueue_9_deq_bits_writeData_mask = writeQueue_dataOut_9_writeData_mask;
  wire [4:0]         writeQueue_9_deq_bits_writeData_groupCounter = writeQueue_dataOut_9_writeData_groupCounter;
  wire [4:0]         writeQueue_9_deq_bits_writeData_vd = writeQueue_dataOut_9_writeData_vd;
  wire [2:0]         writeQueue_9_deq_bits_index = writeQueue_dataOut_9_index;
  wire               writeQueue_9_enq_ready = ~_writeQueue_fifo_9_full;
  wire               writeQueue_9_enq_valid;
  assign writeQueue_10_deq_valid = ~_writeQueue_fifo_10_empty;
  wire               exeResp_10_valid_0 = writeQueue_10_deq_valid;
  wire               writeQueue_dataOut_10_ffoByOther;
  wire [31:0]        writeQueue_dataOut_10_writeData_data;
  wire [31:0]        exeResp_10_bits_data_0 = writeQueue_10_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_10_writeData_mask;
  wire [3:0]         exeResp_10_bits_mask_0 = writeQueue_10_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_10_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_10_writeData_vd;
  wire [2:0]         writeQueue_dataOut_10_index;
  wire [4:0]         writeQueue_10_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_10_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_10 = {writeQueue_10_enq_bits_writeData_groupCounter, writeQueue_10_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_10_enq_bits_writeData_data;
  wire [3:0]         writeQueue_10_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_20 = {writeQueue_10_enq_bits_writeData_data, writeQueue_10_enq_bits_writeData_mask};
  wire               writeQueue_10_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_21 = {writeQueue_10_enq_bits_ffoByOther, writeQueue_dataIn_hi_20, writeQueue_dataIn_lo_10};
  wire [49:0]        writeQueue_dataIn_10 = {writeQueue_dataIn_hi_21, writeQueue_10_enq_bits_index};
  assign writeQueue_dataOut_10_index = _writeQueue_fifo_10_data_out[2:0];
  assign writeQueue_dataOut_10_writeData_vd = _writeQueue_fifo_10_data_out[7:3];
  assign writeQueue_dataOut_10_writeData_groupCounter = _writeQueue_fifo_10_data_out[12:8];
  assign writeQueue_dataOut_10_writeData_mask = _writeQueue_fifo_10_data_out[16:13];
  assign writeQueue_dataOut_10_writeData_data = _writeQueue_fifo_10_data_out[48:17];
  assign writeQueue_dataOut_10_ffoByOther = _writeQueue_fifo_10_data_out[49];
  wire               writeQueue_10_deq_bits_ffoByOther = writeQueue_dataOut_10_ffoByOther;
  assign writeQueue_10_deq_bits_writeData_data = writeQueue_dataOut_10_writeData_data;
  assign writeQueue_10_deq_bits_writeData_mask = writeQueue_dataOut_10_writeData_mask;
  wire [4:0]         writeQueue_10_deq_bits_writeData_groupCounter = writeQueue_dataOut_10_writeData_groupCounter;
  wire [4:0]         writeQueue_10_deq_bits_writeData_vd = writeQueue_dataOut_10_writeData_vd;
  wire [2:0]         writeQueue_10_deq_bits_index = writeQueue_dataOut_10_index;
  wire               writeQueue_10_enq_ready = ~_writeQueue_fifo_10_full;
  wire               writeQueue_10_enq_valid;
  assign writeQueue_11_deq_valid = ~_writeQueue_fifo_11_empty;
  wire               exeResp_11_valid_0 = writeQueue_11_deq_valid;
  wire               writeQueue_dataOut_11_ffoByOther;
  wire [31:0]        writeQueue_dataOut_11_writeData_data;
  wire [31:0]        exeResp_11_bits_data_0 = writeQueue_11_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_11_writeData_mask;
  wire [3:0]         exeResp_11_bits_mask_0 = writeQueue_11_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_11_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_11_writeData_vd;
  wire [2:0]         writeQueue_dataOut_11_index;
  wire [4:0]         writeQueue_11_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_11_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_11 = {writeQueue_11_enq_bits_writeData_groupCounter, writeQueue_11_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_11_enq_bits_writeData_data;
  wire [3:0]         writeQueue_11_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_22 = {writeQueue_11_enq_bits_writeData_data, writeQueue_11_enq_bits_writeData_mask};
  wire               writeQueue_11_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_23 = {writeQueue_11_enq_bits_ffoByOther, writeQueue_dataIn_hi_22, writeQueue_dataIn_lo_11};
  wire [49:0]        writeQueue_dataIn_11 = {writeQueue_dataIn_hi_23, writeQueue_11_enq_bits_index};
  assign writeQueue_dataOut_11_index = _writeQueue_fifo_11_data_out[2:0];
  assign writeQueue_dataOut_11_writeData_vd = _writeQueue_fifo_11_data_out[7:3];
  assign writeQueue_dataOut_11_writeData_groupCounter = _writeQueue_fifo_11_data_out[12:8];
  assign writeQueue_dataOut_11_writeData_mask = _writeQueue_fifo_11_data_out[16:13];
  assign writeQueue_dataOut_11_writeData_data = _writeQueue_fifo_11_data_out[48:17];
  assign writeQueue_dataOut_11_ffoByOther = _writeQueue_fifo_11_data_out[49];
  wire               writeQueue_11_deq_bits_ffoByOther = writeQueue_dataOut_11_ffoByOther;
  assign writeQueue_11_deq_bits_writeData_data = writeQueue_dataOut_11_writeData_data;
  assign writeQueue_11_deq_bits_writeData_mask = writeQueue_dataOut_11_writeData_mask;
  wire [4:0]         writeQueue_11_deq_bits_writeData_groupCounter = writeQueue_dataOut_11_writeData_groupCounter;
  wire [4:0]         writeQueue_11_deq_bits_writeData_vd = writeQueue_dataOut_11_writeData_vd;
  wire [2:0]         writeQueue_11_deq_bits_index = writeQueue_dataOut_11_index;
  wire               writeQueue_11_enq_ready = ~_writeQueue_fifo_11_full;
  wire               writeQueue_11_enq_valid;
  assign writeQueue_12_deq_valid = ~_writeQueue_fifo_12_empty;
  wire               exeResp_12_valid_0 = writeQueue_12_deq_valid;
  wire               writeQueue_dataOut_12_ffoByOther;
  wire [31:0]        writeQueue_dataOut_12_writeData_data;
  wire [31:0]        exeResp_12_bits_data_0 = writeQueue_12_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_12_writeData_mask;
  wire [3:0]         exeResp_12_bits_mask_0 = writeQueue_12_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_12_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_12_writeData_vd;
  wire [2:0]         writeQueue_dataOut_12_index;
  wire [4:0]         writeQueue_12_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_12_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_12 = {writeQueue_12_enq_bits_writeData_groupCounter, writeQueue_12_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_12_enq_bits_writeData_data;
  wire [3:0]         writeQueue_12_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_24 = {writeQueue_12_enq_bits_writeData_data, writeQueue_12_enq_bits_writeData_mask};
  wire               writeQueue_12_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_25 = {writeQueue_12_enq_bits_ffoByOther, writeQueue_dataIn_hi_24, writeQueue_dataIn_lo_12};
  wire [49:0]        writeQueue_dataIn_12 = {writeQueue_dataIn_hi_25, writeQueue_12_enq_bits_index};
  assign writeQueue_dataOut_12_index = _writeQueue_fifo_12_data_out[2:0];
  assign writeQueue_dataOut_12_writeData_vd = _writeQueue_fifo_12_data_out[7:3];
  assign writeQueue_dataOut_12_writeData_groupCounter = _writeQueue_fifo_12_data_out[12:8];
  assign writeQueue_dataOut_12_writeData_mask = _writeQueue_fifo_12_data_out[16:13];
  assign writeQueue_dataOut_12_writeData_data = _writeQueue_fifo_12_data_out[48:17];
  assign writeQueue_dataOut_12_ffoByOther = _writeQueue_fifo_12_data_out[49];
  wire               writeQueue_12_deq_bits_ffoByOther = writeQueue_dataOut_12_ffoByOther;
  assign writeQueue_12_deq_bits_writeData_data = writeQueue_dataOut_12_writeData_data;
  assign writeQueue_12_deq_bits_writeData_mask = writeQueue_dataOut_12_writeData_mask;
  wire [4:0]         writeQueue_12_deq_bits_writeData_groupCounter = writeQueue_dataOut_12_writeData_groupCounter;
  wire [4:0]         writeQueue_12_deq_bits_writeData_vd = writeQueue_dataOut_12_writeData_vd;
  wire [2:0]         writeQueue_12_deq_bits_index = writeQueue_dataOut_12_index;
  wire               writeQueue_12_enq_ready = ~_writeQueue_fifo_12_full;
  wire               writeQueue_12_enq_valid;
  assign writeQueue_13_deq_valid = ~_writeQueue_fifo_13_empty;
  wire               exeResp_13_valid_0 = writeQueue_13_deq_valid;
  wire               writeQueue_dataOut_13_ffoByOther;
  wire [31:0]        writeQueue_dataOut_13_writeData_data;
  wire [31:0]        exeResp_13_bits_data_0 = writeQueue_13_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_13_writeData_mask;
  wire [3:0]         exeResp_13_bits_mask_0 = writeQueue_13_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_13_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_13_writeData_vd;
  wire [2:0]         writeQueue_dataOut_13_index;
  wire [4:0]         writeQueue_13_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_13_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_13 = {writeQueue_13_enq_bits_writeData_groupCounter, writeQueue_13_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_13_enq_bits_writeData_data;
  wire [3:0]         writeQueue_13_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_26 = {writeQueue_13_enq_bits_writeData_data, writeQueue_13_enq_bits_writeData_mask};
  wire               writeQueue_13_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_27 = {writeQueue_13_enq_bits_ffoByOther, writeQueue_dataIn_hi_26, writeQueue_dataIn_lo_13};
  wire [49:0]        writeQueue_dataIn_13 = {writeQueue_dataIn_hi_27, writeQueue_13_enq_bits_index};
  assign writeQueue_dataOut_13_index = _writeQueue_fifo_13_data_out[2:0];
  assign writeQueue_dataOut_13_writeData_vd = _writeQueue_fifo_13_data_out[7:3];
  assign writeQueue_dataOut_13_writeData_groupCounter = _writeQueue_fifo_13_data_out[12:8];
  assign writeQueue_dataOut_13_writeData_mask = _writeQueue_fifo_13_data_out[16:13];
  assign writeQueue_dataOut_13_writeData_data = _writeQueue_fifo_13_data_out[48:17];
  assign writeQueue_dataOut_13_ffoByOther = _writeQueue_fifo_13_data_out[49];
  wire               writeQueue_13_deq_bits_ffoByOther = writeQueue_dataOut_13_ffoByOther;
  assign writeQueue_13_deq_bits_writeData_data = writeQueue_dataOut_13_writeData_data;
  assign writeQueue_13_deq_bits_writeData_mask = writeQueue_dataOut_13_writeData_mask;
  wire [4:0]         writeQueue_13_deq_bits_writeData_groupCounter = writeQueue_dataOut_13_writeData_groupCounter;
  wire [4:0]         writeQueue_13_deq_bits_writeData_vd = writeQueue_dataOut_13_writeData_vd;
  wire [2:0]         writeQueue_13_deq_bits_index = writeQueue_dataOut_13_index;
  wire               writeQueue_13_enq_ready = ~_writeQueue_fifo_13_full;
  wire               writeQueue_13_enq_valid;
  assign writeQueue_14_deq_valid = ~_writeQueue_fifo_14_empty;
  wire               exeResp_14_valid_0 = writeQueue_14_deq_valid;
  wire               writeQueue_dataOut_14_ffoByOther;
  wire [31:0]        writeQueue_dataOut_14_writeData_data;
  wire [31:0]        exeResp_14_bits_data_0 = writeQueue_14_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_14_writeData_mask;
  wire [3:0]         exeResp_14_bits_mask_0 = writeQueue_14_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_14_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_14_writeData_vd;
  wire [2:0]         writeQueue_dataOut_14_index;
  wire [4:0]         writeQueue_14_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_14_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_14 = {writeQueue_14_enq_bits_writeData_groupCounter, writeQueue_14_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_14_enq_bits_writeData_data;
  wire [3:0]         writeQueue_14_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_28 = {writeQueue_14_enq_bits_writeData_data, writeQueue_14_enq_bits_writeData_mask};
  wire               writeQueue_14_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_29 = {writeQueue_14_enq_bits_ffoByOther, writeQueue_dataIn_hi_28, writeQueue_dataIn_lo_14};
  wire [49:0]        writeQueue_dataIn_14 = {writeQueue_dataIn_hi_29, writeQueue_14_enq_bits_index};
  assign writeQueue_dataOut_14_index = _writeQueue_fifo_14_data_out[2:0];
  assign writeQueue_dataOut_14_writeData_vd = _writeQueue_fifo_14_data_out[7:3];
  assign writeQueue_dataOut_14_writeData_groupCounter = _writeQueue_fifo_14_data_out[12:8];
  assign writeQueue_dataOut_14_writeData_mask = _writeQueue_fifo_14_data_out[16:13];
  assign writeQueue_dataOut_14_writeData_data = _writeQueue_fifo_14_data_out[48:17];
  assign writeQueue_dataOut_14_ffoByOther = _writeQueue_fifo_14_data_out[49];
  wire               writeQueue_14_deq_bits_ffoByOther = writeQueue_dataOut_14_ffoByOther;
  assign writeQueue_14_deq_bits_writeData_data = writeQueue_dataOut_14_writeData_data;
  assign writeQueue_14_deq_bits_writeData_mask = writeQueue_dataOut_14_writeData_mask;
  wire [4:0]         writeQueue_14_deq_bits_writeData_groupCounter = writeQueue_dataOut_14_writeData_groupCounter;
  wire [4:0]         writeQueue_14_deq_bits_writeData_vd = writeQueue_dataOut_14_writeData_vd;
  wire [2:0]         writeQueue_14_deq_bits_index = writeQueue_dataOut_14_index;
  wire               writeQueue_14_enq_ready = ~_writeQueue_fifo_14_full;
  wire               writeQueue_14_enq_valid;
  assign writeQueue_15_deq_valid = ~_writeQueue_fifo_15_empty;
  wire               exeResp_15_valid_0 = writeQueue_15_deq_valid;
  wire               writeQueue_dataOut_15_ffoByOther;
  wire [31:0]        writeQueue_dataOut_15_writeData_data;
  wire [31:0]        exeResp_15_bits_data_0 = writeQueue_15_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_15_writeData_mask;
  wire [3:0]         exeResp_15_bits_mask_0 = writeQueue_15_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_15_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_15_writeData_vd;
  wire [2:0]         writeQueue_dataOut_15_index;
  wire [4:0]         writeQueue_15_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_15_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_15 = {writeQueue_15_enq_bits_writeData_groupCounter, writeQueue_15_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_15_enq_bits_writeData_data;
  wire [3:0]         writeQueue_15_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_30 = {writeQueue_15_enq_bits_writeData_data, writeQueue_15_enq_bits_writeData_mask};
  wire               writeQueue_15_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_31 = {writeQueue_15_enq_bits_ffoByOther, writeQueue_dataIn_hi_30, writeQueue_dataIn_lo_15};
  wire [49:0]        writeQueue_dataIn_15 = {writeQueue_dataIn_hi_31, writeQueue_15_enq_bits_index};
  assign writeQueue_dataOut_15_index = _writeQueue_fifo_15_data_out[2:0];
  assign writeQueue_dataOut_15_writeData_vd = _writeQueue_fifo_15_data_out[7:3];
  assign writeQueue_dataOut_15_writeData_groupCounter = _writeQueue_fifo_15_data_out[12:8];
  assign writeQueue_dataOut_15_writeData_mask = _writeQueue_fifo_15_data_out[16:13];
  assign writeQueue_dataOut_15_writeData_data = _writeQueue_fifo_15_data_out[48:17];
  assign writeQueue_dataOut_15_ffoByOther = _writeQueue_fifo_15_data_out[49];
  wire               writeQueue_15_deq_bits_ffoByOther = writeQueue_dataOut_15_ffoByOther;
  assign writeQueue_15_deq_bits_writeData_data = writeQueue_dataOut_15_writeData_data;
  assign writeQueue_15_deq_bits_writeData_mask = writeQueue_dataOut_15_writeData_mask;
  wire [4:0]         writeQueue_15_deq_bits_writeData_groupCounter = writeQueue_dataOut_15_writeData_groupCounter;
  wire [4:0]         writeQueue_15_deq_bits_writeData_vd = writeQueue_dataOut_15_writeData_vd;
  wire [2:0]         writeQueue_15_deq_bits_index = writeQueue_dataOut_15_index;
  wire               writeQueue_15_enq_ready = ~_writeQueue_fifo_15_full;
  wire               writeQueue_15_enq_valid;
  assign writeQueue_16_deq_valid = ~_writeQueue_fifo_16_empty;
  wire               exeResp_16_valid_0 = writeQueue_16_deq_valid;
  wire               writeQueue_dataOut_16_ffoByOther;
  wire [31:0]        writeQueue_dataOut_16_writeData_data;
  wire [31:0]        exeResp_16_bits_data_0 = writeQueue_16_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_16_writeData_mask;
  wire [3:0]         exeResp_16_bits_mask_0 = writeQueue_16_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_16_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_16_writeData_vd;
  wire [2:0]         writeQueue_dataOut_16_index;
  wire [4:0]         writeQueue_16_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_16_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_16 = {writeQueue_16_enq_bits_writeData_groupCounter, writeQueue_16_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_16_enq_bits_writeData_data;
  wire [3:0]         writeQueue_16_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_32 = {writeQueue_16_enq_bits_writeData_data, writeQueue_16_enq_bits_writeData_mask};
  wire               writeQueue_16_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_33 = {writeQueue_16_enq_bits_ffoByOther, writeQueue_dataIn_hi_32, writeQueue_dataIn_lo_16};
  wire [49:0]        writeQueue_dataIn_16 = {writeQueue_dataIn_hi_33, writeQueue_16_enq_bits_index};
  assign writeQueue_dataOut_16_index = _writeQueue_fifo_16_data_out[2:0];
  assign writeQueue_dataOut_16_writeData_vd = _writeQueue_fifo_16_data_out[7:3];
  assign writeQueue_dataOut_16_writeData_groupCounter = _writeQueue_fifo_16_data_out[12:8];
  assign writeQueue_dataOut_16_writeData_mask = _writeQueue_fifo_16_data_out[16:13];
  assign writeQueue_dataOut_16_writeData_data = _writeQueue_fifo_16_data_out[48:17];
  assign writeQueue_dataOut_16_ffoByOther = _writeQueue_fifo_16_data_out[49];
  wire               writeQueue_16_deq_bits_ffoByOther = writeQueue_dataOut_16_ffoByOther;
  assign writeQueue_16_deq_bits_writeData_data = writeQueue_dataOut_16_writeData_data;
  assign writeQueue_16_deq_bits_writeData_mask = writeQueue_dataOut_16_writeData_mask;
  wire [4:0]         writeQueue_16_deq_bits_writeData_groupCounter = writeQueue_dataOut_16_writeData_groupCounter;
  wire [4:0]         writeQueue_16_deq_bits_writeData_vd = writeQueue_dataOut_16_writeData_vd;
  wire [2:0]         writeQueue_16_deq_bits_index = writeQueue_dataOut_16_index;
  wire               writeQueue_16_enq_ready = ~_writeQueue_fifo_16_full;
  wire               writeQueue_16_enq_valid;
  assign writeQueue_17_deq_valid = ~_writeQueue_fifo_17_empty;
  wire               exeResp_17_valid_0 = writeQueue_17_deq_valid;
  wire               writeQueue_dataOut_17_ffoByOther;
  wire [31:0]        writeQueue_dataOut_17_writeData_data;
  wire [31:0]        exeResp_17_bits_data_0 = writeQueue_17_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_17_writeData_mask;
  wire [3:0]         exeResp_17_bits_mask_0 = writeQueue_17_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_17_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_17_writeData_vd;
  wire [2:0]         writeQueue_dataOut_17_index;
  wire [4:0]         writeQueue_17_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_17_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_17 = {writeQueue_17_enq_bits_writeData_groupCounter, writeQueue_17_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_17_enq_bits_writeData_data;
  wire [3:0]         writeQueue_17_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_34 = {writeQueue_17_enq_bits_writeData_data, writeQueue_17_enq_bits_writeData_mask};
  wire               writeQueue_17_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_35 = {writeQueue_17_enq_bits_ffoByOther, writeQueue_dataIn_hi_34, writeQueue_dataIn_lo_17};
  wire [49:0]        writeQueue_dataIn_17 = {writeQueue_dataIn_hi_35, writeQueue_17_enq_bits_index};
  assign writeQueue_dataOut_17_index = _writeQueue_fifo_17_data_out[2:0];
  assign writeQueue_dataOut_17_writeData_vd = _writeQueue_fifo_17_data_out[7:3];
  assign writeQueue_dataOut_17_writeData_groupCounter = _writeQueue_fifo_17_data_out[12:8];
  assign writeQueue_dataOut_17_writeData_mask = _writeQueue_fifo_17_data_out[16:13];
  assign writeQueue_dataOut_17_writeData_data = _writeQueue_fifo_17_data_out[48:17];
  assign writeQueue_dataOut_17_ffoByOther = _writeQueue_fifo_17_data_out[49];
  wire               writeQueue_17_deq_bits_ffoByOther = writeQueue_dataOut_17_ffoByOther;
  assign writeQueue_17_deq_bits_writeData_data = writeQueue_dataOut_17_writeData_data;
  assign writeQueue_17_deq_bits_writeData_mask = writeQueue_dataOut_17_writeData_mask;
  wire [4:0]         writeQueue_17_deq_bits_writeData_groupCounter = writeQueue_dataOut_17_writeData_groupCounter;
  wire [4:0]         writeQueue_17_deq_bits_writeData_vd = writeQueue_dataOut_17_writeData_vd;
  wire [2:0]         writeQueue_17_deq_bits_index = writeQueue_dataOut_17_index;
  wire               writeQueue_17_enq_ready = ~_writeQueue_fifo_17_full;
  wire               writeQueue_17_enq_valid;
  assign writeQueue_18_deq_valid = ~_writeQueue_fifo_18_empty;
  wire               exeResp_18_valid_0 = writeQueue_18_deq_valid;
  wire               writeQueue_dataOut_18_ffoByOther;
  wire [31:0]        writeQueue_dataOut_18_writeData_data;
  wire [31:0]        exeResp_18_bits_data_0 = writeQueue_18_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_18_writeData_mask;
  wire [3:0]         exeResp_18_bits_mask_0 = writeQueue_18_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_18_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_18_writeData_vd;
  wire [2:0]         writeQueue_dataOut_18_index;
  wire [4:0]         writeQueue_18_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_18_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_18 = {writeQueue_18_enq_bits_writeData_groupCounter, writeQueue_18_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_18_enq_bits_writeData_data;
  wire [3:0]         writeQueue_18_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_36 = {writeQueue_18_enq_bits_writeData_data, writeQueue_18_enq_bits_writeData_mask};
  wire               writeQueue_18_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_37 = {writeQueue_18_enq_bits_ffoByOther, writeQueue_dataIn_hi_36, writeQueue_dataIn_lo_18};
  wire [49:0]        writeQueue_dataIn_18 = {writeQueue_dataIn_hi_37, writeQueue_18_enq_bits_index};
  assign writeQueue_dataOut_18_index = _writeQueue_fifo_18_data_out[2:0];
  assign writeQueue_dataOut_18_writeData_vd = _writeQueue_fifo_18_data_out[7:3];
  assign writeQueue_dataOut_18_writeData_groupCounter = _writeQueue_fifo_18_data_out[12:8];
  assign writeQueue_dataOut_18_writeData_mask = _writeQueue_fifo_18_data_out[16:13];
  assign writeQueue_dataOut_18_writeData_data = _writeQueue_fifo_18_data_out[48:17];
  assign writeQueue_dataOut_18_ffoByOther = _writeQueue_fifo_18_data_out[49];
  wire               writeQueue_18_deq_bits_ffoByOther = writeQueue_dataOut_18_ffoByOther;
  assign writeQueue_18_deq_bits_writeData_data = writeQueue_dataOut_18_writeData_data;
  assign writeQueue_18_deq_bits_writeData_mask = writeQueue_dataOut_18_writeData_mask;
  wire [4:0]         writeQueue_18_deq_bits_writeData_groupCounter = writeQueue_dataOut_18_writeData_groupCounter;
  wire [4:0]         writeQueue_18_deq_bits_writeData_vd = writeQueue_dataOut_18_writeData_vd;
  wire [2:0]         writeQueue_18_deq_bits_index = writeQueue_dataOut_18_index;
  wire               writeQueue_18_enq_ready = ~_writeQueue_fifo_18_full;
  wire               writeQueue_18_enq_valid;
  assign writeQueue_19_deq_valid = ~_writeQueue_fifo_19_empty;
  wire               exeResp_19_valid_0 = writeQueue_19_deq_valid;
  wire               writeQueue_dataOut_19_ffoByOther;
  wire [31:0]        writeQueue_dataOut_19_writeData_data;
  wire [31:0]        exeResp_19_bits_data_0 = writeQueue_19_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_19_writeData_mask;
  wire [3:0]         exeResp_19_bits_mask_0 = writeQueue_19_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_19_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_19_writeData_vd;
  wire [2:0]         writeQueue_dataOut_19_index;
  wire [4:0]         writeQueue_19_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_19_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_19 = {writeQueue_19_enq_bits_writeData_groupCounter, writeQueue_19_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_19_enq_bits_writeData_data;
  wire [3:0]         writeQueue_19_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_38 = {writeQueue_19_enq_bits_writeData_data, writeQueue_19_enq_bits_writeData_mask};
  wire               writeQueue_19_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_39 = {writeQueue_19_enq_bits_ffoByOther, writeQueue_dataIn_hi_38, writeQueue_dataIn_lo_19};
  wire [49:0]        writeQueue_dataIn_19 = {writeQueue_dataIn_hi_39, writeQueue_19_enq_bits_index};
  assign writeQueue_dataOut_19_index = _writeQueue_fifo_19_data_out[2:0];
  assign writeQueue_dataOut_19_writeData_vd = _writeQueue_fifo_19_data_out[7:3];
  assign writeQueue_dataOut_19_writeData_groupCounter = _writeQueue_fifo_19_data_out[12:8];
  assign writeQueue_dataOut_19_writeData_mask = _writeQueue_fifo_19_data_out[16:13];
  assign writeQueue_dataOut_19_writeData_data = _writeQueue_fifo_19_data_out[48:17];
  assign writeQueue_dataOut_19_ffoByOther = _writeQueue_fifo_19_data_out[49];
  wire               writeQueue_19_deq_bits_ffoByOther = writeQueue_dataOut_19_ffoByOther;
  assign writeQueue_19_deq_bits_writeData_data = writeQueue_dataOut_19_writeData_data;
  assign writeQueue_19_deq_bits_writeData_mask = writeQueue_dataOut_19_writeData_mask;
  wire [4:0]         writeQueue_19_deq_bits_writeData_groupCounter = writeQueue_dataOut_19_writeData_groupCounter;
  wire [4:0]         writeQueue_19_deq_bits_writeData_vd = writeQueue_dataOut_19_writeData_vd;
  wire [2:0]         writeQueue_19_deq_bits_index = writeQueue_dataOut_19_index;
  wire               writeQueue_19_enq_ready = ~_writeQueue_fifo_19_full;
  wire               writeQueue_19_enq_valid;
  assign writeQueue_20_deq_valid = ~_writeQueue_fifo_20_empty;
  wire               exeResp_20_valid_0 = writeQueue_20_deq_valid;
  wire               writeQueue_dataOut_20_ffoByOther;
  wire [31:0]        writeQueue_dataOut_20_writeData_data;
  wire [31:0]        exeResp_20_bits_data_0 = writeQueue_20_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_20_writeData_mask;
  wire [3:0]         exeResp_20_bits_mask_0 = writeQueue_20_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_20_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_20_writeData_vd;
  wire [2:0]         writeQueue_dataOut_20_index;
  wire [4:0]         writeQueue_20_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_20_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_20 = {writeQueue_20_enq_bits_writeData_groupCounter, writeQueue_20_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_20_enq_bits_writeData_data;
  wire [3:0]         writeQueue_20_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_40 = {writeQueue_20_enq_bits_writeData_data, writeQueue_20_enq_bits_writeData_mask};
  wire               writeQueue_20_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_41 = {writeQueue_20_enq_bits_ffoByOther, writeQueue_dataIn_hi_40, writeQueue_dataIn_lo_20};
  wire [49:0]        writeQueue_dataIn_20 = {writeQueue_dataIn_hi_41, writeQueue_20_enq_bits_index};
  assign writeQueue_dataOut_20_index = _writeQueue_fifo_20_data_out[2:0];
  assign writeQueue_dataOut_20_writeData_vd = _writeQueue_fifo_20_data_out[7:3];
  assign writeQueue_dataOut_20_writeData_groupCounter = _writeQueue_fifo_20_data_out[12:8];
  assign writeQueue_dataOut_20_writeData_mask = _writeQueue_fifo_20_data_out[16:13];
  assign writeQueue_dataOut_20_writeData_data = _writeQueue_fifo_20_data_out[48:17];
  assign writeQueue_dataOut_20_ffoByOther = _writeQueue_fifo_20_data_out[49];
  wire               writeQueue_20_deq_bits_ffoByOther = writeQueue_dataOut_20_ffoByOther;
  assign writeQueue_20_deq_bits_writeData_data = writeQueue_dataOut_20_writeData_data;
  assign writeQueue_20_deq_bits_writeData_mask = writeQueue_dataOut_20_writeData_mask;
  wire [4:0]         writeQueue_20_deq_bits_writeData_groupCounter = writeQueue_dataOut_20_writeData_groupCounter;
  wire [4:0]         writeQueue_20_deq_bits_writeData_vd = writeQueue_dataOut_20_writeData_vd;
  wire [2:0]         writeQueue_20_deq_bits_index = writeQueue_dataOut_20_index;
  wire               writeQueue_20_enq_ready = ~_writeQueue_fifo_20_full;
  wire               writeQueue_20_enq_valid;
  assign writeQueue_21_deq_valid = ~_writeQueue_fifo_21_empty;
  wire               exeResp_21_valid_0 = writeQueue_21_deq_valid;
  wire               writeQueue_dataOut_21_ffoByOther;
  wire [31:0]        writeQueue_dataOut_21_writeData_data;
  wire [31:0]        exeResp_21_bits_data_0 = writeQueue_21_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_21_writeData_mask;
  wire [3:0]         exeResp_21_bits_mask_0 = writeQueue_21_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_21_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_21_writeData_vd;
  wire [2:0]         writeQueue_dataOut_21_index;
  wire [4:0]         writeQueue_21_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_21_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_21 = {writeQueue_21_enq_bits_writeData_groupCounter, writeQueue_21_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_21_enq_bits_writeData_data;
  wire [3:0]         writeQueue_21_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_42 = {writeQueue_21_enq_bits_writeData_data, writeQueue_21_enq_bits_writeData_mask};
  wire               writeQueue_21_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_43 = {writeQueue_21_enq_bits_ffoByOther, writeQueue_dataIn_hi_42, writeQueue_dataIn_lo_21};
  wire [49:0]        writeQueue_dataIn_21 = {writeQueue_dataIn_hi_43, writeQueue_21_enq_bits_index};
  assign writeQueue_dataOut_21_index = _writeQueue_fifo_21_data_out[2:0];
  assign writeQueue_dataOut_21_writeData_vd = _writeQueue_fifo_21_data_out[7:3];
  assign writeQueue_dataOut_21_writeData_groupCounter = _writeQueue_fifo_21_data_out[12:8];
  assign writeQueue_dataOut_21_writeData_mask = _writeQueue_fifo_21_data_out[16:13];
  assign writeQueue_dataOut_21_writeData_data = _writeQueue_fifo_21_data_out[48:17];
  assign writeQueue_dataOut_21_ffoByOther = _writeQueue_fifo_21_data_out[49];
  wire               writeQueue_21_deq_bits_ffoByOther = writeQueue_dataOut_21_ffoByOther;
  assign writeQueue_21_deq_bits_writeData_data = writeQueue_dataOut_21_writeData_data;
  assign writeQueue_21_deq_bits_writeData_mask = writeQueue_dataOut_21_writeData_mask;
  wire [4:0]         writeQueue_21_deq_bits_writeData_groupCounter = writeQueue_dataOut_21_writeData_groupCounter;
  wire [4:0]         writeQueue_21_deq_bits_writeData_vd = writeQueue_dataOut_21_writeData_vd;
  wire [2:0]         writeQueue_21_deq_bits_index = writeQueue_dataOut_21_index;
  wire               writeQueue_21_enq_ready = ~_writeQueue_fifo_21_full;
  wire               writeQueue_21_enq_valid;
  assign writeQueue_22_deq_valid = ~_writeQueue_fifo_22_empty;
  wire               exeResp_22_valid_0 = writeQueue_22_deq_valid;
  wire               writeQueue_dataOut_22_ffoByOther;
  wire [31:0]        writeQueue_dataOut_22_writeData_data;
  wire [31:0]        exeResp_22_bits_data_0 = writeQueue_22_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_22_writeData_mask;
  wire [3:0]         exeResp_22_bits_mask_0 = writeQueue_22_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_22_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_22_writeData_vd;
  wire [2:0]         writeQueue_dataOut_22_index;
  wire [4:0]         writeQueue_22_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_22_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_22 = {writeQueue_22_enq_bits_writeData_groupCounter, writeQueue_22_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_22_enq_bits_writeData_data;
  wire [3:0]         writeQueue_22_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_44 = {writeQueue_22_enq_bits_writeData_data, writeQueue_22_enq_bits_writeData_mask};
  wire               writeQueue_22_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_45 = {writeQueue_22_enq_bits_ffoByOther, writeQueue_dataIn_hi_44, writeQueue_dataIn_lo_22};
  wire [49:0]        writeQueue_dataIn_22 = {writeQueue_dataIn_hi_45, writeQueue_22_enq_bits_index};
  assign writeQueue_dataOut_22_index = _writeQueue_fifo_22_data_out[2:0];
  assign writeQueue_dataOut_22_writeData_vd = _writeQueue_fifo_22_data_out[7:3];
  assign writeQueue_dataOut_22_writeData_groupCounter = _writeQueue_fifo_22_data_out[12:8];
  assign writeQueue_dataOut_22_writeData_mask = _writeQueue_fifo_22_data_out[16:13];
  assign writeQueue_dataOut_22_writeData_data = _writeQueue_fifo_22_data_out[48:17];
  assign writeQueue_dataOut_22_ffoByOther = _writeQueue_fifo_22_data_out[49];
  wire               writeQueue_22_deq_bits_ffoByOther = writeQueue_dataOut_22_ffoByOther;
  assign writeQueue_22_deq_bits_writeData_data = writeQueue_dataOut_22_writeData_data;
  assign writeQueue_22_deq_bits_writeData_mask = writeQueue_dataOut_22_writeData_mask;
  wire [4:0]         writeQueue_22_deq_bits_writeData_groupCounter = writeQueue_dataOut_22_writeData_groupCounter;
  wire [4:0]         writeQueue_22_deq_bits_writeData_vd = writeQueue_dataOut_22_writeData_vd;
  wire [2:0]         writeQueue_22_deq_bits_index = writeQueue_dataOut_22_index;
  wire               writeQueue_22_enq_ready = ~_writeQueue_fifo_22_full;
  wire               writeQueue_22_enq_valid;
  assign writeQueue_23_deq_valid = ~_writeQueue_fifo_23_empty;
  wire               exeResp_23_valid_0 = writeQueue_23_deq_valid;
  wire               writeQueue_dataOut_23_ffoByOther;
  wire [31:0]        writeQueue_dataOut_23_writeData_data;
  wire [31:0]        exeResp_23_bits_data_0 = writeQueue_23_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_23_writeData_mask;
  wire [3:0]         exeResp_23_bits_mask_0 = writeQueue_23_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_23_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_23_writeData_vd;
  wire [2:0]         writeQueue_dataOut_23_index;
  wire [4:0]         writeQueue_23_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_23_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_23 = {writeQueue_23_enq_bits_writeData_groupCounter, writeQueue_23_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_23_enq_bits_writeData_data;
  wire [3:0]         writeQueue_23_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_46 = {writeQueue_23_enq_bits_writeData_data, writeQueue_23_enq_bits_writeData_mask};
  wire               writeQueue_23_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_47 = {writeQueue_23_enq_bits_ffoByOther, writeQueue_dataIn_hi_46, writeQueue_dataIn_lo_23};
  wire [49:0]        writeQueue_dataIn_23 = {writeQueue_dataIn_hi_47, writeQueue_23_enq_bits_index};
  assign writeQueue_dataOut_23_index = _writeQueue_fifo_23_data_out[2:0];
  assign writeQueue_dataOut_23_writeData_vd = _writeQueue_fifo_23_data_out[7:3];
  assign writeQueue_dataOut_23_writeData_groupCounter = _writeQueue_fifo_23_data_out[12:8];
  assign writeQueue_dataOut_23_writeData_mask = _writeQueue_fifo_23_data_out[16:13];
  assign writeQueue_dataOut_23_writeData_data = _writeQueue_fifo_23_data_out[48:17];
  assign writeQueue_dataOut_23_ffoByOther = _writeQueue_fifo_23_data_out[49];
  wire               writeQueue_23_deq_bits_ffoByOther = writeQueue_dataOut_23_ffoByOther;
  assign writeQueue_23_deq_bits_writeData_data = writeQueue_dataOut_23_writeData_data;
  assign writeQueue_23_deq_bits_writeData_mask = writeQueue_dataOut_23_writeData_mask;
  wire [4:0]         writeQueue_23_deq_bits_writeData_groupCounter = writeQueue_dataOut_23_writeData_groupCounter;
  wire [4:0]         writeQueue_23_deq_bits_writeData_vd = writeQueue_dataOut_23_writeData_vd;
  wire [2:0]         writeQueue_23_deq_bits_index = writeQueue_dataOut_23_index;
  wire               writeQueue_23_enq_ready = ~_writeQueue_fifo_23_full;
  wire               writeQueue_23_enq_valid;
  assign writeQueue_24_deq_valid = ~_writeQueue_fifo_24_empty;
  wire               exeResp_24_valid_0 = writeQueue_24_deq_valid;
  wire               writeQueue_dataOut_24_ffoByOther;
  wire [31:0]        writeQueue_dataOut_24_writeData_data;
  wire [31:0]        exeResp_24_bits_data_0 = writeQueue_24_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_24_writeData_mask;
  wire [3:0]         exeResp_24_bits_mask_0 = writeQueue_24_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_24_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_24_writeData_vd;
  wire [2:0]         writeQueue_dataOut_24_index;
  wire [4:0]         writeQueue_24_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_24_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_24 = {writeQueue_24_enq_bits_writeData_groupCounter, writeQueue_24_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_24_enq_bits_writeData_data;
  wire [3:0]         writeQueue_24_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_48 = {writeQueue_24_enq_bits_writeData_data, writeQueue_24_enq_bits_writeData_mask};
  wire               writeQueue_24_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_49 = {writeQueue_24_enq_bits_ffoByOther, writeQueue_dataIn_hi_48, writeQueue_dataIn_lo_24};
  wire [49:0]        writeQueue_dataIn_24 = {writeQueue_dataIn_hi_49, writeQueue_24_enq_bits_index};
  assign writeQueue_dataOut_24_index = _writeQueue_fifo_24_data_out[2:0];
  assign writeQueue_dataOut_24_writeData_vd = _writeQueue_fifo_24_data_out[7:3];
  assign writeQueue_dataOut_24_writeData_groupCounter = _writeQueue_fifo_24_data_out[12:8];
  assign writeQueue_dataOut_24_writeData_mask = _writeQueue_fifo_24_data_out[16:13];
  assign writeQueue_dataOut_24_writeData_data = _writeQueue_fifo_24_data_out[48:17];
  assign writeQueue_dataOut_24_ffoByOther = _writeQueue_fifo_24_data_out[49];
  wire               writeQueue_24_deq_bits_ffoByOther = writeQueue_dataOut_24_ffoByOther;
  assign writeQueue_24_deq_bits_writeData_data = writeQueue_dataOut_24_writeData_data;
  assign writeQueue_24_deq_bits_writeData_mask = writeQueue_dataOut_24_writeData_mask;
  wire [4:0]         writeQueue_24_deq_bits_writeData_groupCounter = writeQueue_dataOut_24_writeData_groupCounter;
  wire [4:0]         writeQueue_24_deq_bits_writeData_vd = writeQueue_dataOut_24_writeData_vd;
  wire [2:0]         writeQueue_24_deq_bits_index = writeQueue_dataOut_24_index;
  wire               writeQueue_24_enq_ready = ~_writeQueue_fifo_24_full;
  wire               writeQueue_24_enq_valid;
  assign writeQueue_25_deq_valid = ~_writeQueue_fifo_25_empty;
  wire               exeResp_25_valid_0 = writeQueue_25_deq_valid;
  wire               writeQueue_dataOut_25_ffoByOther;
  wire [31:0]        writeQueue_dataOut_25_writeData_data;
  wire [31:0]        exeResp_25_bits_data_0 = writeQueue_25_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_25_writeData_mask;
  wire [3:0]         exeResp_25_bits_mask_0 = writeQueue_25_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_25_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_25_writeData_vd;
  wire [2:0]         writeQueue_dataOut_25_index;
  wire [4:0]         writeQueue_25_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_25_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_25 = {writeQueue_25_enq_bits_writeData_groupCounter, writeQueue_25_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_25_enq_bits_writeData_data;
  wire [3:0]         writeQueue_25_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_50 = {writeQueue_25_enq_bits_writeData_data, writeQueue_25_enq_bits_writeData_mask};
  wire               writeQueue_25_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_51 = {writeQueue_25_enq_bits_ffoByOther, writeQueue_dataIn_hi_50, writeQueue_dataIn_lo_25};
  wire [49:0]        writeQueue_dataIn_25 = {writeQueue_dataIn_hi_51, writeQueue_25_enq_bits_index};
  assign writeQueue_dataOut_25_index = _writeQueue_fifo_25_data_out[2:0];
  assign writeQueue_dataOut_25_writeData_vd = _writeQueue_fifo_25_data_out[7:3];
  assign writeQueue_dataOut_25_writeData_groupCounter = _writeQueue_fifo_25_data_out[12:8];
  assign writeQueue_dataOut_25_writeData_mask = _writeQueue_fifo_25_data_out[16:13];
  assign writeQueue_dataOut_25_writeData_data = _writeQueue_fifo_25_data_out[48:17];
  assign writeQueue_dataOut_25_ffoByOther = _writeQueue_fifo_25_data_out[49];
  wire               writeQueue_25_deq_bits_ffoByOther = writeQueue_dataOut_25_ffoByOther;
  assign writeQueue_25_deq_bits_writeData_data = writeQueue_dataOut_25_writeData_data;
  assign writeQueue_25_deq_bits_writeData_mask = writeQueue_dataOut_25_writeData_mask;
  wire [4:0]         writeQueue_25_deq_bits_writeData_groupCounter = writeQueue_dataOut_25_writeData_groupCounter;
  wire [4:0]         writeQueue_25_deq_bits_writeData_vd = writeQueue_dataOut_25_writeData_vd;
  wire [2:0]         writeQueue_25_deq_bits_index = writeQueue_dataOut_25_index;
  wire               writeQueue_25_enq_ready = ~_writeQueue_fifo_25_full;
  wire               writeQueue_25_enq_valid;
  assign writeQueue_26_deq_valid = ~_writeQueue_fifo_26_empty;
  wire               exeResp_26_valid_0 = writeQueue_26_deq_valid;
  wire               writeQueue_dataOut_26_ffoByOther;
  wire [31:0]        writeQueue_dataOut_26_writeData_data;
  wire [31:0]        exeResp_26_bits_data_0 = writeQueue_26_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_26_writeData_mask;
  wire [3:0]         exeResp_26_bits_mask_0 = writeQueue_26_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_26_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_26_writeData_vd;
  wire [2:0]         writeQueue_dataOut_26_index;
  wire [4:0]         writeQueue_26_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_26_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_26 = {writeQueue_26_enq_bits_writeData_groupCounter, writeQueue_26_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_26_enq_bits_writeData_data;
  wire [3:0]         writeQueue_26_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_52 = {writeQueue_26_enq_bits_writeData_data, writeQueue_26_enq_bits_writeData_mask};
  wire               writeQueue_26_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_53 = {writeQueue_26_enq_bits_ffoByOther, writeQueue_dataIn_hi_52, writeQueue_dataIn_lo_26};
  wire [49:0]        writeQueue_dataIn_26 = {writeQueue_dataIn_hi_53, writeQueue_26_enq_bits_index};
  assign writeQueue_dataOut_26_index = _writeQueue_fifo_26_data_out[2:0];
  assign writeQueue_dataOut_26_writeData_vd = _writeQueue_fifo_26_data_out[7:3];
  assign writeQueue_dataOut_26_writeData_groupCounter = _writeQueue_fifo_26_data_out[12:8];
  assign writeQueue_dataOut_26_writeData_mask = _writeQueue_fifo_26_data_out[16:13];
  assign writeQueue_dataOut_26_writeData_data = _writeQueue_fifo_26_data_out[48:17];
  assign writeQueue_dataOut_26_ffoByOther = _writeQueue_fifo_26_data_out[49];
  wire               writeQueue_26_deq_bits_ffoByOther = writeQueue_dataOut_26_ffoByOther;
  assign writeQueue_26_deq_bits_writeData_data = writeQueue_dataOut_26_writeData_data;
  assign writeQueue_26_deq_bits_writeData_mask = writeQueue_dataOut_26_writeData_mask;
  wire [4:0]         writeQueue_26_deq_bits_writeData_groupCounter = writeQueue_dataOut_26_writeData_groupCounter;
  wire [4:0]         writeQueue_26_deq_bits_writeData_vd = writeQueue_dataOut_26_writeData_vd;
  wire [2:0]         writeQueue_26_deq_bits_index = writeQueue_dataOut_26_index;
  wire               writeQueue_26_enq_ready = ~_writeQueue_fifo_26_full;
  wire               writeQueue_26_enq_valid;
  assign writeQueue_27_deq_valid = ~_writeQueue_fifo_27_empty;
  wire               exeResp_27_valid_0 = writeQueue_27_deq_valid;
  wire               writeQueue_dataOut_27_ffoByOther;
  wire [31:0]        writeQueue_dataOut_27_writeData_data;
  wire [31:0]        exeResp_27_bits_data_0 = writeQueue_27_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_27_writeData_mask;
  wire [3:0]         exeResp_27_bits_mask_0 = writeQueue_27_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_27_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_27_writeData_vd;
  wire [2:0]         writeQueue_dataOut_27_index;
  wire [4:0]         writeQueue_27_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_27_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_27 = {writeQueue_27_enq_bits_writeData_groupCounter, writeQueue_27_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_27_enq_bits_writeData_data;
  wire [3:0]         writeQueue_27_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_54 = {writeQueue_27_enq_bits_writeData_data, writeQueue_27_enq_bits_writeData_mask};
  wire               writeQueue_27_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_55 = {writeQueue_27_enq_bits_ffoByOther, writeQueue_dataIn_hi_54, writeQueue_dataIn_lo_27};
  wire [49:0]        writeQueue_dataIn_27 = {writeQueue_dataIn_hi_55, writeQueue_27_enq_bits_index};
  assign writeQueue_dataOut_27_index = _writeQueue_fifo_27_data_out[2:0];
  assign writeQueue_dataOut_27_writeData_vd = _writeQueue_fifo_27_data_out[7:3];
  assign writeQueue_dataOut_27_writeData_groupCounter = _writeQueue_fifo_27_data_out[12:8];
  assign writeQueue_dataOut_27_writeData_mask = _writeQueue_fifo_27_data_out[16:13];
  assign writeQueue_dataOut_27_writeData_data = _writeQueue_fifo_27_data_out[48:17];
  assign writeQueue_dataOut_27_ffoByOther = _writeQueue_fifo_27_data_out[49];
  wire               writeQueue_27_deq_bits_ffoByOther = writeQueue_dataOut_27_ffoByOther;
  assign writeQueue_27_deq_bits_writeData_data = writeQueue_dataOut_27_writeData_data;
  assign writeQueue_27_deq_bits_writeData_mask = writeQueue_dataOut_27_writeData_mask;
  wire [4:0]         writeQueue_27_deq_bits_writeData_groupCounter = writeQueue_dataOut_27_writeData_groupCounter;
  wire [4:0]         writeQueue_27_deq_bits_writeData_vd = writeQueue_dataOut_27_writeData_vd;
  wire [2:0]         writeQueue_27_deq_bits_index = writeQueue_dataOut_27_index;
  wire               writeQueue_27_enq_ready = ~_writeQueue_fifo_27_full;
  wire               writeQueue_27_enq_valid;
  assign writeQueue_28_deq_valid = ~_writeQueue_fifo_28_empty;
  wire               exeResp_28_valid_0 = writeQueue_28_deq_valid;
  wire               writeQueue_dataOut_28_ffoByOther;
  wire [31:0]        writeQueue_dataOut_28_writeData_data;
  wire [31:0]        exeResp_28_bits_data_0 = writeQueue_28_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_28_writeData_mask;
  wire [3:0]         exeResp_28_bits_mask_0 = writeQueue_28_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_28_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_28_writeData_vd;
  wire [2:0]         writeQueue_dataOut_28_index;
  wire [4:0]         writeQueue_28_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_28_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_28 = {writeQueue_28_enq_bits_writeData_groupCounter, writeQueue_28_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_28_enq_bits_writeData_data;
  wire [3:0]         writeQueue_28_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_56 = {writeQueue_28_enq_bits_writeData_data, writeQueue_28_enq_bits_writeData_mask};
  wire               writeQueue_28_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_57 = {writeQueue_28_enq_bits_ffoByOther, writeQueue_dataIn_hi_56, writeQueue_dataIn_lo_28};
  wire [49:0]        writeQueue_dataIn_28 = {writeQueue_dataIn_hi_57, writeQueue_28_enq_bits_index};
  assign writeQueue_dataOut_28_index = _writeQueue_fifo_28_data_out[2:0];
  assign writeQueue_dataOut_28_writeData_vd = _writeQueue_fifo_28_data_out[7:3];
  assign writeQueue_dataOut_28_writeData_groupCounter = _writeQueue_fifo_28_data_out[12:8];
  assign writeQueue_dataOut_28_writeData_mask = _writeQueue_fifo_28_data_out[16:13];
  assign writeQueue_dataOut_28_writeData_data = _writeQueue_fifo_28_data_out[48:17];
  assign writeQueue_dataOut_28_ffoByOther = _writeQueue_fifo_28_data_out[49];
  wire               writeQueue_28_deq_bits_ffoByOther = writeQueue_dataOut_28_ffoByOther;
  assign writeQueue_28_deq_bits_writeData_data = writeQueue_dataOut_28_writeData_data;
  assign writeQueue_28_deq_bits_writeData_mask = writeQueue_dataOut_28_writeData_mask;
  wire [4:0]         writeQueue_28_deq_bits_writeData_groupCounter = writeQueue_dataOut_28_writeData_groupCounter;
  wire [4:0]         writeQueue_28_deq_bits_writeData_vd = writeQueue_dataOut_28_writeData_vd;
  wire [2:0]         writeQueue_28_deq_bits_index = writeQueue_dataOut_28_index;
  wire               writeQueue_28_enq_ready = ~_writeQueue_fifo_28_full;
  wire               writeQueue_28_enq_valid;
  assign writeQueue_29_deq_valid = ~_writeQueue_fifo_29_empty;
  wire               exeResp_29_valid_0 = writeQueue_29_deq_valid;
  wire               writeQueue_dataOut_29_ffoByOther;
  wire [31:0]        writeQueue_dataOut_29_writeData_data;
  wire [31:0]        exeResp_29_bits_data_0 = writeQueue_29_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_29_writeData_mask;
  wire [3:0]         exeResp_29_bits_mask_0 = writeQueue_29_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_29_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_29_writeData_vd;
  wire [2:0]         writeQueue_dataOut_29_index;
  wire [4:0]         writeQueue_29_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_29_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_29 = {writeQueue_29_enq_bits_writeData_groupCounter, writeQueue_29_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_29_enq_bits_writeData_data;
  wire [3:0]         writeQueue_29_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_58 = {writeQueue_29_enq_bits_writeData_data, writeQueue_29_enq_bits_writeData_mask};
  wire               writeQueue_29_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_59 = {writeQueue_29_enq_bits_ffoByOther, writeQueue_dataIn_hi_58, writeQueue_dataIn_lo_29};
  wire [49:0]        writeQueue_dataIn_29 = {writeQueue_dataIn_hi_59, writeQueue_29_enq_bits_index};
  assign writeQueue_dataOut_29_index = _writeQueue_fifo_29_data_out[2:0];
  assign writeQueue_dataOut_29_writeData_vd = _writeQueue_fifo_29_data_out[7:3];
  assign writeQueue_dataOut_29_writeData_groupCounter = _writeQueue_fifo_29_data_out[12:8];
  assign writeQueue_dataOut_29_writeData_mask = _writeQueue_fifo_29_data_out[16:13];
  assign writeQueue_dataOut_29_writeData_data = _writeQueue_fifo_29_data_out[48:17];
  assign writeQueue_dataOut_29_ffoByOther = _writeQueue_fifo_29_data_out[49];
  wire               writeQueue_29_deq_bits_ffoByOther = writeQueue_dataOut_29_ffoByOther;
  assign writeQueue_29_deq_bits_writeData_data = writeQueue_dataOut_29_writeData_data;
  assign writeQueue_29_deq_bits_writeData_mask = writeQueue_dataOut_29_writeData_mask;
  wire [4:0]         writeQueue_29_deq_bits_writeData_groupCounter = writeQueue_dataOut_29_writeData_groupCounter;
  wire [4:0]         writeQueue_29_deq_bits_writeData_vd = writeQueue_dataOut_29_writeData_vd;
  wire [2:0]         writeQueue_29_deq_bits_index = writeQueue_dataOut_29_index;
  wire               writeQueue_29_enq_ready = ~_writeQueue_fifo_29_full;
  wire               writeQueue_29_enq_valid;
  assign writeQueue_30_deq_valid = ~_writeQueue_fifo_30_empty;
  wire               exeResp_30_valid_0 = writeQueue_30_deq_valid;
  wire               writeQueue_dataOut_30_ffoByOther;
  wire [31:0]        writeQueue_dataOut_30_writeData_data;
  wire [31:0]        exeResp_30_bits_data_0 = writeQueue_30_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_30_writeData_mask;
  wire [3:0]         exeResp_30_bits_mask_0 = writeQueue_30_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_30_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_30_writeData_vd;
  wire [2:0]         writeQueue_dataOut_30_index;
  wire [4:0]         writeQueue_30_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_30_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_30 = {writeQueue_30_enq_bits_writeData_groupCounter, writeQueue_30_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_30_enq_bits_writeData_data;
  wire [3:0]         writeQueue_30_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_60 = {writeQueue_30_enq_bits_writeData_data, writeQueue_30_enq_bits_writeData_mask};
  wire               writeQueue_30_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_61 = {writeQueue_30_enq_bits_ffoByOther, writeQueue_dataIn_hi_60, writeQueue_dataIn_lo_30};
  wire [49:0]        writeQueue_dataIn_30 = {writeQueue_dataIn_hi_61, writeQueue_30_enq_bits_index};
  assign writeQueue_dataOut_30_index = _writeQueue_fifo_30_data_out[2:0];
  assign writeQueue_dataOut_30_writeData_vd = _writeQueue_fifo_30_data_out[7:3];
  assign writeQueue_dataOut_30_writeData_groupCounter = _writeQueue_fifo_30_data_out[12:8];
  assign writeQueue_dataOut_30_writeData_mask = _writeQueue_fifo_30_data_out[16:13];
  assign writeQueue_dataOut_30_writeData_data = _writeQueue_fifo_30_data_out[48:17];
  assign writeQueue_dataOut_30_ffoByOther = _writeQueue_fifo_30_data_out[49];
  wire               writeQueue_30_deq_bits_ffoByOther = writeQueue_dataOut_30_ffoByOther;
  assign writeQueue_30_deq_bits_writeData_data = writeQueue_dataOut_30_writeData_data;
  assign writeQueue_30_deq_bits_writeData_mask = writeQueue_dataOut_30_writeData_mask;
  wire [4:0]         writeQueue_30_deq_bits_writeData_groupCounter = writeQueue_dataOut_30_writeData_groupCounter;
  wire [4:0]         writeQueue_30_deq_bits_writeData_vd = writeQueue_dataOut_30_writeData_vd;
  wire [2:0]         writeQueue_30_deq_bits_index = writeQueue_dataOut_30_index;
  wire               writeQueue_30_enq_ready = ~_writeQueue_fifo_30_full;
  wire               writeQueue_30_enq_valid;
  assign writeQueue_31_deq_valid = ~_writeQueue_fifo_31_empty;
  wire               exeResp_31_valid_0 = writeQueue_31_deq_valid;
  wire               writeQueue_dataOut_31_ffoByOther;
  wire [31:0]        writeQueue_dataOut_31_writeData_data;
  wire [31:0]        exeResp_31_bits_data_0 = writeQueue_31_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_31_writeData_mask;
  wire [3:0]         exeResp_31_bits_mask_0 = writeQueue_31_deq_bits_writeData_mask;
  wire [4:0]         writeQueue_dataOut_31_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_31_writeData_vd;
  wire [2:0]         writeQueue_dataOut_31_index;
  wire [4:0]         writeQueue_31_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_31_enq_bits_writeData_vd;
  wire [9:0]         writeQueue_dataIn_lo_31 = {writeQueue_31_enq_bits_writeData_groupCounter, writeQueue_31_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_31_enq_bits_writeData_data;
  wire [3:0]         writeQueue_31_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_62 = {writeQueue_31_enq_bits_writeData_data, writeQueue_31_enq_bits_writeData_mask};
  wire               writeQueue_31_enq_bits_ffoByOther;
  wire [46:0]        writeQueue_dataIn_hi_63 = {writeQueue_31_enq_bits_ffoByOther, writeQueue_dataIn_hi_62, writeQueue_dataIn_lo_31};
  wire [49:0]        writeQueue_dataIn_31 = {writeQueue_dataIn_hi_63, writeQueue_31_enq_bits_index};
  assign writeQueue_dataOut_31_index = _writeQueue_fifo_31_data_out[2:0];
  assign writeQueue_dataOut_31_writeData_vd = _writeQueue_fifo_31_data_out[7:3];
  assign writeQueue_dataOut_31_writeData_groupCounter = _writeQueue_fifo_31_data_out[12:8];
  assign writeQueue_dataOut_31_writeData_mask = _writeQueue_fifo_31_data_out[16:13];
  assign writeQueue_dataOut_31_writeData_data = _writeQueue_fifo_31_data_out[48:17];
  assign writeQueue_dataOut_31_ffoByOther = _writeQueue_fifo_31_data_out[49];
  wire               writeQueue_31_deq_bits_ffoByOther = writeQueue_dataOut_31_ffoByOther;
  assign writeQueue_31_deq_bits_writeData_data = writeQueue_dataOut_31_writeData_data;
  assign writeQueue_31_deq_bits_writeData_mask = writeQueue_dataOut_31_writeData_mask;
  wire [4:0]         writeQueue_31_deq_bits_writeData_groupCounter = writeQueue_dataOut_31_writeData_groupCounter;
  wire [4:0]         writeQueue_31_deq_bits_writeData_vd = writeQueue_dataOut_31_writeData_vd;
  wire [2:0]         writeQueue_31_deq_bits_index = writeQueue_dataOut_31_index;
  wire               writeQueue_31_enq_ready = ~_writeQueue_fifo_31_full;
  wire               writeQueue_31_enq_valid;
  wire               dataNotInShifter_readTypeWriteVrf = waiteStageDeqFire & WillWriteLane[0];
  assign writeQueue_0_enq_valid = _maskedWrite_out_0_valid | dataNotInShifter_readTypeWriteVrf;
  assign writeQueue_0_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_vd : 5'h0;
  assign writeQueue_0_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_groupCounter : _maskedWrite_out_0_bits_writeData_groupCounter;
  assign writeQueue_0_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_mask : _maskedWrite_out_0_bits_writeData_mask;
  assign writeQueue_0_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_data : _maskedWrite_out_0_bits_writeData_data;
  assign writeQueue_0_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf & _maskedWrite_out_0_bits_ffoByOther;
  wire [4:0]         exeResp_0_bits_vd_0 = instReg_vd + {1'h0, writeQueue_0_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_0_bits_offset_0 = writeQueue_0_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter;
  wire               _dataNotInShifter_T = exeResp_0_ready_0 & exeResp_0_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange = _dataNotInShifter_T ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_1 = waiteStageDeqFire & WillWriteLane[1];
  assign writeQueue_1_enq_valid = _maskedWrite_out_1_valid | dataNotInShifter_readTypeWriteVrf_1;
  assign writeQueue_1_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_vd : 5'h0;
  assign writeQueue_1_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_groupCounter : _maskedWrite_out_1_bits_writeData_groupCounter;
  assign writeQueue_1_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_mask : _maskedWrite_out_1_bits_writeData_mask;
  assign writeQueue_1_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_data : _maskedWrite_out_1_bits_writeData_data;
  assign writeQueue_1_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_1 & _maskedWrite_out_1_bits_ffoByOther;
  wire [4:0]         exeResp_1_bits_vd_0 = instReg_vd + {1'h0, writeQueue_1_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_1_bits_offset_0 = writeQueue_1_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_1;
  wire               _dataNotInShifter_T_3 = exeResp_1_ready_0 & exeResp_1_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_1 = _dataNotInShifter_T_3 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_2 = waiteStageDeqFire & WillWriteLane[2];
  assign writeQueue_2_enq_valid = _maskedWrite_out_2_valid | dataNotInShifter_readTypeWriteVrf_2;
  assign writeQueue_2_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_vd : 5'h0;
  assign writeQueue_2_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_groupCounter : _maskedWrite_out_2_bits_writeData_groupCounter;
  assign writeQueue_2_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_mask : _maskedWrite_out_2_bits_writeData_mask;
  assign writeQueue_2_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_data : _maskedWrite_out_2_bits_writeData_data;
  assign writeQueue_2_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_2 & _maskedWrite_out_2_bits_ffoByOther;
  wire [4:0]         exeResp_2_bits_vd_0 = instReg_vd + {1'h0, writeQueue_2_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_2_bits_offset_0 = writeQueue_2_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_2;
  wire               _dataNotInShifter_T_6 = exeResp_2_ready_0 & exeResp_2_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_2 = _dataNotInShifter_T_6 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_3 = waiteStageDeqFire & WillWriteLane[3];
  assign writeQueue_3_enq_valid = _maskedWrite_out_3_valid | dataNotInShifter_readTypeWriteVrf_3;
  assign writeQueue_3_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_vd : 5'h0;
  assign writeQueue_3_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_groupCounter : _maskedWrite_out_3_bits_writeData_groupCounter;
  assign writeQueue_3_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_mask : _maskedWrite_out_3_bits_writeData_mask;
  assign writeQueue_3_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_data : _maskedWrite_out_3_bits_writeData_data;
  assign writeQueue_3_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_3 & _maskedWrite_out_3_bits_ffoByOther;
  wire [4:0]         exeResp_3_bits_vd_0 = instReg_vd + {1'h0, writeQueue_3_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_3_bits_offset_0 = writeQueue_3_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_3;
  wire               _dataNotInShifter_T_9 = exeResp_3_ready_0 & exeResp_3_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_3 = _dataNotInShifter_T_9 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_4 = waiteStageDeqFire & WillWriteLane[4];
  assign writeQueue_4_enq_valid = _maskedWrite_out_4_valid | dataNotInShifter_readTypeWriteVrf_4;
  assign writeQueue_4_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_4 ? writeRequest_4_writeData_vd : 5'h0;
  assign writeQueue_4_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_4 ? writeRequest_4_writeData_groupCounter : _maskedWrite_out_4_bits_writeData_groupCounter;
  assign writeQueue_4_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_4 ? writeRequest_4_writeData_mask : _maskedWrite_out_4_bits_writeData_mask;
  assign writeQueue_4_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_4 ? writeRequest_4_writeData_data : _maskedWrite_out_4_bits_writeData_data;
  assign writeQueue_4_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_4 & _maskedWrite_out_4_bits_ffoByOther;
  wire [4:0]         exeResp_4_bits_vd_0 = instReg_vd + {1'h0, writeQueue_4_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_4_bits_offset_0 = writeQueue_4_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_4;
  wire               _dataNotInShifter_T_12 = exeResp_4_ready_0 & exeResp_4_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_4 = _dataNotInShifter_T_12 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_5 = waiteStageDeqFire & WillWriteLane[5];
  assign writeQueue_5_enq_valid = _maskedWrite_out_5_valid | dataNotInShifter_readTypeWriteVrf_5;
  assign writeQueue_5_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_5 ? writeRequest_5_writeData_vd : 5'h0;
  assign writeQueue_5_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_5 ? writeRequest_5_writeData_groupCounter : _maskedWrite_out_5_bits_writeData_groupCounter;
  assign writeQueue_5_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_5 ? writeRequest_5_writeData_mask : _maskedWrite_out_5_bits_writeData_mask;
  assign writeQueue_5_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_5 ? writeRequest_5_writeData_data : _maskedWrite_out_5_bits_writeData_data;
  assign writeQueue_5_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_5 & _maskedWrite_out_5_bits_ffoByOther;
  wire [4:0]         exeResp_5_bits_vd_0 = instReg_vd + {1'h0, writeQueue_5_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_5_bits_offset_0 = writeQueue_5_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_5;
  wire               _dataNotInShifter_T_15 = exeResp_5_ready_0 & exeResp_5_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_5 = _dataNotInShifter_T_15 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_6 = waiteStageDeqFire & WillWriteLane[6];
  assign writeQueue_6_enq_valid = _maskedWrite_out_6_valid | dataNotInShifter_readTypeWriteVrf_6;
  assign writeQueue_6_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_6 ? writeRequest_6_writeData_vd : 5'h0;
  assign writeQueue_6_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_6 ? writeRequest_6_writeData_groupCounter : _maskedWrite_out_6_bits_writeData_groupCounter;
  assign writeQueue_6_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_6 ? writeRequest_6_writeData_mask : _maskedWrite_out_6_bits_writeData_mask;
  assign writeQueue_6_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_6 ? writeRequest_6_writeData_data : _maskedWrite_out_6_bits_writeData_data;
  assign writeQueue_6_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_6 & _maskedWrite_out_6_bits_ffoByOther;
  wire [4:0]         exeResp_6_bits_vd_0 = instReg_vd + {1'h0, writeQueue_6_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_6_bits_offset_0 = writeQueue_6_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_6;
  wire               _dataNotInShifter_T_18 = exeResp_6_ready_0 & exeResp_6_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_6 = _dataNotInShifter_T_18 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_7 = waiteStageDeqFire & WillWriteLane[7];
  assign writeQueue_7_enq_valid = _maskedWrite_out_7_valid | dataNotInShifter_readTypeWriteVrf_7;
  assign writeQueue_7_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_7 ? writeRequest_7_writeData_vd : 5'h0;
  assign writeQueue_7_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_7 ? writeRequest_7_writeData_groupCounter : _maskedWrite_out_7_bits_writeData_groupCounter;
  assign writeQueue_7_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_7 ? writeRequest_7_writeData_mask : _maskedWrite_out_7_bits_writeData_mask;
  assign writeQueue_7_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_7 ? writeRequest_7_writeData_data : _maskedWrite_out_7_bits_writeData_data;
  assign writeQueue_7_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_7 & _maskedWrite_out_7_bits_ffoByOther;
  wire [4:0]         exeResp_7_bits_vd_0 = instReg_vd + {1'h0, writeQueue_7_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_7_bits_offset_0 = writeQueue_7_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_7;
  wire               _dataNotInShifter_T_21 = exeResp_7_ready_0 & exeResp_7_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_7 = _dataNotInShifter_T_21 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_8 = waiteStageDeqFire & WillWriteLane[8];
  assign writeQueue_8_enq_valid = _maskedWrite_out_8_valid | dataNotInShifter_readTypeWriteVrf_8;
  assign writeQueue_8_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_8 ? writeRequest_8_writeData_vd : 5'h0;
  assign writeQueue_8_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_8 ? writeRequest_8_writeData_groupCounter : _maskedWrite_out_8_bits_writeData_groupCounter;
  assign writeQueue_8_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_8 ? writeRequest_8_writeData_mask : _maskedWrite_out_8_bits_writeData_mask;
  assign writeQueue_8_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_8 ? writeRequest_8_writeData_data : _maskedWrite_out_8_bits_writeData_data;
  assign writeQueue_8_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_8 & _maskedWrite_out_8_bits_ffoByOther;
  wire [4:0]         exeResp_8_bits_vd_0 = instReg_vd + {1'h0, writeQueue_8_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_8_bits_offset_0 = writeQueue_8_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_8;
  wire               _dataNotInShifter_T_24 = exeResp_8_ready_0 & exeResp_8_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_8 = _dataNotInShifter_T_24 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_9 = waiteStageDeqFire & WillWriteLane[9];
  assign writeQueue_9_enq_valid = _maskedWrite_out_9_valid | dataNotInShifter_readTypeWriteVrf_9;
  assign writeQueue_9_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_9 ? writeRequest_9_writeData_vd : 5'h0;
  assign writeQueue_9_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_9 ? writeRequest_9_writeData_groupCounter : _maskedWrite_out_9_bits_writeData_groupCounter;
  assign writeQueue_9_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_9 ? writeRequest_9_writeData_mask : _maskedWrite_out_9_bits_writeData_mask;
  assign writeQueue_9_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_9 ? writeRequest_9_writeData_data : _maskedWrite_out_9_bits_writeData_data;
  assign writeQueue_9_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_9 & _maskedWrite_out_9_bits_ffoByOther;
  wire [4:0]         exeResp_9_bits_vd_0 = instReg_vd + {1'h0, writeQueue_9_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_9_bits_offset_0 = writeQueue_9_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_9;
  wire               _dataNotInShifter_T_27 = exeResp_9_ready_0 & exeResp_9_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_9 = _dataNotInShifter_T_27 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_10 = waiteStageDeqFire & WillWriteLane[10];
  assign writeQueue_10_enq_valid = _maskedWrite_out_10_valid | dataNotInShifter_readTypeWriteVrf_10;
  assign writeQueue_10_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_10 ? writeRequest_10_writeData_vd : 5'h0;
  assign writeQueue_10_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_10 ? writeRequest_10_writeData_groupCounter : _maskedWrite_out_10_bits_writeData_groupCounter;
  assign writeQueue_10_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_10 ? writeRequest_10_writeData_mask : _maskedWrite_out_10_bits_writeData_mask;
  assign writeQueue_10_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_10 ? writeRequest_10_writeData_data : _maskedWrite_out_10_bits_writeData_data;
  assign writeQueue_10_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_10 & _maskedWrite_out_10_bits_ffoByOther;
  wire [4:0]         exeResp_10_bits_vd_0 = instReg_vd + {1'h0, writeQueue_10_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_10_bits_offset_0 = writeQueue_10_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_10;
  wire               _dataNotInShifter_T_30 = exeResp_10_ready_0 & exeResp_10_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_10 = _dataNotInShifter_T_30 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_11 = waiteStageDeqFire & WillWriteLane[11];
  assign writeQueue_11_enq_valid = _maskedWrite_out_11_valid | dataNotInShifter_readTypeWriteVrf_11;
  assign writeQueue_11_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_11 ? writeRequest_11_writeData_vd : 5'h0;
  assign writeQueue_11_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_11 ? writeRequest_11_writeData_groupCounter : _maskedWrite_out_11_bits_writeData_groupCounter;
  assign writeQueue_11_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_11 ? writeRequest_11_writeData_mask : _maskedWrite_out_11_bits_writeData_mask;
  assign writeQueue_11_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_11 ? writeRequest_11_writeData_data : _maskedWrite_out_11_bits_writeData_data;
  assign writeQueue_11_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_11 & _maskedWrite_out_11_bits_ffoByOther;
  wire [4:0]         exeResp_11_bits_vd_0 = instReg_vd + {1'h0, writeQueue_11_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_11_bits_offset_0 = writeQueue_11_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_11;
  wire               _dataNotInShifter_T_33 = exeResp_11_ready_0 & exeResp_11_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_11 = _dataNotInShifter_T_33 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_12 = waiteStageDeqFire & WillWriteLane[12];
  assign writeQueue_12_enq_valid = _maskedWrite_out_12_valid | dataNotInShifter_readTypeWriteVrf_12;
  assign writeQueue_12_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_12 ? writeRequest_12_writeData_vd : 5'h0;
  assign writeQueue_12_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_12 ? writeRequest_12_writeData_groupCounter : _maskedWrite_out_12_bits_writeData_groupCounter;
  assign writeQueue_12_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_12 ? writeRequest_12_writeData_mask : _maskedWrite_out_12_bits_writeData_mask;
  assign writeQueue_12_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_12 ? writeRequest_12_writeData_data : _maskedWrite_out_12_bits_writeData_data;
  assign writeQueue_12_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_12 & _maskedWrite_out_12_bits_ffoByOther;
  wire [4:0]         exeResp_12_bits_vd_0 = instReg_vd + {1'h0, writeQueue_12_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_12_bits_offset_0 = writeQueue_12_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_12;
  wire               _dataNotInShifter_T_36 = exeResp_12_ready_0 & exeResp_12_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_12 = _dataNotInShifter_T_36 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_13 = waiteStageDeqFire & WillWriteLane[13];
  assign writeQueue_13_enq_valid = _maskedWrite_out_13_valid | dataNotInShifter_readTypeWriteVrf_13;
  assign writeQueue_13_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_13 ? writeRequest_13_writeData_vd : 5'h0;
  assign writeQueue_13_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_13 ? writeRequest_13_writeData_groupCounter : _maskedWrite_out_13_bits_writeData_groupCounter;
  assign writeQueue_13_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_13 ? writeRequest_13_writeData_mask : _maskedWrite_out_13_bits_writeData_mask;
  assign writeQueue_13_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_13 ? writeRequest_13_writeData_data : _maskedWrite_out_13_bits_writeData_data;
  assign writeQueue_13_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_13 & _maskedWrite_out_13_bits_ffoByOther;
  wire [4:0]         exeResp_13_bits_vd_0 = instReg_vd + {1'h0, writeQueue_13_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_13_bits_offset_0 = writeQueue_13_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_13;
  wire               _dataNotInShifter_T_39 = exeResp_13_ready_0 & exeResp_13_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_13 = _dataNotInShifter_T_39 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_14 = waiteStageDeqFire & WillWriteLane[14];
  assign writeQueue_14_enq_valid = _maskedWrite_out_14_valid | dataNotInShifter_readTypeWriteVrf_14;
  assign writeQueue_14_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_14 ? writeRequest_14_writeData_vd : 5'h0;
  assign writeQueue_14_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_14 ? writeRequest_14_writeData_groupCounter : _maskedWrite_out_14_bits_writeData_groupCounter;
  assign writeQueue_14_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_14 ? writeRequest_14_writeData_mask : _maskedWrite_out_14_bits_writeData_mask;
  assign writeQueue_14_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_14 ? writeRequest_14_writeData_data : _maskedWrite_out_14_bits_writeData_data;
  assign writeQueue_14_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_14 & _maskedWrite_out_14_bits_ffoByOther;
  wire [4:0]         exeResp_14_bits_vd_0 = instReg_vd + {1'h0, writeQueue_14_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_14_bits_offset_0 = writeQueue_14_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_14;
  wire               _dataNotInShifter_T_42 = exeResp_14_ready_0 & exeResp_14_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_14 = _dataNotInShifter_T_42 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_15 = waiteStageDeqFire & WillWriteLane[15];
  assign writeQueue_15_enq_valid = _maskedWrite_out_15_valid | dataNotInShifter_readTypeWriteVrf_15;
  assign writeQueue_15_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_15 ? writeRequest_15_writeData_vd : 5'h0;
  assign writeQueue_15_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_15 ? writeRequest_15_writeData_groupCounter : _maskedWrite_out_15_bits_writeData_groupCounter;
  assign writeQueue_15_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_15 ? writeRequest_15_writeData_mask : _maskedWrite_out_15_bits_writeData_mask;
  assign writeQueue_15_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_15 ? writeRequest_15_writeData_data : _maskedWrite_out_15_bits_writeData_data;
  assign writeQueue_15_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_15 & _maskedWrite_out_15_bits_ffoByOther;
  wire [4:0]         exeResp_15_bits_vd_0 = instReg_vd + {1'h0, writeQueue_15_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_15_bits_offset_0 = writeQueue_15_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_15;
  wire               _dataNotInShifter_T_45 = exeResp_15_ready_0 & exeResp_15_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_15 = _dataNotInShifter_T_45 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_16 = waiteStageDeqFire & WillWriteLane[16];
  assign writeQueue_16_enq_valid = _maskedWrite_out_16_valid | dataNotInShifter_readTypeWriteVrf_16;
  assign writeQueue_16_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_16 ? writeRequest_16_writeData_vd : 5'h0;
  assign writeQueue_16_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_16 ? writeRequest_16_writeData_groupCounter : _maskedWrite_out_16_bits_writeData_groupCounter;
  assign writeQueue_16_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_16 ? writeRequest_16_writeData_mask : _maskedWrite_out_16_bits_writeData_mask;
  assign writeQueue_16_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_16 ? writeRequest_16_writeData_data : _maskedWrite_out_16_bits_writeData_data;
  assign writeQueue_16_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_16 & _maskedWrite_out_16_bits_ffoByOther;
  wire [4:0]         exeResp_16_bits_vd_0 = instReg_vd + {1'h0, writeQueue_16_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_16_bits_offset_0 = writeQueue_16_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_16;
  wire               _dataNotInShifter_T_48 = exeResp_16_ready_0 & exeResp_16_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_16 = _dataNotInShifter_T_48 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_17 = waiteStageDeqFire & WillWriteLane[17];
  assign writeQueue_17_enq_valid = _maskedWrite_out_17_valid | dataNotInShifter_readTypeWriteVrf_17;
  assign writeQueue_17_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_17 ? writeRequest_17_writeData_vd : 5'h0;
  assign writeQueue_17_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_17 ? writeRequest_17_writeData_groupCounter : _maskedWrite_out_17_bits_writeData_groupCounter;
  assign writeQueue_17_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_17 ? writeRequest_17_writeData_mask : _maskedWrite_out_17_bits_writeData_mask;
  assign writeQueue_17_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_17 ? writeRequest_17_writeData_data : _maskedWrite_out_17_bits_writeData_data;
  assign writeQueue_17_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_17 & _maskedWrite_out_17_bits_ffoByOther;
  wire [4:0]         exeResp_17_bits_vd_0 = instReg_vd + {1'h0, writeQueue_17_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_17_bits_offset_0 = writeQueue_17_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_17;
  wire               _dataNotInShifter_T_51 = exeResp_17_ready_0 & exeResp_17_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_17 = _dataNotInShifter_T_51 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_18 = waiteStageDeqFire & WillWriteLane[18];
  assign writeQueue_18_enq_valid = _maskedWrite_out_18_valid | dataNotInShifter_readTypeWriteVrf_18;
  assign writeQueue_18_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_18 ? writeRequest_18_writeData_vd : 5'h0;
  assign writeQueue_18_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_18 ? writeRequest_18_writeData_groupCounter : _maskedWrite_out_18_bits_writeData_groupCounter;
  assign writeQueue_18_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_18 ? writeRequest_18_writeData_mask : _maskedWrite_out_18_bits_writeData_mask;
  assign writeQueue_18_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_18 ? writeRequest_18_writeData_data : _maskedWrite_out_18_bits_writeData_data;
  assign writeQueue_18_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_18 & _maskedWrite_out_18_bits_ffoByOther;
  wire [4:0]         exeResp_18_bits_vd_0 = instReg_vd + {1'h0, writeQueue_18_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_18_bits_offset_0 = writeQueue_18_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_18;
  wire               _dataNotInShifter_T_54 = exeResp_18_ready_0 & exeResp_18_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_18 = _dataNotInShifter_T_54 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_19 = waiteStageDeqFire & WillWriteLane[19];
  assign writeQueue_19_enq_valid = _maskedWrite_out_19_valid | dataNotInShifter_readTypeWriteVrf_19;
  assign writeQueue_19_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_19 ? writeRequest_19_writeData_vd : 5'h0;
  assign writeQueue_19_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_19 ? writeRequest_19_writeData_groupCounter : _maskedWrite_out_19_bits_writeData_groupCounter;
  assign writeQueue_19_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_19 ? writeRequest_19_writeData_mask : _maskedWrite_out_19_bits_writeData_mask;
  assign writeQueue_19_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_19 ? writeRequest_19_writeData_data : _maskedWrite_out_19_bits_writeData_data;
  assign writeQueue_19_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_19 & _maskedWrite_out_19_bits_ffoByOther;
  wire [4:0]         exeResp_19_bits_vd_0 = instReg_vd + {1'h0, writeQueue_19_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_19_bits_offset_0 = writeQueue_19_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_19;
  wire               _dataNotInShifter_T_57 = exeResp_19_ready_0 & exeResp_19_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_19 = _dataNotInShifter_T_57 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_20 = waiteStageDeqFire & WillWriteLane[20];
  assign writeQueue_20_enq_valid = _maskedWrite_out_20_valid | dataNotInShifter_readTypeWriteVrf_20;
  assign writeQueue_20_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_20 ? writeRequest_20_writeData_vd : 5'h0;
  assign writeQueue_20_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_20 ? writeRequest_20_writeData_groupCounter : _maskedWrite_out_20_bits_writeData_groupCounter;
  assign writeQueue_20_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_20 ? writeRequest_20_writeData_mask : _maskedWrite_out_20_bits_writeData_mask;
  assign writeQueue_20_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_20 ? writeRequest_20_writeData_data : _maskedWrite_out_20_bits_writeData_data;
  assign writeQueue_20_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_20 & _maskedWrite_out_20_bits_ffoByOther;
  wire [4:0]         exeResp_20_bits_vd_0 = instReg_vd + {1'h0, writeQueue_20_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_20_bits_offset_0 = writeQueue_20_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_20;
  wire               _dataNotInShifter_T_60 = exeResp_20_ready_0 & exeResp_20_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_20 = _dataNotInShifter_T_60 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_21 = waiteStageDeqFire & WillWriteLane[21];
  assign writeQueue_21_enq_valid = _maskedWrite_out_21_valid | dataNotInShifter_readTypeWriteVrf_21;
  assign writeQueue_21_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_21 ? writeRequest_21_writeData_vd : 5'h0;
  assign writeQueue_21_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_21 ? writeRequest_21_writeData_groupCounter : _maskedWrite_out_21_bits_writeData_groupCounter;
  assign writeQueue_21_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_21 ? writeRequest_21_writeData_mask : _maskedWrite_out_21_bits_writeData_mask;
  assign writeQueue_21_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_21 ? writeRequest_21_writeData_data : _maskedWrite_out_21_bits_writeData_data;
  assign writeQueue_21_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_21 & _maskedWrite_out_21_bits_ffoByOther;
  wire [4:0]         exeResp_21_bits_vd_0 = instReg_vd + {1'h0, writeQueue_21_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_21_bits_offset_0 = writeQueue_21_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_21;
  wire               _dataNotInShifter_T_63 = exeResp_21_ready_0 & exeResp_21_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_21 = _dataNotInShifter_T_63 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_22 = waiteStageDeqFire & WillWriteLane[22];
  assign writeQueue_22_enq_valid = _maskedWrite_out_22_valid | dataNotInShifter_readTypeWriteVrf_22;
  assign writeQueue_22_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_22 ? writeRequest_22_writeData_vd : 5'h0;
  assign writeQueue_22_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_22 ? writeRequest_22_writeData_groupCounter : _maskedWrite_out_22_bits_writeData_groupCounter;
  assign writeQueue_22_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_22 ? writeRequest_22_writeData_mask : _maskedWrite_out_22_bits_writeData_mask;
  assign writeQueue_22_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_22 ? writeRequest_22_writeData_data : _maskedWrite_out_22_bits_writeData_data;
  assign writeQueue_22_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_22 & _maskedWrite_out_22_bits_ffoByOther;
  wire [4:0]         exeResp_22_bits_vd_0 = instReg_vd + {1'h0, writeQueue_22_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_22_bits_offset_0 = writeQueue_22_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_22;
  wire               _dataNotInShifter_T_66 = exeResp_22_ready_0 & exeResp_22_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_22 = _dataNotInShifter_T_66 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_23 = waiteStageDeqFire & WillWriteLane[23];
  assign writeQueue_23_enq_valid = _maskedWrite_out_23_valid | dataNotInShifter_readTypeWriteVrf_23;
  assign writeQueue_23_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_23 ? writeRequest_23_writeData_vd : 5'h0;
  assign writeQueue_23_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_23 ? writeRequest_23_writeData_groupCounter : _maskedWrite_out_23_bits_writeData_groupCounter;
  assign writeQueue_23_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_23 ? writeRequest_23_writeData_mask : _maskedWrite_out_23_bits_writeData_mask;
  assign writeQueue_23_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_23 ? writeRequest_23_writeData_data : _maskedWrite_out_23_bits_writeData_data;
  assign writeQueue_23_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_23 & _maskedWrite_out_23_bits_ffoByOther;
  wire [4:0]         exeResp_23_bits_vd_0 = instReg_vd + {1'h0, writeQueue_23_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_23_bits_offset_0 = writeQueue_23_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_23;
  wire               _dataNotInShifter_T_69 = exeResp_23_ready_0 & exeResp_23_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_23 = _dataNotInShifter_T_69 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_24 = waiteStageDeqFire & WillWriteLane[24];
  assign writeQueue_24_enq_valid = _maskedWrite_out_24_valid | dataNotInShifter_readTypeWriteVrf_24;
  assign writeQueue_24_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_24 ? writeRequest_24_writeData_vd : 5'h0;
  assign writeQueue_24_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_24 ? writeRequest_24_writeData_groupCounter : _maskedWrite_out_24_bits_writeData_groupCounter;
  assign writeQueue_24_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_24 ? writeRequest_24_writeData_mask : _maskedWrite_out_24_bits_writeData_mask;
  assign writeQueue_24_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_24 ? writeRequest_24_writeData_data : _maskedWrite_out_24_bits_writeData_data;
  assign writeQueue_24_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_24 & _maskedWrite_out_24_bits_ffoByOther;
  wire [4:0]         exeResp_24_bits_vd_0 = instReg_vd + {1'h0, writeQueue_24_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_24_bits_offset_0 = writeQueue_24_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_24;
  wire               _dataNotInShifter_T_72 = exeResp_24_ready_0 & exeResp_24_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_24 = _dataNotInShifter_T_72 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_25 = waiteStageDeqFire & WillWriteLane[25];
  assign writeQueue_25_enq_valid = _maskedWrite_out_25_valid | dataNotInShifter_readTypeWriteVrf_25;
  assign writeQueue_25_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_25 ? writeRequest_25_writeData_vd : 5'h0;
  assign writeQueue_25_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_25 ? writeRequest_25_writeData_groupCounter : _maskedWrite_out_25_bits_writeData_groupCounter;
  assign writeQueue_25_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_25 ? writeRequest_25_writeData_mask : _maskedWrite_out_25_bits_writeData_mask;
  assign writeQueue_25_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_25 ? writeRequest_25_writeData_data : _maskedWrite_out_25_bits_writeData_data;
  assign writeQueue_25_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_25 & _maskedWrite_out_25_bits_ffoByOther;
  wire [4:0]         exeResp_25_bits_vd_0 = instReg_vd + {1'h0, writeQueue_25_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_25_bits_offset_0 = writeQueue_25_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_25;
  wire               _dataNotInShifter_T_75 = exeResp_25_ready_0 & exeResp_25_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_25 = _dataNotInShifter_T_75 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_26 = waiteStageDeqFire & WillWriteLane[26];
  assign writeQueue_26_enq_valid = _maskedWrite_out_26_valid | dataNotInShifter_readTypeWriteVrf_26;
  assign writeQueue_26_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_26 ? writeRequest_26_writeData_vd : 5'h0;
  assign writeQueue_26_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_26 ? writeRequest_26_writeData_groupCounter : _maskedWrite_out_26_bits_writeData_groupCounter;
  assign writeQueue_26_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_26 ? writeRequest_26_writeData_mask : _maskedWrite_out_26_bits_writeData_mask;
  assign writeQueue_26_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_26 ? writeRequest_26_writeData_data : _maskedWrite_out_26_bits_writeData_data;
  assign writeQueue_26_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_26 & _maskedWrite_out_26_bits_ffoByOther;
  wire [4:0]         exeResp_26_bits_vd_0 = instReg_vd + {1'h0, writeQueue_26_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_26_bits_offset_0 = writeQueue_26_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_26;
  wire               _dataNotInShifter_T_78 = exeResp_26_ready_0 & exeResp_26_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_26 = _dataNotInShifter_T_78 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_27 = waiteStageDeqFire & WillWriteLane[27];
  assign writeQueue_27_enq_valid = _maskedWrite_out_27_valid | dataNotInShifter_readTypeWriteVrf_27;
  assign writeQueue_27_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_27 ? writeRequest_27_writeData_vd : 5'h0;
  assign writeQueue_27_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_27 ? writeRequest_27_writeData_groupCounter : _maskedWrite_out_27_bits_writeData_groupCounter;
  assign writeQueue_27_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_27 ? writeRequest_27_writeData_mask : _maskedWrite_out_27_bits_writeData_mask;
  assign writeQueue_27_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_27 ? writeRequest_27_writeData_data : _maskedWrite_out_27_bits_writeData_data;
  assign writeQueue_27_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_27 & _maskedWrite_out_27_bits_ffoByOther;
  wire [4:0]         exeResp_27_bits_vd_0 = instReg_vd + {1'h0, writeQueue_27_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_27_bits_offset_0 = writeQueue_27_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_27;
  wire               _dataNotInShifter_T_81 = exeResp_27_ready_0 & exeResp_27_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_27 = _dataNotInShifter_T_81 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_28 = waiteStageDeqFire & WillWriteLane[28];
  assign writeQueue_28_enq_valid = _maskedWrite_out_28_valid | dataNotInShifter_readTypeWriteVrf_28;
  assign writeQueue_28_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_28 ? writeRequest_28_writeData_vd : 5'h0;
  assign writeQueue_28_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_28 ? writeRequest_28_writeData_groupCounter : _maskedWrite_out_28_bits_writeData_groupCounter;
  assign writeQueue_28_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_28 ? writeRequest_28_writeData_mask : _maskedWrite_out_28_bits_writeData_mask;
  assign writeQueue_28_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_28 ? writeRequest_28_writeData_data : _maskedWrite_out_28_bits_writeData_data;
  assign writeQueue_28_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_28 & _maskedWrite_out_28_bits_ffoByOther;
  wire [4:0]         exeResp_28_bits_vd_0 = instReg_vd + {1'h0, writeQueue_28_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_28_bits_offset_0 = writeQueue_28_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_28;
  wire               _dataNotInShifter_T_84 = exeResp_28_ready_0 & exeResp_28_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_28 = _dataNotInShifter_T_84 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_29 = waiteStageDeqFire & WillWriteLane[29];
  assign writeQueue_29_enq_valid = _maskedWrite_out_29_valid | dataNotInShifter_readTypeWriteVrf_29;
  assign writeQueue_29_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_29 ? writeRequest_29_writeData_vd : 5'h0;
  assign writeQueue_29_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_29 ? writeRequest_29_writeData_groupCounter : _maskedWrite_out_29_bits_writeData_groupCounter;
  assign writeQueue_29_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_29 ? writeRequest_29_writeData_mask : _maskedWrite_out_29_bits_writeData_mask;
  assign writeQueue_29_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_29 ? writeRequest_29_writeData_data : _maskedWrite_out_29_bits_writeData_data;
  assign writeQueue_29_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_29 & _maskedWrite_out_29_bits_ffoByOther;
  wire [4:0]         exeResp_29_bits_vd_0 = instReg_vd + {1'h0, writeQueue_29_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_29_bits_offset_0 = writeQueue_29_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_29;
  wire               _dataNotInShifter_T_87 = exeResp_29_ready_0 & exeResp_29_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_29 = _dataNotInShifter_T_87 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_30 = waiteStageDeqFire & WillWriteLane[30];
  assign writeQueue_30_enq_valid = _maskedWrite_out_30_valid | dataNotInShifter_readTypeWriteVrf_30;
  assign writeQueue_30_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_30 ? writeRequest_30_writeData_vd : 5'h0;
  assign writeQueue_30_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_30 ? writeRequest_30_writeData_groupCounter : _maskedWrite_out_30_bits_writeData_groupCounter;
  assign writeQueue_30_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_30 ? writeRequest_30_writeData_mask : _maskedWrite_out_30_bits_writeData_mask;
  assign writeQueue_30_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_30 ? writeRequest_30_writeData_data : _maskedWrite_out_30_bits_writeData_data;
  assign writeQueue_30_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_30 & _maskedWrite_out_30_bits_ffoByOther;
  wire [4:0]         exeResp_30_bits_vd_0 = instReg_vd + {1'h0, writeQueue_30_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_30_bits_offset_0 = writeQueue_30_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_30;
  wire               _dataNotInShifter_T_90 = exeResp_30_ready_0 & exeResp_30_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_30 = _dataNotInShifter_T_90 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_31 = waiteStageDeqFire & WillWriteLane[31];
  assign writeQueue_31_enq_valid = _maskedWrite_out_31_valid | dataNotInShifter_readTypeWriteVrf_31;
  assign writeQueue_31_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_31 ? writeRequest_31_writeData_vd : 5'h0;
  assign writeQueue_31_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_31 ? writeRequest_31_writeData_groupCounter : _maskedWrite_out_31_bits_writeData_groupCounter;
  assign writeQueue_31_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_31 ? writeRequest_31_writeData_mask : _maskedWrite_out_31_bits_writeData_mask;
  assign writeQueue_31_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_31 ? writeRequest_31_writeData_data : _maskedWrite_out_31_bits_writeData_data;
  assign writeQueue_31_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_31 & _maskedWrite_out_31_bits_ffoByOther;
  wire [4:0]         exeResp_31_bits_vd_0 = instReg_vd + {1'h0, writeQueue_31_deq_bits_writeData_groupCounter[4:1]};
  wire               exeResp_31_bits_offset_0 = writeQueue_31_deq_bits_writeData_groupCounter[0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_31;
  wire               _dataNotInShifter_T_93 = exeResp_31_ready_0 & exeResp_31_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_31 = _dataNotInShifter_T_93 ? 3'h1 : 3'h7;
  wire               dataNotInShifter =
    dataNotInShifter_writeTokenCounter == 3'h0 & dataNotInShifter_writeTokenCounter_1 == 3'h0 & dataNotInShifter_writeTokenCounter_2 == 3'h0 & dataNotInShifter_writeTokenCounter_3 == 3'h0 & dataNotInShifter_writeTokenCounter_4 == 3'h0
    & dataNotInShifter_writeTokenCounter_5 == 3'h0 & dataNotInShifter_writeTokenCounter_6 == 3'h0 & dataNotInShifter_writeTokenCounter_7 == 3'h0 & dataNotInShifter_writeTokenCounter_8 == 3'h0 & dataNotInShifter_writeTokenCounter_9 == 3'h0
    & dataNotInShifter_writeTokenCounter_10 == 3'h0 & dataNotInShifter_writeTokenCounter_11 == 3'h0 & dataNotInShifter_writeTokenCounter_12 == 3'h0 & dataNotInShifter_writeTokenCounter_13 == 3'h0
    & dataNotInShifter_writeTokenCounter_14 == 3'h0 & dataNotInShifter_writeTokenCounter_15 == 3'h0 & dataNotInShifter_writeTokenCounter_16 == 3'h0 & dataNotInShifter_writeTokenCounter_17 == 3'h0
    & dataNotInShifter_writeTokenCounter_18 == 3'h0 & dataNotInShifter_writeTokenCounter_19 == 3'h0 & dataNotInShifter_writeTokenCounter_20 == 3'h0 & dataNotInShifter_writeTokenCounter_21 == 3'h0
    & dataNotInShifter_writeTokenCounter_22 == 3'h0 & dataNotInShifter_writeTokenCounter_23 == 3'h0 & dataNotInShifter_writeTokenCounter_24 == 3'h0 & dataNotInShifter_writeTokenCounter_25 == 3'h0
    & dataNotInShifter_writeTokenCounter_26 == 3'h0 & dataNotInShifter_writeTokenCounter_27 == 3'h0 & dataNotInShifter_writeTokenCounter_28 == 3'h0 & dataNotInShifter_writeTokenCounter_29 == 3'h0
    & dataNotInShifter_writeTokenCounter_30 == 3'h0 & dataNotInShifter_writeTokenCounter_31 == 3'h0;
  assign waiteStageDeqReady =
    (~(WillWriteLane[0]) | writeQueue_0_enq_ready) & (~(WillWriteLane[1]) | writeQueue_1_enq_ready) & (~(WillWriteLane[2]) | writeQueue_2_enq_ready) & (~(WillWriteLane[3]) | writeQueue_3_enq_ready)
    & (~(WillWriteLane[4]) | writeQueue_4_enq_ready) & (~(WillWriteLane[5]) | writeQueue_5_enq_ready) & (~(WillWriteLane[6]) | writeQueue_6_enq_ready) & (~(WillWriteLane[7]) | writeQueue_7_enq_ready)
    & (~(WillWriteLane[8]) | writeQueue_8_enq_ready) & (~(WillWriteLane[9]) | writeQueue_9_enq_ready) & (~(WillWriteLane[10]) | writeQueue_10_enq_ready) & (~(WillWriteLane[11]) | writeQueue_11_enq_ready)
    & (~(WillWriteLane[12]) | writeQueue_12_enq_ready) & (~(WillWriteLane[13]) | writeQueue_13_enq_ready) & (~(WillWriteLane[14]) | writeQueue_14_enq_ready) & (~(WillWriteLane[15]) | writeQueue_15_enq_ready)
    & (~(WillWriteLane[16]) | writeQueue_16_enq_ready) & (~(WillWriteLane[17]) | writeQueue_17_enq_ready) & (~(WillWriteLane[18]) | writeQueue_18_enq_ready) & (~(WillWriteLane[19]) | writeQueue_19_enq_ready)
    & (~(WillWriteLane[20]) | writeQueue_20_enq_ready) & (~(WillWriteLane[21]) | writeQueue_21_enq_ready) & (~(WillWriteLane[22]) | writeQueue_22_enq_ready) & (~(WillWriteLane[23]) | writeQueue_23_enq_ready)
    & (~(WillWriteLane[24]) | writeQueue_24_enq_ready) & (~(WillWriteLane[25]) | writeQueue_25_enq_ready) & (~(WillWriteLane[26]) | writeQueue_26_enq_ready) & (~(WillWriteLane[27]) | writeQueue_27_enq_ready)
    & (~(WillWriteLane[28]) | writeQueue_28_enq_ready) & (~(WillWriteLane[29]) | writeQueue_29_enq_ready) & (~(WillWriteLane[30]) | writeQueue_30_enq_ready) & (~(WillWriteLane[31]) | writeQueue_31_enq_ready);
  reg                waiteLastRequest;
  reg                waitQueueClear;
  wire               lastReportValid =
    waitQueueClear
    & ~(writeQueue_0_deq_valid | writeQueue_1_deq_valid | writeQueue_2_deq_valid | writeQueue_3_deq_valid | writeQueue_4_deq_valid | writeQueue_5_deq_valid | writeQueue_6_deq_valid | writeQueue_7_deq_valid | writeQueue_8_deq_valid
        | writeQueue_9_deq_valid | writeQueue_10_deq_valid | writeQueue_11_deq_valid | writeQueue_12_deq_valid | writeQueue_13_deq_valid | writeQueue_14_deq_valid | writeQueue_15_deq_valid | writeQueue_16_deq_valid | writeQueue_17_deq_valid
        | writeQueue_18_deq_valid | writeQueue_19_deq_valid | writeQueue_20_deq_valid | writeQueue_21_deq_valid | writeQueue_22_deq_valid | writeQueue_23_deq_valid | writeQueue_24_deq_valid | writeQueue_25_deq_valid
        | writeQueue_26_deq_valid | writeQueue_27_deq_valid | writeQueue_28_deq_valid | writeQueue_29_deq_valid | writeQueue_30_deq_valid | writeQueue_31_deq_valid) & dataNotInShifter;
  wire               executeStageInvalid = unitType[1] & ~compressUnitResultQueue_deq_valid & ~_compressUnit_stageValid | unitType[2] & _reduceUnit_in_ready | unitType[3];
  wire               executeStageClean = readType ? waiteStageDeqFire & waiteReadDataPipeReg_last : waiteLastRequest & _maskedWrite_stageClear & executeStageInvalid;
  wire               invalidEnq = instReq_valid & instReq_bits_vl == 12'h0 & ~enqMvRD;
  wire [7:0]         _lastReport_output = lastReportValid ? 8'h1 << instReg_instructionIndex : 8'h0;
  wire [31:0]        gatherData_bits_0 = readVS1Reg_dataValid ? readVS1Reg_data : 32'h0;
  always @(posedge clock) begin
    if (reset) begin
      v0_0 <= 32'h0;
      v0_1 <= 32'h0;
      v0_2 <= 32'h0;
      v0_3 <= 32'h0;
      v0_4 <= 32'h0;
      v0_5 <= 32'h0;
      v0_6 <= 32'h0;
      v0_7 <= 32'h0;
      v0_8 <= 32'h0;
      v0_9 <= 32'h0;
      v0_10 <= 32'h0;
      v0_11 <= 32'h0;
      v0_12 <= 32'h0;
      v0_13 <= 32'h0;
      v0_14 <= 32'h0;
      v0_15 <= 32'h0;
      v0_16 <= 32'h0;
      v0_17 <= 32'h0;
      v0_18 <= 32'h0;
      v0_19 <= 32'h0;
      v0_20 <= 32'h0;
      v0_21 <= 32'h0;
      v0_22 <= 32'h0;
      v0_23 <= 32'h0;
      v0_24 <= 32'h0;
      v0_25 <= 32'h0;
      v0_26 <= 32'h0;
      v0_27 <= 32'h0;
      v0_28 <= 32'h0;
      v0_29 <= 32'h0;
      v0_30 <= 32'h0;
      v0_31 <= 32'h0;
      v0_32 <= 32'h0;
      v0_33 <= 32'h0;
      v0_34 <= 32'h0;
      v0_35 <= 32'h0;
      v0_36 <= 32'h0;
      v0_37 <= 32'h0;
      v0_38 <= 32'h0;
      v0_39 <= 32'h0;
      v0_40 <= 32'h0;
      v0_41 <= 32'h0;
      v0_42 <= 32'h0;
      v0_43 <= 32'h0;
      v0_44 <= 32'h0;
      v0_45 <= 32'h0;
      v0_46 <= 32'h0;
      v0_47 <= 32'h0;
      v0_48 <= 32'h0;
      v0_49 <= 32'h0;
      v0_50 <= 32'h0;
      v0_51 <= 32'h0;
      v0_52 <= 32'h0;
      v0_53 <= 32'h0;
      v0_54 <= 32'h0;
      v0_55 <= 32'h0;
      v0_56 <= 32'h0;
      v0_57 <= 32'h0;
      v0_58 <= 32'h0;
      v0_59 <= 32'h0;
      v0_60 <= 32'h0;
      v0_61 <= 32'h0;
      v0_62 <= 32'h0;
      v0_63 <= 32'h0;
      gatherReadState <= 2'h0;
      gatherDatOffset <= 2'h0;
      gatherLane <= 5'h0;
      gatherOffset <= 1'h0;
      gatherGrowth <= 3'h0;
      instReg_instructionIndex <= 3'h0;
      instReg_decodeResult_specialSlot <= 1'h0;
      instReg_decodeResult_topUop <= 5'h0;
      instReg_decodeResult_popCount <= 1'h0;
      instReg_decodeResult_ffo <= 1'h0;
      instReg_decodeResult_average <= 1'h0;
      instReg_decodeResult_reverse <= 1'h0;
      instReg_decodeResult_dontNeedExecuteInLane <= 1'h0;
      instReg_decodeResult_scheduler <= 1'h0;
      instReg_decodeResult_sReadVD <= 1'h0;
      instReg_decodeResult_vtype <= 1'h0;
      instReg_decodeResult_sWrite <= 1'h0;
      instReg_decodeResult_crossRead <= 1'h0;
      instReg_decodeResult_crossWrite <= 1'h0;
      instReg_decodeResult_maskUnit <= 1'h0;
      instReg_decodeResult_special <= 1'h0;
      instReg_decodeResult_saturate <= 1'h0;
      instReg_decodeResult_vwmacc <= 1'h0;
      instReg_decodeResult_readOnly <= 1'h0;
      instReg_decodeResult_maskSource <= 1'h0;
      instReg_decodeResult_maskDestination <= 1'h0;
      instReg_decodeResult_maskLogic <= 1'h0;
      instReg_decodeResult_uop <= 4'h0;
      instReg_decodeResult_iota <= 1'h0;
      instReg_decodeResult_mv <= 1'h0;
      instReg_decodeResult_extend <= 1'h0;
      instReg_decodeResult_unOrderWrite <= 1'h0;
      instReg_decodeResult_compress <= 1'h0;
      instReg_decodeResult_gather16 <= 1'h0;
      instReg_decodeResult_gather <= 1'h0;
      instReg_decodeResult_slid <= 1'h0;
      instReg_decodeResult_targetRd <= 1'h0;
      instReg_decodeResult_widenReduce <= 1'h0;
      instReg_decodeResult_red <= 1'h0;
      instReg_decodeResult_nr <= 1'h0;
      instReg_decodeResult_itype <= 1'h0;
      instReg_decodeResult_unsigned1 <= 1'h0;
      instReg_decodeResult_unsigned0 <= 1'h0;
      instReg_decodeResult_other <= 1'h0;
      instReg_decodeResult_multiCycle <= 1'h0;
      instReg_decodeResult_divider <= 1'h0;
      instReg_decodeResult_multiplier <= 1'h0;
      instReg_decodeResult_shift <= 1'h0;
      instReg_decodeResult_adder <= 1'h0;
      instReg_decodeResult_logic <= 1'h0;
      instReg_readFromScala <= 32'h0;
      instReg_sew <= 2'h0;
      instReg_vlmul <= 3'h0;
      instReg_maskType <= 1'h0;
      instReg_vxrm <= 3'h0;
      instReg_vs2 <= 5'h0;
      instReg_vs1 <= 5'h0;
      instReg_vd <= 5'h0;
      instReg_vl <= 12'h0;
      instVlValid <= 1'h0;
      readVS1Reg_dataValid <= 1'h0;
      readVS1Reg_requestSend <= 1'h0;
      readVS1Reg_sendToExecution <= 1'h0;
      readVS1Reg_data <= 32'h0;
      readVS1Reg_readIndex <= 4'h0;
      exeReqReg_0_valid <= 1'h0;
      exeReqReg_0_bits_source1 <= 32'h0;
      exeReqReg_0_bits_source2 <= 32'h0;
      exeReqReg_0_bits_index <= 3'h0;
      exeReqReg_0_bits_ffo <= 1'h0;
      exeReqReg_1_valid <= 1'h0;
      exeReqReg_1_bits_source1 <= 32'h0;
      exeReqReg_1_bits_source2 <= 32'h0;
      exeReqReg_1_bits_index <= 3'h0;
      exeReqReg_1_bits_ffo <= 1'h0;
      exeReqReg_2_valid <= 1'h0;
      exeReqReg_2_bits_source1 <= 32'h0;
      exeReqReg_2_bits_source2 <= 32'h0;
      exeReqReg_2_bits_index <= 3'h0;
      exeReqReg_2_bits_ffo <= 1'h0;
      exeReqReg_3_valid <= 1'h0;
      exeReqReg_3_bits_source1 <= 32'h0;
      exeReqReg_3_bits_source2 <= 32'h0;
      exeReqReg_3_bits_index <= 3'h0;
      exeReqReg_3_bits_ffo <= 1'h0;
      exeReqReg_4_valid <= 1'h0;
      exeReqReg_4_bits_source1 <= 32'h0;
      exeReqReg_4_bits_source2 <= 32'h0;
      exeReqReg_4_bits_index <= 3'h0;
      exeReqReg_4_bits_ffo <= 1'h0;
      exeReqReg_5_valid <= 1'h0;
      exeReqReg_5_bits_source1 <= 32'h0;
      exeReqReg_5_bits_source2 <= 32'h0;
      exeReqReg_5_bits_index <= 3'h0;
      exeReqReg_5_bits_ffo <= 1'h0;
      exeReqReg_6_valid <= 1'h0;
      exeReqReg_6_bits_source1 <= 32'h0;
      exeReqReg_6_bits_source2 <= 32'h0;
      exeReqReg_6_bits_index <= 3'h0;
      exeReqReg_6_bits_ffo <= 1'h0;
      exeReqReg_7_valid <= 1'h0;
      exeReqReg_7_bits_source1 <= 32'h0;
      exeReqReg_7_bits_source2 <= 32'h0;
      exeReqReg_7_bits_index <= 3'h0;
      exeReqReg_7_bits_ffo <= 1'h0;
      exeReqReg_8_valid <= 1'h0;
      exeReqReg_8_bits_source1 <= 32'h0;
      exeReqReg_8_bits_source2 <= 32'h0;
      exeReqReg_8_bits_index <= 3'h0;
      exeReqReg_8_bits_ffo <= 1'h0;
      exeReqReg_9_valid <= 1'h0;
      exeReqReg_9_bits_source1 <= 32'h0;
      exeReqReg_9_bits_source2 <= 32'h0;
      exeReqReg_9_bits_index <= 3'h0;
      exeReqReg_9_bits_ffo <= 1'h0;
      exeReqReg_10_valid <= 1'h0;
      exeReqReg_10_bits_source1 <= 32'h0;
      exeReqReg_10_bits_source2 <= 32'h0;
      exeReqReg_10_bits_index <= 3'h0;
      exeReqReg_10_bits_ffo <= 1'h0;
      exeReqReg_11_valid <= 1'h0;
      exeReqReg_11_bits_source1 <= 32'h0;
      exeReqReg_11_bits_source2 <= 32'h0;
      exeReqReg_11_bits_index <= 3'h0;
      exeReqReg_11_bits_ffo <= 1'h0;
      exeReqReg_12_valid <= 1'h0;
      exeReqReg_12_bits_source1 <= 32'h0;
      exeReqReg_12_bits_source2 <= 32'h0;
      exeReqReg_12_bits_index <= 3'h0;
      exeReqReg_12_bits_ffo <= 1'h0;
      exeReqReg_13_valid <= 1'h0;
      exeReqReg_13_bits_source1 <= 32'h0;
      exeReqReg_13_bits_source2 <= 32'h0;
      exeReqReg_13_bits_index <= 3'h0;
      exeReqReg_13_bits_ffo <= 1'h0;
      exeReqReg_14_valid <= 1'h0;
      exeReqReg_14_bits_source1 <= 32'h0;
      exeReqReg_14_bits_source2 <= 32'h0;
      exeReqReg_14_bits_index <= 3'h0;
      exeReqReg_14_bits_ffo <= 1'h0;
      exeReqReg_15_valid <= 1'h0;
      exeReqReg_15_bits_source1 <= 32'h0;
      exeReqReg_15_bits_source2 <= 32'h0;
      exeReqReg_15_bits_index <= 3'h0;
      exeReqReg_15_bits_ffo <= 1'h0;
      exeReqReg_16_valid <= 1'h0;
      exeReqReg_16_bits_source1 <= 32'h0;
      exeReqReg_16_bits_source2 <= 32'h0;
      exeReqReg_16_bits_index <= 3'h0;
      exeReqReg_16_bits_ffo <= 1'h0;
      exeReqReg_17_valid <= 1'h0;
      exeReqReg_17_bits_source1 <= 32'h0;
      exeReqReg_17_bits_source2 <= 32'h0;
      exeReqReg_17_bits_index <= 3'h0;
      exeReqReg_17_bits_ffo <= 1'h0;
      exeReqReg_18_valid <= 1'h0;
      exeReqReg_18_bits_source1 <= 32'h0;
      exeReqReg_18_bits_source2 <= 32'h0;
      exeReqReg_18_bits_index <= 3'h0;
      exeReqReg_18_bits_ffo <= 1'h0;
      exeReqReg_19_valid <= 1'h0;
      exeReqReg_19_bits_source1 <= 32'h0;
      exeReqReg_19_bits_source2 <= 32'h0;
      exeReqReg_19_bits_index <= 3'h0;
      exeReqReg_19_bits_ffo <= 1'h0;
      exeReqReg_20_valid <= 1'h0;
      exeReqReg_20_bits_source1 <= 32'h0;
      exeReqReg_20_bits_source2 <= 32'h0;
      exeReqReg_20_bits_index <= 3'h0;
      exeReqReg_20_bits_ffo <= 1'h0;
      exeReqReg_21_valid <= 1'h0;
      exeReqReg_21_bits_source1 <= 32'h0;
      exeReqReg_21_bits_source2 <= 32'h0;
      exeReqReg_21_bits_index <= 3'h0;
      exeReqReg_21_bits_ffo <= 1'h0;
      exeReqReg_22_valid <= 1'h0;
      exeReqReg_22_bits_source1 <= 32'h0;
      exeReqReg_22_bits_source2 <= 32'h0;
      exeReqReg_22_bits_index <= 3'h0;
      exeReqReg_22_bits_ffo <= 1'h0;
      exeReqReg_23_valid <= 1'h0;
      exeReqReg_23_bits_source1 <= 32'h0;
      exeReqReg_23_bits_source2 <= 32'h0;
      exeReqReg_23_bits_index <= 3'h0;
      exeReqReg_23_bits_ffo <= 1'h0;
      exeReqReg_24_valid <= 1'h0;
      exeReqReg_24_bits_source1 <= 32'h0;
      exeReqReg_24_bits_source2 <= 32'h0;
      exeReqReg_24_bits_index <= 3'h0;
      exeReqReg_24_bits_ffo <= 1'h0;
      exeReqReg_25_valid <= 1'h0;
      exeReqReg_25_bits_source1 <= 32'h0;
      exeReqReg_25_bits_source2 <= 32'h0;
      exeReqReg_25_bits_index <= 3'h0;
      exeReqReg_25_bits_ffo <= 1'h0;
      exeReqReg_26_valid <= 1'h0;
      exeReqReg_26_bits_source1 <= 32'h0;
      exeReqReg_26_bits_source2 <= 32'h0;
      exeReqReg_26_bits_index <= 3'h0;
      exeReqReg_26_bits_ffo <= 1'h0;
      exeReqReg_27_valid <= 1'h0;
      exeReqReg_27_bits_source1 <= 32'h0;
      exeReqReg_27_bits_source2 <= 32'h0;
      exeReqReg_27_bits_index <= 3'h0;
      exeReqReg_27_bits_ffo <= 1'h0;
      exeReqReg_28_valid <= 1'h0;
      exeReqReg_28_bits_source1 <= 32'h0;
      exeReqReg_28_bits_source2 <= 32'h0;
      exeReqReg_28_bits_index <= 3'h0;
      exeReqReg_28_bits_ffo <= 1'h0;
      exeReqReg_29_valid <= 1'h0;
      exeReqReg_29_bits_source1 <= 32'h0;
      exeReqReg_29_bits_source2 <= 32'h0;
      exeReqReg_29_bits_index <= 3'h0;
      exeReqReg_29_bits_ffo <= 1'h0;
      exeReqReg_30_valid <= 1'h0;
      exeReqReg_30_bits_source1 <= 32'h0;
      exeReqReg_30_bits_source2 <= 32'h0;
      exeReqReg_30_bits_index <= 3'h0;
      exeReqReg_30_bits_ffo <= 1'h0;
      exeReqReg_31_valid <= 1'h0;
      exeReqReg_31_bits_source1 <= 32'h0;
      exeReqReg_31_bits_source2 <= 32'h0;
      exeReqReg_31_bits_index <= 3'h0;
      exeReqReg_31_bits_ffo <= 1'h0;
      requestCounter <= 5'h0;
      executeIndex <= 2'h0;
      readIssueStageState_groupReadState <= 32'h0;
      readIssueStageState_needRead <= 32'h0;
      readIssueStageState_elementValid <= 32'h0;
      readIssueStageState_replaceVs1 <= 32'h0;
      readIssueStageState_readOffset <= 32'h0;
      readIssueStageState_accessLane_0 <= 5'h0;
      readIssueStageState_accessLane_1 <= 5'h0;
      readIssueStageState_accessLane_2 <= 5'h0;
      readIssueStageState_accessLane_3 <= 5'h0;
      readIssueStageState_accessLane_4 <= 5'h0;
      readIssueStageState_accessLane_5 <= 5'h0;
      readIssueStageState_accessLane_6 <= 5'h0;
      readIssueStageState_accessLane_7 <= 5'h0;
      readIssueStageState_accessLane_8 <= 5'h0;
      readIssueStageState_accessLane_9 <= 5'h0;
      readIssueStageState_accessLane_10 <= 5'h0;
      readIssueStageState_accessLane_11 <= 5'h0;
      readIssueStageState_accessLane_12 <= 5'h0;
      readIssueStageState_accessLane_13 <= 5'h0;
      readIssueStageState_accessLane_14 <= 5'h0;
      readIssueStageState_accessLane_15 <= 5'h0;
      readIssueStageState_accessLane_16 <= 5'h0;
      readIssueStageState_accessLane_17 <= 5'h0;
      readIssueStageState_accessLane_18 <= 5'h0;
      readIssueStageState_accessLane_19 <= 5'h0;
      readIssueStageState_accessLane_20 <= 5'h0;
      readIssueStageState_accessLane_21 <= 5'h0;
      readIssueStageState_accessLane_22 <= 5'h0;
      readIssueStageState_accessLane_23 <= 5'h0;
      readIssueStageState_accessLane_24 <= 5'h0;
      readIssueStageState_accessLane_25 <= 5'h0;
      readIssueStageState_accessLane_26 <= 5'h0;
      readIssueStageState_accessLane_27 <= 5'h0;
      readIssueStageState_accessLane_28 <= 5'h0;
      readIssueStageState_accessLane_29 <= 5'h0;
      readIssueStageState_accessLane_30 <= 5'h0;
      readIssueStageState_accessLane_31 <= 5'h0;
      readIssueStageState_vsGrowth_0 <= 3'h0;
      readIssueStageState_vsGrowth_1 <= 3'h0;
      readIssueStageState_vsGrowth_2 <= 3'h0;
      readIssueStageState_vsGrowth_3 <= 3'h0;
      readIssueStageState_vsGrowth_4 <= 3'h0;
      readIssueStageState_vsGrowth_5 <= 3'h0;
      readIssueStageState_vsGrowth_6 <= 3'h0;
      readIssueStageState_vsGrowth_7 <= 3'h0;
      readIssueStageState_vsGrowth_8 <= 3'h0;
      readIssueStageState_vsGrowth_9 <= 3'h0;
      readIssueStageState_vsGrowth_10 <= 3'h0;
      readIssueStageState_vsGrowth_11 <= 3'h0;
      readIssueStageState_vsGrowth_12 <= 3'h0;
      readIssueStageState_vsGrowth_13 <= 3'h0;
      readIssueStageState_vsGrowth_14 <= 3'h0;
      readIssueStageState_vsGrowth_15 <= 3'h0;
      readIssueStageState_vsGrowth_16 <= 3'h0;
      readIssueStageState_vsGrowth_17 <= 3'h0;
      readIssueStageState_vsGrowth_18 <= 3'h0;
      readIssueStageState_vsGrowth_19 <= 3'h0;
      readIssueStageState_vsGrowth_20 <= 3'h0;
      readIssueStageState_vsGrowth_21 <= 3'h0;
      readIssueStageState_vsGrowth_22 <= 3'h0;
      readIssueStageState_vsGrowth_23 <= 3'h0;
      readIssueStageState_vsGrowth_24 <= 3'h0;
      readIssueStageState_vsGrowth_25 <= 3'h0;
      readIssueStageState_vsGrowth_26 <= 3'h0;
      readIssueStageState_vsGrowth_27 <= 3'h0;
      readIssueStageState_vsGrowth_28 <= 3'h0;
      readIssueStageState_vsGrowth_29 <= 3'h0;
      readIssueStageState_vsGrowth_30 <= 3'h0;
      readIssueStageState_vsGrowth_31 <= 3'h0;
      readIssueStageState_executeGroup <= 7'h0;
      readIssueStageState_readDataOffset <= 64'h0;
      readIssueStageState_last <= 1'h0;
      readIssueStageValid <= 1'h0;
      tokenCheck_counter <= 4'h0;
      tokenCheck_counter_1 <= 4'h0;
      tokenCheck_counter_2 <= 4'h0;
      tokenCheck_counter_3 <= 4'h0;
      tokenCheck_counter_4 <= 4'h0;
      tokenCheck_counter_5 <= 4'h0;
      tokenCheck_counter_6 <= 4'h0;
      tokenCheck_counter_7 <= 4'h0;
      tokenCheck_counter_8 <= 4'h0;
      tokenCheck_counter_9 <= 4'h0;
      tokenCheck_counter_10 <= 4'h0;
      tokenCheck_counter_11 <= 4'h0;
      tokenCheck_counter_12 <= 4'h0;
      tokenCheck_counter_13 <= 4'h0;
      tokenCheck_counter_14 <= 4'h0;
      tokenCheck_counter_15 <= 4'h0;
      tokenCheck_counter_16 <= 4'h0;
      tokenCheck_counter_17 <= 4'h0;
      tokenCheck_counter_18 <= 4'h0;
      tokenCheck_counter_19 <= 4'h0;
      tokenCheck_counter_20 <= 4'h0;
      tokenCheck_counter_21 <= 4'h0;
      tokenCheck_counter_22 <= 4'h0;
      tokenCheck_counter_23 <= 4'h0;
      tokenCheck_counter_24 <= 4'h0;
      tokenCheck_counter_25 <= 4'h0;
      tokenCheck_counter_26 <= 4'h0;
      tokenCheck_counter_27 <= 4'h0;
      tokenCheck_counter_28 <= 4'h0;
      tokenCheck_counter_29 <= 4'h0;
      tokenCheck_counter_30 <= 4'h0;
      tokenCheck_counter_31 <= 4'h0;
      reorderQueueAllocate_counter <= 7'h0;
      reorderQueueAllocate_counterWillUpdate <= 7'h0;
      reorderQueueAllocate_counter_1 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_1 <= 7'h0;
      reorderQueueAllocate_counter_2 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_2 <= 7'h0;
      reorderQueueAllocate_counter_3 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_3 <= 7'h0;
      reorderQueueAllocate_counter_4 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_4 <= 7'h0;
      reorderQueueAllocate_counter_5 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_5 <= 7'h0;
      reorderQueueAllocate_counter_6 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_6 <= 7'h0;
      reorderQueueAllocate_counter_7 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_7 <= 7'h0;
      reorderQueueAllocate_counter_8 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_8 <= 7'h0;
      reorderQueueAllocate_counter_9 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_9 <= 7'h0;
      reorderQueueAllocate_counter_10 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_10 <= 7'h0;
      reorderQueueAllocate_counter_11 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_11 <= 7'h0;
      reorderQueueAllocate_counter_12 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_12 <= 7'h0;
      reorderQueueAllocate_counter_13 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_13 <= 7'h0;
      reorderQueueAllocate_counter_14 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_14 <= 7'h0;
      reorderQueueAllocate_counter_15 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_15 <= 7'h0;
      reorderQueueAllocate_counter_16 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_16 <= 7'h0;
      reorderQueueAllocate_counter_17 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_17 <= 7'h0;
      reorderQueueAllocate_counter_18 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_18 <= 7'h0;
      reorderQueueAllocate_counter_19 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_19 <= 7'h0;
      reorderQueueAllocate_counter_20 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_20 <= 7'h0;
      reorderQueueAllocate_counter_21 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_21 <= 7'h0;
      reorderQueueAllocate_counter_22 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_22 <= 7'h0;
      reorderQueueAllocate_counter_23 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_23 <= 7'h0;
      reorderQueueAllocate_counter_24 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_24 <= 7'h0;
      reorderQueueAllocate_counter_25 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_25 <= 7'h0;
      reorderQueueAllocate_counter_26 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_26 <= 7'h0;
      reorderQueueAllocate_counter_27 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_27 <= 7'h0;
      reorderQueueAllocate_counter_28 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_28 <= 7'h0;
      reorderQueueAllocate_counter_29 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_29 <= 7'h0;
      reorderQueueAllocate_counter_30 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_30 <= 7'h0;
      reorderQueueAllocate_counter_31 <= 7'h0;
      reorderQueueAllocate_counterWillUpdate_31 <= 7'h0;
      reorderStageValid <= 1'h0;
      reorderStageState_0 <= 6'h0;
      reorderStageState_1 <= 6'h0;
      reorderStageState_2 <= 6'h0;
      reorderStageState_3 <= 6'h0;
      reorderStageState_4 <= 6'h0;
      reorderStageState_5 <= 6'h0;
      reorderStageState_6 <= 6'h0;
      reorderStageState_7 <= 6'h0;
      reorderStageState_8 <= 6'h0;
      reorderStageState_9 <= 6'h0;
      reorderStageState_10 <= 6'h0;
      reorderStageState_11 <= 6'h0;
      reorderStageState_12 <= 6'h0;
      reorderStageState_13 <= 6'h0;
      reorderStageState_14 <= 6'h0;
      reorderStageState_15 <= 6'h0;
      reorderStageState_16 <= 6'h0;
      reorderStageState_17 <= 6'h0;
      reorderStageState_18 <= 6'h0;
      reorderStageState_19 <= 6'h0;
      reorderStageState_20 <= 6'h0;
      reorderStageState_21 <= 6'h0;
      reorderStageState_22 <= 6'h0;
      reorderStageState_23 <= 6'h0;
      reorderStageState_24 <= 6'h0;
      reorderStageState_25 <= 6'h0;
      reorderStageState_26 <= 6'h0;
      reorderStageState_27 <= 6'h0;
      reorderStageState_28 <= 6'h0;
      reorderStageState_29 <= 6'h0;
      reorderStageState_30 <= 6'h0;
      reorderStageState_31 <= 6'h0;
      reorderStageNeed_0 <= 6'h0;
      reorderStageNeed_1 <= 6'h0;
      reorderStageNeed_2 <= 6'h0;
      reorderStageNeed_3 <= 6'h0;
      reorderStageNeed_4 <= 6'h0;
      reorderStageNeed_5 <= 6'h0;
      reorderStageNeed_6 <= 6'h0;
      reorderStageNeed_7 <= 6'h0;
      reorderStageNeed_8 <= 6'h0;
      reorderStageNeed_9 <= 6'h0;
      reorderStageNeed_10 <= 6'h0;
      reorderStageNeed_11 <= 6'h0;
      reorderStageNeed_12 <= 6'h0;
      reorderStageNeed_13 <= 6'h0;
      reorderStageNeed_14 <= 6'h0;
      reorderStageNeed_15 <= 6'h0;
      reorderStageNeed_16 <= 6'h0;
      reorderStageNeed_17 <= 6'h0;
      reorderStageNeed_18 <= 6'h0;
      reorderStageNeed_19 <= 6'h0;
      reorderStageNeed_20 <= 6'h0;
      reorderStageNeed_21 <= 6'h0;
      reorderStageNeed_22 <= 6'h0;
      reorderStageNeed_23 <= 6'h0;
      reorderStageNeed_24 <= 6'h0;
      reorderStageNeed_25 <= 6'h0;
      reorderStageNeed_26 <= 6'h0;
      reorderStageNeed_27 <= 6'h0;
      reorderStageNeed_28 <= 6'h0;
      reorderStageNeed_29 <= 6'h0;
      reorderStageNeed_30 <= 6'h0;
      reorderStageNeed_31 <= 6'h0;
      waiteReadDataPipeReg_executeGroup <= 7'h0;
      waiteReadDataPipeReg_sourceValid <= 32'h0;
      waiteReadDataPipeReg_replaceVs1 <= 32'h0;
      waiteReadDataPipeReg_needRead <= 32'h0;
      waiteReadDataPipeReg_last <= 1'h0;
      waiteReadData_0 <= 32'h0;
      waiteReadData_1 <= 32'h0;
      waiteReadData_2 <= 32'h0;
      waiteReadData_3 <= 32'h0;
      waiteReadData_4 <= 32'h0;
      waiteReadData_5 <= 32'h0;
      waiteReadData_6 <= 32'h0;
      waiteReadData_7 <= 32'h0;
      waiteReadData_8 <= 32'h0;
      waiteReadData_9 <= 32'h0;
      waiteReadData_10 <= 32'h0;
      waiteReadData_11 <= 32'h0;
      waiteReadData_12 <= 32'h0;
      waiteReadData_13 <= 32'h0;
      waiteReadData_14 <= 32'h0;
      waiteReadData_15 <= 32'h0;
      waiteReadData_16 <= 32'h0;
      waiteReadData_17 <= 32'h0;
      waiteReadData_18 <= 32'h0;
      waiteReadData_19 <= 32'h0;
      waiteReadData_20 <= 32'h0;
      waiteReadData_21 <= 32'h0;
      waiteReadData_22 <= 32'h0;
      waiteReadData_23 <= 32'h0;
      waiteReadData_24 <= 32'h0;
      waiteReadData_25 <= 32'h0;
      waiteReadData_26 <= 32'h0;
      waiteReadData_27 <= 32'h0;
      waiteReadData_28 <= 32'h0;
      waiteReadData_29 <= 32'h0;
      waiteReadData_30 <= 32'h0;
      waiteReadData_31 <= 32'h0;
      waiteReadSate <= 32'h0;
      waiteReadStageValid <= 1'h0;
      dataNotInShifter_writeTokenCounter <= 3'h0;
      dataNotInShifter_writeTokenCounter_1 <= 3'h0;
      dataNotInShifter_writeTokenCounter_2 <= 3'h0;
      dataNotInShifter_writeTokenCounter_3 <= 3'h0;
      dataNotInShifter_writeTokenCounter_4 <= 3'h0;
      dataNotInShifter_writeTokenCounter_5 <= 3'h0;
      dataNotInShifter_writeTokenCounter_6 <= 3'h0;
      dataNotInShifter_writeTokenCounter_7 <= 3'h0;
      dataNotInShifter_writeTokenCounter_8 <= 3'h0;
      dataNotInShifter_writeTokenCounter_9 <= 3'h0;
      dataNotInShifter_writeTokenCounter_10 <= 3'h0;
      dataNotInShifter_writeTokenCounter_11 <= 3'h0;
      dataNotInShifter_writeTokenCounter_12 <= 3'h0;
      dataNotInShifter_writeTokenCounter_13 <= 3'h0;
      dataNotInShifter_writeTokenCounter_14 <= 3'h0;
      dataNotInShifter_writeTokenCounter_15 <= 3'h0;
      dataNotInShifter_writeTokenCounter_16 <= 3'h0;
      dataNotInShifter_writeTokenCounter_17 <= 3'h0;
      dataNotInShifter_writeTokenCounter_18 <= 3'h0;
      dataNotInShifter_writeTokenCounter_19 <= 3'h0;
      dataNotInShifter_writeTokenCounter_20 <= 3'h0;
      dataNotInShifter_writeTokenCounter_21 <= 3'h0;
      dataNotInShifter_writeTokenCounter_22 <= 3'h0;
      dataNotInShifter_writeTokenCounter_23 <= 3'h0;
      dataNotInShifter_writeTokenCounter_24 <= 3'h0;
      dataNotInShifter_writeTokenCounter_25 <= 3'h0;
      dataNotInShifter_writeTokenCounter_26 <= 3'h0;
      dataNotInShifter_writeTokenCounter_27 <= 3'h0;
      dataNotInShifter_writeTokenCounter_28 <= 3'h0;
      dataNotInShifter_writeTokenCounter_29 <= 3'h0;
      dataNotInShifter_writeTokenCounter_30 <= 3'h0;
      dataNotInShifter_writeTokenCounter_31 <= 3'h0;
      waiteLastRequest <= 1'h0;
      waitQueueClear <= 1'h0;
    end
    else begin
      automatic logic _GEN_171 = instReq_valid & (viotaReq | enqMvRD) | gatherRequestFire;
      automatic logic _GEN_172;
      automatic logic _GEN_173 = source1Change & viotaCounterAdd;
      _GEN_172 = instReq_valid | gatherRequestFire;
      if (v0UpdateVec_0_valid & ~v0UpdateVec_0_bits_offset)
        v0_0 <= v0_0 & ~maskExt | maskExt & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & ~v0UpdateVec_1_bits_offset)
        v0_1 <= v0_1 & ~maskExt_1 | maskExt_1 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & ~v0UpdateVec_2_bits_offset)
        v0_2 <= v0_2 & ~maskExt_2 | maskExt_2 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & ~v0UpdateVec_3_bits_offset)
        v0_3 <= v0_3 & ~maskExt_3 | maskExt_3 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_4_valid & ~v0UpdateVec_4_bits_offset)
        v0_4 <= v0_4 & ~maskExt_4 | maskExt_4 & v0UpdateVec_4_bits_data;
      if (v0UpdateVec_5_valid & ~v0UpdateVec_5_bits_offset)
        v0_5 <= v0_5 & ~maskExt_5 | maskExt_5 & v0UpdateVec_5_bits_data;
      if (v0UpdateVec_6_valid & ~v0UpdateVec_6_bits_offset)
        v0_6 <= v0_6 & ~maskExt_6 | maskExt_6 & v0UpdateVec_6_bits_data;
      if (v0UpdateVec_7_valid & ~v0UpdateVec_7_bits_offset)
        v0_7 <= v0_7 & ~maskExt_7 | maskExt_7 & v0UpdateVec_7_bits_data;
      if (v0UpdateVec_8_valid & ~v0UpdateVec_8_bits_offset)
        v0_8 <= v0_8 & ~maskExt_8 | maskExt_8 & v0UpdateVec_8_bits_data;
      if (v0UpdateVec_9_valid & ~v0UpdateVec_9_bits_offset)
        v0_9 <= v0_9 & ~maskExt_9 | maskExt_9 & v0UpdateVec_9_bits_data;
      if (v0UpdateVec_10_valid & ~v0UpdateVec_10_bits_offset)
        v0_10 <= v0_10 & ~maskExt_10 | maskExt_10 & v0UpdateVec_10_bits_data;
      if (v0UpdateVec_11_valid & ~v0UpdateVec_11_bits_offset)
        v0_11 <= v0_11 & ~maskExt_11 | maskExt_11 & v0UpdateVec_11_bits_data;
      if (v0UpdateVec_12_valid & ~v0UpdateVec_12_bits_offset)
        v0_12 <= v0_12 & ~maskExt_12 | maskExt_12 & v0UpdateVec_12_bits_data;
      if (v0UpdateVec_13_valid & ~v0UpdateVec_13_bits_offset)
        v0_13 <= v0_13 & ~maskExt_13 | maskExt_13 & v0UpdateVec_13_bits_data;
      if (v0UpdateVec_14_valid & ~v0UpdateVec_14_bits_offset)
        v0_14 <= v0_14 & ~maskExt_14 | maskExt_14 & v0UpdateVec_14_bits_data;
      if (v0UpdateVec_15_valid & ~v0UpdateVec_15_bits_offset)
        v0_15 <= v0_15 & ~maskExt_15 | maskExt_15 & v0UpdateVec_15_bits_data;
      if (v0UpdateVec_16_valid & ~v0UpdateVec_16_bits_offset)
        v0_16 <= v0_16 & ~maskExt_16 | maskExt_16 & v0UpdateVec_16_bits_data;
      if (v0UpdateVec_17_valid & ~v0UpdateVec_17_bits_offset)
        v0_17 <= v0_17 & ~maskExt_17 | maskExt_17 & v0UpdateVec_17_bits_data;
      if (v0UpdateVec_18_valid & ~v0UpdateVec_18_bits_offset)
        v0_18 <= v0_18 & ~maskExt_18 | maskExt_18 & v0UpdateVec_18_bits_data;
      if (v0UpdateVec_19_valid & ~v0UpdateVec_19_bits_offset)
        v0_19 <= v0_19 & ~maskExt_19 | maskExt_19 & v0UpdateVec_19_bits_data;
      if (v0UpdateVec_20_valid & ~v0UpdateVec_20_bits_offset)
        v0_20 <= v0_20 & ~maskExt_20 | maskExt_20 & v0UpdateVec_20_bits_data;
      if (v0UpdateVec_21_valid & ~v0UpdateVec_21_bits_offset)
        v0_21 <= v0_21 & ~maskExt_21 | maskExt_21 & v0UpdateVec_21_bits_data;
      if (v0UpdateVec_22_valid & ~v0UpdateVec_22_bits_offset)
        v0_22 <= v0_22 & ~maskExt_22 | maskExt_22 & v0UpdateVec_22_bits_data;
      if (v0UpdateVec_23_valid & ~v0UpdateVec_23_bits_offset)
        v0_23 <= v0_23 & ~maskExt_23 | maskExt_23 & v0UpdateVec_23_bits_data;
      if (v0UpdateVec_24_valid & ~v0UpdateVec_24_bits_offset)
        v0_24 <= v0_24 & ~maskExt_24 | maskExt_24 & v0UpdateVec_24_bits_data;
      if (v0UpdateVec_25_valid & ~v0UpdateVec_25_bits_offset)
        v0_25 <= v0_25 & ~maskExt_25 | maskExt_25 & v0UpdateVec_25_bits_data;
      if (v0UpdateVec_26_valid & ~v0UpdateVec_26_bits_offset)
        v0_26 <= v0_26 & ~maskExt_26 | maskExt_26 & v0UpdateVec_26_bits_data;
      if (v0UpdateVec_27_valid & ~v0UpdateVec_27_bits_offset)
        v0_27 <= v0_27 & ~maskExt_27 | maskExt_27 & v0UpdateVec_27_bits_data;
      if (v0UpdateVec_28_valid & ~v0UpdateVec_28_bits_offset)
        v0_28 <= v0_28 & ~maskExt_28 | maskExt_28 & v0UpdateVec_28_bits_data;
      if (v0UpdateVec_29_valid & ~v0UpdateVec_29_bits_offset)
        v0_29 <= v0_29 & ~maskExt_29 | maskExt_29 & v0UpdateVec_29_bits_data;
      if (v0UpdateVec_30_valid & ~v0UpdateVec_30_bits_offset)
        v0_30 <= v0_30 & ~maskExt_30 | maskExt_30 & v0UpdateVec_30_bits_data;
      if (v0UpdateVec_31_valid & ~v0UpdateVec_31_bits_offset)
        v0_31 <= v0_31 & ~maskExt_31 | maskExt_31 & v0UpdateVec_31_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset)
        v0_32 <= v0_32 & ~maskExt_32 | maskExt_32 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset)
        v0_33 <= v0_33 & ~maskExt_33 | maskExt_33 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset)
        v0_34 <= v0_34 & ~maskExt_34 | maskExt_34 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset)
        v0_35 <= v0_35 & ~maskExt_35 | maskExt_35 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_4_valid & v0UpdateVec_4_bits_offset)
        v0_36 <= v0_36 & ~maskExt_36 | maskExt_36 & v0UpdateVec_4_bits_data;
      if (v0UpdateVec_5_valid & v0UpdateVec_5_bits_offset)
        v0_37 <= v0_37 & ~maskExt_37 | maskExt_37 & v0UpdateVec_5_bits_data;
      if (v0UpdateVec_6_valid & v0UpdateVec_6_bits_offset)
        v0_38 <= v0_38 & ~maskExt_38 | maskExt_38 & v0UpdateVec_6_bits_data;
      if (v0UpdateVec_7_valid & v0UpdateVec_7_bits_offset)
        v0_39 <= v0_39 & ~maskExt_39 | maskExt_39 & v0UpdateVec_7_bits_data;
      if (v0UpdateVec_8_valid & v0UpdateVec_8_bits_offset)
        v0_40 <= v0_40 & ~maskExt_40 | maskExt_40 & v0UpdateVec_8_bits_data;
      if (v0UpdateVec_9_valid & v0UpdateVec_9_bits_offset)
        v0_41 <= v0_41 & ~maskExt_41 | maskExt_41 & v0UpdateVec_9_bits_data;
      if (v0UpdateVec_10_valid & v0UpdateVec_10_bits_offset)
        v0_42 <= v0_42 & ~maskExt_42 | maskExt_42 & v0UpdateVec_10_bits_data;
      if (v0UpdateVec_11_valid & v0UpdateVec_11_bits_offset)
        v0_43 <= v0_43 & ~maskExt_43 | maskExt_43 & v0UpdateVec_11_bits_data;
      if (v0UpdateVec_12_valid & v0UpdateVec_12_bits_offset)
        v0_44 <= v0_44 & ~maskExt_44 | maskExt_44 & v0UpdateVec_12_bits_data;
      if (v0UpdateVec_13_valid & v0UpdateVec_13_bits_offset)
        v0_45 <= v0_45 & ~maskExt_45 | maskExt_45 & v0UpdateVec_13_bits_data;
      if (v0UpdateVec_14_valid & v0UpdateVec_14_bits_offset)
        v0_46 <= v0_46 & ~maskExt_46 | maskExt_46 & v0UpdateVec_14_bits_data;
      if (v0UpdateVec_15_valid & v0UpdateVec_15_bits_offset)
        v0_47 <= v0_47 & ~maskExt_47 | maskExt_47 & v0UpdateVec_15_bits_data;
      if (v0UpdateVec_16_valid & v0UpdateVec_16_bits_offset)
        v0_48 <= v0_48 & ~maskExt_48 | maskExt_48 & v0UpdateVec_16_bits_data;
      if (v0UpdateVec_17_valid & v0UpdateVec_17_bits_offset)
        v0_49 <= v0_49 & ~maskExt_49 | maskExt_49 & v0UpdateVec_17_bits_data;
      if (v0UpdateVec_18_valid & v0UpdateVec_18_bits_offset)
        v0_50 <= v0_50 & ~maskExt_50 | maskExt_50 & v0UpdateVec_18_bits_data;
      if (v0UpdateVec_19_valid & v0UpdateVec_19_bits_offset)
        v0_51 <= v0_51 & ~maskExt_51 | maskExt_51 & v0UpdateVec_19_bits_data;
      if (v0UpdateVec_20_valid & v0UpdateVec_20_bits_offset)
        v0_52 <= v0_52 & ~maskExt_52 | maskExt_52 & v0UpdateVec_20_bits_data;
      if (v0UpdateVec_21_valid & v0UpdateVec_21_bits_offset)
        v0_53 <= v0_53 & ~maskExt_53 | maskExt_53 & v0UpdateVec_21_bits_data;
      if (v0UpdateVec_22_valid & v0UpdateVec_22_bits_offset)
        v0_54 <= v0_54 & ~maskExt_54 | maskExt_54 & v0UpdateVec_22_bits_data;
      if (v0UpdateVec_23_valid & v0UpdateVec_23_bits_offset)
        v0_55 <= v0_55 & ~maskExt_55 | maskExt_55 & v0UpdateVec_23_bits_data;
      if (v0UpdateVec_24_valid & v0UpdateVec_24_bits_offset)
        v0_56 <= v0_56 & ~maskExt_56 | maskExt_56 & v0UpdateVec_24_bits_data;
      if (v0UpdateVec_25_valid & v0UpdateVec_25_bits_offset)
        v0_57 <= v0_57 & ~maskExt_57 | maskExt_57 & v0UpdateVec_25_bits_data;
      if (v0UpdateVec_26_valid & v0UpdateVec_26_bits_offset)
        v0_58 <= v0_58 & ~maskExt_58 | maskExt_58 & v0UpdateVec_26_bits_data;
      if (v0UpdateVec_27_valid & v0UpdateVec_27_bits_offset)
        v0_59 <= v0_59 & ~maskExt_59 | maskExt_59 & v0UpdateVec_27_bits_data;
      if (v0UpdateVec_28_valid & v0UpdateVec_28_bits_offset)
        v0_60 <= v0_60 & ~maskExt_60 | maskExt_60 & v0UpdateVec_28_bits_data;
      if (v0UpdateVec_29_valid & v0UpdateVec_29_bits_offset)
        v0_61 <= v0_61 & ~maskExt_61 | maskExt_61 & v0UpdateVec_29_bits_data;
      if (v0UpdateVec_30_valid & v0UpdateVec_30_bits_offset)
        v0_62 <= v0_62 & ~maskExt_62 | maskExt_62 & v0UpdateVec_30_bits_data;
      if (v0UpdateVec_31_valid & v0UpdateVec_31_bits_offset)
        v0_63 <= v0_63 & ~maskExt_63 | maskExt_63 & v0UpdateVec_31_bits_data;
      if (gatherData_ready_0 & gatherData_valid_0)
        gatherReadState <= 2'h0;
      else if (_tokenCheck_T & gatherSRead)
        gatherReadState <= 2'h2;
      else if (gatherRequestFire)
        gatherReadState <= {notNeedRead, 1'h1};
      else if (readTokenRelease_0 & gatherWaiteRead)
        gatherReadState <= 2'h3;
      if (gatherRequestFire) begin
        gatherDatOffset <= dataOffset;
        gatherLane <= accessLane;
        gatherOffset <= offset;
        gatherGrowth <= reallyGrowth;
      end
      if (_GEN_171 | instReq_valid)
        instReg_instructionIndex <= instReq_bits_instructionIndex;
      if (instReq_valid) begin
        instReg_decodeResult_specialSlot <= instReq_bits_decodeResult_specialSlot;
        instReg_decodeResult_topUop <= instReq_bits_decodeResult_topUop;
        instReg_decodeResult_popCount <= instReq_bits_decodeResult_popCount;
        instReg_decodeResult_ffo <= instReq_bits_decodeResult_ffo;
        instReg_decodeResult_average <= instReq_bits_decodeResult_average;
        instReg_decodeResult_reverse <= instReq_bits_decodeResult_reverse;
        instReg_decodeResult_dontNeedExecuteInLane <= instReq_bits_decodeResult_dontNeedExecuteInLane;
        instReg_decodeResult_scheduler <= instReq_bits_decodeResult_scheduler;
        instReg_decodeResult_sReadVD <= instReq_bits_decodeResult_sReadVD;
        instReg_decodeResult_vtype <= instReq_bits_decodeResult_vtype;
        instReg_decodeResult_sWrite <= instReq_bits_decodeResult_sWrite;
        instReg_decodeResult_crossRead <= instReq_bits_decodeResult_crossRead;
        instReg_decodeResult_crossWrite <= instReq_bits_decodeResult_crossWrite;
        instReg_decodeResult_maskUnit <= instReq_bits_decodeResult_maskUnit;
        instReg_decodeResult_special <= instReq_bits_decodeResult_special;
        instReg_decodeResult_saturate <= instReq_bits_decodeResult_saturate;
        instReg_decodeResult_vwmacc <= instReq_bits_decodeResult_vwmacc;
        instReg_decodeResult_readOnly <= instReq_bits_decodeResult_readOnly;
        instReg_decodeResult_maskSource <= instReq_bits_decodeResult_maskSource;
        instReg_decodeResult_maskDestination <= instReq_bits_decodeResult_maskDestination;
        instReg_decodeResult_maskLogic <= instReq_bits_decodeResult_maskLogic;
        instReg_decodeResult_uop <= instReq_bits_decodeResult_uop;
        instReg_decodeResult_iota <= instReq_bits_decodeResult_iota;
        instReg_decodeResult_mv <= instReq_bits_decodeResult_mv;
        instReg_decodeResult_extend <= instReq_bits_decodeResult_extend;
        instReg_decodeResult_unOrderWrite <= instReq_bits_decodeResult_unOrderWrite;
        instReg_decodeResult_compress <= instReq_bits_decodeResult_compress;
        instReg_decodeResult_gather16 <= instReq_bits_decodeResult_gather16;
        instReg_decodeResult_gather <= instReq_bits_decodeResult_gather;
        instReg_decodeResult_slid <= instReq_bits_decodeResult_slid;
        instReg_decodeResult_targetRd <= instReq_bits_decodeResult_targetRd;
        instReg_decodeResult_widenReduce <= instReq_bits_decodeResult_widenReduce;
        instReg_decodeResult_red <= instReq_bits_decodeResult_red;
        instReg_decodeResult_nr <= instReq_bits_decodeResult_nr;
        instReg_decodeResult_itype <= instReq_bits_decodeResult_itype;
        instReg_decodeResult_unsigned1 <= instReq_bits_decodeResult_unsigned1;
        instReg_decodeResult_unsigned0 <= instReq_bits_decodeResult_unsigned0;
        instReg_decodeResult_other <= instReq_bits_decodeResult_other;
        instReg_decodeResult_multiCycle <= instReq_bits_decodeResult_multiCycle;
        instReg_decodeResult_divider <= instReq_bits_decodeResult_divider;
        instReg_decodeResult_multiplier <= instReq_bits_decodeResult_multiplier;
        instReg_decodeResult_shift <= instReq_bits_decodeResult_shift;
        instReg_decodeResult_adder <= instReq_bits_decodeResult_adder;
        instReg_decodeResult_logic <= instReq_bits_decodeResult_logic;
        instReg_readFromScala <= instReq_bits_readFromScala;
        instReg_sew <= instReq_bits_sew;
        instReg_vlmul <= instReq_bits_vlmul;
        instReg_maskType <= instReq_bits_maskType;
        instReg_vxrm <= instReq_bits_vxrm;
        instReg_vs2 <= instReq_bits_vs2;
        instReg_vd <= instReq_bits_vd;
        instReg_vl <= instReq_bits_vl;
      end
      if (_GEN_171)
        instReg_vs1 <= instReq_bits_vs2;
      else if (instReq_valid)
        instReg_vs1 <= instReq_bits_vs1;
      if (|{instReq_valid, _lastReport_output})
        instVlValid <= ((|instReq_bits_vl) | enqMvRD) & instReq_valid;
      readVS1Reg_dataValid <= ~_GEN_173 & (readTokenRelease_0 | ~_GEN_172 & readVS1Reg_dataValid);
      readVS1Reg_requestSend <= ~_GEN_173 & (_tokenCheck_T | ~_GEN_172 & readVS1Reg_requestSend);
      readVS1Reg_sendToExecution <= _view__firstGroup_T_1 | viotaCounterAdd | ~_GEN_172 & readVS1Reg_sendToExecution;
      if (readTokenRelease_0) begin
        readVS1Reg_data <= readData_readDataQueue_deq_bits;
        waiteReadData_0 <= readData_readDataQueue_deq_bits;
      end
      if (_GEN_173)
        readVS1Reg_readIndex <= readVS1Reg_readIndex + 4'h1;
      else if (_GEN_172)
        readVS1Reg_readIndex <= 4'h0;
      if (tokenIO_0_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_0_valid <= tokenIO_0_maskRequestRelease_0 & ~viota;
      if (tokenIO_0_maskRequestRelease_0) begin
        exeReqReg_0_bits_source1 <= exeRequestQueue_0_deq_bits_source1;
        exeReqReg_0_bits_source2 <= exeRequestQueue_0_deq_bits_source2;
        exeReqReg_0_bits_index <= exeRequestQueue_0_deq_bits_index;
        exeReqReg_0_bits_ffo <= exeRequestQueue_0_deq_bits_ffo;
      end
      if (tokenIO_1_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_1_valid <= tokenIO_1_maskRequestRelease_0 & ~viota;
      if (tokenIO_1_maskRequestRelease_0) begin
        exeReqReg_1_bits_source1 <= exeRequestQueue_1_deq_bits_source1;
        exeReqReg_1_bits_source2 <= exeRequestQueue_1_deq_bits_source2;
        exeReqReg_1_bits_index <= exeRequestQueue_1_deq_bits_index;
        exeReqReg_1_bits_ffo <= exeRequestQueue_1_deq_bits_ffo;
      end
      if (tokenIO_2_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_2_valid <= tokenIO_2_maskRequestRelease_0 & ~viota;
      if (tokenIO_2_maskRequestRelease_0) begin
        exeReqReg_2_bits_source1 <= exeRequestQueue_2_deq_bits_source1;
        exeReqReg_2_bits_source2 <= exeRequestQueue_2_deq_bits_source2;
        exeReqReg_2_bits_index <= exeRequestQueue_2_deq_bits_index;
        exeReqReg_2_bits_ffo <= exeRequestQueue_2_deq_bits_ffo;
      end
      if (tokenIO_3_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_3_valid <= tokenIO_3_maskRequestRelease_0 & ~viota;
      if (tokenIO_3_maskRequestRelease_0) begin
        exeReqReg_3_bits_source1 <= exeRequestQueue_3_deq_bits_source1;
        exeReqReg_3_bits_source2 <= exeRequestQueue_3_deq_bits_source2;
        exeReqReg_3_bits_index <= exeRequestQueue_3_deq_bits_index;
        exeReqReg_3_bits_ffo <= exeRequestQueue_3_deq_bits_ffo;
      end
      if (tokenIO_4_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_4_valid <= tokenIO_4_maskRequestRelease_0 & ~viota;
      if (tokenIO_4_maskRequestRelease_0) begin
        exeReqReg_4_bits_source1 <= exeRequestQueue_4_deq_bits_source1;
        exeReqReg_4_bits_source2 <= exeRequestQueue_4_deq_bits_source2;
        exeReqReg_4_bits_index <= exeRequestQueue_4_deq_bits_index;
        exeReqReg_4_bits_ffo <= exeRequestQueue_4_deq_bits_ffo;
      end
      if (tokenIO_5_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_5_valid <= tokenIO_5_maskRequestRelease_0 & ~viota;
      if (tokenIO_5_maskRequestRelease_0) begin
        exeReqReg_5_bits_source1 <= exeRequestQueue_5_deq_bits_source1;
        exeReqReg_5_bits_source2 <= exeRequestQueue_5_deq_bits_source2;
        exeReqReg_5_bits_index <= exeRequestQueue_5_deq_bits_index;
        exeReqReg_5_bits_ffo <= exeRequestQueue_5_deq_bits_ffo;
      end
      if (tokenIO_6_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_6_valid <= tokenIO_6_maskRequestRelease_0 & ~viota;
      if (tokenIO_6_maskRequestRelease_0) begin
        exeReqReg_6_bits_source1 <= exeRequestQueue_6_deq_bits_source1;
        exeReqReg_6_bits_source2 <= exeRequestQueue_6_deq_bits_source2;
        exeReqReg_6_bits_index <= exeRequestQueue_6_deq_bits_index;
        exeReqReg_6_bits_ffo <= exeRequestQueue_6_deq_bits_ffo;
      end
      if (tokenIO_7_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_7_valid <= tokenIO_7_maskRequestRelease_0 & ~viota;
      if (tokenIO_7_maskRequestRelease_0) begin
        exeReqReg_7_bits_source1 <= exeRequestQueue_7_deq_bits_source1;
        exeReqReg_7_bits_source2 <= exeRequestQueue_7_deq_bits_source2;
        exeReqReg_7_bits_index <= exeRequestQueue_7_deq_bits_index;
        exeReqReg_7_bits_ffo <= exeRequestQueue_7_deq_bits_ffo;
      end
      if (tokenIO_8_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_8_valid <= tokenIO_8_maskRequestRelease_0 & ~viota;
      if (tokenIO_8_maskRequestRelease_0) begin
        exeReqReg_8_bits_source1 <= exeRequestQueue_8_deq_bits_source1;
        exeReqReg_8_bits_source2 <= exeRequestQueue_8_deq_bits_source2;
        exeReqReg_8_bits_index <= exeRequestQueue_8_deq_bits_index;
        exeReqReg_8_bits_ffo <= exeRequestQueue_8_deq_bits_ffo;
      end
      if (tokenIO_9_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_9_valid <= tokenIO_9_maskRequestRelease_0 & ~viota;
      if (tokenIO_9_maskRequestRelease_0) begin
        exeReqReg_9_bits_source1 <= exeRequestQueue_9_deq_bits_source1;
        exeReqReg_9_bits_source2 <= exeRequestQueue_9_deq_bits_source2;
        exeReqReg_9_bits_index <= exeRequestQueue_9_deq_bits_index;
        exeReqReg_9_bits_ffo <= exeRequestQueue_9_deq_bits_ffo;
      end
      if (tokenIO_10_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_10_valid <= tokenIO_10_maskRequestRelease_0 & ~viota;
      if (tokenIO_10_maskRequestRelease_0) begin
        exeReqReg_10_bits_source1 <= exeRequestQueue_10_deq_bits_source1;
        exeReqReg_10_bits_source2 <= exeRequestQueue_10_deq_bits_source2;
        exeReqReg_10_bits_index <= exeRequestQueue_10_deq_bits_index;
        exeReqReg_10_bits_ffo <= exeRequestQueue_10_deq_bits_ffo;
      end
      if (tokenIO_11_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_11_valid <= tokenIO_11_maskRequestRelease_0 & ~viota;
      if (tokenIO_11_maskRequestRelease_0) begin
        exeReqReg_11_bits_source1 <= exeRequestQueue_11_deq_bits_source1;
        exeReqReg_11_bits_source2 <= exeRequestQueue_11_deq_bits_source2;
        exeReqReg_11_bits_index <= exeRequestQueue_11_deq_bits_index;
        exeReqReg_11_bits_ffo <= exeRequestQueue_11_deq_bits_ffo;
      end
      if (tokenIO_12_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_12_valid <= tokenIO_12_maskRequestRelease_0 & ~viota;
      if (tokenIO_12_maskRequestRelease_0) begin
        exeReqReg_12_bits_source1 <= exeRequestQueue_12_deq_bits_source1;
        exeReqReg_12_bits_source2 <= exeRequestQueue_12_deq_bits_source2;
        exeReqReg_12_bits_index <= exeRequestQueue_12_deq_bits_index;
        exeReqReg_12_bits_ffo <= exeRequestQueue_12_deq_bits_ffo;
      end
      if (tokenIO_13_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_13_valid <= tokenIO_13_maskRequestRelease_0 & ~viota;
      if (tokenIO_13_maskRequestRelease_0) begin
        exeReqReg_13_bits_source1 <= exeRequestQueue_13_deq_bits_source1;
        exeReqReg_13_bits_source2 <= exeRequestQueue_13_deq_bits_source2;
        exeReqReg_13_bits_index <= exeRequestQueue_13_deq_bits_index;
        exeReqReg_13_bits_ffo <= exeRequestQueue_13_deq_bits_ffo;
      end
      if (tokenIO_14_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_14_valid <= tokenIO_14_maskRequestRelease_0 & ~viota;
      if (tokenIO_14_maskRequestRelease_0) begin
        exeReqReg_14_bits_source1 <= exeRequestQueue_14_deq_bits_source1;
        exeReqReg_14_bits_source2 <= exeRequestQueue_14_deq_bits_source2;
        exeReqReg_14_bits_index <= exeRequestQueue_14_deq_bits_index;
        exeReqReg_14_bits_ffo <= exeRequestQueue_14_deq_bits_ffo;
      end
      if (tokenIO_15_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_15_valid <= tokenIO_15_maskRequestRelease_0 & ~viota;
      if (tokenIO_15_maskRequestRelease_0) begin
        exeReqReg_15_bits_source1 <= exeRequestQueue_15_deq_bits_source1;
        exeReqReg_15_bits_source2 <= exeRequestQueue_15_deq_bits_source2;
        exeReqReg_15_bits_index <= exeRequestQueue_15_deq_bits_index;
        exeReqReg_15_bits_ffo <= exeRequestQueue_15_deq_bits_ffo;
      end
      if (tokenIO_16_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_16_valid <= tokenIO_16_maskRequestRelease_0 & ~viota;
      if (tokenIO_16_maskRequestRelease_0) begin
        exeReqReg_16_bits_source1 <= exeRequestQueue_16_deq_bits_source1;
        exeReqReg_16_bits_source2 <= exeRequestQueue_16_deq_bits_source2;
        exeReqReg_16_bits_index <= exeRequestQueue_16_deq_bits_index;
        exeReqReg_16_bits_ffo <= exeRequestQueue_16_deq_bits_ffo;
      end
      if (tokenIO_17_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_17_valid <= tokenIO_17_maskRequestRelease_0 & ~viota;
      if (tokenIO_17_maskRequestRelease_0) begin
        exeReqReg_17_bits_source1 <= exeRequestQueue_17_deq_bits_source1;
        exeReqReg_17_bits_source2 <= exeRequestQueue_17_deq_bits_source2;
        exeReqReg_17_bits_index <= exeRequestQueue_17_deq_bits_index;
        exeReqReg_17_bits_ffo <= exeRequestQueue_17_deq_bits_ffo;
      end
      if (tokenIO_18_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_18_valid <= tokenIO_18_maskRequestRelease_0 & ~viota;
      if (tokenIO_18_maskRequestRelease_0) begin
        exeReqReg_18_bits_source1 <= exeRequestQueue_18_deq_bits_source1;
        exeReqReg_18_bits_source2 <= exeRequestQueue_18_deq_bits_source2;
        exeReqReg_18_bits_index <= exeRequestQueue_18_deq_bits_index;
        exeReqReg_18_bits_ffo <= exeRequestQueue_18_deq_bits_ffo;
      end
      if (tokenIO_19_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_19_valid <= tokenIO_19_maskRequestRelease_0 & ~viota;
      if (tokenIO_19_maskRequestRelease_0) begin
        exeReqReg_19_bits_source1 <= exeRequestQueue_19_deq_bits_source1;
        exeReqReg_19_bits_source2 <= exeRequestQueue_19_deq_bits_source2;
        exeReqReg_19_bits_index <= exeRequestQueue_19_deq_bits_index;
        exeReqReg_19_bits_ffo <= exeRequestQueue_19_deq_bits_ffo;
      end
      if (tokenIO_20_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_20_valid <= tokenIO_20_maskRequestRelease_0 & ~viota;
      if (tokenIO_20_maskRequestRelease_0) begin
        exeReqReg_20_bits_source1 <= exeRequestQueue_20_deq_bits_source1;
        exeReqReg_20_bits_source2 <= exeRequestQueue_20_deq_bits_source2;
        exeReqReg_20_bits_index <= exeRequestQueue_20_deq_bits_index;
        exeReqReg_20_bits_ffo <= exeRequestQueue_20_deq_bits_ffo;
      end
      if (tokenIO_21_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_21_valid <= tokenIO_21_maskRequestRelease_0 & ~viota;
      if (tokenIO_21_maskRequestRelease_0) begin
        exeReqReg_21_bits_source1 <= exeRequestQueue_21_deq_bits_source1;
        exeReqReg_21_bits_source2 <= exeRequestQueue_21_deq_bits_source2;
        exeReqReg_21_bits_index <= exeRequestQueue_21_deq_bits_index;
        exeReqReg_21_bits_ffo <= exeRequestQueue_21_deq_bits_ffo;
      end
      if (tokenIO_22_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_22_valid <= tokenIO_22_maskRequestRelease_0 & ~viota;
      if (tokenIO_22_maskRequestRelease_0) begin
        exeReqReg_22_bits_source1 <= exeRequestQueue_22_deq_bits_source1;
        exeReqReg_22_bits_source2 <= exeRequestQueue_22_deq_bits_source2;
        exeReqReg_22_bits_index <= exeRequestQueue_22_deq_bits_index;
        exeReqReg_22_bits_ffo <= exeRequestQueue_22_deq_bits_ffo;
      end
      if (tokenIO_23_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_23_valid <= tokenIO_23_maskRequestRelease_0 & ~viota;
      if (tokenIO_23_maskRequestRelease_0) begin
        exeReqReg_23_bits_source1 <= exeRequestQueue_23_deq_bits_source1;
        exeReqReg_23_bits_source2 <= exeRequestQueue_23_deq_bits_source2;
        exeReqReg_23_bits_index <= exeRequestQueue_23_deq_bits_index;
        exeReqReg_23_bits_ffo <= exeRequestQueue_23_deq_bits_ffo;
      end
      if (tokenIO_24_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_24_valid <= tokenIO_24_maskRequestRelease_0 & ~viota;
      if (tokenIO_24_maskRequestRelease_0) begin
        exeReqReg_24_bits_source1 <= exeRequestQueue_24_deq_bits_source1;
        exeReqReg_24_bits_source2 <= exeRequestQueue_24_deq_bits_source2;
        exeReqReg_24_bits_index <= exeRequestQueue_24_deq_bits_index;
        exeReqReg_24_bits_ffo <= exeRequestQueue_24_deq_bits_ffo;
      end
      if (tokenIO_25_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_25_valid <= tokenIO_25_maskRequestRelease_0 & ~viota;
      if (tokenIO_25_maskRequestRelease_0) begin
        exeReqReg_25_bits_source1 <= exeRequestQueue_25_deq_bits_source1;
        exeReqReg_25_bits_source2 <= exeRequestQueue_25_deq_bits_source2;
        exeReqReg_25_bits_index <= exeRequestQueue_25_deq_bits_index;
        exeReqReg_25_bits_ffo <= exeRequestQueue_25_deq_bits_ffo;
      end
      if (tokenIO_26_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_26_valid <= tokenIO_26_maskRequestRelease_0 & ~viota;
      if (tokenIO_26_maskRequestRelease_0) begin
        exeReqReg_26_bits_source1 <= exeRequestQueue_26_deq_bits_source1;
        exeReqReg_26_bits_source2 <= exeRequestQueue_26_deq_bits_source2;
        exeReqReg_26_bits_index <= exeRequestQueue_26_deq_bits_index;
        exeReqReg_26_bits_ffo <= exeRequestQueue_26_deq_bits_ffo;
      end
      if (tokenIO_27_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_27_valid <= tokenIO_27_maskRequestRelease_0 & ~viota;
      if (tokenIO_27_maskRequestRelease_0) begin
        exeReqReg_27_bits_source1 <= exeRequestQueue_27_deq_bits_source1;
        exeReqReg_27_bits_source2 <= exeRequestQueue_27_deq_bits_source2;
        exeReqReg_27_bits_index <= exeRequestQueue_27_deq_bits_index;
        exeReqReg_27_bits_ffo <= exeRequestQueue_27_deq_bits_ffo;
      end
      if (tokenIO_28_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_28_valid <= tokenIO_28_maskRequestRelease_0 & ~viota;
      if (tokenIO_28_maskRequestRelease_0) begin
        exeReqReg_28_bits_source1 <= exeRequestQueue_28_deq_bits_source1;
        exeReqReg_28_bits_source2 <= exeRequestQueue_28_deq_bits_source2;
        exeReqReg_28_bits_index <= exeRequestQueue_28_deq_bits_index;
        exeReqReg_28_bits_ffo <= exeRequestQueue_28_deq_bits_ffo;
      end
      if (tokenIO_29_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_29_valid <= tokenIO_29_maskRequestRelease_0 & ~viota;
      if (tokenIO_29_maskRequestRelease_0) begin
        exeReqReg_29_bits_source1 <= exeRequestQueue_29_deq_bits_source1;
        exeReqReg_29_bits_source2 <= exeRequestQueue_29_deq_bits_source2;
        exeReqReg_29_bits_index <= exeRequestQueue_29_deq_bits_index;
        exeReqReg_29_bits_ffo <= exeRequestQueue_29_deq_bits_ffo;
      end
      if (tokenIO_30_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_30_valid <= tokenIO_30_maskRequestRelease_0 & ~viota;
      if (tokenIO_30_maskRequestRelease_0) begin
        exeReqReg_30_bits_source1 <= exeRequestQueue_30_deq_bits_source1;
        exeReqReg_30_bits_source2 <= exeRequestQueue_30_deq_bits_source2;
        exeReqReg_30_bits_index <= exeRequestQueue_30_deq_bits_index;
        exeReqReg_30_bits_ffo <= exeRequestQueue_30_deq_bits_ffo;
      end
      if (tokenIO_31_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_31_valid <= tokenIO_31_maskRequestRelease_0 & ~viota;
      if (tokenIO_31_maskRequestRelease_0) begin
        exeReqReg_31_bits_source1 <= exeRequestQueue_31_deq_bits_source1;
        exeReqReg_31_bits_source2 <= exeRequestQueue_31_deq_bits_source2;
        exeReqReg_31_bits_index <= exeRequestQueue_31_deq_bits_index;
        exeReqReg_31_bits_ffo <= exeRequestQueue_31_deq_bits_ffo;
      end
      if (instReq_valid | groupCounterAdd)
        requestCounter <= instReq_valid ? 5'h0 : requestCounter + 5'h1;
      if (requestStageDeq & anyDataValid)
        executeIndex <= executeIndex + executeIndexGrowth[1:0];
      if (readIssueStageEnq) begin
        readIssueStageState_groupReadState <= 32'h0;
        readIssueStageState_needRead <= _GEN_139 ? _slideAddressGen_indexDeq_bits_needRead : ~notReadSelect;
        readIssueStageState_elementValid <= _GEN_139 ? _slideAddressGen_indexDeq_bits_elementValid : elementValidSelect;
        readIssueStageState_replaceVs1 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_replaceVs1 : 32'h0;
        readIssueStageState_readOffset <= _GEN_139 ? _slideAddressGen_indexDeq_bits_readOffset : offsetSelect;
        readIssueStageState_accessLane_0 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_0 : accessLaneSelect[4:0];
        readIssueStageState_accessLane_1 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_1 : accessLaneSelect[9:5];
        readIssueStageState_accessLane_2 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_2 : accessLaneSelect[14:10];
        readIssueStageState_accessLane_3 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_3 : accessLaneSelect[19:15];
        readIssueStageState_accessLane_4 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_4 : accessLaneSelect[24:20];
        readIssueStageState_accessLane_5 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_5 : accessLaneSelect[29:25];
        readIssueStageState_accessLane_6 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_6 : accessLaneSelect[34:30];
        readIssueStageState_accessLane_7 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_7 : accessLaneSelect[39:35];
        readIssueStageState_accessLane_8 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_8 : accessLaneSelect[44:40];
        readIssueStageState_accessLane_9 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_9 : accessLaneSelect[49:45];
        readIssueStageState_accessLane_10 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_10 : accessLaneSelect[54:50];
        readIssueStageState_accessLane_11 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_11 : accessLaneSelect[59:55];
        readIssueStageState_accessLane_12 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_12 : accessLaneSelect[64:60];
        readIssueStageState_accessLane_13 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_13 : accessLaneSelect[69:65];
        readIssueStageState_accessLane_14 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_14 : accessLaneSelect[74:70];
        readIssueStageState_accessLane_15 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_15 : accessLaneSelect[79:75];
        readIssueStageState_accessLane_16 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_16 : accessLaneSelect[84:80];
        readIssueStageState_accessLane_17 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_17 : accessLaneSelect[89:85];
        readIssueStageState_accessLane_18 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_18 : accessLaneSelect[94:90];
        readIssueStageState_accessLane_19 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_19 : accessLaneSelect[99:95];
        readIssueStageState_accessLane_20 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_20 : accessLaneSelect[104:100];
        readIssueStageState_accessLane_21 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_21 : accessLaneSelect[109:105];
        readIssueStageState_accessLane_22 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_22 : accessLaneSelect[114:110];
        readIssueStageState_accessLane_23 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_23 : accessLaneSelect[119:115];
        readIssueStageState_accessLane_24 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_24 : accessLaneSelect[124:120];
        readIssueStageState_accessLane_25 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_25 : accessLaneSelect[129:125];
        readIssueStageState_accessLane_26 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_26 : accessLaneSelect[134:130];
        readIssueStageState_accessLane_27 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_27 : accessLaneSelect[139:135];
        readIssueStageState_accessLane_28 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_28 : accessLaneSelect[144:140];
        readIssueStageState_accessLane_29 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_29 : accessLaneSelect[149:145];
        readIssueStageState_accessLane_30 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_30 : accessLaneSelect[154:150];
        readIssueStageState_accessLane_31 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_accessLane_31 : accessLaneSelect[159:155];
        readIssueStageState_vsGrowth_0 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_0 : growthSelect[2:0];
        readIssueStageState_vsGrowth_1 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_1 : growthSelect[5:3];
        readIssueStageState_vsGrowth_2 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_2 : growthSelect[8:6];
        readIssueStageState_vsGrowth_3 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_3 : growthSelect[11:9];
        readIssueStageState_vsGrowth_4 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_4 : growthSelect[14:12];
        readIssueStageState_vsGrowth_5 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_5 : growthSelect[17:15];
        readIssueStageState_vsGrowth_6 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_6 : growthSelect[20:18];
        readIssueStageState_vsGrowth_7 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_7 : growthSelect[23:21];
        readIssueStageState_vsGrowth_8 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_8 : growthSelect[26:24];
        readIssueStageState_vsGrowth_9 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_9 : growthSelect[29:27];
        readIssueStageState_vsGrowth_10 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_10 : growthSelect[32:30];
        readIssueStageState_vsGrowth_11 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_11 : growthSelect[35:33];
        readIssueStageState_vsGrowth_12 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_12 : growthSelect[38:36];
        readIssueStageState_vsGrowth_13 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_13 : growthSelect[41:39];
        readIssueStageState_vsGrowth_14 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_14 : growthSelect[44:42];
        readIssueStageState_vsGrowth_15 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_15 : growthSelect[47:45];
        readIssueStageState_vsGrowth_16 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_16 : growthSelect[50:48];
        readIssueStageState_vsGrowth_17 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_17 : growthSelect[53:51];
        readIssueStageState_vsGrowth_18 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_18 : growthSelect[56:54];
        readIssueStageState_vsGrowth_19 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_19 : growthSelect[59:57];
        readIssueStageState_vsGrowth_20 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_20 : growthSelect[62:60];
        readIssueStageState_vsGrowth_21 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_21 : growthSelect[65:63];
        readIssueStageState_vsGrowth_22 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_22 : growthSelect[68:66];
        readIssueStageState_vsGrowth_23 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_23 : growthSelect[71:69];
        readIssueStageState_vsGrowth_24 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_24 : growthSelect[74:72];
        readIssueStageState_vsGrowth_25 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_25 : growthSelect[77:75];
        readIssueStageState_vsGrowth_26 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_26 : growthSelect[80:78];
        readIssueStageState_vsGrowth_27 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_27 : growthSelect[83:81];
        readIssueStageState_vsGrowth_28 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_28 : growthSelect[86:84];
        readIssueStageState_vsGrowth_29 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_29 : growthSelect[89:87];
        readIssueStageState_vsGrowth_30 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_30 : growthSelect[92:90];
        readIssueStageState_vsGrowth_31 <= _GEN_139 ? _slideAddressGen_indexDeq_bits_vsGrowth_31 : growthSelect[95:93];
        readIssueStageState_executeGroup <= _GEN_139 ? _slideAddressGen_indexDeq_bits_executeGroup : executeGroup;
        readIssueStageState_readDataOffset <= _GEN_139 ? _slideAddressGen_indexDeq_bits_readDataOffset : dataOffsetSelect;
        readIssueStageState_last <= _GEN_139 ? _slideAddressGen_indexDeq_bits_last : isVlBoundary;
      end
      else if (anyReadFire)
        readIssueStageState_groupReadState <= readStateUpdate;
      if (readTypeRequestDeq ^ readIssueStageEnq)
        readIssueStageValid <= readIssueStageEnq;
      if (_tokenCheck_T ^ readTokenRelease_0)
        tokenCheck_counter <= tokenCheck_counter + tokenCheck_counterChange;
      if (pipeReadFire_1 ^ readTokenRelease_1)
        tokenCheck_counter_1 <= tokenCheck_counter_1 + tokenCheck_counterChange_1;
      if (pipeReadFire_2 ^ readTokenRelease_2)
        tokenCheck_counter_2 <= tokenCheck_counter_2 + tokenCheck_counterChange_2;
      if (pipeReadFire_3 ^ readTokenRelease_3)
        tokenCheck_counter_3 <= tokenCheck_counter_3 + tokenCheck_counterChange_3;
      if (pipeReadFire_4 ^ readTokenRelease_4)
        tokenCheck_counter_4 <= tokenCheck_counter_4 + tokenCheck_counterChange_4;
      if (pipeReadFire_5 ^ readTokenRelease_5)
        tokenCheck_counter_5 <= tokenCheck_counter_5 + tokenCheck_counterChange_5;
      if (pipeReadFire_6 ^ readTokenRelease_6)
        tokenCheck_counter_6 <= tokenCheck_counter_6 + tokenCheck_counterChange_6;
      if (pipeReadFire_7 ^ readTokenRelease_7)
        tokenCheck_counter_7 <= tokenCheck_counter_7 + tokenCheck_counterChange_7;
      if (pipeReadFire_8 ^ readTokenRelease_8)
        tokenCheck_counter_8 <= tokenCheck_counter_8 + tokenCheck_counterChange_8;
      if (pipeReadFire_9 ^ readTokenRelease_9)
        tokenCheck_counter_9 <= tokenCheck_counter_9 + tokenCheck_counterChange_9;
      if (pipeReadFire_10 ^ readTokenRelease_10)
        tokenCheck_counter_10 <= tokenCheck_counter_10 + tokenCheck_counterChange_10;
      if (pipeReadFire_11 ^ readTokenRelease_11)
        tokenCheck_counter_11 <= tokenCheck_counter_11 + tokenCheck_counterChange_11;
      if (pipeReadFire_12 ^ readTokenRelease_12)
        tokenCheck_counter_12 <= tokenCheck_counter_12 + tokenCheck_counterChange_12;
      if (pipeReadFire_13 ^ readTokenRelease_13)
        tokenCheck_counter_13 <= tokenCheck_counter_13 + tokenCheck_counterChange_13;
      if (pipeReadFire_14 ^ readTokenRelease_14)
        tokenCheck_counter_14 <= tokenCheck_counter_14 + tokenCheck_counterChange_14;
      if (pipeReadFire_15 ^ readTokenRelease_15)
        tokenCheck_counter_15 <= tokenCheck_counter_15 + tokenCheck_counterChange_15;
      if (pipeReadFire_16 ^ readTokenRelease_16)
        tokenCheck_counter_16 <= tokenCheck_counter_16 + tokenCheck_counterChange_16;
      if (pipeReadFire_17 ^ readTokenRelease_17)
        tokenCheck_counter_17 <= tokenCheck_counter_17 + tokenCheck_counterChange_17;
      if (pipeReadFire_18 ^ readTokenRelease_18)
        tokenCheck_counter_18 <= tokenCheck_counter_18 + tokenCheck_counterChange_18;
      if (pipeReadFire_19 ^ readTokenRelease_19)
        tokenCheck_counter_19 <= tokenCheck_counter_19 + tokenCheck_counterChange_19;
      if (pipeReadFire_20 ^ readTokenRelease_20)
        tokenCheck_counter_20 <= tokenCheck_counter_20 + tokenCheck_counterChange_20;
      if (pipeReadFire_21 ^ readTokenRelease_21)
        tokenCheck_counter_21 <= tokenCheck_counter_21 + tokenCheck_counterChange_21;
      if (pipeReadFire_22 ^ readTokenRelease_22)
        tokenCheck_counter_22 <= tokenCheck_counter_22 + tokenCheck_counterChange_22;
      if (pipeReadFire_23 ^ readTokenRelease_23)
        tokenCheck_counter_23 <= tokenCheck_counter_23 + tokenCheck_counterChange_23;
      if (pipeReadFire_24 ^ readTokenRelease_24)
        tokenCheck_counter_24 <= tokenCheck_counter_24 + tokenCheck_counterChange_24;
      if (pipeReadFire_25 ^ readTokenRelease_25)
        tokenCheck_counter_25 <= tokenCheck_counter_25 + tokenCheck_counterChange_25;
      if (pipeReadFire_26 ^ readTokenRelease_26)
        tokenCheck_counter_26 <= tokenCheck_counter_26 + tokenCheck_counterChange_26;
      if (pipeReadFire_27 ^ readTokenRelease_27)
        tokenCheck_counter_27 <= tokenCheck_counter_27 + tokenCheck_counterChange_27;
      if (pipeReadFire_28 ^ readTokenRelease_28)
        tokenCheck_counter_28 <= tokenCheck_counter_28 + tokenCheck_counterChange_28;
      if (pipeReadFire_29 ^ readTokenRelease_29)
        tokenCheck_counter_29 <= tokenCheck_counter_29 + tokenCheck_counterChange_29;
      if (pipeReadFire_30 ^ readTokenRelease_30)
        tokenCheck_counter_30 <= tokenCheck_counter_30 + tokenCheck_counterChange_30;
      if (pipeReadFire_31 ^ readTokenRelease_31)
        tokenCheck_counter_31 <= tokenCheck_counter_31 + tokenCheck_counterChange_31;
      if (reorderQueueAllocate_release | readIssueStageEnq) begin
        reorderQueueAllocate_counter <= reorderQueueAllocate_counterUpdate;
        reorderQueueAllocate_counterWillUpdate <= reorderQueueAllocate_counterUpdate + 7'h20;
      end
      if (reorderQueueAllocate_release_1 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_1 <= reorderQueueAllocate_counterUpdate_1;
        reorderQueueAllocate_counterWillUpdate_1 <= reorderQueueAllocate_counterUpdate_1 + 7'h20;
      end
      if (reorderQueueAllocate_release_2 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_2 <= reorderQueueAllocate_counterUpdate_2;
        reorderQueueAllocate_counterWillUpdate_2 <= reorderQueueAllocate_counterUpdate_2 + 7'h20;
      end
      if (reorderQueueAllocate_release_3 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_3 <= reorderQueueAllocate_counterUpdate_3;
        reorderQueueAllocate_counterWillUpdate_3 <= reorderQueueAllocate_counterUpdate_3 + 7'h20;
      end
      if (reorderQueueAllocate_release_4 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_4 <= reorderQueueAllocate_counterUpdate_4;
        reorderQueueAllocate_counterWillUpdate_4 <= reorderQueueAllocate_counterUpdate_4 + 7'h20;
      end
      if (reorderQueueAllocate_release_5 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_5 <= reorderQueueAllocate_counterUpdate_5;
        reorderQueueAllocate_counterWillUpdate_5 <= reorderQueueAllocate_counterUpdate_5 + 7'h20;
      end
      if (reorderQueueAllocate_release_6 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_6 <= reorderQueueAllocate_counterUpdate_6;
        reorderQueueAllocate_counterWillUpdate_6 <= reorderQueueAllocate_counterUpdate_6 + 7'h20;
      end
      if (reorderQueueAllocate_release_7 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_7 <= reorderQueueAllocate_counterUpdate_7;
        reorderQueueAllocate_counterWillUpdate_7 <= reorderQueueAllocate_counterUpdate_7 + 7'h20;
      end
      if (reorderQueueAllocate_release_8 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_8 <= reorderQueueAllocate_counterUpdate_8;
        reorderQueueAllocate_counterWillUpdate_8 <= reorderQueueAllocate_counterUpdate_8 + 7'h20;
      end
      if (reorderQueueAllocate_release_9 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_9 <= reorderQueueAllocate_counterUpdate_9;
        reorderQueueAllocate_counterWillUpdate_9 <= reorderQueueAllocate_counterUpdate_9 + 7'h20;
      end
      if (reorderQueueAllocate_release_10 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_10 <= reorderQueueAllocate_counterUpdate_10;
        reorderQueueAllocate_counterWillUpdate_10 <= reorderQueueAllocate_counterUpdate_10 + 7'h20;
      end
      if (reorderQueueAllocate_release_11 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_11 <= reorderQueueAllocate_counterUpdate_11;
        reorderQueueAllocate_counterWillUpdate_11 <= reorderQueueAllocate_counterUpdate_11 + 7'h20;
      end
      if (reorderQueueAllocate_release_12 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_12 <= reorderQueueAllocate_counterUpdate_12;
        reorderQueueAllocate_counterWillUpdate_12 <= reorderQueueAllocate_counterUpdate_12 + 7'h20;
      end
      if (reorderQueueAllocate_release_13 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_13 <= reorderQueueAllocate_counterUpdate_13;
        reorderQueueAllocate_counterWillUpdate_13 <= reorderQueueAllocate_counterUpdate_13 + 7'h20;
      end
      if (reorderQueueAllocate_release_14 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_14 <= reorderQueueAllocate_counterUpdate_14;
        reorderQueueAllocate_counterWillUpdate_14 <= reorderQueueAllocate_counterUpdate_14 + 7'h20;
      end
      if (reorderQueueAllocate_release_15 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_15 <= reorderQueueAllocate_counterUpdate_15;
        reorderQueueAllocate_counterWillUpdate_15 <= reorderQueueAllocate_counterUpdate_15 + 7'h20;
      end
      if (reorderQueueAllocate_release_16 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_16 <= reorderQueueAllocate_counterUpdate_16;
        reorderQueueAllocate_counterWillUpdate_16 <= reorderQueueAllocate_counterUpdate_16 + 7'h20;
      end
      if (reorderQueueAllocate_release_17 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_17 <= reorderQueueAllocate_counterUpdate_17;
        reorderQueueAllocate_counterWillUpdate_17 <= reorderQueueAllocate_counterUpdate_17 + 7'h20;
      end
      if (reorderQueueAllocate_release_18 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_18 <= reorderQueueAllocate_counterUpdate_18;
        reorderQueueAllocate_counterWillUpdate_18 <= reorderQueueAllocate_counterUpdate_18 + 7'h20;
      end
      if (reorderQueueAllocate_release_19 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_19 <= reorderQueueAllocate_counterUpdate_19;
        reorderQueueAllocate_counterWillUpdate_19 <= reorderQueueAllocate_counterUpdate_19 + 7'h20;
      end
      if (reorderQueueAllocate_release_20 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_20 <= reorderQueueAllocate_counterUpdate_20;
        reorderQueueAllocate_counterWillUpdate_20 <= reorderQueueAllocate_counterUpdate_20 + 7'h20;
      end
      if (reorderQueueAllocate_release_21 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_21 <= reorderQueueAllocate_counterUpdate_21;
        reorderQueueAllocate_counterWillUpdate_21 <= reorderQueueAllocate_counterUpdate_21 + 7'h20;
      end
      if (reorderQueueAllocate_release_22 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_22 <= reorderQueueAllocate_counterUpdate_22;
        reorderQueueAllocate_counterWillUpdate_22 <= reorderQueueAllocate_counterUpdate_22 + 7'h20;
      end
      if (reorderQueueAllocate_release_23 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_23 <= reorderQueueAllocate_counterUpdate_23;
        reorderQueueAllocate_counterWillUpdate_23 <= reorderQueueAllocate_counterUpdate_23 + 7'h20;
      end
      if (reorderQueueAllocate_release_24 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_24 <= reorderQueueAllocate_counterUpdate_24;
        reorderQueueAllocate_counterWillUpdate_24 <= reorderQueueAllocate_counterUpdate_24 + 7'h20;
      end
      if (reorderQueueAllocate_release_25 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_25 <= reorderQueueAllocate_counterUpdate_25;
        reorderQueueAllocate_counterWillUpdate_25 <= reorderQueueAllocate_counterUpdate_25 + 7'h20;
      end
      if (reorderQueueAllocate_release_26 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_26 <= reorderQueueAllocate_counterUpdate_26;
        reorderQueueAllocate_counterWillUpdate_26 <= reorderQueueAllocate_counterUpdate_26 + 7'h20;
      end
      if (reorderQueueAllocate_release_27 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_27 <= reorderQueueAllocate_counterUpdate_27;
        reorderQueueAllocate_counterWillUpdate_27 <= reorderQueueAllocate_counterUpdate_27 + 7'h20;
      end
      if (reorderQueueAllocate_release_28 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_28 <= reorderQueueAllocate_counterUpdate_28;
        reorderQueueAllocate_counterWillUpdate_28 <= reorderQueueAllocate_counterUpdate_28 + 7'h20;
      end
      if (reorderQueueAllocate_release_29 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_29 <= reorderQueueAllocate_counterUpdate_29;
        reorderQueueAllocate_counterWillUpdate_29 <= reorderQueueAllocate_counterUpdate_29 + 7'h20;
      end
      if (reorderQueueAllocate_release_30 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_30 <= reorderQueueAllocate_counterUpdate_30;
        reorderQueueAllocate_counterWillUpdate_30 <= reorderQueueAllocate_counterUpdate_30 + 7'h20;
      end
      if (reorderQueueAllocate_release_31 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_31 <= reorderQueueAllocate_counterUpdate_31;
        reorderQueueAllocate_counterWillUpdate_31 <= reorderQueueAllocate_counterUpdate_31 + 7'h20;
      end
      if (reorderStageEnqFire ^ reorderStageDeqFire)
        reorderStageValid <= reorderStageEnqFire;
      if (_write1HPipe_0_T & readType)
        reorderStageState_0 <= reorderStageState_0 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_0 <= 6'h0;
      if (_write1HPipe_1_T & readType)
        reorderStageState_1 <= reorderStageState_1 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_1 <= 6'h0;
      if (_write1HPipe_2_T & readType)
        reorderStageState_2 <= reorderStageState_2 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_2 <= 6'h0;
      if (_write1HPipe_3_T & readType)
        reorderStageState_3 <= reorderStageState_3 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_3 <= 6'h0;
      if (_write1HPipe_4_T & readType)
        reorderStageState_4 <= reorderStageState_4 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_4 <= 6'h0;
      if (_write1HPipe_5_T & readType)
        reorderStageState_5 <= reorderStageState_5 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_5 <= 6'h0;
      if (_write1HPipe_6_T & readType)
        reorderStageState_6 <= reorderStageState_6 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_6 <= 6'h0;
      if (_write1HPipe_7_T & readType)
        reorderStageState_7 <= reorderStageState_7 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_7 <= 6'h0;
      if (_write1HPipe_8_T & readType)
        reorderStageState_8 <= reorderStageState_8 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_8 <= 6'h0;
      if (_write1HPipe_9_T & readType)
        reorderStageState_9 <= reorderStageState_9 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_9 <= 6'h0;
      if (_write1HPipe_10_T & readType)
        reorderStageState_10 <= reorderStageState_10 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_10 <= 6'h0;
      if (_write1HPipe_11_T & readType)
        reorderStageState_11 <= reorderStageState_11 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_11 <= 6'h0;
      if (_write1HPipe_12_T & readType)
        reorderStageState_12 <= reorderStageState_12 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_12 <= 6'h0;
      if (_write1HPipe_13_T & readType)
        reorderStageState_13 <= reorderStageState_13 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_13 <= 6'h0;
      if (_write1HPipe_14_T & readType)
        reorderStageState_14 <= reorderStageState_14 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_14 <= 6'h0;
      if (_write1HPipe_15_T & readType)
        reorderStageState_15 <= reorderStageState_15 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_15 <= 6'h0;
      if (_write1HPipe_16_T & readType)
        reorderStageState_16 <= reorderStageState_16 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_16 <= 6'h0;
      if (_write1HPipe_17_T & readType)
        reorderStageState_17 <= reorderStageState_17 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_17 <= 6'h0;
      if (_write1HPipe_18_T & readType)
        reorderStageState_18 <= reorderStageState_18 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_18 <= 6'h0;
      if (_write1HPipe_19_T & readType)
        reorderStageState_19 <= reorderStageState_19 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_19 <= 6'h0;
      if (_write1HPipe_20_T & readType)
        reorderStageState_20 <= reorderStageState_20 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_20 <= 6'h0;
      if (_write1HPipe_21_T & readType)
        reorderStageState_21 <= reorderStageState_21 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_21 <= 6'h0;
      if (_write1HPipe_22_T & readType)
        reorderStageState_22 <= reorderStageState_22 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_22 <= 6'h0;
      if (_write1HPipe_23_T & readType)
        reorderStageState_23 <= reorderStageState_23 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_23 <= 6'h0;
      if (_write1HPipe_24_T & readType)
        reorderStageState_24 <= reorderStageState_24 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_24 <= 6'h0;
      if (_write1HPipe_25_T & readType)
        reorderStageState_25 <= reorderStageState_25 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_25 <= 6'h0;
      if (_write1HPipe_26_T & readType)
        reorderStageState_26 <= reorderStageState_26 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_26 <= 6'h0;
      if (_write1HPipe_27_T & readType)
        reorderStageState_27 <= reorderStageState_27 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_27 <= 6'h0;
      if (_write1HPipe_28_T & readType)
        reorderStageState_28 <= reorderStageState_28 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_28 <= 6'h0;
      if (_write1HPipe_29_T & readType)
        reorderStageState_29 <= reorderStageState_29 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_29 <= 6'h0;
      if (_write1HPipe_30_T & readType)
        reorderStageState_30 <= reorderStageState_30 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_30 <= 6'h0;
      if (_write1HPipe_31_T & readType)
        reorderStageState_31 <= reorderStageState_31 + 6'h1;
      else if (reorderStageEnqFire)
        reorderStageState_31 <= 6'h0;
      if (reorderStageEnqFire) begin
        reorderStageNeed_0 <= accessCountQueue_deq_bits_0;
        reorderStageNeed_1 <= accessCountQueue_deq_bits_1;
        reorderStageNeed_2 <= accessCountQueue_deq_bits_2;
        reorderStageNeed_3 <= accessCountQueue_deq_bits_3;
        reorderStageNeed_4 <= accessCountQueue_deq_bits_4;
        reorderStageNeed_5 <= accessCountQueue_deq_bits_5;
        reorderStageNeed_6 <= accessCountQueue_deq_bits_6;
        reorderStageNeed_7 <= accessCountQueue_deq_bits_7;
        reorderStageNeed_8 <= accessCountQueue_deq_bits_8;
        reorderStageNeed_9 <= accessCountQueue_deq_bits_9;
        reorderStageNeed_10 <= accessCountQueue_deq_bits_10;
        reorderStageNeed_11 <= accessCountQueue_deq_bits_11;
        reorderStageNeed_12 <= accessCountQueue_deq_bits_12;
        reorderStageNeed_13 <= accessCountQueue_deq_bits_13;
        reorderStageNeed_14 <= accessCountQueue_deq_bits_14;
        reorderStageNeed_15 <= accessCountQueue_deq_bits_15;
        reorderStageNeed_16 <= accessCountQueue_deq_bits_16;
        reorderStageNeed_17 <= accessCountQueue_deq_bits_17;
        reorderStageNeed_18 <= accessCountQueue_deq_bits_18;
        reorderStageNeed_19 <= accessCountQueue_deq_bits_19;
        reorderStageNeed_20 <= accessCountQueue_deq_bits_20;
        reorderStageNeed_21 <= accessCountQueue_deq_bits_21;
        reorderStageNeed_22 <= accessCountQueue_deq_bits_22;
        reorderStageNeed_23 <= accessCountQueue_deq_bits_23;
        reorderStageNeed_24 <= accessCountQueue_deq_bits_24;
        reorderStageNeed_25 <= accessCountQueue_deq_bits_25;
        reorderStageNeed_26 <= accessCountQueue_deq_bits_26;
        reorderStageNeed_27 <= accessCountQueue_deq_bits_27;
        reorderStageNeed_28 <= accessCountQueue_deq_bits_28;
        reorderStageNeed_29 <= accessCountQueue_deq_bits_29;
        reorderStageNeed_30 <= accessCountQueue_deq_bits_30;
        reorderStageNeed_31 <= accessCountQueue_deq_bits_31;
      end
      if (waiteStageEnqFire) begin
        waiteReadDataPipeReg_executeGroup <= readWaitQueue_deq_bits_executeGroup;
        waiteReadDataPipeReg_sourceValid <= readWaitQueue_deq_bits_sourceValid;
        waiteReadDataPipeReg_replaceVs1 <= readWaitQueue_deq_bits_replaceVs1;
        waiteReadDataPipeReg_needRead <= readWaitQueue_deq_bits_needRead;
        waiteReadDataPipeReg_last <= readWaitQueue_deq_bits_last;
      end
      if (readTokenRelease_1)
        waiteReadData_1 <= readData_readDataQueue_1_deq_bits;
      if (readTokenRelease_2)
        waiteReadData_2 <= readData_readDataQueue_2_deq_bits;
      if (readTokenRelease_3)
        waiteReadData_3 <= readData_readDataQueue_3_deq_bits;
      if (readTokenRelease_4)
        waiteReadData_4 <= readData_readDataQueue_4_deq_bits;
      if (readTokenRelease_5)
        waiteReadData_5 <= readData_readDataQueue_5_deq_bits;
      if (readTokenRelease_6)
        waiteReadData_6 <= readData_readDataQueue_6_deq_bits;
      if (readTokenRelease_7)
        waiteReadData_7 <= readData_readDataQueue_7_deq_bits;
      if (readTokenRelease_8)
        waiteReadData_8 <= readData_readDataQueue_8_deq_bits;
      if (readTokenRelease_9)
        waiteReadData_9 <= readData_readDataQueue_9_deq_bits;
      if (readTokenRelease_10)
        waiteReadData_10 <= readData_readDataQueue_10_deq_bits;
      if (readTokenRelease_11)
        waiteReadData_11 <= readData_readDataQueue_11_deq_bits;
      if (readTokenRelease_12)
        waiteReadData_12 <= readData_readDataQueue_12_deq_bits;
      if (readTokenRelease_13)
        waiteReadData_13 <= readData_readDataQueue_13_deq_bits;
      if (readTokenRelease_14)
        waiteReadData_14 <= readData_readDataQueue_14_deq_bits;
      if (readTokenRelease_15)
        waiteReadData_15 <= readData_readDataQueue_15_deq_bits;
      if (readTokenRelease_16)
        waiteReadData_16 <= readData_readDataQueue_16_deq_bits;
      if (readTokenRelease_17)
        waiteReadData_17 <= readData_readDataQueue_17_deq_bits;
      if (readTokenRelease_18)
        waiteReadData_18 <= readData_readDataQueue_18_deq_bits;
      if (readTokenRelease_19)
        waiteReadData_19 <= readData_readDataQueue_19_deq_bits;
      if (readTokenRelease_20)
        waiteReadData_20 <= readData_readDataQueue_20_deq_bits;
      if (readTokenRelease_21)
        waiteReadData_21 <= readData_readDataQueue_21_deq_bits;
      if (readTokenRelease_22)
        waiteReadData_22 <= readData_readDataQueue_22_deq_bits;
      if (readTokenRelease_23)
        waiteReadData_23 <= readData_readDataQueue_23_deq_bits;
      if (readTokenRelease_24)
        waiteReadData_24 <= readData_readDataQueue_24_deq_bits;
      if (readTokenRelease_25)
        waiteReadData_25 <= readData_readDataQueue_25_deq_bits;
      if (readTokenRelease_26)
        waiteReadData_26 <= readData_readDataQueue_26_deq_bits;
      if (readTokenRelease_27)
        waiteReadData_27 <= readData_readDataQueue_27_deq_bits;
      if (readTokenRelease_28)
        waiteReadData_28 <= readData_readDataQueue_28_deq_bits;
      if (readTokenRelease_29)
        waiteReadData_29 <= readData_readDataQueue_29_deq_bits;
      if (readTokenRelease_30)
        waiteReadData_30 <= readData_readDataQueue_30_deq_bits;
      if (readTokenRelease_31)
        waiteReadData_31 <= readData_readDataQueue_31_deq_bits;
      if (waiteStageEnqFire & (|readResultValid))
        waiteReadSate <= readResultValid;
      else if (|readResultValid)
        waiteReadSate <= waiteReadSate | readResultValid;
      else if (waiteStageEnqFire)
        waiteReadSate <= 32'h0;
      if (waiteStageDeqFire ^ waiteStageEnqFire)
        waiteReadStageValid <= waiteStageEnqFire;
      if (_dataNotInShifter_T ^ writeRelease_0)
        dataNotInShifter_writeTokenCounter <= dataNotInShifter_writeTokenCounter + dataNotInShifter_writeTokenChange;
      if (_dataNotInShifter_T_3 ^ writeRelease_1)
        dataNotInShifter_writeTokenCounter_1 <= dataNotInShifter_writeTokenCounter_1 + dataNotInShifter_writeTokenChange_1;
      if (_dataNotInShifter_T_6 ^ writeRelease_2)
        dataNotInShifter_writeTokenCounter_2 <= dataNotInShifter_writeTokenCounter_2 + dataNotInShifter_writeTokenChange_2;
      if (_dataNotInShifter_T_9 ^ writeRelease_3)
        dataNotInShifter_writeTokenCounter_3 <= dataNotInShifter_writeTokenCounter_3 + dataNotInShifter_writeTokenChange_3;
      if (_dataNotInShifter_T_12 ^ writeRelease_4)
        dataNotInShifter_writeTokenCounter_4 <= dataNotInShifter_writeTokenCounter_4 + dataNotInShifter_writeTokenChange_4;
      if (_dataNotInShifter_T_15 ^ writeRelease_5)
        dataNotInShifter_writeTokenCounter_5 <= dataNotInShifter_writeTokenCounter_5 + dataNotInShifter_writeTokenChange_5;
      if (_dataNotInShifter_T_18 ^ writeRelease_6)
        dataNotInShifter_writeTokenCounter_6 <= dataNotInShifter_writeTokenCounter_6 + dataNotInShifter_writeTokenChange_6;
      if (_dataNotInShifter_T_21 ^ writeRelease_7)
        dataNotInShifter_writeTokenCounter_7 <= dataNotInShifter_writeTokenCounter_7 + dataNotInShifter_writeTokenChange_7;
      if (_dataNotInShifter_T_24 ^ writeRelease_8)
        dataNotInShifter_writeTokenCounter_8 <= dataNotInShifter_writeTokenCounter_8 + dataNotInShifter_writeTokenChange_8;
      if (_dataNotInShifter_T_27 ^ writeRelease_9)
        dataNotInShifter_writeTokenCounter_9 <= dataNotInShifter_writeTokenCounter_9 + dataNotInShifter_writeTokenChange_9;
      if (_dataNotInShifter_T_30 ^ writeRelease_10)
        dataNotInShifter_writeTokenCounter_10 <= dataNotInShifter_writeTokenCounter_10 + dataNotInShifter_writeTokenChange_10;
      if (_dataNotInShifter_T_33 ^ writeRelease_11)
        dataNotInShifter_writeTokenCounter_11 <= dataNotInShifter_writeTokenCounter_11 + dataNotInShifter_writeTokenChange_11;
      if (_dataNotInShifter_T_36 ^ writeRelease_12)
        dataNotInShifter_writeTokenCounter_12 <= dataNotInShifter_writeTokenCounter_12 + dataNotInShifter_writeTokenChange_12;
      if (_dataNotInShifter_T_39 ^ writeRelease_13)
        dataNotInShifter_writeTokenCounter_13 <= dataNotInShifter_writeTokenCounter_13 + dataNotInShifter_writeTokenChange_13;
      if (_dataNotInShifter_T_42 ^ writeRelease_14)
        dataNotInShifter_writeTokenCounter_14 <= dataNotInShifter_writeTokenCounter_14 + dataNotInShifter_writeTokenChange_14;
      if (_dataNotInShifter_T_45 ^ writeRelease_15)
        dataNotInShifter_writeTokenCounter_15 <= dataNotInShifter_writeTokenCounter_15 + dataNotInShifter_writeTokenChange_15;
      if (_dataNotInShifter_T_48 ^ writeRelease_16)
        dataNotInShifter_writeTokenCounter_16 <= dataNotInShifter_writeTokenCounter_16 + dataNotInShifter_writeTokenChange_16;
      if (_dataNotInShifter_T_51 ^ writeRelease_17)
        dataNotInShifter_writeTokenCounter_17 <= dataNotInShifter_writeTokenCounter_17 + dataNotInShifter_writeTokenChange_17;
      if (_dataNotInShifter_T_54 ^ writeRelease_18)
        dataNotInShifter_writeTokenCounter_18 <= dataNotInShifter_writeTokenCounter_18 + dataNotInShifter_writeTokenChange_18;
      if (_dataNotInShifter_T_57 ^ writeRelease_19)
        dataNotInShifter_writeTokenCounter_19 <= dataNotInShifter_writeTokenCounter_19 + dataNotInShifter_writeTokenChange_19;
      if (_dataNotInShifter_T_60 ^ writeRelease_20)
        dataNotInShifter_writeTokenCounter_20 <= dataNotInShifter_writeTokenCounter_20 + dataNotInShifter_writeTokenChange_20;
      if (_dataNotInShifter_T_63 ^ writeRelease_21)
        dataNotInShifter_writeTokenCounter_21 <= dataNotInShifter_writeTokenCounter_21 + dataNotInShifter_writeTokenChange_21;
      if (_dataNotInShifter_T_66 ^ writeRelease_22)
        dataNotInShifter_writeTokenCounter_22 <= dataNotInShifter_writeTokenCounter_22 + dataNotInShifter_writeTokenChange_22;
      if (_dataNotInShifter_T_69 ^ writeRelease_23)
        dataNotInShifter_writeTokenCounter_23 <= dataNotInShifter_writeTokenCounter_23 + dataNotInShifter_writeTokenChange_23;
      if (_dataNotInShifter_T_72 ^ writeRelease_24)
        dataNotInShifter_writeTokenCounter_24 <= dataNotInShifter_writeTokenCounter_24 + dataNotInShifter_writeTokenChange_24;
      if (_dataNotInShifter_T_75 ^ writeRelease_25)
        dataNotInShifter_writeTokenCounter_25 <= dataNotInShifter_writeTokenCounter_25 + dataNotInShifter_writeTokenChange_25;
      if (_dataNotInShifter_T_78 ^ writeRelease_26)
        dataNotInShifter_writeTokenCounter_26 <= dataNotInShifter_writeTokenCounter_26 + dataNotInShifter_writeTokenChange_26;
      if (_dataNotInShifter_T_81 ^ writeRelease_27)
        dataNotInShifter_writeTokenCounter_27 <= dataNotInShifter_writeTokenCounter_27 + dataNotInShifter_writeTokenChange_27;
      if (_dataNotInShifter_T_84 ^ writeRelease_28)
        dataNotInShifter_writeTokenCounter_28 <= dataNotInShifter_writeTokenCounter_28 + dataNotInShifter_writeTokenChange_28;
      if (_dataNotInShifter_T_87 ^ writeRelease_29)
        dataNotInShifter_writeTokenCounter_29 <= dataNotInShifter_writeTokenCounter_29 + dataNotInShifter_writeTokenChange_29;
      if (_dataNotInShifter_T_90 ^ writeRelease_30)
        dataNotInShifter_writeTokenCounter_30 <= dataNotInShifter_writeTokenCounter_30 + dataNotInShifter_writeTokenChange_30;
      if (_dataNotInShifter_T_93 ^ writeRelease_31)
        dataNotInShifter_writeTokenCounter_31 <= dataNotInShifter_writeTokenCounter_31 + dataNotInShifter_writeTokenChange_31;
      waiteLastRequest <= ~readType & requestStageDeq & lastGroup | ~lastReportValid & waiteLastRequest;
      waitQueueClear <= executeStageClean | invalidEnq | ~lastReportValid & waitQueueClear;
    end
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:224];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [7:0] i = 8'h0; i < 8'hE1; i += 8'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        v0_0 = _RANDOM[8'h0];
        v0_1 = _RANDOM[8'h1];
        v0_2 = _RANDOM[8'h2];
        v0_3 = _RANDOM[8'h3];
        v0_4 = _RANDOM[8'h4];
        v0_5 = _RANDOM[8'h5];
        v0_6 = _RANDOM[8'h6];
        v0_7 = _RANDOM[8'h7];
        v0_8 = _RANDOM[8'h8];
        v0_9 = _RANDOM[8'h9];
        v0_10 = _RANDOM[8'hA];
        v0_11 = _RANDOM[8'hB];
        v0_12 = _RANDOM[8'hC];
        v0_13 = _RANDOM[8'hD];
        v0_14 = _RANDOM[8'hE];
        v0_15 = _RANDOM[8'hF];
        v0_16 = _RANDOM[8'h10];
        v0_17 = _RANDOM[8'h11];
        v0_18 = _RANDOM[8'h12];
        v0_19 = _RANDOM[8'h13];
        v0_20 = _RANDOM[8'h14];
        v0_21 = _RANDOM[8'h15];
        v0_22 = _RANDOM[8'h16];
        v0_23 = _RANDOM[8'h17];
        v0_24 = _RANDOM[8'h18];
        v0_25 = _RANDOM[8'h19];
        v0_26 = _RANDOM[8'h1A];
        v0_27 = _RANDOM[8'h1B];
        v0_28 = _RANDOM[8'h1C];
        v0_29 = _RANDOM[8'h1D];
        v0_30 = _RANDOM[8'h1E];
        v0_31 = _RANDOM[8'h1F];
        v0_32 = _RANDOM[8'h20];
        v0_33 = _RANDOM[8'h21];
        v0_34 = _RANDOM[8'h22];
        v0_35 = _RANDOM[8'h23];
        v0_36 = _RANDOM[8'h24];
        v0_37 = _RANDOM[8'h25];
        v0_38 = _RANDOM[8'h26];
        v0_39 = _RANDOM[8'h27];
        v0_40 = _RANDOM[8'h28];
        v0_41 = _RANDOM[8'h29];
        v0_42 = _RANDOM[8'h2A];
        v0_43 = _RANDOM[8'h2B];
        v0_44 = _RANDOM[8'h2C];
        v0_45 = _RANDOM[8'h2D];
        v0_46 = _RANDOM[8'h2E];
        v0_47 = _RANDOM[8'h2F];
        v0_48 = _RANDOM[8'h30];
        v0_49 = _RANDOM[8'h31];
        v0_50 = _RANDOM[8'h32];
        v0_51 = _RANDOM[8'h33];
        v0_52 = _RANDOM[8'h34];
        v0_53 = _RANDOM[8'h35];
        v0_54 = _RANDOM[8'h36];
        v0_55 = _RANDOM[8'h37];
        v0_56 = _RANDOM[8'h38];
        v0_57 = _RANDOM[8'h39];
        v0_58 = _RANDOM[8'h3A];
        v0_59 = _RANDOM[8'h3B];
        v0_60 = _RANDOM[8'h3C];
        v0_61 = _RANDOM[8'h3D];
        v0_62 = _RANDOM[8'h3E];
        v0_63 = _RANDOM[8'h3F];
        gatherReadState = _RANDOM[8'h40][1:0];
        gatherDatOffset = _RANDOM[8'h40][3:2];
        gatherLane = _RANDOM[8'h40][8:4];
        gatherOffset = _RANDOM[8'h40][9];
        gatherGrowth = _RANDOM[8'h40][12:10];
        instReg_instructionIndex = _RANDOM[8'h40][15:13];
        instReg_decodeResult_specialSlot = _RANDOM[8'h40][16];
        instReg_decodeResult_topUop = _RANDOM[8'h40][21:17];
        instReg_decodeResult_popCount = _RANDOM[8'h40][22];
        instReg_decodeResult_ffo = _RANDOM[8'h40][23];
        instReg_decodeResult_average = _RANDOM[8'h40][24];
        instReg_decodeResult_reverse = _RANDOM[8'h40][25];
        instReg_decodeResult_dontNeedExecuteInLane = _RANDOM[8'h40][26];
        instReg_decodeResult_scheduler = _RANDOM[8'h40][27];
        instReg_decodeResult_sReadVD = _RANDOM[8'h40][28];
        instReg_decodeResult_vtype = _RANDOM[8'h40][29];
        instReg_decodeResult_sWrite = _RANDOM[8'h40][30];
        instReg_decodeResult_crossRead = _RANDOM[8'h40][31];
        instReg_decodeResult_crossWrite = _RANDOM[8'h41][0];
        instReg_decodeResult_maskUnit = _RANDOM[8'h41][1];
        instReg_decodeResult_special = _RANDOM[8'h41][2];
        instReg_decodeResult_saturate = _RANDOM[8'h41][3];
        instReg_decodeResult_vwmacc = _RANDOM[8'h41][4];
        instReg_decodeResult_readOnly = _RANDOM[8'h41][5];
        instReg_decodeResult_maskSource = _RANDOM[8'h41][6];
        instReg_decodeResult_maskDestination = _RANDOM[8'h41][7];
        instReg_decodeResult_maskLogic = _RANDOM[8'h41][8];
        instReg_decodeResult_uop = _RANDOM[8'h41][12:9];
        instReg_decodeResult_iota = _RANDOM[8'h41][13];
        instReg_decodeResult_mv = _RANDOM[8'h41][14];
        instReg_decodeResult_extend = _RANDOM[8'h41][15];
        instReg_decodeResult_unOrderWrite = _RANDOM[8'h41][16];
        instReg_decodeResult_compress = _RANDOM[8'h41][17];
        instReg_decodeResult_gather16 = _RANDOM[8'h41][18];
        instReg_decodeResult_gather = _RANDOM[8'h41][19];
        instReg_decodeResult_slid = _RANDOM[8'h41][20];
        instReg_decodeResult_targetRd = _RANDOM[8'h41][21];
        instReg_decodeResult_widenReduce = _RANDOM[8'h41][22];
        instReg_decodeResult_red = _RANDOM[8'h41][23];
        instReg_decodeResult_nr = _RANDOM[8'h41][24];
        instReg_decodeResult_itype = _RANDOM[8'h41][25];
        instReg_decodeResult_unsigned1 = _RANDOM[8'h41][26];
        instReg_decodeResult_unsigned0 = _RANDOM[8'h41][27];
        instReg_decodeResult_other = _RANDOM[8'h41][28];
        instReg_decodeResult_multiCycle = _RANDOM[8'h41][29];
        instReg_decodeResult_divider = _RANDOM[8'h41][30];
        instReg_decodeResult_multiplier = _RANDOM[8'h41][31];
        instReg_decodeResult_shift = _RANDOM[8'h42][0];
        instReg_decodeResult_adder = _RANDOM[8'h42][1];
        instReg_decodeResult_logic = _RANDOM[8'h42][2];
        instReg_readFromScala = {_RANDOM[8'h42][31:3], _RANDOM[8'h43][2:0]};
        instReg_sew = _RANDOM[8'h43][4:3];
        instReg_vlmul = _RANDOM[8'h43][7:5];
        instReg_maskType = _RANDOM[8'h43][8];
        instReg_vxrm = _RANDOM[8'h43][11:9];
        instReg_vs2 = _RANDOM[8'h43][16:12];
        instReg_vs1 = _RANDOM[8'h43][21:17];
        instReg_vd = _RANDOM[8'h43][26:22];
        instReg_vl = {_RANDOM[8'h43][31:27], _RANDOM[8'h44][6:0]};
        instVlValid = _RANDOM[8'h44][7];
        readVS1Reg_dataValid = _RANDOM[8'h44][8];
        readVS1Reg_requestSend = _RANDOM[8'h44][9];
        readVS1Reg_sendToExecution = _RANDOM[8'h44][10];
        readVS1Reg_data = {_RANDOM[8'h44][31:11], _RANDOM[8'h45][10:0]};
        readVS1Reg_readIndex = _RANDOM[8'h45][14:11];
        exeReqReg_0_valid = _RANDOM[8'h46][15];
        exeReqReg_0_bits_source1 = {_RANDOM[8'h46][31:16], _RANDOM[8'h47][15:0]};
        exeReqReg_0_bits_source2 = {_RANDOM[8'h47][31:16], _RANDOM[8'h48][15:0]};
        exeReqReg_0_bits_index = _RANDOM[8'h48][18:16];
        exeReqReg_0_bits_ffo = _RANDOM[8'h48][19];
        exeReqReg_1_valid = _RANDOM[8'h48][20];
        exeReqReg_1_bits_source1 = {_RANDOM[8'h48][31:21], _RANDOM[8'h49][20:0]};
        exeReqReg_1_bits_source2 = {_RANDOM[8'h49][31:21], _RANDOM[8'h4A][20:0]};
        exeReqReg_1_bits_index = _RANDOM[8'h4A][23:21];
        exeReqReg_1_bits_ffo = _RANDOM[8'h4A][24];
        exeReqReg_2_valid = _RANDOM[8'h4A][25];
        exeReqReg_2_bits_source1 = {_RANDOM[8'h4A][31:26], _RANDOM[8'h4B][25:0]};
        exeReqReg_2_bits_source2 = {_RANDOM[8'h4B][31:26], _RANDOM[8'h4C][25:0]};
        exeReqReg_2_bits_index = _RANDOM[8'h4C][28:26];
        exeReqReg_2_bits_ffo = _RANDOM[8'h4C][29];
        exeReqReg_3_valid = _RANDOM[8'h4C][30];
        exeReqReg_3_bits_source1 = {_RANDOM[8'h4C][31], _RANDOM[8'h4D][30:0]};
        exeReqReg_3_bits_source2 = {_RANDOM[8'h4D][31], _RANDOM[8'h4E][30:0]};
        exeReqReg_3_bits_index = {_RANDOM[8'h4E][31], _RANDOM[8'h4F][1:0]};
        exeReqReg_3_bits_ffo = _RANDOM[8'h4F][2];
        exeReqReg_4_valid = _RANDOM[8'h4F][3];
        exeReqReg_4_bits_source1 = {_RANDOM[8'h4F][31:4], _RANDOM[8'h50][3:0]};
        exeReqReg_4_bits_source2 = {_RANDOM[8'h50][31:4], _RANDOM[8'h51][3:0]};
        exeReqReg_4_bits_index = _RANDOM[8'h51][6:4];
        exeReqReg_4_bits_ffo = _RANDOM[8'h51][7];
        exeReqReg_5_valid = _RANDOM[8'h51][8];
        exeReqReg_5_bits_source1 = {_RANDOM[8'h51][31:9], _RANDOM[8'h52][8:0]};
        exeReqReg_5_bits_source2 = {_RANDOM[8'h52][31:9], _RANDOM[8'h53][8:0]};
        exeReqReg_5_bits_index = _RANDOM[8'h53][11:9];
        exeReqReg_5_bits_ffo = _RANDOM[8'h53][12];
        exeReqReg_6_valid = _RANDOM[8'h53][13];
        exeReqReg_6_bits_source1 = {_RANDOM[8'h53][31:14], _RANDOM[8'h54][13:0]};
        exeReqReg_6_bits_source2 = {_RANDOM[8'h54][31:14], _RANDOM[8'h55][13:0]};
        exeReqReg_6_bits_index = _RANDOM[8'h55][16:14];
        exeReqReg_6_bits_ffo = _RANDOM[8'h55][17];
        exeReqReg_7_valid = _RANDOM[8'h55][18];
        exeReqReg_7_bits_source1 = {_RANDOM[8'h55][31:19], _RANDOM[8'h56][18:0]};
        exeReqReg_7_bits_source2 = {_RANDOM[8'h56][31:19], _RANDOM[8'h57][18:0]};
        exeReqReg_7_bits_index = _RANDOM[8'h57][21:19];
        exeReqReg_7_bits_ffo = _RANDOM[8'h57][22];
        exeReqReg_8_valid = _RANDOM[8'h57][23];
        exeReqReg_8_bits_source1 = {_RANDOM[8'h57][31:24], _RANDOM[8'h58][23:0]};
        exeReqReg_8_bits_source2 = {_RANDOM[8'h58][31:24], _RANDOM[8'h59][23:0]};
        exeReqReg_8_bits_index = _RANDOM[8'h59][26:24];
        exeReqReg_8_bits_ffo = _RANDOM[8'h59][27];
        exeReqReg_9_valid = _RANDOM[8'h59][28];
        exeReqReg_9_bits_source1 = {_RANDOM[8'h59][31:29], _RANDOM[8'h5A][28:0]};
        exeReqReg_9_bits_source2 = {_RANDOM[8'h5A][31:29], _RANDOM[8'h5B][28:0]};
        exeReqReg_9_bits_index = _RANDOM[8'h5B][31:29];
        exeReqReg_9_bits_ffo = _RANDOM[8'h5C][0];
        exeReqReg_10_valid = _RANDOM[8'h5C][1];
        exeReqReg_10_bits_source1 = {_RANDOM[8'h5C][31:2], _RANDOM[8'h5D][1:0]};
        exeReqReg_10_bits_source2 = {_RANDOM[8'h5D][31:2], _RANDOM[8'h5E][1:0]};
        exeReqReg_10_bits_index = _RANDOM[8'h5E][4:2];
        exeReqReg_10_bits_ffo = _RANDOM[8'h5E][5];
        exeReqReg_11_valid = _RANDOM[8'h5E][6];
        exeReqReg_11_bits_source1 = {_RANDOM[8'h5E][31:7], _RANDOM[8'h5F][6:0]};
        exeReqReg_11_bits_source2 = {_RANDOM[8'h5F][31:7], _RANDOM[8'h60][6:0]};
        exeReqReg_11_bits_index = _RANDOM[8'h60][9:7];
        exeReqReg_11_bits_ffo = _RANDOM[8'h60][10];
        exeReqReg_12_valid = _RANDOM[8'h60][11];
        exeReqReg_12_bits_source1 = {_RANDOM[8'h60][31:12], _RANDOM[8'h61][11:0]};
        exeReqReg_12_bits_source2 = {_RANDOM[8'h61][31:12], _RANDOM[8'h62][11:0]};
        exeReqReg_12_bits_index = _RANDOM[8'h62][14:12];
        exeReqReg_12_bits_ffo = _RANDOM[8'h62][15];
        exeReqReg_13_valid = _RANDOM[8'h62][16];
        exeReqReg_13_bits_source1 = {_RANDOM[8'h62][31:17], _RANDOM[8'h63][16:0]};
        exeReqReg_13_bits_source2 = {_RANDOM[8'h63][31:17], _RANDOM[8'h64][16:0]};
        exeReqReg_13_bits_index = _RANDOM[8'h64][19:17];
        exeReqReg_13_bits_ffo = _RANDOM[8'h64][20];
        exeReqReg_14_valid = _RANDOM[8'h64][21];
        exeReqReg_14_bits_source1 = {_RANDOM[8'h64][31:22], _RANDOM[8'h65][21:0]};
        exeReqReg_14_bits_source2 = {_RANDOM[8'h65][31:22], _RANDOM[8'h66][21:0]};
        exeReqReg_14_bits_index = _RANDOM[8'h66][24:22];
        exeReqReg_14_bits_ffo = _RANDOM[8'h66][25];
        exeReqReg_15_valid = _RANDOM[8'h66][26];
        exeReqReg_15_bits_source1 = {_RANDOM[8'h66][31:27], _RANDOM[8'h67][26:0]};
        exeReqReg_15_bits_source2 = {_RANDOM[8'h67][31:27], _RANDOM[8'h68][26:0]};
        exeReqReg_15_bits_index = _RANDOM[8'h68][29:27];
        exeReqReg_15_bits_ffo = _RANDOM[8'h68][30];
        exeReqReg_16_valid = _RANDOM[8'h68][31];
        exeReqReg_16_bits_source1 = _RANDOM[8'h69];
        exeReqReg_16_bits_source2 = _RANDOM[8'h6A];
        exeReqReg_16_bits_index = _RANDOM[8'h6B][2:0];
        exeReqReg_16_bits_ffo = _RANDOM[8'h6B][3];
        exeReqReg_17_valid = _RANDOM[8'h6B][4];
        exeReqReg_17_bits_source1 = {_RANDOM[8'h6B][31:5], _RANDOM[8'h6C][4:0]};
        exeReqReg_17_bits_source2 = {_RANDOM[8'h6C][31:5], _RANDOM[8'h6D][4:0]};
        exeReqReg_17_bits_index = _RANDOM[8'h6D][7:5];
        exeReqReg_17_bits_ffo = _RANDOM[8'h6D][8];
        exeReqReg_18_valid = _RANDOM[8'h6D][9];
        exeReqReg_18_bits_source1 = {_RANDOM[8'h6D][31:10], _RANDOM[8'h6E][9:0]};
        exeReqReg_18_bits_source2 = {_RANDOM[8'h6E][31:10], _RANDOM[8'h6F][9:0]};
        exeReqReg_18_bits_index = _RANDOM[8'h6F][12:10];
        exeReqReg_18_bits_ffo = _RANDOM[8'h6F][13];
        exeReqReg_19_valid = _RANDOM[8'h6F][14];
        exeReqReg_19_bits_source1 = {_RANDOM[8'h6F][31:15], _RANDOM[8'h70][14:0]};
        exeReqReg_19_bits_source2 = {_RANDOM[8'h70][31:15], _RANDOM[8'h71][14:0]};
        exeReqReg_19_bits_index = _RANDOM[8'h71][17:15];
        exeReqReg_19_bits_ffo = _RANDOM[8'h71][18];
        exeReqReg_20_valid = _RANDOM[8'h71][19];
        exeReqReg_20_bits_source1 = {_RANDOM[8'h71][31:20], _RANDOM[8'h72][19:0]};
        exeReqReg_20_bits_source2 = {_RANDOM[8'h72][31:20], _RANDOM[8'h73][19:0]};
        exeReqReg_20_bits_index = _RANDOM[8'h73][22:20];
        exeReqReg_20_bits_ffo = _RANDOM[8'h73][23];
        exeReqReg_21_valid = _RANDOM[8'h73][24];
        exeReqReg_21_bits_source1 = {_RANDOM[8'h73][31:25], _RANDOM[8'h74][24:0]};
        exeReqReg_21_bits_source2 = {_RANDOM[8'h74][31:25], _RANDOM[8'h75][24:0]};
        exeReqReg_21_bits_index = _RANDOM[8'h75][27:25];
        exeReqReg_21_bits_ffo = _RANDOM[8'h75][28];
        exeReqReg_22_valid = _RANDOM[8'h75][29];
        exeReqReg_22_bits_source1 = {_RANDOM[8'h75][31:30], _RANDOM[8'h76][29:0]};
        exeReqReg_22_bits_source2 = {_RANDOM[8'h76][31:30], _RANDOM[8'h77][29:0]};
        exeReqReg_22_bits_index = {_RANDOM[8'h77][31:30], _RANDOM[8'h78][0]};
        exeReqReg_22_bits_ffo = _RANDOM[8'h78][1];
        exeReqReg_23_valid = _RANDOM[8'h78][2];
        exeReqReg_23_bits_source1 = {_RANDOM[8'h78][31:3], _RANDOM[8'h79][2:0]};
        exeReqReg_23_bits_source2 = {_RANDOM[8'h79][31:3], _RANDOM[8'h7A][2:0]};
        exeReqReg_23_bits_index = _RANDOM[8'h7A][5:3];
        exeReqReg_23_bits_ffo = _RANDOM[8'h7A][6];
        exeReqReg_24_valid = _RANDOM[8'h7A][7];
        exeReqReg_24_bits_source1 = {_RANDOM[8'h7A][31:8], _RANDOM[8'h7B][7:0]};
        exeReqReg_24_bits_source2 = {_RANDOM[8'h7B][31:8], _RANDOM[8'h7C][7:0]};
        exeReqReg_24_bits_index = _RANDOM[8'h7C][10:8];
        exeReqReg_24_bits_ffo = _RANDOM[8'h7C][11];
        exeReqReg_25_valid = _RANDOM[8'h7C][12];
        exeReqReg_25_bits_source1 = {_RANDOM[8'h7C][31:13], _RANDOM[8'h7D][12:0]};
        exeReqReg_25_bits_source2 = {_RANDOM[8'h7D][31:13], _RANDOM[8'h7E][12:0]};
        exeReqReg_25_bits_index = _RANDOM[8'h7E][15:13];
        exeReqReg_25_bits_ffo = _RANDOM[8'h7E][16];
        exeReqReg_26_valid = _RANDOM[8'h7E][17];
        exeReqReg_26_bits_source1 = {_RANDOM[8'h7E][31:18], _RANDOM[8'h7F][17:0]};
        exeReqReg_26_bits_source2 = {_RANDOM[8'h7F][31:18], _RANDOM[8'h80][17:0]};
        exeReqReg_26_bits_index = _RANDOM[8'h80][20:18];
        exeReqReg_26_bits_ffo = _RANDOM[8'h80][21];
        exeReqReg_27_valid = _RANDOM[8'h80][22];
        exeReqReg_27_bits_source1 = {_RANDOM[8'h80][31:23], _RANDOM[8'h81][22:0]};
        exeReqReg_27_bits_source2 = {_RANDOM[8'h81][31:23], _RANDOM[8'h82][22:0]};
        exeReqReg_27_bits_index = _RANDOM[8'h82][25:23];
        exeReqReg_27_bits_ffo = _RANDOM[8'h82][26];
        exeReqReg_28_valid = _RANDOM[8'h82][27];
        exeReqReg_28_bits_source1 = {_RANDOM[8'h82][31:28], _RANDOM[8'h83][27:0]};
        exeReqReg_28_bits_source2 = {_RANDOM[8'h83][31:28], _RANDOM[8'h84][27:0]};
        exeReqReg_28_bits_index = _RANDOM[8'h84][30:28];
        exeReqReg_28_bits_ffo = _RANDOM[8'h84][31];
        exeReqReg_29_valid = _RANDOM[8'h85][0];
        exeReqReg_29_bits_source1 = {_RANDOM[8'h85][31:1], _RANDOM[8'h86][0]};
        exeReqReg_29_bits_source2 = {_RANDOM[8'h86][31:1], _RANDOM[8'h87][0]};
        exeReqReg_29_bits_index = _RANDOM[8'h87][3:1];
        exeReqReg_29_bits_ffo = _RANDOM[8'h87][4];
        exeReqReg_30_valid = _RANDOM[8'h87][5];
        exeReqReg_30_bits_source1 = {_RANDOM[8'h87][31:6], _RANDOM[8'h88][5:0]};
        exeReqReg_30_bits_source2 = {_RANDOM[8'h88][31:6], _RANDOM[8'h89][5:0]};
        exeReqReg_30_bits_index = _RANDOM[8'h89][8:6];
        exeReqReg_30_bits_ffo = _RANDOM[8'h89][9];
        exeReqReg_31_valid = _RANDOM[8'h89][10];
        exeReqReg_31_bits_source1 = {_RANDOM[8'h89][31:11], _RANDOM[8'h8A][10:0]};
        exeReqReg_31_bits_source2 = {_RANDOM[8'h8A][31:11], _RANDOM[8'h8B][10:0]};
        exeReqReg_31_bits_index = _RANDOM[8'h8B][13:11];
        exeReqReg_31_bits_ffo = _RANDOM[8'h8B][14];
        requestCounter = _RANDOM[8'h8B][19:15];
        executeIndex = _RANDOM[8'h8B][21:20];
        readIssueStageState_groupReadState = {_RANDOM[8'h8B][31:22], _RANDOM[8'h8C][21:0]};
        readIssueStageState_needRead = {_RANDOM[8'h8C][31:22], _RANDOM[8'h8D][21:0]};
        readIssueStageState_elementValid = {_RANDOM[8'h8D][31:22], _RANDOM[8'h8E][21:0]};
        readIssueStageState_replaceVs1 = {_RANDOM[8'h8E][31:22], _RANDOM[8'h8F][21:0]};
        readIssueStageState_readOffset = {_RANDOM[8'h8F][31:22], _RANDOM[8'h90][21:0]};
        readIssueStageState_accessLane_0 = _RANDOM[8'h90][26:22];
        readIssueStageState_accessLane_1 = _RANDOM[8'h90][31:27];
        readIssueStageState_accessLane_2 = _RANDOM[8'h91][4:0];
        readIssueStageState_accessLane_3 = _RANDOM[8'h91][9:5];
        readIssueStageState_accessLane_4 = _RANDOM[8'h91][14:10];
        readIssueStageState_accessLane_5 = _RANDOM[8'h91][19:15];
        readIssueStageState_accessLane_6 = _RANDOM[8'h91][24:20];
        readIssueStageState_accessLane_7 = _RANDOM[8'h91][29:25];
        readIssueStageState_accessLane_8 = {_RANDOM[8'h91][31:30], _RANDOM[8'h92][2:0]};
        readIssueStageState_accessLane_9 = _RANDOM[8'h92][7:3];
        readIssueStageState_accessLane_10 = _RANDOM[8'h92][12:8];
        readIssueStageState_accessLane_11 = _RANDOM[8'h92][17:13];
        readIssueStageState_accessLane_12 = _RANDOM[8'h92][22:18];
        readIssueStageState_accessLane_13 = _RANDOM[8'h92][27:23];
        readIssueStageState_accessLane_14 = {_RANDOM[8'h92][31:28], _RANDOM[8'h93][0]};
        readIssueStageState_accessLane_15 = _RANDOM[8'h93][5:1];
        readIssueStageState_accessLane_16 = _RANDOM[8'h93][10:6];
        readIssueStageState_accessLane_17 = _RANDOM[8'h93][15:11];
        readIssueStageState_accessLane_18 = _RANDOM[8'h93][20:16];
        readIssueStageState_accessLane_19 = _RANDOM[8'h93][25:21];
        readIssueStageState_accessLane_20 = _RANDOM[8'h93][30:26];
        readIssueStageState_accessLane_21 = {_RANDOM[8'h93][31], _RANDOM[8'h94][3:0]};
        readIssueStageState_accessLane_22 = _RANDOM[8'h94][8:4];
        readIssueStageState_accessLane_23 = _RANDOM[8'h94][13:9];
        readIssueStageState_accessLane_24 = _RANDOM[8'h94][18:14];
        readIssueStageState_accessLane_25 = _RANDOM[8'h94][23:19];
        readIssueStageState_accessLane_26 = _RANDOM[8'h94][28:24];
        readIssueStageState_accessLane_27 = {_RANDOM[8'h94][31:29], _RANDOM[8'h95][1:0]};
        readIssueStageState_accessLane_28 = _RANDOM[8'h95][6:2];
        readIssueStageState_accessLane_29 = _RANDOM[8'h95][11:7];
        readIssueStageState_accessLane_30 = _RANDOM[8'h95][16:12];
        readIssueStageState_accessLane_31 = _RANDOM[8'h95][21:17];
        readIssueStageState_vsGrowth_0 = _RANDOM[8'h95][24:22];
        readIssueStageState_vsGrowth_1 = _RANDOM[8'h95][27:25];
        readIssueStageState_vsGrowth_2 = _RANDOM[8'h95][30:28];
        readIssueStageState_vsGrowth_3 = {_RANDOM[8'h95][31], _RANDOM[8'h96][1:0]};
        readIssueStageState_vsGrowth_4 = _RANDOM[8'h96][4:2];
        readIssueStageState_vsGrowth_5 = _RANDOM[8'h96][7:5];
        readIssueStageState_vsGrowth_6 = _RANDOM[8'h96][10:8];
        readIssueStageState_vsGrowth_7 = _RANDOM[8'h96][13:11];
        readIssueStageState_vsGrowth_8 = _RANDOM[8'h96][16:14];
        readIssueStageState_vsGrowth_9 = _RANDOM[8'h96][19:17];
        readIssueStageState_vsGrowth_10 = _RANDOM[8'h96][22:20];
        readIssueStageState_vsGrowth_11 = _RANDOM[8'h96][25:23];
        readIssueStageState_vsGrowth_12 = _RANDOM[8'h96][28:26];
        readIssueStageState_vsGrowth_13 = _RANDOM[8'h96][31:29];
        readIssueStageState_vsGrowth_14 = _RANDOM[8'h97][2:0];
        readIssueStageState_vsGrowth_15 = _RANDOM[8'h97][5:3];
        readIssueStageState_vsGrowth_16 = _RANDOM[8'h97][8:6];
        readIssueStageState_vsGrowth_17 = _RANDOM[8'h97][11:9];
        readIssueStageState_vsGrowth_18 = _RANDOM[8'h97][14:12];
        readIssueStageState_vsGrowth_19 = _RANDOM[8'h97][17:15];
        readIssueStageState_vsGrowth_20 = _RANDOM[8'h97][20:18];
        readIssueStageState_vsGrowth_21 = _RANDOM[8'h97][23:21];
        readIssueStageState_vsGrowth_22 = _RANDOM[8'h97][26:24];
        readIssueStageState_vsGrowth_23 = _RANDOM[8'h97][29:27];
        readIssueStageState_vsGrowth_24 = {_RANDOM[8'h97][31:30], _RANDOM[8'h98][0]};
        readIssueStageState_vsGrowth_25 = _RANDOM[8'h98][3:1];
        readIssueStageState_vsGrowth_26 = _RANDOM[8'h98][6:4];
        readIssueStageState_vsGrowth_27 = _RANDOM[8'h98][9:7];
        readIssueStageState_vsGrowth_28 = _RANDOM[8'h98][12:10];
        readIssueStageState_vsGrowth_29 = _RANDOM[8'h98][15:13];
        readIssueStageState_vsGrowth_30 = _RANDOM[8'h98][18:16];
        readIssueStageState_vsGrowth_31 = _RANDOM[8'h98][21:19];
        readIssueStageState_executeGroup = _RANDOM[8'h98][28:22];
        readIssueStageState_readDataOffset = {_RANDOM[8'h98][31:29], _RANDOM[8'h99], _RANDOM[8'h9A][28:0]};
        readIssueStageState_last = _RANDOM[8'h9A][29];
        readIssueStageValid = _RANDOM[8'h9A][30];
        tokenCheck_counter = {_RANDOM[8'h9A][31], _RANDOM[8'h9B][2:0]};
        tokenCheck_counter_1 = _RANDOM[8'h9B][6:3];
        tokenCheck_counter_2 = _RANDOM[8'h9B][10:7];
        tokenCheck_counter_3 = _RANDOM[8'h9B][14:11];
        tokenCheck_counter_4 = _RANDOM[8'h9B][18:15];
        tokenCheck_counter_5 = _RANDOM[8'h9B][22:19];
        tokenCheck_counter_6 = _RANDOM[8'h9B][26:23];
        tokenCheck_counter_7 = _RANDOM[8'h9B][30:27];
        tokenCheck_counter_8 = {_RANDOM[8'h9B][31], _RANDOM[8'h9C][2:0]};
        tokenCheck_counter_9 = _RANDOM[8'h9C][6:3];
        tokenCheck_counter_10 = _RANDOM[8'h9C][10:7];
        tokenCheck_counter_11 = _RANDOM[8'h9C][14:11];
        tokenCheck_counter_12 = _RANDOM[8'h9C][18:15];
        tokenCheck_counter_13 = _RANDOM[8'h9C][22:19];
        tokenCheck_counter_14 = _RANDOM[8'h9C][26:23];
        tokenCheck_counter_15 = _RANDOM[8'h9C][30:27];
        tokenCheck_counter_16 = {_RANDOM[8'h9C][31], _RANDOM[8'h9D][2:0]};
        tokenCheck_counter_17 = _RANDOM[8'h9D][6:3];
        tokenCheck_counter_18 = _RANDOM[8'h9D][10:7];
        tokenCheck_counter_19 = _RANDOM[8'h9D][14:11];
        tokenCheck_counter_20 = _RANDOM[8'h9D][18:15];
        tokenCheck_counter_21 = _RANDOM[8'h9D][22:19];
        tokenCheck_counter_22 = _RANDOM[8'h9D][26:23];
        tokenCheck_counter_23 = _RANDOM[8'h9D][30:27];
        tokenCheck_counter_24 = {_RANDOM[8'h9D][31], _RANDOM[8'h9E][2:0]};
        tokenCheck_counter_25 = _RANDOM[8'h9E][6:3];
        tokenCheck_counter_26 = _RANDOM[8'h9E][10:7];
        tokenCheck_counter_27 = _RANDOM[8'h9E][14:11];
        tokenCheck_counter_28 = _RANDOM[8'h9E][18:15];
        tokenCheck_counter_29 = _RANDOM[8'h9E][22:19];
        tokenCheck_counter_30 = _RANDOM[8'h9E][26:23];
        tokenCheck_counter_31 = _RANDOM[8'h9E][30:27];
        reorderQueueAllocate_counter = {_RANDOM[8'h9E][31], _RANDOM[8'h9F][5:0]};
        reorderQueueAllocate_counterWillUpdate = _RANDOM[8'h9F][12:6];
        reorderQueueAllocate_counter_1 = _RANDOM[8'h9F][19:13];
        reorderQueueAllocate_counterWillUpdate_1 = _RANDOM[8'h9F][26:20];
        reorderQueueAllocate_counter_2 = {_RANDOM[8'h9F][31:27], _RANDOM[8'hA0][1:0]};
        reorderQueueAllocate_counterWillUpdate_2 = _RANDOM[8'hA0][8:2];
        reorderQueueAllocate_counter_3 = _RANDOM[8'hA0][15:9];
        reorderQueueAllocate_counterWillUpdate_3 = _RANDOM[8'hA0][22:16];
        reorderQueueAllocate_counter_4 = _RANDOM[8'hA0][29:23];
        reorderQueueAllocate_counterWillUpdate_4 = {_RANDOM[8'hA0][31:30], _RANDOM[8'hA1][4:0]};
        reorderQueueAllocate_counter_5 = _RANDOM[8'hA1][11:5];
        reorderQueueAllocate_counterWillUpdate_5 = _RANDOM[8'hA1][18:12];
        reorderQueueAllocate_counter_6 = _RANDOM[8'hA1][25:19];
        reorderQueueAllocate_counterWillUpdate_6 = {_RANDOM[8'hA1][31:26], _RANDOM[8'hA2][0]};
        reorderQueueAllocate_counter_7 = _RANDOM[8'hA2][7:1];
        reorderQueueAllocate_counterWillUpdate_7 = _RANDOM[8'hA2][14:8];
        reorderQueueAllocate_counter_8 = _RANDOM[8'hA2][21:15];
        reorderQueueAllocate_counterWillUpdate_8 = _RANDOM[8'hA2][28:22];
        reorderQueueAllocate_counter_9 = {_RANDOM[8'hA2][31:29], _RANDOM[8'hA3][3:0]};
        reorderQueueAllocate_counterWillUpdate_9 = _RANDOM[8'hA3][10:4];
        reorderQueueAllocate_counter_10 = _RANDOM[8'hA3][17:11];
        reorderQueueAllocate_counterWillUpdate_10 = _RANDOM[8'hA3][24:18];
        reorderQueueAllocate_counter_11 = _RANDOM[8'hA3][31:25];
        reorderQueueAllocate_counterWillUpdate_11 = _RANDOM[8'hA4][6:0];
        reorderQueueAllocate_counter_12 = _RANDOM[8'hA4][13:7];
        reorderQueueAllocate_counterWillUpdate_12 = _RANDOM[8'hA4][20:14];
        reorderQueueAllocate_counter_13 = _RANDOM[8'hA4][27:21];
        reorderQueueAllocate_counterWillUpdate_13 = {_RANDOM[8'hA4][31:28], _RANDOM[8'hA5][2:0]};
        reorderQueueAllocate_counter_14 = _RANDOM[8'hA5][9:3];
        reorderQueueAllocate_counterWillUpdate_14 = _RANDOM[8'hA5][16:10];
        reorderQueueAllocate_counter_15 = _RANDOM[8'hA5][23:17];
        reorderQueueAllocate_counterWillUpdate_15 = _RANDOM[8'hA5][30:24];
        reorderQueueAllocate_counter_16 = {_RANDOM[8'hA5][31], _RANDOM[8'hA6][5:0]};
        reorderQueueAllocate_counterWillUpdate_16 = _RANDOM[8'hA6][12:6];
        reorderQueueAllocate_counter_17 = _RANDOM[8'hA6][19:13];
        reorderQueueAllocate_counterWillUpdate_17 = _RANDOM[8'hA6][26:20];
        reorderQueueAllocate_counter_18 = {_RANDOM[8'hA6][31:27], _RANDOM[8'hA7][1:0]};
        reorderQueueAllocate_counterWillUpdate_18 = _RANDOM[8'hA7][8:2];
        reorderQueueAllocate_counter_19 = _RANDOM[8'hA7][15:9];
        reorderQueueAllocate_counterWillUpdate_19 = _RANDOM[8'hA7][22:16];
        reorderQueueAllocate_counter_20 = _RANDOM[8'hA7][29:23];
        reorderQueueAllocate_counterWillUpdate_20 = {_RANDOM[8'hA7][31:30], _RANDOM[8'hA8][4:0]};
        reorderQueueAllocate_counter_21 = _RANDOM[8'hA8][11:5];
        reorderQueueAllocate_counterWillUpdate_21 = _RANDOM[8'hA8][18:12];
        reorderQueueAllocate_counter_22 = _RANDOM[8'hA8][25:19];
        reorderQueueAllocate_counterWillUpdate_22 = {_RANDOM[8'hA8][31:26], _RANDOM[8'hA9][0]};
        reorderQueueAllocate_counter_23 = _RANDOM[8'hA9][7:1];
        reorderQueueAllocate_counterWillUpdate_23 = _RANDOM[8'hA9][14:8];
        reorderQueueAllocate_counter_24 = _RANDOM[8'hA9][21:15];
        reorderQueueAllocate_counterWillUpdate_24 = _RANDOM[8'hA9][28:22];
        reorderQueueAllocate_counter_25 = {_RANDOM[8'hA9][31:29], _RANDOM[8'hAA][3:0]};
        reorderQueueAllocate_counterWillUpdate_25 = _RANDOM[8'hAA][10:4];
        reorderQueueAllocate_counter_26 = _RANDOM[8'hAA][17:11];
        reorderQueueAllocate_counterWillUpdate_26 = _RANDOM[8'hAA][24:18];
        reorderQueueAllocate_counter_27 = _RANDOM[8'hAA][31:25];
        reorderQueueAllocate_counterWillUpdate_27 = _RANDOM[8'hAB][6:0];
        reorderQueueAllocate_counter_28 = _RANDOM[8'hAB][13:7];
        reorderQueueAllocate_counterWillUpdate_28 = _RANDOM[8'hAB][20:14];
        reorderQueueAllocate_counter_29 = _RANDOM[8'hAB][27:21];
        reorderQueueAllocate_counterWillUpdate_29 = {_RANDOM[8'hAB][31:28], _RANDOM[8'hAC][2:0]};
        reorderQueueAllocate_counter_30 = _RANDOM[8'hAC][9:3];
        reorderQueueAllocate_counterWillUpdate_30 = _RANDOM[8'hAC][16:10];
        reorderQueueAllocate_counter_31 = _RANDOM[8'hAC][23:17];
        reorderQueueAllocate_counterWillUpdate_31 = _RANDOM[8'hAC][30:24];
        reorderStageValid = _RANDOM[8'hAC][31];
        reorderStageState_0 = _RANDOM[8'hAD][5:0];
        reorderStageState_1 = _RANDOM[8'hAD][11:6];
        reorderStageState_2 = _RANDOM[8'hAD][17:12];
        reorderStageState_3 = _RANDOM[8'hAD][23:18];
        reorderStageState_4 = _RANDOM[8'hAD][29:24];
        reorderStageState_5 = {_RANDOM[8'hAD][31:30], _RANDOM[8'hAE][3:0]};
        reorderStageState_6 = _RANDOM[8'hAE][9:4];
        reorderStageState_7 = _RANDOM[8'hAE][15:10];
        reorderStageState_8 = _RANDOM[8'hAE][21:16];
        reorderStageState_9 = _RANDOM[8'hAE][27:22];
        reorderStageState_10 = {_RANDOM[8'hAE][31:28], _RANDOM[8'hAF][1:0]};
        reorderStageState_11 = _RANDOM[8'hAF][7:2];
        reorderStageState_12 = _RANDOM[8'hAF][13:8];
        reorderStageState_13 = _RANDOM[8'hAF][19:14];
        reorderStageState_14 = _RANDOM[8'hAF][25:20];
        reorderStageState_15 = _RANDOM[8'hAF][31:26];
        reorderStageState_16 = _RANDOM[8'hB0][5:0];
        reorderStageState_17 = _RANDOM[8'hB0][11:6];
        reorderStageState_18 = _RANDOM[8'hB0][17:12];
        reorderStageState_19 = _RANDOM[8'hB0][23:18];
        reorderStageState_20 = _RANDOM[8'hB0][29:24];
        reorderStageState_21 = {_RANDOM[8'hB0][31:30], _RANDOM[8'hB1][3:0]};
        reorderStageState_22 = _RANDOM[8'hB1][9:4];
        reorderStageState_23 = _RANDOM[8'hB1][15:10];
        reorderStageState_24 = _RANDOM[8'hB1][21:16];
        reorderStageState_25 = _RANDOM[8'hB1][27:22];
        reorderStageState_26 = {_RANDOM[8'hB1][31:28], _RANDOM[8'hB2][1:0]};
        reorderStageState_27 = _RANDOM[8'hB2][7:2];
        reorderStageState_28 = _RANDOM[8'hB2][13:8];
        reorderStageState_29 = _RANDOM[8'hB2][19:14];
        reorderStageState_30 = _RANDOM[8'hB2][25:20];
        reorderStageState_31 = _RANDOM[8'hB2][31:26];
        reorderStageNeed_0 = _RANDOM[8'hB3][5:0];
        reorderStageNeed_1 = _RANDOM[8'hB3][11:6];
        reorderStageNeed_2 = _RANDOM[8'hB3][17:12];
        reorderStageNeed_3 = _RANDOM[8'hB3][23:18];
        reorderStageNeed_4 = _RANDOM[8'hB3][29:24];
        reorderStageNeed_5 = {_RANDOM[8'hB3][31:30], _RANDOM[8'hB4][3:0]};
        reorderStageNeed_6 = _RANDOM[8'hB4][9:4];
        reorderStageNeed_7 = _RANDOM[8'hB4][15:10];
        reorderStageNeed_8 = _RANDOM[8'hB4][21:16];
        reorderStageNeed_9 = _RANDOM[8'hB4][27:22];
        reorderStageNeed_10 = {_RANDOM[8'hB4][31:28], _RANDOM[8'hB5][1:0]};
        reorderStageNeed_11 = _RANDOM[8'hB5][7:2];
        reorderStageNeed_12 = _RANDOM[8'hB5][13:8];
        reorderStageNeed_13 = _RANDOM[8'hB5][19:14];
        reorderStageNeed_14 = _RANDOM[8'hB5][25:20];
        reorderStageNeed_15 = _RANDOM[8'hB5][31:26];
        reorderStageNeed_16 = _RANDOM[8'hB6][5:0];
        reorderStageNeed_17 = _RANDOM[8'hB6][11:6];
        reorderStageNeed_18 = _RANDOM[8'hB6][17:12];
        reorderStageNeed_19 = _RANDOM[8'hB6][23:18];
        reorderStageNeed_20 = _RANDOM[8'hB6][29:24];
        reorderStageNeed_21 = {_RANDOM[8'hB6][31:30], _RANDOM[8'hB7][3:0]};
        reorderStageNeed_22 = _RANDOM[8'hB7][9:4];
        reorderStageNeed_23 = _RANDOM[8'hB7][15:10];
        reorderStageNeed_24 = _RANDOM[8'hB7][21:16];
        reorderStageNeed_25 = _RANDOM[8'hB7][27:22];
        reorderStageNeed_26 = {_RANDOM[8'hB7][31:28], _RANDOM[8'hB8][1:0]};
        reorderStageNeed_27 = _RANDOM[8'hB8][7:2];
        reorderStageNeed_28 = _RANDOM[8'hB8][13:8];
        reorderStageNeed_29 = _RANDOM[8'hB8][19:14];
        reorderStageNeed_30 = _RANDOM[8'hB8][25:20];
        reorderStageNeed_31 = _RANDOM[8'hB8][31:26];
        waiteReadDataPipeReg_executeGroup = _RANDOM[8'hB9][6:0];
        waiteReadDataPipeReg_sourceValid = {_RANDOM[8'hB9][31:7], _RANDOM[8'hBA][6:0]};
        waiteReadDataPipeReg_replaceVs1 = {_RANDOM[8'hBA][31:7], _RANDOM[8'hBB][6:0]};
        waiteReadDataPipeReg_needRead = {_RANDOM[8'hBB][31:7], _RANDOM[8'hBC][6:0]};
        waiteReadDataPipeReg_last = _RANDOM[8'hBC][7];
        waiteReadData_0 = {_RANDOM[8'hBC][31:8], _RANDOM[8'hBD][7:0]};
        waiteReadData_1 = {_RANDOM[8'hBD][31:8], _RANDOM[8'hBE][7:0]};
        waiteReadData_2 = {_RANDOM[8'hBE][31:8], _RANDOM[8'hBF][7:0]};
        waiteReadData_3 = {_RANDOM[8'hBF][31:8], _RANDOM[8'hC0][7:0]};
        waiteReadData_4 = {_RANDOM[8'hC0][31:8], _RANDOM[8'hC1][7:0]};
        waiteReadData_5 = {_RANDOM[8'hC1][31:8], _RANDOM[8'hC2][7:0]};
        waiteReadData_6 = {_RANDOM[8'hC2][31:8], _RANDOM[8'hC3][7:0]};
        waiteReadData_7 = {_RANDOM[8'hC3][31:8], _RANDOM[8'hC4][7:0]};
        waiteReadData_8 = {_RANDOM[8'hC4][31:8], _RANDOM[8'hC5][7:0]};
        waiteReadData_9 = {_RANDOM[8'hC5][31:8], _RANDOM[8'hC6][7:0]};
        waiteReadData_10 = {_RANDOM[8'hC6][31:8], _RANDOM[8'hC7][7:0]};
        waiteReadData_11 = {_RANDOM[8'hC7][31:8], _RANDOM[8'hC8][7:0]};
        waiteReadData_12 = {_RANDOM[8'hC8][31:8], _RANDOM[8'hC9][7:0]};
        waiteReadData_13 = {_RANDOM[8'hC9][31:8], _RANDOM[8'hCA][7:0]};
        waiteReadData_14 = {_RANDOM[8'hCA][31:8], _RANDOM[8'hCB][7:0]};
        waiteReadData_15 = {_RANDOM[8'hCB][31:8], _RANDOM[8'hCC][7:0]};
        waiteReadData_16 = {_RANDOM[8'hCC][31:8], _RANDOM[8'hCD][7:0]};
        waiteReadData_17 = {_RANDOM[8'hCD][31:8], _RANDOM[8'hCE][7:0]};
        waiteReadData_18 = {_RANDOM[8'hCE][31:8], _RANDOM[8'hCF][7:0]};
        waiteReadData_19 = {_RANDOM[8'hCF][31:8], _RANDOM[8'hD0][7:0]};
        waiteReadData_20 = {_RANDOM[8'hD0][31:8], _RANDOM[8'hD1][7:0]};
        waiteReadData_21 = {_RANDOM[8'hD1][31:8], _RANDOM[8'hD2][7:0]};
        waiteReadData_22 = {_RANDOM[8'hD2][31:8], _RANDOM[8'hD3][7:0]};
        waiteReadData_23 = {_RANDOM[8'hD3][31:8], _RANDOM[8'hD4][7:0]};
        waiteReadData_24 = {_RANDOM[8'hD4][31:8], _RANDOM[8'hD5][7:0]};
        waiteReadData_25 = {_RANDOM[8'hD5][31:8], _RANDOM[8'hD6][7:0]};
        waiteReadData_26 = {_RANDOM[8'hD6][31:8], _RANDOM[8'hD7][7:0]};
        waiteReadData_27 = {_RANDOM[8'hD7][31:8], _RANDOM[8'hD8][7:0]};
        waiteReadData_28 = {_RANDOM[8'hD8][31:8], _RANDOM[8'hD9][7:0]};
        waiteReadData_29 = {_RANDOM[8'hD9][31:8], _RANDOM[8'hDA][7:0]};
        waiteReadData_30 = {_RANDOM[8'hDA][31:8], _RANDOM[8'hDB][7:0]};
        waiteReadData_31 = {_RANDOM[8'hDB][31:8], _RANDOM[8'hDC][7:0]};
        waiteReadSate = {_RANDOM[8'hDC][31:8], _RANDOM[8'hDD][7:0]};
        waiteReadStageValid = _RANDOM[8'hDD][8];
        dataNotInShifter_writeTokenCounter = _RANDOM[8'hDD][11:9];
        dataNotInShifter_writeTokenCounter_1 = _RANDOM[8'hDD][14:12];
        dataNotInShifter_writeTokenCounter_2 = _RANDOM[8'hDD][17:15];
        dataNotInShifter_writeTokenCounter_3 = _RANDOM[8'hDD][20:18];
        dataNotInShifter_writeTokenCounter_4 = _RANDOM[8'hDD][23:21];
        dataNotInShifter_writeTokenCounter_5 = _RANDOM[8'hDD][26:24];
        dataNotInShifter_writeTokenCounter_6 = _RANDOM[8'hDD][29:27];
        dataNotInShifter_writeTokenCounter_7 = {_RANDOM[8'hDD][31:30], _RANDOM[8'hDE][0]};
        dataNotInShifter_writeTokenCounter_8 = _RANDOM[8'hDE][3:1];
        dataNotInShifter_writeTokenCounter_9 = _RANDOM[8'hDE][6:4];
        dataNotInShifter_writeTokenCounter_10 = _RANDOM[8'hDE][9:7];
        dataNotInShifter_writeTokenCounter_11 = _RANDOM[8'hDE][12:10];
        dataNotInShifter_writeTokenCounter_12 = _RANDOM[8'hDE][15:13];
        dataNotInShifter_writeTokenCounter_13 = _RANDOM[8'hDE][18:16];
        dataNotInShifter_writeTokenCounter_14 = _RANDOM[8'hDE][21:19];
        dataNotInShifter_writeTokenCounter_15 = _RANDOM[8'hDE][24:22];
        dataNotInShifter_writeTokenCounter_16 = _RANDOM[8'hDE][27:25];
        dataNotInShifter_writeTokenCounter_17 = _RANDOM[8'hDE][30:28];
        dataNotInShifter_writeTokenCounter_18 = {_RANDOM[8'hDE][31], _RANDOM[8'hDF][1:0]};
        dataNotInShifter_writeTokenCounter_19 = _RANDOM[8'hDF][4:2];
        dataNotInShifter_writeTokenCounter_20 = _RANDOM[8'hDF][7:5];
        dataNotInShifter_writeTokenCounter_21 = _RANDOM[8'hDF][10:8];
        dataNotInShifter_writeTokenCounter_22 = _RANDOM[8'hDF][13:11];
        dataNotInShifter_writeTokenCounter_23 = _RANDOM[8'hDF][16:14];
        dataNotInShifter_writeTokenCounter_24 = _RANDOM[8'hDF][19:17];
        dataNotInShifter_writeTokenCounter_25 = _RANDOM[8'hDF][22:20];
        dataNotInShifter_writeTokenCounter_26 = _RANDOM[8'hDF][25:23];
        dataNotInShifter_writeTokenCounter_27 = _RANDOM[8'hDF][28:26];
        dataNotInShifter_writeTokenCounter_28 = _RANDOM[8'hDF][31:29];
        dataNotInShifter_writeTokenCounter_29 = _RANDOM[8'hE0][2:0];
        dataNotInShifter_writeTokenCounter_30 = _RANDOM[8'hE0][5:3];
        dataNotInShifter_writeTokenCounter_31 = _RANDOM[8'hE0][8:6];
        waiteLastRequest = _RANDOM[8'hE0][9];
        waitQueueClear = _RANDOM[8'hE0][10];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  wire               exeRequestQueue_0_empty;
  assign exeRequestQueue_0_empty = _exeRequestQueue_queue_fifo_empty;
  wire               exeRequestQueue_0_full;
  assign exeRequestQueue_0_full = _exeRequestQueue_queue_fifo_full;
  wire               exeRequestQueue_1_empty;
  assign exeRequestQueue_1_empty = _exeRequestQueue_queue_fifo_1_empty;
  wire               exeRequestQueue_1_full;
  assign exeRequestQueue_1_full = _exeRequestQueue_queue_fifo_1_full;
  wire               exeRequestQueue_2_empty;
  assign exeRequestQueue_2_empty = _exeRequestQueue_queue_fifo_2_empty;
  wire               exeRequestQueue_2_full;
  assign exeRequestQueue_2_full = _exeRequestQueue_queue_fifo_2_full;
  wire               exeRequestQueue_3_empty;
  assign exeRequestQueue_3_empty = _exeRequestQueue_queue_fifo_3_empty;
  wire               exeRequestQueue_3_full;
  assign exeRequestQueue_3_full = _exeRequestQueue_queue_fifo_3_full;
  wire               exeRequestQueue_4_empty;
  assign exeRequestQueue_4_empty = _exeRequestQueue_queue_fifo_4_empty;
  wire               exeRequestQueue_4_full;
  assign exeRequestQueue_4_full = _exeRequestQueue_queue_fifo_4_full;
  wire               exeRequestQueue_5_empty;
  assign exeRequestQueue_5_empty = _exeRequestQueue_queue_fifo_5_empty;
  wire               exeRequestQueue_5_full;
  assign exeRequestQueue_5_full = _exeRequestQueue_queue_fifo_5_full;
  wire               exeRequestQueue_6_empty;
  assign exeRequestQueue_6_empty = _exeRequestQueue_queue_fifo_6_empty;
  wire               exeRequestQueue_6_full;
  assign exeRequestQueue_6_full = _exeRequestQueue_queue_fifo_6_full;
  wire               exeRequestQueue_7_empty;
  assign exeRequestQueue_7_empty = _exeRequestQueue_queue_fifo_7_empty;
  wire               exeRequestQueue_7_full;
  assign exeRequestQueue_7_full = _exeRequestQueue_queue_fifo_7_full;
  wire               exeRequestQueue_8_empty;
  assign exeRequestQueue_8_empty = _exeRequestQueue_queue_fifo_8_empty;
  wire               exeRequestQueue_8_full;
  assign exeRequestQueue_8_full = _exeRequestQueue_queue_fifo_8_full;
  wire               exeRequestQueue_9_empty;
  assign exeRequestQueue_9_empty = _exeRequestQueue_queue_fifo_9_empty;
  wire               exeRequestQueue_9_full;
  assign exeRequestQueue_9_full = _exeRequestQueue_queue_fifo_9_full;
  wire               exeRequestQueue_10_empty;
  assign exeRequestQueue_10_empty = _exeRequestQueue_queue_fifo_10_empty;
  wire               exeRequestQueue_10_full;
  assign exeRequestQueue_10_full = _exeRequestQueue_queue_fifo_10_full;
  wire               exeRequestQueue_11_empty;
  assign exeRequestQueue_11_empty = _exeRequestQueue_queue_fifo_11_empty;
  wire               exeRequestQueue_11_full;
  assign exeRequestQueue_11_full = _exeRequestQueue_queue_fifo_11_full;
  wire               exeRequestQueue_12_empty;
  assign exeRequestQueue_12_empty = _exeRequestQueue_queue_fifo_12_empty;
  wire               exeRequestQueue_12_full;
  assign exeRequestQueue_12_full = _exeRequestQueue_queue_fifo_12_full;
  wire               exeRequestQueue_13_empty;
  assign exeRequestQueue_13_empty = _exeRequestQueue_queue_fifo_13_empty;
  wire               exeRequestQueue_13_full;
  assign exeRequestQueue_13_full = _exeRequestQueue_queue_fifo_13_full;
  wire               exeRequestQueue_14_empty;
  assign exeRequestQueue_14_empty = _exeRequestQueue_queue_fifo_14_empty;
  wire               exeRequestQueue_14_full;
  assign exeRequestQueue_14_full = _exeRequestQueue_queue_fifo_14_full;
  wire               exeRequestQueue_15_empty;
  assign exeRequestQueue_15_empty = _exeRequestQueue_queue_fifo_15_empty;
  wire               exeRequestQueue_15_full;
  assign exeRequestQueue_15_full = _exeRequestQueue_queue_fifo_15_full;
  wire               exeRequestQueue_16_empty;
  assign exeRequestQueue_16_empty = _exeRequestQueue_queue_fifo_16_empty;
  wire               exeRequestQueue_16_full;
  assign exeRequestQueue_16_full = _exeRequestQueue_queue_fifo_16_full;
  wire               exeRequestQueue_17_empty;
  assign exeRequestQueue_17_empty = _exeRequestQueue_queue_fifo_17_empty;
  wire               exeRequestQueue_17_full;
  assign exeRequestQueue_17_full = _exeRequestQueue_queue_fifo_17_full;
  wire               exeRequestQueue_18_empty;
  assign exeRequestQueue_18_empty = _exeRequestQueue_queue_fifo_18_empty;
  wire               exeRequestQueue_18_full;
  assign exeRequestQueue_18_full = _exeRequestQueue_queue_fifo_18_full;
  wire               exeRequestQueue_19_empty;
  assign exeRequestQueue_19_empty = _exeRequestQueue_queue_fifo_19_empty;
  wire               exeRequestQueue_19_full;
  assign exeRequestQueue_19_full = _exeRequestQueue_queue_fifo_19_full;
  wire               exeRequestQueue_20_empty;
  assign exeRequestQueue_20_empty = _exeRequestQueue_queue_fifo_20_empty;
  wire               exeRequestQueue_20_full;
  assign exeRequestQueue_20_full = _exeRequestQueue_queue_fifo_20_full;
  wire               exeRequestQueue_21_empty;
  assign exeRequestQueue_21_empty = _exeRequestQueue_queue_fifo_21_empty;
  wire               exeRequestQueue_21_full;
  assign exeRequestQueue_21_full = _exeRequestQueue_queue_fifo_21_full;
  wire               exeRequestQueue_22_empty;
  assign exeRequestQueue_22_empty = _exeRequestQueue_queue_fifo_22_empty;
  wire               exeRequestQueue_22_full;
  assign exeRequestQueue_22_full = _exeRequestQueue_queue_fifo_22_full;
  wire               exeRequestQueue_23_empty;
  assign exeRequestQueue_23_empty = _exeRequestQueue_queue_fifo_23_empty;
  wire               exeRequestQueue_23_full;
  assign exeRequestQueue_23_full = _exeRequestQueue_queue_fifo_23_full;
  wire               exeRequestQueue_24_empty;
  assign exeRequestQueue_24_empty = _exeRequestQueue_queue_fifo_24_empty;
  wire               exeRequestQueue_24_full;
  assign exeRequestQueue_24_full = _exeRequestQueue_queue_fifo_24_full;
  wire               exeRequestQueue_25_empty;
  assign exeRequestQueue_25_empty = _exeRequestQueue_queue_fifo_25_empty;
  wire               exeRequestQueue_25_full;
  assign exeRequestQueue_25_full = _exeRequestQueue_queue_fifo_25_full;
  wire               exeRequestQueue_26_empty;
  assign exeRequestQueue_26_empty = _exeRequestQueue_queue_fifo_26_empty;
  wire               exeRequestQueue_26_full;
  assign exeRequestQueue_26_full = _exeRequestQueue_queue_fifo_26_full;
  wire               exeRequestQueue_27_empty;
  assign exeRequestQueue_27_empty = _exeRequestQueue_queue_fifo_27_empty;
  wire               exeRequestQueue_27_full;
  assign exeRequestQueue_27_full = _exeRequestQueue_queue_fifo_27_full;
  wire               exeRequestQueue_28_empty;
  assign exeRequestQueue_28_empty = _exeRequestQueue_queue_fifo_28_empty;
  wire               exeRequestQueue_28_full;
  assign exeRequestQueue_28_full = _exeRequestQueue_queue_fifo_28_full;
  wire               exeRequestQueue_29_empty;
  assign exeRequestQueue_29_empty = _exeRequestQueue_queue_fifo_29_empty;
  wire               exeRequestQueue_29_full;
  assign exeRequestQueue_29_full = _exeRequestQueue_queue_fifo_29_full;
  wire               exeRequestQueue_30_empty;
  assign exeRequestQueue_30_empty = _exeRequestQueue_queue_fifo_30_empty;
  wire               exeRequestQueue_30_full;
  assign exeRequestQueue_30_full = _exeRequestQueue_queue_fifo_30_full;
  wire               exeRequestQueue_31_empty;
  assign exeRequestQueue_31_empty = _exeRequestQueue_queue_fifo_31_empty;
  wire               exeRequestQueue_31_full;
  assign exeRequestQueue_31_full = _exeRequestQueue_queue_fifo_31_full;
  wire               accessCountQueue_empty;
  assign accessCountQueue_empty = _accessCountQueue_fifo_empty;
  wire               accessCountQueue_full;
  assign accessCountQueue_full = _accessCountQueue_fifo_full;
  wire               readWaitQueue_empty;
  assign readWaitQueue_empty = _readWaitQueue_fifo_empty;
  wire               readWaitQueue_full;
  assign readWaitQueue_full = _readWaitQueue_fifo_full;
  assign compressUnitResultQueue_empty = _compressUnitResultQueue_fifo_empty;
  wire               compressUnitResultQueue_full;
  assign compressUnitResultQueue_full = _compressUnitResultQueue_fifo_full;
  wire               reorderQueueVec_0_empty;
  assign reorderQueueVec_0_empty = _reorderQueueVec_fifo_empty;
  wire               reorderQueueVec_0_full;
  assign reorderQueueVec_0_full = _reorderQueueVec_fifo_full;
  wire               reorderQueueVec_1_empty;
  assign reorderQueueVec_1_empty = _reorderQueueVec_fifo_1_empty;
  wire               reorderQueueVec_1_full;
  assign reorderQueueVec_1_full = _reorderQueueVec_fifo_1_full;
  wire               reorderQueueVec_2_empty;
  assign reorderQueueVec_2_empty = _reorderQueueVec_fifo_2_empty;
  wire               reorderQueueVec_2_full;
  assign reorderQueueVec_2_full = _reorderQueueVec_fifo_2_full;
  wire               reorderQueueVec_3_empty;
  assign reorderQueueVec_3_empty = _reorderQueueVec_fifo_3_empty;
  wire               reorderQueueVec_3_full;
  assign reorderQueueVec_3_full = _reorderQueueVec_fifo_3_full;
  wire               reorderQueueVec_4_empty;
  assign reorderQueueVec_4_empty = _reorderQueueVec_fifo_4_empty;
  wire               reorderQueueVec_4_full;
  assign reorderQueueVec_4_full = _reorderQueueVec_fifo_4_full;
  wire               reorderQueueVec_5_empty;
  assign reorderQueueVec_5_empty = _reorderQueueVec_fifo_5_empty;
  wire               reorderQueueVec_5_full;
  assign reorderQueueVec_5_full = _reorderQueueVec_fifo_5_full;
  wire               reorderQueueVec_6_empty;
  assign reorderQueueVec_6_empty = _reorderQueueVec_fifo_6_empty;
  wire               reorderQueueVec_6_full;
  assign reorderQueueVec_6_full = _reorderQueueVec_fifo_6_full;
  wire               reorderQueueVec_7_empty;
  assign reorderQueueVec_7_empty = _reorderQueueVec_fifo_7_empty;
  wire               reorderQueueVec_7_full;
  assign reorderQueueVec_7_full = _reorderQueueVec_fifo_7_full;
  wire               reorderQueueVec_8_empty;
  assign reorderQueueVec_8_empty = _reorderQueueVec_fifo_8_empty;
  wire               reorderQueueVec_8_full;
  assign reorderQueueVec_8_full = _reorderQueueVec_fifo_8_full;
  wire               reorderQueueVec_9_empty;
  assign reorderQueueVec_9_empty = _reorderQueueVec_fifo_9_empty;
  wire               reorderQueueVec_9_full;
  assign reorderQueueVec_9_full = _reorderQueueVec_fifo_9_full;
  wire               reorderQueueVec_10_empty;
  assign reorderQueueVec_10_empty = _reorderQueueVec_fifo_10_empty;
  wire               reorderQueueVec_10_full;
  assign reorderQueueVec_10_full = _reorderQueueVec_fifo_10_full;
  wire               reorderQueueVec_11_empty;
  assign reorderQueueVec_11_empty = _reorderQueueVec_fifo_11_empty;
  wire               reorderQueueVec_11_full;
  assign reorderQueueVec_11_full = _reorderQueueVec_fifo_11_full;
  wire               reorderQueueVec_12_empty;
  assign reorderQueueVec_12_empty = _reorderQueueVec_fifo_12_empty;
  wire               reorderQueueVec_12_full;
  assign reorderQueueVec_12_full = _reorderQueueVec_fifo_12_full;
  wire               reorderQueueVec_13_empty;
  assign reorderQueueVec_13_empty = _reorderQueueVec_fifo_13_empty;
  wire               reorderQueueVec_13_full;
  assign reorderQueueVec_13_full = _reorderQueueVec_fifo_13_full;
  wire               reorderQueueVec_14_empty;
  assign reorderQueueVec_14_empty = _reorderQueueVec_fifo_14_empty;
  wire               reorderQueueVec_14_full;
  assign reorderQueueVec_14_full = _reorderQueueVec_fifo_14_full;
  wire               reorderQueueVec_15_empty;
  assign reorderQueueVec_15_empty = _reorderQueueVec_fifo_15_empty;
  wire               reorderQueueVec_15_full;
  assign reorderQueueVec_15_full = _reorderQueueVec_fifo_15_full;
  wire               reorderQueueVec_16_empty;
  assign reorderQueueVec_16_empty = _reorderQueueVec_fifo_16_empty;
  wire               reorderQueueVec_16_full;
  assign reorderQueueVec_16_full = _reorderQueueVec_fifo_16_full;
  wire               reorderQueueVec_17_empty;
  assign reorderQueueVec_17_empty = _reorderQueueVec_fifo_17_empty;
  wire               reorderQueueVec_17_full;
  assign reorderQueueVec_17_full = _reorderQueueVec_fifo_17_full;
  wire               reorderQueueVec_18_empty;
  assign reorderQueueVec_18_empty = _reorderQueueVec_fifo_18_empty;
  wire               reorderQueueVec_18_full;
  assign reorderQueueVec_18_full = _reorderQueueVec_fifo_18_full;
  wire               reorderQueueVec_19_empty;
  assign reorderQueueVec_19_empty = _reorderQueueVec_fifo_19_empty;
  wire               reorderQueueVec_19_full;
  assign reorderQueueVec_19_full = _reorderQueueVec_fifo_19_full;
  wire               reorderQueueVec_20_empty;
  assign reorderQueueVec_20_empty = _reorderQueueVec_fifo_20_empty;
  wire               reorderQueueVec_20_full;
  assign reorderQueueVec_20_full = _reorderQueueVec_fifo_20_full;
  wire               reorderQueueVec_21_empty;
  assign reorderQueueVec_21_empty = _reorderQueueVec_fifo_21_empty;
  wire               reorderQueueVec_21_full;
  assign reorderQueueVec_21_full = _reorderQueueVec_fifo_21_full;
  wire               reorderQueueVec_22_empty;
  assign reorderQueueVec_22_empty = _reorderQueueVec_fifo_22_empty;
  wire               reorderQueueVec_22_full;
  assign reorderQueueVec_22_full = _reorderQueueVec_fifo_22_full;
  wire               reorderQueueVec_23_empty;
  assign reorderQueueVec_23_empty = _reorderQueueVec_fifo_23_empty;
  wire               reorderQueueVec_23_full;
  assign reorderQueueVec_23_full = _reorderQueueVec_fifo_23_full;
  wire               reorderQueueVec_24_empty;
  assign reorderQueueVec_24_empty = _reorderQueueVec_fifo_24_empty;
  wire               reorderQueueVec_24_full;
  assign reorderQueueVec_24_full = _reorderQueueVec_fifo_24_full;
  wire               reorderQueueVec_25_empty;
  assign reorderQueueVec_25_empty = _reorderQueueVec_fifo_25_empty;
  wire               reorderQueueVec_25_full;
  assign reorderQueueVec_25_full = _reorderQueueVec_fifo_25_full;
  wire               reorderQueueVec_26_empty;
  assign reorderQueueVec_26_empty = _reorderQueueVec_fifo_26_empty;
  wire               reorderQueueVec_26_full;
  assign reorderQueueVec_26_full = _reorderQueueVec_fifo_26_full;
  wire               reorderQueueVec_27_empty;
  assign reorderQueueVec_27_empty = _reorderQueueVec_fifo_27_empty;
  wire               reorderQueueVec_27_full;
  assign reorderQueueVec_27_full = _reorderQueueVec_fifo_27_full;
  wire               reorderQueueVec_28_empty;
  assign reorderQueueVec_28_empty = _reorderQueueVec_fifo_28_empty;
  wire               reorderQueueVec_28_full;
  assign reorderQueueVec_28_full = _reorderQueueVec_fifo_28_full;
  wire               reorderQueueVec_29_empty;
  assign reorderQueueVec_29_empty = _reorderQueueVec_fifo_29_empty;
  wire               reorderQueueVec_29_full;
  assign reorderQueueVec_29_full = _reorderQueueVec_fifo_29_full;
  wire               reorderQueueVec_30_empty;
  assign reorderQueueVec_30_empty = _reorderQueueVec_fifo_30_empty;
  wire               reorderQueueVec_30_full;
  assign reorderQueueVec_30_full = _reorderQueueVec_fifo_30_full;
  wire               reorderQueueVec_31_empty;
  assign reorderQueueVec_31_empty = _reorderQueueVec_fifo_31_empty;
  wire               reorderQueueVec_31_full;
  assign reorderQueueVec_31_full = _reorderQueueVec_fifo_31_full;
  wire               readMessageQueue_empty;
  assign readMessageQueue_empty = _readMessageQueue_fifo_empty;
  wire               readMessageQueue_full;
  assign readMessageQueue_full = _readMessageQueue_fifo_full;
  wire               readMessageQueue_1_empty;
  assign readMessageQueue_1_empty = _readMessageQueue_fifo_1_empty;
  wire               readMessageQueue_1_full;
  assign readMessageQueue_1_full = _readMessageQueue_fifo_1_full;
  wire               readMessageQueue_2_empty;
  assign readMessageQueue_2_empty = _readMessageQueue_fifo_2_empty;
  wire               readMessageQueue_2_full;
  assign readMessageQueue_2_full = _readMessageQueue_fifo_2_full;
  wire               readMessageQueue_3_empty;
  assign readMessageQueue_3_empty = _readMessageQueue_fifo_3_empty;
  wire               readMessageQueue_3_full;
  assign readMessageQueue_3_full = _readMessageQueue_fifo_3_full;
  wire               readMessageQueue_4_empty;
  assign readMessageQueue_4_empty = _readMessageQueue_fifo_4_empty;
  wire               readMessageQueue_4_full;
  assign readMessageQueue_4_full = _readMessageQueue_fifo_4_full;
  wire               readMessageQueue_5_empty;
  assign readMessageQueue_5_empty = _readMessageQueue_fifo_5_empty;
  wire               readMessageQueue_5_full;
  assign readMessageQueue_5_full = _readMessageQueue_fifo_5_full;
  wire               readMessageQueue_6_empty;
  assign readMessageQueue_6_empty = _readMessageQueue_fifo_6_empty;
  wire               readMessageQueue_6_full;
  assign readMessageQueue_6_full = _readMessageQueue_fifo_6_full;
  wire               readMessageQueue_7_empty;
  assign readMessageQueue_7_empty = _readMessageQueue_fifo_7_empty;
  wire               readMessageQueue_7_full;
  assign readMessageQueue_7_full = _readMessageQueue_fifo_7_full;
  wire               readMessageQueue_8_empty;
  assign readMessageQueue_8_empty = _readMessageQueue_fifo_8_empty;
  wire               readMessageQueue_8_full;
  assign readMessageQueue_8_full = _readMessageQueue_fifo_8_full;
  wire               readMessageQueue_9_empty;
  assign readMessageQueue_9_empty = _readMessageQueue_fifo_9_empty;
  wire               readMessageQueue_9_full;
  assign readMessageQueue_9_full = _readMessageQueue_fifo_9_full;
  wire               readMessageQueue_10_empty;
  assign readMessageQueue_10_empty = _readMessageQueue_fifo_10_empty;
  wire               readMessageQueue_10_full;
  assign readMessageQueue_10_full = _readMessageQueue_fifo_10_full;
  wire               readMessageQueue_11_empty;
  assign readMessageQueue_11_empty = _readMessageQueue_fifo_11_empty;
  wire               readMessageQueue_11_full;
  assign readMessageQueue_11_full = _readMessageQueue_fifo_11_full;
  wire               readMessageQueue_12_empty;
  assign readMessageQueue_12_empty = _readMessageQueue_fifo_12_empty;
  wire               readMessageQueue_12_full;
  assign readMessageQueue_12_full = _readMessageQueue_fifo_12_full;
  wire               readMessageQueue_13_empty;
  assign readMessageQueue_13_empty = _readMessageQueue_fifo_13_empty;
  wire               readMessageQueue_13_full;
  assign readMessageQueue_13_full = _readMessageQueue_fifo_13_full;
  wire               readMessageQueue_14_empty;
  assign readMessageQueue_14_empty = _readMessageQueue_fifo_14_empty;
  wire               readMessageQueue_14_full;
  assign readMessageQueue_14_full = _readMessageQueue_fifo_14_full;
  wire               readMessageQueue_15_empty;
  assign readMessageQueue_15_empty = _readMessageQueue_fifo_15_empty;
  wire               readMessageQueue_15_full;
  assign readMessageQueue_15_full = _readMessageQueue_fifo_15_full;
  wire               readMessageQueue_16_empty;
  assign readMessageQueue_16_empty = _readMessageQueue_fifo_16_empty;
  wire               readMessageQueue_16_full;
  assign readMessageQueue_16_full = _readMessageQueue_fifo_16_full;
  wire               readMessageQueue_17_empty;
  assign readMessageQueue_17_empty = _readMessageQueue_fifo_17_empty;
  wire               readMessageQueue_17_full;
  assign readMessageQueue_17_full = _readMessageQueue_fifo_17_full;
  wire               readMessageQueue_18_empty;
  assign readMessageQueue_18_empty = _readMessageQueue_fifo_18_empty;
  wire               readMessageQueue_18_full;
  assign readMessageQueue_18_full = _readMessageQueue_fifo_18_full;
  wire               readMessageQueue_19_empty;
  assign readMessageQueue_19_empty = _readMessageQueue_fifo_19_empty;
  wire               readMessageQueue_19_full;
  assign readMessageQueue_19_full = _readMessageQueue_fifo_19_full;
  wire               readMessageQueue_20_empty;
  assign readMessageQueue_20_empty = _readMessageQueue_fifo_20_empty;
  wire               readMessageQueue_20_full;
  assign readMessageQueue_20_full = _readMessageQueue_fifo_20_full;
  wire               readMessageQueue_21_empty;
  assign readMessageQueue_21_empty = _readMessageQueue_fifo_21_empty;
  wire               readMessageQueue_21_full;
  assign readMessageQueue_21_full = _readMessageQueue_fifo_21_full;
  wire               readMessageQueue_22_empty;
  assign readMessageQueue_22_empty = _readMessageQueue_fifo_22_empty;
  wire               readMessageQueue_22_full;
  assign readMessageQueue_22_full = _readMessageQueue_fifo_22_full;
  wire               readMessageQueue_23_empty;
  assign readMessageQueue_23_empty = _readMessageQueue_fifo_23_empty;
  wire               readMessageQueue_23_full;
  assign readMessageQueue_23_full = _readMessageQueue_fifo_23_full;
  wire               readMessageQueue_24_empty;
  assign readMessageQueue_24_empty = _readMessageQueue_fifo_24_empty;
  wire               readMessageQueue_24_full;
  assign readMessageQueue_24_full = _readMessageQueue_fifo_24_full;
  wire               readMessageQueue_25_empty;
  assign readMessageQueue_25_empty = _readMessageQueue_fifo_25_empty;
  wire               readMessageQueue_25_full;
  assign readMessageQueue_25_full = _readMessageQueue_fifo_25_full;
  wire               readMessageQueue_26_empty;
  assign readMessageQueue_26_empty = _readMessageQueue_fifo_26_empty;
  wire               readMessageQueue_26_full;
  assign readMessageQueue_26_full = _readMessageQueue_fifo_26_full;
  wire               readMessageQueue_27_empty;
  assign readMessageQueue_27_empty = _readMessageQueue_fifo_27_empty;
  wire               readMessageQueue_27_full;
  assign readMessageQueue_27_full = _readMessageQueue_fifo_27_full;
  wire               readMessageQueue_28_empty;
  assign readMessageQueue_28_empty = _readMessageQueue_fifo_28_empty;
  wire               readMessageQueue_28_full;
  assign readMessageQueue_28_full = _readMessageQueue_fifo_28_full;
  wire               readMessageQueue_29_empty;
  assign readMessageQueue_29_empty = _readMessageQueue_fifo_29_empty;
  wire               readMessageQueue_29_full;
  assign readMessageQueue_29_full = _readMessageQueue_fifo_29_full;
  wire               readMessageQueue_30_empty;
  assign readMessageQueue_30_empty = _readMessageQueue_fifo_30_empty;
  wire               readMessageQueue_30_full;
  assign readMessageQueue_30_full = _readMessageQueue_fifo_30_full;
  wire               readMessageQueue_31_empty;
  assign readMessageQueue_31_empty = _readMessageQueue_fifo_31_empty;
  wire               readMessageQueue_31_full;
  assign readMessageQueue_31_full = _readMessageQueue_fifo_31_full;
  wire               readData_readDataQueue_empty;
  assign readData_readDataQueue_empty = _readData_readDataQueue_fifo_empty;
  wire               readData_readDataQueue_full;
  assign readData_readDataQueue_full = _readData_readDataQueue_fifo_full;
  wire               readData_readDataQueue_1_empty;
  assign readData_readDataQueue_1_empty = _readData_readDataQueue_fifo_1_empty;
  wire               readData_readDataQueue_1_full;
  assign readData_readDataQueue_1_full = _readData_readDataQueue_fifo_1_full;
  wire               readData_readDataQueue_2_empty;
  assign readData_readDataQueue_2_empty = _readData_readDataQueue_fifo_2_empty;
  wire               readData_readDataQueue_2_full;
  assign readData_readDataQueue_2_full = _readData_readDataQueue_fifo_2_full;
  wire               readData_readDataQueue_3_empty;
  assign readData_readDataQueue_3_empty = _readData_readDataQueue_fifo_3_empty;
  wire               readData_readDataQueue_3_full;
  assign readData_readDataQueue_3_full = _readData_readDataQueue_fifo_3_full;
  wire               readData_readDataQueue_4_empty;
  assign readData_readDataQueue_4_empty = _readData_readDataQueue_fifo_4_empty;
  wire               readData_readDataQueue_4_full;
  assign readData_readDataQueue_4_full = _readData_readDataQueue_fifo_4_full;
  wire               readData_readDataQueue_5_empty;
  assign readData_readDataQueue_5_empty = _readData_readDataQueue_fifo_5_empty;
  wire               readData_readDataQueue_5_full;
  assign readData_readDataQueue_5_full = _readData_readDataQueue_fifo_5_full;
  wire               readData_readDataQueue_6_empty;
  assign readData_readDataQueue_6_empty = _readData_readDataQueue_fifo_6_empty;
  wire               readData_readDataQueue_6_full;
  assign readData_readDataQueue_6_full = _readData_readDataQueue_fifo_6_full;
  wire               readData_readDataQueue_7_empty;
  assign readData_readDataQueue_7_empty = _readData_readDataQueue_fifo_7_empty;
  wire               readData_readDataQueue_7_full;
  assign readData_readDataQueue_7_full = _readData_readDataQueue_fifo_7_full;
  wire               readData_readDataQueue_8_empty;
  assign readData_readDataQueue_8_empty = _readData_readDataQueue_fifo_8_empty;
  wire               readData_readDataQueue_8_full;
  assign readData_readDataQueue_8_full = _readData_readDataQueue_fifo_8_full;
  wire               readData_readDataQueue_9_empty;
  assign readData_readDataQueue_9_empty = _readData_readDataQueue_fifo_9_empty;
  wire               readData_readDataQueue_9_full;
  assign readData_readDataQueue_9_full = _readData_readDataQueue_fifo_9_full;
  wire               readData_readDataQueue_10_empty;
  assign readData_readDataQueue_10_empty = _readData_readDataQueue_fifo_10_empty;
  wire               readData_readDataQueue_10_full;
  assign readData_readDataQueue_10_full = _readData_readDataQueue_fifo_10_full;
  wire               readData_readDataQueue_11_empty;
  assign readData_readDataQueue_11_empty = _readData_readDataQueue_fifo_11_empty;
  wire               readData_readDataQueue_11_full;
  assign readData_readDataQueue_11_full = _readData_readDataQueue_fifo_11_full;
  wire               readData_readDataQueue_12_empty;
  assign readData_readDataQueue_12_empty = _readData_readDataQueue_fifo_12_empty;
  wire               readData_readDataQueue_12_full;
  assign readData_readDataQueue_12_full = _readData_readDataQueue_fifo_12_full;
  wire               readData_readDataQueue_13_empty;
  assign readData_readDataQueue_13_empty = _readData_readDataQueue_fifo_13_empty;
  wire               readData_readDataQueue_13_full;
  assign readData_readDataQueue_13_full = _readData_readDataQueue_fifo_13_full;
  wire               readData_readDataQueue_14_empty;
  assign readData_readDataQueue_14_empty = _readData_readDataQueue_fifo_14_empty;
  wire               readData_readDataQueue_14_full;
  assign readData_readDataQueue_14_full = _readData_readDataQueue_fifo_14_full;
  wire               readData_readDataQueue_15_empty;
  assign readData_readDataQueue_15_empty = _readData_readDataQueue_fifo_15_empty;
  wire               readData_readDataQueue_15_full;
  assign readData_readDataQueue_15_full = _readData_readDataQueue_fifo_15_full;
  wire               readData_readDataQueue_16_empty;
  assign readData_readDataQueue_16_empty = _readData_readDataQueue_fifo_16_empty;
  wire               readData_readDataQueue_16_full;
  assign readData_readDataQueue_16_full = _readData_readDataQueue_fifo_16_full;
  wire               readData_readDataQueue_17_empty;
  assign readData_readDataQueue_17_empty = _readData_readDataQueue_fifo_17_empty;
  wire               readData_readDataQueue_17_full;
  assign readData_readDataQueue_17_full = _readData_readDataQueue_fifo_17_full;
  wire               readData_readDataQueue_18_empty;
  assign readData_readDataQueue_18_empty = _readData_readDataQueue_fifo_18_empty;
  wire               readData_readDataQueue_18_full;
  assign readData_readDataQueue_18_full = _readData_readDataQueue_fifo_18_full;
  wire               readData_readDataQueue_19_empty;
  assign readData_readDataQueue_19_empty = _readData_readDataQueue_fifo_19_empty;
  wire               readData_readDataQueue_19_full;
  assign readData_readDataQueue_19_full = _readData_readDataQueue_fifo_19_full;
  wire               readData_readDataQueue_20_empty;
  assign readData_readDataQueue_20_empty = _readData_readDataQueue_fifo_20_empty;
  wire               readData_readDataQueue_20_full;
  assign readData_readDataQueue_20_full = _readData_readDataQueue_fifo_20_full;
  wire               readData_readDataQueue_21_empty;
  assign readData_readDataQueue_21_empty = _readData_readDataQueue_fifo_21_empty;
  wire               readData_readDataQueue_21_full;
  assign readData_readDataQueue_21_full = _readData_readDataQueue_fifo_21_full;
  wire               readData_readDataQueue_22_empty;
  assign readData_readDataQueue_22_empty = _readData_readDataQueue_fifo_22_empty;
  wire               readData_readDataQueue_22_full;
  assign readData_readDataQueue_22_full = _readData_readDataQueue_fifo_22_full;
  wire               readData_readDataQueue_23_empty;
  assign readData_readDataQueue_23_empty = _readData_readDataQueue_fifo_23_empty;
  wire               readData_readDataQueue_23_full;
  assign readData_readDataQueue_23_full = _readData_readDataQueue_fifo_23_full;
  wire               readData_readDataQueue_24_empty;
  assign readData_readDataQueue_24_empty = _readData_readDataQueue_fifo_24_empty;
  wire               readData_readDataQueue_24_full;
  assign readData_readDataQueue_24_full = _readData_readDataQueue_fifo_24_full;
  wire               readData_readDataQueue_25_empty;
  assign readData_readDataQueue_25_empty = _readData_readDataQueue_fifo_25_empty;
  wire               readData_readDataQueue_25_full;
  assign readData_readDataQueue_25_full = _readData_readDataQueue_fifo_25_full;
  wire               readData_readDataQueue_26_empty;
  assign readData_readDataQueue_26_empty = _readData_readDataQueue_fifo_26_empty;
  wire               readData_readDataQueue_26_full;
  assign readData_readDataQueue_26_full = _readData_readDataQueue_fifo_26_full;
  wire               readData_readDataQueue_27_empty;
  assign readData_readDataQueue_27_empty = _readData_readDataQueue_fifo_27_empty;
  wire               readData_readDataQueue_27_full;
  assign readData_readDataQueue_27_full = _readData_readDataQueue_fifo_27_full;
  wire               readData_readDataQueue_28_empty;
  assign readData_readDataQueue_28_empty = _readData_readDataQueue_fifo_28_empty;
  wire               readData_readDataQueue_28_full;
  assign readData_readDataQueue_28_full = _readData_readDataQueue_fifo_28_full;
  wire               readData_readDataQueue_29_empty;
  assign readData_readDataQueue_29_empty = _readData_readDataQueue_fifo_29_empty;
  wire               readData_readDataQueue_29_full;
  assign readData_readDataQueue_29_full = _readData_readDataQueue_fifo_29_full;
  wire               readData_readDataQueue_30_empty;
  assign readData_readDataQueue_30_empty = _readData_readDataQueue_fifo_30_empty;
  wire               readData_readDataQueue_30_full;
  assign readData_readDataQueue_30_full = _readData_readDataQueue_fifo_30_full;
  wire               readData_readDataQueue_31_empty;
  assign readData_readDataQueue_31_empty = _readData_readDataQueue_fifo_31_empty;
  wire               readData_readDataQueue_31_full;
  assign readData_readDataQueue_31_full = _readData_readDataQueue_fifo_31_full;
  assign compressUnitResultQueue_enq_valid = _compressUnit_out_compressValid;
  assign compressUnitResultQueue_enq_bits_compressValid = _compressUnit_out_compressValid;
  wire               writeQueue_0_empty;
  assign writeQueue_0_empty = _writeQueue_fifo_empty;
  wire               writeQueue_0_full;
  assign writeQueue_0_full = _writeQueue_fifo_full;
  wire               writeQueue_1_empty;
  assign writeQueue_1_empty = _writeQueue_fifo_1_empty;
  wire               writeQueue_1_full;
  assign writeQueue_1_full = _writeQueue_fifo_1_full;
  wire               writeQueue_2_empty;
  assign writeQueue_2_empty = _writeQueue_fifo_2_empty;
  wire               writeQueue_2_full;
  assign writeQueue_2_full = _writeQueue_fifo_2_full;
  wire               writeQueue_3_empty;
  assign writeQueue_3_empty = _writeQueue_fifo_3_empty;
  wire               writeQueue_3_full;
  assign writeQueue_3_full = _writeQueue_fifo_3_full;
  wire               writeQueue_4_empty;
  assign writeQueue_4_empty = _writeQueue_fifo_4_empty;
  wire               writeQueue_4_full;
  assign writeQueue_4_full = _writeQueue_fifo_4_full;
  wire               writeQueue_5_empty;
  assign writeQueue_5_empty = _writeQueue_fifo_5_empty;
  wire               writeQueue_5_full;
  assign writeQueue_5_full = _writeQueue_fifo_5_full;
  wire               writeQueue_6_empty;
  assign writeQueue_6_empty = _writeQueue_fifo_6_empty;
  wire               writeQueue_6_full;
  assign writeQueue_6_full = _writeQueue_fifo_6_full;
  wire               writeQueue_7_empty;
  assign writeQueue_7_empty = _writeQueue_fifo_7_empty;
  wire               writeQueue_7_full;
  assign writeQueue_7_full = _writeQueue_fifo_7_full;
  wire               writeQueue_8_empty;
  assign writeQueue_8_empty = _writeQueue_fifo_8_empty;
  wire               writeQueue_8_full;
  assign writeQueue_8_full = _writeQueue_fifo_8_full;
  wire               writeQueue_9_empty;
  assign writeQueue_9_empty = _writeQueue_fifo_9_empty;
  wire               writeQueue_9_full;
  assign writeQueue_9_full = _writeQueue_fifo_9_full;
  wire               writeQueue_10_empty;
  assign writeQueue_10_empty = _writeQueue_fifo_10_empty;
  wire               writeQueue_10_full;
  assign writeQueue_10_full = _writeQueue_fifo_10_full;
  wire               writeQueue_11_empty;
  assign writeQueue_11_empty = _writeQueue_fifo_11_empty;
  wire               writeQueue_11_full;
  assign writeQueue_11_full = _writeQueue_fifo_11_full;
  wire               writeQueue_12_empty;
  assign writeQueue_12_empty = _writeQueue_fifo_12_empty;
  wire               writeQueue_12_full;
  assign writeQueue_12_full = _writeQueue_fifo_12_full;
  wire               writeQueue_13_empty;
  assign writeQueue_13_empty = _writeQueue_fifo_13_empty;
  wire               writeQueue_13_full;
  assign writeQueue_13_full = _writeQueue_fifo_13_full;
  wire               writeQueue_14_empty;
  assign writeQueue_14_empty = _writeQueue_fifo_14_empty;
  wire               writeQueue_14_full;
  assign writeQueue_14_full = _writeQueue_fifo_14_full;
  wire               writeQueue_15_empty;
  assign writeQueue_15_empty = _writeQueue_fifo_15_empty;
  wire               writeQueue_15_full;
  assign writeQueue_15_full = _writeQueue_fifo_15_full;
  wire               writeQueue_16_empty;
  assign writeQueue_16_empty = _writeQueue_fifo_16_empty;
  wire               writeQueue_16_full;
  assign writeQueue_16_full = _writeQueue_fifo_16_full;
  wire               writeQueue_17_empty;
  assign writeQueue_17_empty = _writeQueue_fifo_17_empty;
  wire               writeQueue_17_full;
  assign writeQueue_17_full = _writeQueue_fifo_17_full;
  wire               writeQueue_18_empty;
  assign writeQueue_18_empty = _writeQueue_fifo_18_empty;
  wire               writeQueue_18_full;
  assign writeQueue_18_full = _writeQueue_fifo_18_full;
  wire               writeQueue_19_empty;
  assign writeQueue_19_empty = _writeQueue_fifo_19_empty;
  wire               writeQueue_19_full;
  assign writeQueue_19_full = _writeQueue_fifo_19_full;
  wire               writeQueue_20_empty;
  assign writeQueue_20_empty = _writeQueue_fifo_20_empty;
  wire               writeQueue_20_full;
  assign writeQueue_20_full = _writeQueue_fifo_20_full;
  wire               writeQueue_21_empty;
  assign writeQueue_21_empty = _writeQueue_fifo_21_empty;
  wire               writeQueue_21_full;
  assign writeQueue_21_full = _writeQueue_fifo_21_full;
  wire               writeQueue_22_empty;
  assign writeQueue_22_empty = _writeQueue_fifo_22_empty;
  wire               writeQueue_22_full;
  assign writeQueue_22_full = _writeQueue_fifo_22_full;
  wire               writeQueue_23_empty;
  assign writeQueue_23_empty = _writeQueue_fifo_23_empty;
  wire               writeQueue_23_full;
  assign writeQueue_23_full = _writeQueue_fifo_23_full;
  wire               writeQueue_24_empty;
  assign writeQueue_24_empty = _writeQueue_fifo_24_empty;
  wire               writeQueue_24_full;
  assign writeQueue_24_full = _writeQueue_fifo_24_full;
  wire               writeQueue_25_empty;
  assign writeQueue_25_empty = _writeQueue_fifo_25_empty;
  wire               writeQueue_25_full;
  assign writeQueue_25_full = _writeQueue_fifo_25_full;
  wire               writeQueue_26_empty;
  assign writeQueue_26_empty = _writeQueue_fifo_26_empty;
  wire               writeQueue_26_full;
  assign writeQueue_26_full = _writeQueue_fifo_26_full;
  wire               writeQueue_27_empty;
  assign writeQueue_27_empty = _writeQueue_fifo_27_empty;
  wire               writeQueue_27_full;
  assign writeQueue_27_full = _writeQueue_fifo_27_full;
  wire               writeQueue_28_empty;
  assign writeQueue_28_empty = _writeQueue_fifo_28_empty;
  wire               writeQueue_28_full;
  assign writeQueue_28_full = _writeQueue_fifo_28_full;
  wire               writeQueue_29_empty;
  assign writeQueue_29_empty = _writeQueue_fifo_29_empty;
  wire               writeQueue_29_full;
  assign writeQueue_29_full = _writeQueue_fifo_29_full;
  wire               writeQueue_30_empty;
  assign writeQueue_30_empty = _writeQueue_fifo_30_empty;
  wire               writeQueue_30_full;
  assign writeQueue_30_full = _writeQueue_fifo_30_full;
  wire               writeQueue_31_empty;
  assign writeQueue_31_empty = _writeQueue_fifo_31_empty;
  wire               writeQueue_31_full;
  assign writeQueue_31_full = _writeQueue_fifo_31_full;
  BitLevelMaskWrite maskedWrite (
    .clock                              (clock),
    .reset                              (reset),
    .needWAR                            (maskDestinationType),
    .vd                                 (instReg_vd),
    .in_0_ready                         (_maskedWrite_in_0_ready),
    .in_0_valid                         (unitType[2] ? _reduceUnit_out_valid : executeValid & maskFilter),
    .in_0_bits_data                     (unitType[2] ? _reduceUnit_out_bits_data : executeResult[31:0]),
    .in_0_bits_bitMask                  (currentMaskGroupForDestination[31:0]),
    .in_0_bits_mask                     (unitType[2] ? _reduceUnit_out_bits_mask : executeWriteByteMask[3:0]),
    .in_0_bits_groupCounter             (unitType[2] ? 5'h0 : executeDeqGroupCounter[4:0]),
    .in_0_bits_ffoByOther               (compressUnitResultQueue_deq_bits_ffoOutput[0] & ffo),
    .in_1_ready                         (_maskedWrite_in_1_ready),
    .in_1_valid                         (executeValid & maskFilter_1),
    .in_1_bits_data                     (executeResult[63:32]),
    .in_1_bits_bitMask                  (currentMaskGroupForDestination[63:32]),
    .in_1_bits_mask                     (executeWriteByteMask[7:4]),
    .in_1_bits_groupCounter             (executeDeqGroupCounter[4:0]),
    .in_1_bits_ffoByOther               (compressUnitResultQueue_deq_bits_ffoOutput[1] & ffo),
    .in_2_ready                         (_maskedWrite_in_2_ready),
    .in_2_valid                         (executeValid & maskFilter_2),
    .in_2_bits_data                     (executeResult[95:64]),
    .in_2_bits_bitMask                  (currentMaskGroupForDestination[95:64]),
    .in_2_bits_mask                     (executeWriteByteMask[11:8]),
    .in_2_bits_groupCounter             (executeDeqGroupCounter[4:0]),
    .in_2_bits_ffoByOther               (compressUnitResultQueue_deq_bits_ffoOutput[2] & ffo),
    .in_3_ready                         (_maskedWrite_in_3_ready),
    .in_3_valid                         (executeValid & maskFilter_3),
    .in_3_bits_data                     (executeResult[127:96]),
    .in_3_bits_bitMask                  (currentMaskGroupForDestination[127:96]),
    .in_3_bits_mask                     (executeWriteByteMask[15:12]),
    .in_3_bits_groupCounter             (executeDeqGroupCounter[4:0]),
    .in_3_bits_ffoByOther               (compressUnitResultQueue_deq_bits_ffoOutput[3] & ffo),
    .in_4_ready                         (_maskedWrite_in_4_ready),
    .in_4_valid                         (executeValid & maskFilter_4),
    .in_4_bits_data                     (executeResult[159:128]),
    .in_4_bits_bitMask                  (currentMaskGroupForDestination[159:128]),
    .in_4_bits_mask                     (executeWriteByteMask[19:16]),
    .in_4_bits_groupCounter             (executeDeqGroupCounter[4:0]),
    .in_4_bits_ffoByOther               (compressUnitResultQueue_deq_bits_ffoOutput[4] & ffo),
    .in_5_ready                         (_maskedWrite_in_5_ready),
    .in_5_valid                         (executeValid & maskFilter_5),
    .in_5_bits_data                     (executeResult[191:160]),
    .in_5_bits_bitMask                  (currentMaskGroupForDestination[191:160]),
    .in_5_bits_mask                     (executeWriteByteMask[23:20]),
    .in_5_bits_groupCounter             (executeDeqGroupCounter[4:0]),
    .in_5_bits_ffoByOther               (compressUnitResultQueue_deq_bits_ffoOutput[5] & ffo),
    .in_6_ready                         (_maskedWrite_in_6_ready),
    .in_6_valid                         (executeValid & maskFilter_6),
    .in_6_bits_data                     (executeResult[223:192]),
    .in_6_bits_bitMask                  (currentMaskGroupForDestination[223:192]),
    .in_6_bits_mask                     (executeWriteByteMask[27:24]),
    .in_6_bits_groupCounter             (executeDeqGroupCounter[4:0]),
    .in_6_bits_ffoByOther               (compressUnitResultQueue_deq_bits_ffoOutput[6] & ffo),
    .in_7_ready                         (_maskedWrite_in_7_ready),
    .in_7_valid                         (executeValid & maskFilter_7),
    .in_7_bits_data                     (executeResult[255:224]),
    .in_7_bits_bitMask                  (currentMaskGroupForDestination[255:224]),
    .in_7_bits_mask                     (executeWriteByteMask[31:28]),
    .in_7_bits_groupCounter             (executeDeqGroupCounter[4:0]),
    .in_7_bits_ffoByOther               (compressUnitResultQueue_deq_bits_ffoOutput[7] & ffo),
    .in_8_ready                         (_maskedWrite_in_8_ready),
    .in_8_valid                         (executeValid & maskFilter_8),
    .in_8_bits_data                     (executeResult[287:256]),
    .in_8_bits_bitMask                  (currentMaskGroupForDestination[287:256]),
    .in_8_bits_mask                     (executeWriteByteMask[35:32]),
    .in_8_bits_groupCounter             (executeDeqGroupCounter[4:0]),
    .in_8_bits_ffoByOther               (compressUnitResultQueue_deq_bits_ffoOutput[8] & ffo),
    .in_9_ready                         (_maskedWrite_in_9_ready),
    .in_9_valid                         (executeValid & maskFilter_9),
    .in_9_bits_data                     (executeResult[319:288]),
    .in_9_bits_bitMask                  (currentMaskGroupForDestination[319:288]),
    .in_9_bits_mask                     (executeWriteByteMask[39:36]),
    .in_9_bits_groupCounter             (executeDeqGroupCounter[4:0]),
    .in_9_bits_ffoByOther               (compressUnitResultQueue_deq_bits_ffoOutput[9] & ffo),
    .in_10_ready                        (_maskedWrite_in_10_ready),
    .in_10_valid                        (executeValid & maskFilter_10),
    .in_10_bits_data                    (executeResult[351:320]),
    .in_10_bits_bitMask                 (currentMaskGroupForDestination[351:320]),
    .in_10_bits_mask                    (executeWriteByteMask[43:40]),
    .in_10_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_10_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[10] & ffo),
    .in_11_ready                        (_maskedWrite_in_11_ready),
    .in_11_valid                        (executeValid & maskFilter_11),
    .in_11_bits_data                    (executeResult[383:352]),
    .in_11_bits_bitMask                 (currentMaskGroupForDestination[383:352]),
    .in_11_bits_mask                    (executeWriteByteMask[47:44]),
    .in_11_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_11_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[11] & ffo),
    .in_12_ready                        (_maskedWrite_in_12_ready),
    .in_12_valid                        (executeValid & maskFilter_12),
    .in_12_bits_data                    (executeResult[415:384]),
    .in_12_bits_bitMask                 (currentMaskGroupForDestination[415:384]),
    .in_12_bits_mask                    (executeWriteByteMask[51:48]),
    .in_12_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_12_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[12] & ffo),
    .in_13_ready                        (_maskedWrite_in_13_ready),
    .in_13_valid                        (executeValid & maskFilter_13),
    .in_13_bits_data                    (executeResult[447:416]),
    .in_13_bits_bitMask                 (currentMaskGroupForDestination[447:416]),
    .in_13_bits_mask                    (executeWriteByteMask[55:52]),
    .in_13_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_13_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[13] & ffo),
    .in_14_ready                        (_maskedWrite_in_14_ready),
    .in_14_valid                        (executeValid & maskFilter_14),
    .in_14_bits_data                    (executeResult[479:448]),
    .in_14_bits_bitMask                 (currentMaskGroupForDestination[479:448]),
    .in_14_bits_mask                    (executeWriteByteMask[59:56]),
    .in_14_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_14_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[14] & ffo),
    .in_15_ready                        (_maskedWrite_in_15_ready),
    .in_15_valid                        (executeValid & maskFilter_15),
    .in_15_bits_data                    (executeResult[511:480]),
    .in_15_bits_bitMask                 (currentMaskGroupForDestination[511:480]),
    .in_15_bits_mask                    (executeWriteByteMask[63:60]),
    .in_15_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_15_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[15] & ffo),
    .in_16_ready                        (_maskedWrite_in_16_ready),
    .in_16_valid                        (executeValid & maskFilter_16),
    .in_16_bits_data                    (executeResult[543:512]),
    .in_16_bits_bitMask                 (currentMaskGroupForDestination[543:512]),
    .in_16_bits_mask                    (executeWriteByteMask[67:64]),
    .in_16_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_16_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[16] & ffo),
    .in_17_ready                        (_maskedWrite_in_17_ready),
    .in_17_valid                        (executeValid & maskFilter_17),
    .in_17_bits_data                    (executeResult[575:544]),
    .in_17_bits_bitMask                 (currentMaskGroupForDestination[575:544]),
    .in_17_bits_mask                    (executeWriteByteMask[71:68]),
    .in_17_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_17_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[17] & ffo),
    .in_18_ready                        (_maskedWrite_in_18_ready),
    .in_18_valid                        (executeValid & maskFilter_18),
    .in_18_bits_data                    (executeResult[607:576]),
    .in_18_bits_bitMask                 (currentMaskGroupForDestination[607:576]),
    .in_18_bits_mask                    (executeWriteByteMask[75:72]),
    .in_18_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_18_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[18] & ffo),
    .in_19_ready                        (_maskedWrite_in_19_ready),
    .in_19_valid                        (executeValid & maskFilter_19),
    .in_19_bits_data                    (executeResult[639:608]),
    .in_19_bits_bitMask                 (currentMaskGroupForDestination[639:608]),
    .in_19_bits_mask                    (executeWriteByteMask[79:76]),
    .in_19_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_19_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[19] & ffo),
    .in_20_ready                        (_maskedWrite_in_20_ready),
    .in_20_valid                        (executeValid & maskFilter_20),
    .in_20_bits_data                    (executeResult[671:640]),
    .in_20_bits_bitMask                 (currentMaskGroupForDestination[671:640]),
    .in_20_bits_mask                    (executeWriteByteMask[83:80]),
    .in_20_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_20_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[20] & ffo),
    .in_21_ready                        (_maskedWrite_in_21_ready),
    .in_21_valid                        (executeValid & maskFilter_21),
    .in_21_bits_data                    (executeResult[703:672]),
    .in_21_bits_bitMask                 (currentMaskGroupForDestination[703:672]),
    .in_21_bits_mask                    (executeWriteByteMask[87:84]),
    .in_21_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_21_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[21] & ffo),
    .in_22_ready                        (_maskedWrite_in_22_ready),
    .in_22_valid                        (executeValid & maskFilter_22),
    .in_22_bits_data                    (executeResult[735:704]),
    .in_22_bits_bitMask                 (currentMaskGroupForDestination[735:704]),
    .in_22_bits_mask                    (executeWriteByteMask[91:88]),
    .in_22_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_22_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[22] & ffo),
    .in_23_ready                        (_maskedWrite_in_23_ready),
    .in_23_valid                        (executeValid & maskFilter_23),
    .in_23_bits_data                    (executeResult[767:736]),
    .in_23_bits_bitMask                 (currentMaskGroupForDestination[767:736]),
    .in_23_bits_mask                    (executeWriteByteMask[95:92]),
    .in_23_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_23_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[23] & ffo),
    .in_24_ready                        (_maskedWrite_in_24_ready),
    .in_24_valid                        (executeValid & maskFilter_24),
    .in_24_bits_data                    (executeResult[799:768]),
    .in_24_bits_bitMask                 (currentMaskGroupForDestination[799:768]),
    .in_24_bits_mask                    (executeWriteByteMask[99:96]),
    .in_24_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_24_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[24] & ffo),
    .in_25_ready                        (_maskedWrite_in_25_ready),
    .in_25_valid                        (executeValid & maskFilter_25),
    .in_25_bits_data                    (executeResult[831:800]),
    .in_25_bits_bitMask                 (currentMaskGroupForDestination[831:800]),
    .in_25_bits_mask                    (executeWriteByteMask[103:100]),
    .in_25_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_25_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[25] & ffo),
    .in_26_ready                        (_maskedWrite_in_26_ready),
    .in_26_valid                        (executeValid & maskFilter_26),
    .in_26_bits_data                    (executeResult[863:832]),
    .in_26_bits_bitMask                 (currentMaskGroupForDestination[863:832]),
    .in_26_bits_mask                    (executeWriteByteMask[107:104]),
    .in_26_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_26_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[26] & ffo),
    .in_27_ready                        (_maskedWrite_in_27_ready),
    .in_27_valid                        (executeValid & maskFilter_27),
    .in_27_bits_data                    (executeResult[895:864]),
    .in_27_bits_bitMask                 (currentMaskGroupForDestination[895:864]),
    .in_27_bits_mask                    (executeWriteByteMask[111:108]),
    .in_27_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_27_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[27] & ffo),
    .in_28_ready                        (_maskedWrite_in_28_ready),
    .in_28_valid                        (executeValid & maskFilter_28),
    .in_28_bits_data                    (executeResult[927:896]),
    .in_28_bits_bitMask                 (currentMaskGroupForDestination[927:896]),
    .in_28_bits_mask                    (executeWriteByteMask[115:112]),
    .in_28_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_28_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[28] & ffo),
    .in_29_ready                        (_maskedWrite_in_29_ready),
    .in_29_valid                        (executeValid & maskFilter_29),
    .in_29_bits_data                    (executeResult[959:928]),
    .in_29_bits_bitMask                 (currentMaskGroupForDestination[959:928]),
    .in_29_bits_mask                    (executeWriteByteMask[119:116]),
    .in_29_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_29_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[29] & ffo),
    .in_30_ready                        (_maskedWrite_in_30_ready),
    .in_30_valid                        (executeValid & maskFilter_30),
    .in_30_bits_data                    (executeResult[991:960]),
    .in_30_bits_bitMask                 (currentMaskGroupForDestination[991:960]),
    .in_30_bits_mask                    (executeWriteByteMask[123:120]),
    .in_30_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_30_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[30] & ffo),
    .in_31_ready                        (_maskedWrite_in_31_ready),
    .in_31_valid                        (executeValid & maskFilter_31),
    .in_31_bits_data                    (executeResult[1023:992]),
    .in_31_bits_bitMask                 (currentMaskGroupForDestination[1023:992]),
    .in_31_bits_mask                    (executeWriteByteMask[127:124]),
    .in_31_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_31_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[31] & ffo),
    .out_0_ready                        (writeQueue_0_enq_ready),
    .out_0_valid                        (_maskedWrite_out_0_valid),
    .out_0_bits_ffoByOther              (_maskedWrite_out_0_bits_ffoByOther),
    .out_0_bits_writeData_data          (_maskedWrite_out_0_bits_writeData_data),
    .out_0_bits_writeData_mask          (_maskedWrite_out_0_bits_writeData_mask),
    .out_0_bits_writeData_groupCounter  (_maskedWrite_out_0_bits_writeData_groupCounter),
    .out_1_ready                        (writeQueue_1_enq_ready),
    .out_1_valid                        (_maskedWrite_out_1_valid),
    .out_1_bits_ffoByOther              (_maskedWrite_out_1_bits_ffoByOther),
    .out_1_bits_writeData_data          (_maskedWrite_out_1_bits_writeData_data),
    .out_1_bits_writeData_mask          (_maskedWrite_out_1_bits_writeData_mask),
    .out_1_bits_writeData_groupCounter  (_maskedWrite_out_1_bits_writeData_groupCounter),
    .out_2_ready                        (writeQueue_2_enq_ready),
    .out_2_valid                        (_maskedWrite_out_2_valid),
    .out_2_bits_ffoByOther              (_maskedWrite_out_2_bits_ffoByOther),
    .out_2_bits_writeData_data          (_maskedWrite_out_2_bits_writeData_data),
    .out_2_bits_writeData_mask          (_maskedWrite_out_2_bits_writeData_mask),
    .out_2_bits_writeData_groupCounter  (_maskedWrite_out_2_bits_writeData_groupCounter),
    .out_3_ready                        (writeQueue_3_enq_ready),
    .out_3_valid                        (_maskedWrite_out_3_valid),
    .out_3_bits_ffoByOther              (_maskedWrite_out_3_bits_ffoByOther),
    .out_3_bits_writeData_data          (_maskedWrite_out_3_bits_writeData_data),
    .out_3_bits_writeData_mask          (_maskedWrite_out_3_bits_writeData_mask),
    .out_3_bits_writeData_groupCounter  (_maskedWrite_out_3_bits_writeData_groupCounter),
    .out_4_ready                        (writeQueue_4_enq_ready),
    .out_4_valid                        (_maskedWrite_out_4_valid),
    .out_4_bits_ffoByOther              (_maskedWrite_out_4_bits_ffoByOther),
    .out_4_bits_writeData_data          (_maskedWrite_out_4_bits_writeData_data),
    .out_4_bits_writeData_mask          (_maskedWrite_out_4_bits_writeData_mask),
    .out_4_bits_writeData_groupCounter  (_maskedWrite_out_4_bits_writeData_groupCounter),
    .out_5_ready                        (writeQueue_5_enq_ready),
    .out_5_valid                        (_maskedWrite_out_5_valid),
    .out_5_bits_ffoByOther              (_maskedWrite_out_5_bits_ffoByOther),
    .out_5_bits_writeData_data          (_maskedWrite_out_5_bits_writeData_data),
    .out_5_bits_writeData_mask          (_maskedWrite_out_5_bits_writeData_mask),
    .out_5_bits_writeData_groupCounter  (_maskedWrite_out_5_bits_writeData_groupCounter),
    .out_6_ready                        (writeQueue_6_enq_ready),
    .out_6_valid                        (_maskedWrite_out_6_valid),
    .out_6_bits_ffoByOther              (_maskedWrite_out_6_bits_ffoByOther),
    .out_6_bits_writeData_data          (_maskedWrite_out_6_bits_writeData_data),
    .out_6_bits_writeData_mask          (_maskedWrite_out_6_bits_writeData_mask),
    .out_6_bits_writeData_groupCounter  (_maskedWrite_out_6_bits_writeData_groupCounter),
    .out_7_ready                        (writeQueue_7_enq_ready),
    .out_7_valid                        (_maskedWrite_out_7_valid),
    .out_7_bits_ffoByOther              (_maskedWrite_out_7_bits_ffoByOther),
    .out_7_bits_writeData_data          (_maskedWrite_out_7_bits_writeData_data),
    .out_7_bits_writeData_mask          (_maskedWrite_out_7_bits_writeData_mask),
    .out_7_bits_writeData_groupCounter  (_maskedWrite_out_7_bits_writeData_groupCounter),
    .out_8_ready                        (writeQueue_8_enq_ready),
    .out_8_valid                        (_maskedWrite_out_8_valid),
    .out_8_bits_ffoByOther              (_maskedWrite_out_8_bits_ffoByOther),
    .out_8_bits_writeData_data          (_maskedWrite_out_8_bits_writeData_data),
    .out_8_bits_writeData_mask          (_maskedWrite_out_8_bits_writeData_mask),
    .out_8_bits_writeData_groupCounter  (_maskedWrite_out_8_bits_writeData_groupCounter),
    .out_9_ready                        (writeQueue_9_enq_ready),
    .out_9_valid                        (_maskedWrite_out_9_valid),
    .out_9_bits_ffoByOther              (_maskedWrite_out_9_bits_ffoByOther),
    .out_9_bits_writeData_data          (_maskedWrite_out_9_bits_writeData_data),
    .out_9_bits_writeData_mask          (_maskedWrite_out_9_bits_writeData_mask),
    .out_9_bits_writeData_groupCounter  (_maskedWrite_out_9_bits_writeData_groupCounter),
    .out_10_ready                       (writeQueue_10_enq_ready),
    .out_10_valid                       (_maskedWrite_out_10_valid),
    .out_10_bits_ffoByOther             (_maskedWrite_out_10_bits_ffoByOther),
    .out_10_bits_writeData_data         (_maskedWrite_out_10_bits_writeData_data),
    .out_10_bits_writeData_mask         (_maskedWrite_out_10_bits_writeData_mask),
    .out_10_bits_writeData_groupCounter (_maskedWrite_out_10_bits_writeData_groupCounter),
    .out_11_ready                       (writeQueue_11_enq_ready),
    .out_11_valid                       (_maskedWrite_out_11_valid),
    .out_11_bits_ffoByOther             (_maskedWrite_out_11_bits_ffoByOther),
    .out_11_bits_writeData_data         (_maskedWrite_out_11_bits_writeData_data),
    .out_11_bits_writeData_mask         (_maskedWrite_out_11_bits_writeData_mask),
    .out_11_bits_writeData_groupCounter (_maskedWrite_out_11_bits_writeData_groupCounter),
    .out_12_ready                       (writeQueue_12_enq_ready),
    .out_12_valid                       (_maskedWrite_out_12_valid),
    .out_12_bits_ffoByOther             (_maskedWrite_out_12_bits_ffoByOther),
    .out_12_bits_writeData_data         (_maskedWrite_out_12_bits_writeData_data),
    .out_12_bits_writeData_mask         (_maskedWrite_out_12_bits_writeData_mask),
    .out_12_bits_writeData_groupCounter (_maskedWrite_out_12_bits_writeData_groupCounter),
    .out_13_ready                       (writeQueue_13_enq_ready),
    .out_13_valid                       (_maskedWrite_out_13_valid),
    .out_13_bits_ffoByOther             (_maskedWrite_out_13_bits_ffoByOther),
    .out_13_bits_writeData_data         (_maskedWrite_out_13_bits_writeData_data),
    .out_13_bits_writeData_mask         (_maskedWrite_out_13_bits_writeData_mask),
    .out_13_bits_writeData_groupCounter (_maskedWrite_out_13_bits_writeData_groupCounter),
    .out_14_ready                       (writeQueue_14_enq_ready),
    .out_14_valid                       (_maskedWrite_out_14_valid),
    .out_14_bits_ffoByOther             (_maskedWrite_out_14_bits_ffoByOther),
    .out_14_bits_writeData_data         (_maskedWrite_out_14_bits_writeData_data),
    .out_14_bits_writeData_mask         (_maskedWrite_out_14_bits_writeData_mask),
    .out_14_bits_writeData_groupCounter (_maskedWrite_out_14_bits_writeData_groupCounter),
    .out_15_ready                       (writeQueue_15_enq_ready),
    .out_15_valid                       (_maskedWrite_out_15_valid),
    .out_15_bits_ffoByOther             (_maskedWrite_out_15_bits_ffoByOther),
    .out_15_bits_writeData_data         (_maskedWrite_out_15_bits_writeData_data),
    .out_15_bits_writeData_mask         (_maskedWrite_out_15_bits_writeData_mask),
    .out_15_bits_writeData_groupCounter (_maskedWrite_out_15_bits_writeData_groupCounter),
    .out_16_ready                       (writeQueue_16_enq_ready),
    .out_16_valid                       (_maskedWrite_out_16_valid),
    .out_16_bits_ffoByOther             (_maskedWrite_out_16_bits_ffoByOther),
    .out_16_bits_writeData_data         (_maskedWrite_out_16_bits_writeData_data),
    .out_16_bits_writeData_mask         (_maskedWrite_out_16_bits_writeData_mask),
    .out_16_bits_writeData_groupCounter (_maskedWrite_out_16_bits_writeData_groupCounter),
    .out_17_ready                       (writeQueue_17_enq_ready),
    .out_17_valid                       (_maskedWrite_out_17_valid),
    .out_17_bits_ffoByOther             (_maskedWrite_out_17_bits_ffoByOther),
    .out_17_bits_writeData_data         (_maskedWrite_out_17_bits_writeData_data),
    .out_17_bits_writeData_mask         (_maskedWrite_out_17_bits_writeData_mask),
    .out_17_bits_writeData_groupCounter (_maskedWrite_out_17_bits_writeData_groupCounter),
    .out_18_ready                       (writeQueue_18_enq_ready),
    .out_18_valid                       (_maskedWrite_out_18_valid),
    .out_18_bits_ffoByOther             (_maskedWrite_out_18_bits_ffoByOther),
    .out_18_bits_writeData_data         (_maskedWrite_out_18_bits_writeData_data),
    .out_18_bits_writeData_mask         (_maskedWrite_out_18_bits_writeData_mask),
    .out_18_bits_writeData_groupCounter (_maskedWrite_out_18_bits_writeData_groupCounter),
    .out_19_ready                       (writeQueue_19_enq_ready),
    .out_19_valid                       (_maskedWrite_out_19_valid),
    .out_19_bits_ffoByOther             (_maskedWrite_out_19_bits_ffoByOther),
    .out_19_bits_writeData_data         (_maskedWrite_out_19_bits_writeData_data),
    .out_19_bits_writeData_mask         (_maskedWrite_out_19_bits_writeData_mask),
    .out_19_bits_writeData_groupCounter (_maskedWrite_out_19_bits_writeData_groupCounter),
    .out_20_ready                       (writeQueue_20_enq_ready),
    .out_20_valid                       (_maskedWrite_out_20_valid),
    .out_20_bits_ffoByOther             (_maskedWrite_out_20_bits_ffoByOther),
    .out_20_bits_writeData_data         (_maskedWrite_out_20_bits_writeData_data),
    .out_20_bits_writeData_mask         (_maskedWrite_out_20_bits_writeData_mask),
    .out_20_bits_writeData_groupCounter (_maskedWrite_out_20_bits_writeData_groupCounter),
    .out_21_ready                       (writeQueue_21_enq_ready),
    .out_21_valid                       (_maskedWrite_out_21_valid),
    .out_21_bits_ffoByOther             (_maskedWrite_out_21_bits_ffoByOther),
    .out_21_bits_writeData_data         (_maskedWrite_out_21_bits_writeData_data),
    .out_21_bits_writeData_mask         (_maskedWrite_out_21_bits_writeData_mask),
    .out_21_bits_writeData_groupCounter (_maskedWrite_out_21_bits_writeData_groupCounter),
    .out_22_ready                       (writeQueue_22_enq_ready),
    .out_22_valid                       (_maskedWrite_out_22_valid),
    .out_22_bits_ffoByOther             (_maskedWrite_out_22_bits_ffoByOther),
    .out_22_bits_writeData_data         (_maskedWrite_out_22_bits_writeData_data),
    .out_22_bits_writeData_mask         (_maskedWrite_out_22_bits_writeData_mask),
    .out_22_bits_writeData_groupCounter (_maskedWrite_out_22_bits_writeData_groupCounter),
    .out_23_ready                       (writeQueue_23_enq_ready),
    .out_23_valid                       (_maskedWrite_out_23_valid),
    .out_23_bits_ffoByOther             (_maskedWrite_out_23_bits_ffoByOther),
    .out_23_bits_writeData_data         (_maskedWrite_out_23_bits_writeData_data),
    .out_23_bits_writeData_mask         (_maskedWrite_out_23_bits_writeData_mask),
    .out_23_bits_writeData_groupCounter (_maskedWrite_out_23_bits_writeData_groupCounter),
    .out_24_ready                       (writeQueue_24_enq_ready),
    .out_24_valid                       (_maskedWrite_out_24_valid),
    .out_24_bits_ffoByOther             (_maskedWrite_out_24_bits_ffoByOther),
    .out_24_bits_writeData_data         (_maskedWrite_out_24_bits_writeData_data),
    .out_24_bits_writeData_mask         (_maskedWrite_out_24_bits_writeData_mask),
    .out_24_bits_writeData_groupCounter (_maskedWrite_out_24_bits_writeData_groupCounter),
    .out_25_ready                       (writeQueue_25_enq_ready),
    .out_25_valid                       (_maskedWrite_out_25_valid),
    .out_25_bits_ffoByOther             (_maskedWrite_out_25_bits_ffoByOther),
    .out_25_bits_writeData_data         (_maskedWrite_out_25_bits_writeData_data),
    .out_25_bits_writeData_mask         (_maskedWrite_out_25_bits_writeData_mask),
    .out_25_bits_writeData_groupCounter (_maskedWrite_out_25_bits_writeData_groupCounter),
    .out_26_ready                       (writeQueue_26_enq_ready),
    .out_26_valid                       (_maskedWrite_out_26_valid),
    .out_26_bits_ffoByOther             (_maskedWrite_out_26_bits_ffoByOther),
    .out_26_bits_writeData_data         (_maskedWrite_out_26_bits_writeData_data),
    .out_26_bits_writeData_mask         (_maskedWrite_out_26_bits_writeData_mask),
    .out_26_bits_writeData_groupCounter (_maskedWrite_out_26_bits_writeData_groupCounter),
    .out_27_ready                       (writeQueue_27_enq_ready),
    .out_27_valid                       (_maskedWrite_out_27_valid),
    .out_27_bits_ffoByOther             (_maskedWrite_out_27_bits_ffoByOther),
    .out_27_bits_writeData_data         (_maskedWrite_out_27_bits_writeData_data),
    .out_27_bits_writeData_mask         (_maskedWrite_out_27_bits_writeData_mask),
    .out_27_bits_writeData_groupCounter (_maskedWrite_out_27_bits_writeData_groupCounter),
    .out_28_ready                       (writeQueue_28_enq_ready),
    .out_28_valid                       (_maskedWrite_out_28_valid),
    .out_28_bits_ffoByOther             (_maskedWrite_out_28_bits_ffoByOther),
    .out_28_bits_writeData_data         (_maskedWrite_out_28_bits_writeData_data),
    .out_28_bits_writeData_mask         (_maskedWrite_out_28_bits_writeData_mask),
    .out_28_bits_writeData_groupCounter (_maskedWrite_out_28_bits_writeData_groupCounter),
    .out_29_ready                       (writeQueue_29_enq_ready),
    .out_29_valid                       (_maskedWrite_out_29_valid),
    .out_29_bits_ffoByOther             (_maskedWrite_out_29_bits_ffoByOther),
    .out_29_bits_writeData_data         (_maskedWrite_out_29_bits_writeData_data),
    .out_29_bits_writeData_mask         (_maskedWrite_out_29_bits_writeData_mask),
    .out_29_bits_writeData_groupCounter (_maskedWrite_out_29_bits_writeData_groupCounter),
    .out_30_ready                       (writeQueue_30_enq_ready),
    .out_30_valid                       (_maskedWrite_out_30_valid),
    .out_30_bits_ffoByOther             (_maskedWrite_out_30_bits_ffoByOther),
    .out_30_bits_writeData_data         (_maskedWrite_out_30_bits_writeData_data),
    .out_30_bits_writeData_mask         (_maskedWrite_out_30_bits_writeData_mask),
    .out_30_bits_writeData_groupCounter (_maskedWrite_out_30_bits_writeData_groupCounter),
    .out_31_ready                       (writeQueue_31_enq_ready),
    .out_31_valid                       (_maskedWrite_out_31_valid),
    .out_31_bits_ffoByOther             (_maskedWrite_out_31_bits_ffoByOther),
    .out_31_bits_writeData_data         (_maskedWrite_out_31_bits_writeData_data),
    .out_31_bits_writeData_mask         (_maskedWrite_out_31_bits_writeData_mask),
    .out_31_bits_writeData_groupCounter (_maskedWrite_out_31_bits_writeData_groupCounter),
    .readChannel_0_ready                (readChannel_0_ready_0),
    .readChannel_0_valid                (_maskedWrite_readChannel_0_valid),
    .readChannel_0_bits_vs              (_maskedWrite_readChannel_0_bits_vs),
    .readChannel_0_bits_offset          (_maskedWrite_readChannel_0_bits_offset),
    .readChannel_1_ready                (readChannel_1_ready_0),
    .readChannel_1_valid                (_maskedWrite_readChannel_1_valid),
    .readChannel_1_bits_vs              (_maskedWrite_readChannel_1_bits_vs),
    .readChannel_1_bits_offset          (_maskedWrite_readChannel_1_bits_offset),
    .readChannel_2_ready                (readChannel_2_ready_0),
    .readChannel_2_valid                (_maskedWrite_readChannel_2_valid),
    .readChannel_2_bits_vs              (_maskedWrite_readChannel_2_bits_vs),
    .readChannel_2_bits_offset          (_maskedWrite_readChannel_2_bits_offset),
    .readChannel_3_ready                (readChannel_3_ready_0),
    .readChannel_3_valid                (_maskedWrite_readChannel_3_valid),
    .readChannel_3_bits_vs              (_maskedWrite_readChannel_3_bits_vs),
    .readChannel_3_bits_offset          (_maskedWrite_readChannel_3_bits_offset),
    .readChannel_4_ready                (readChannel_4_ready_0),
    .readChannel_4_valid                (_maskedWrite_readChannel_4_valid),
    .readChannel_4_bits_vs              (_maskedWrite_readChannel_4_bits_vs),
    .readChannel_4_bits_offset          (_maskedWrite_readChannel_4_bits_offset),
    .readChannel_5_ready                (readChannel_5_ready_0),
    .readChannel_5_valid                (_maskedWrite_readChannel_5_valid),
    .readChannel_5_bits_vs              (_maskedWrite_readChannel_5_bits_vs),
    .readChannel_5_bits_offset          (_maskedWrite_readChannel_5_bits_offset),
    .readChannel_6_ready                (readChannel_6_ready_0),
    .readChannel_6_valid                (_maskedWrite_readChannel_6_valid),
    .readChannel_6_bits_vs              (_maskedWrite_readChannel_6_bits_vs),
    .readChannel_6_bits_offset          (_maskedWrite_readChannel_6_bits_offset),
    .readChannel_7_ready                (readChannel_7_ready_0),
    .readChannel_7_valid                (_maskedWrite_readChannel_7_valid),
    .readChannel_7_bits_vs              (_maskedWrite_readChannel_7_bits_vs),
    .readChannel_7_bits_offset          (_maskedWrite_readChannel_7_bits_offset),
    .readChannel_8_ready                (readChannel_8_ready_0),
    .readChannel_8_valid                (_maskedWrite_readChannel_8_valid),
    .readChannel_8_bits_vs              (_maskedWrite_readChannel_8_bits_vs),
    .readChannel_8_bits_offset          (_maskedWrite_readChannel_8_bits_offset),
    .readChannel_9_ready                (readChannel_9_ready_0),
    .readChannel_9_valid                (_maskedWrite_readChannel_9_valid),
    .readChannel_9_bits_vs              (_maskedWrite_readChannel_9_bits_vs),
    .readChannel_9_bits_offset          (_maskedWrite_readChannel_9_bits_offset),
    .readChannel_10_ready               (readChannel_10_ready_0),
    .readChannel_10_valid               (_maskedWrite_readChannel_10_valid),
    .readChannel_10_bits_vs             (_maskedWrite_readChannel_10_bits_vs),
    .readChannel_10_bits_offset         (_maskedWrite_readChannel_10_bits_offset),
    .readChannel_11_ready               (readChannel_11_ready_0),
    .readChannel_11_valid               (_maskedWrite_readChannel_11_valid),
    .readChannel_11_bits_vs             (_maskedWrite_readChannel_11_bits_vs),
    .readChannel_11_bits_offset         (_maskedWrite_readChannel_11_bits_offset),
    .readChannel_12_ready               (readChannel_12_ready_0),
    .readChannel_12_valid               (_maskedWrite_readChannel_12_valid),
    .readChannel_12_bits_vs             (_maskedWrite_readChannel_12_bits_vs),
    .readChannel_12_bits_offset         (_maskedWrite_readChannel_12_bits_offset),
    .readChannel_13_ready               (readChannel_13_ready_0),
    .readChannel_13_valid               (_maskedWrite_readChannel_13_valid),
    .readChannel_13_bits_vs             (_maskedWrite_readChannel_13_bits_vs),
    .readChannel_13_bits_offset         (_maskedWrite_readChannel_13_bits_offset),
    .readChannel_14_ready               (readChannel_14_ready_0),
    .readChannel_14_valid               (_maskedWrite_readChannel_14_valid),
    .readChannel_14_bits_vs             (_maskedWrite_readChannel_14_bits_vs),
    .readChannel_14_bits_offset         (_maskedWrite_readChannel_14_bits_offset),
    .readChannel_15_ready               (readChannel_15_ready_0),
    .readChannel_15_valid               (_maskedWrite_readChannel_15_valid),
    .readChannel_15_bits_vs             (_maskedWrite_readChannel_15_bits_vs),
    .readChannel_15_bits_offset         (_maskedWrite_readChannel_15_bits_offset),
    .readChannel_16_ready               (readChannel_16_ready_0),
    .readChannel_16_valid               (_maskedWrite_readChannel_16_valid),
    .readChannel_16_bits_vs             (_maskedWrite_readChannel_16_bits_vs),
    .readChannel_16_bits_offset         (_maskedWrite_readChannel_16_bits_offset),
    .readChannel_17_ready               (readChannel_17_ready_0),
    .readChannel_17_valid               (_maskedWrite_readChannel_17_valid),
    .readChannel_17_bits_vs             (_maskedWrite_readChannel_17_bits_vs),
    .readChannel_17_bits_offset         (_maskedWrite_readChannel_17_bits_offset),
    .readChannel_18_ready               (readChannel_18_ready_0),
    .readChannel_18_valid               (_maskedWrite_readChannel_18_valid),
    .readChannel_18_bits_vs             (_maskedWrite_readChannel_18_bits_vs),
    .readChannel_18_bits_offset         (_maskedWrite_readChannel_18_bits_offset),
    .readChannel_19_ready               (readChannel_19_ready_0),
    .readChannel_19_valid               (_maskedWrite_readChannel_19_valid),
    .readChannel_19_bits_vs             (_maskedWrite_readChannel_19_bits_vs),
    .readChannel_19_bits_offset         (_maskedWrite_readChannel_19_bits_offset),
    .readChannel_20_ready               (readChannel_20_ready_0),
    .readChannel_20_valid               (_maskedWrite_readChannel_20_valid),
    .readChannel_20_bits_vs             (_maskedWrite_readChannel_20_bits_vs),
    .readChannel_20_bits_offset         (_maskedWrite_readChannel_20_bits_offset),
    .readChannel_21_ready               (readChannel_21_ready_0),
    .readChannel_21_valid               (_maskedWrite_readChannel_21_valid),
    .readChannel_21_bits_vs             (_maskedWrite_readChannel_21_bits_vs),
    .readChannel_21_bits_offset         (_maskedWrite_readChannel_21_bits_offset),
    .readChannel_22_ready               (readChannel_22_ready_0),
    .readChannel_22_valid               (_maskedWrite_readChannel_22_valid),
    .readChannel_22_bits_vs             (_maskedWrite_readChannel_22_bits_vs),
    .readChannel_22_bits_offset         (_maskedWrite_readChannel_22_bits_offset),
    .readChannel_23_ready               (readChannel_23_ready_0),
    .readChannel_23_valid               (_maskedWrite_readChannel_23_valid),
    .readChannel_23_bits_vs             (_maskedWrite_readChannel_23_bits_vs),
    .readChannel_23_bits_offset         (_maskedWrite_readChannel_23_bits_offset),
    .readChannel_24_ready               (readChannel_24_ready_0),
    .readChannel_24_valid               (_maskedWrite_readChannel_24_valid),
    .readChannel_24_bits_vs             (_maskedWrite_readChannel_24_bits_vs),
    .readChannel_24_bits_offset         (_maskedWrite_readChannel_24_bits_offset),
    .readChannel_25_ready               (readChannel_25_ready_0),
    .readChannel_25_valid               (_maskedWrite_readChannel_25_valid),
    .readChannel_25_bits_vs             (_maskedWrite_readChannel_25_bits_vs),
    .readChannel_25_bits_offset         (_maskedWrite_readChannel_25_bits_offset),
    .readChannel_26_ready               (readChannel_26_ready_0),
    .readChannel_26_valid               (_maskedWrite_readChannel_26_valid),
    .readChannel_26_bits_vs             (_maskedWrite_readChannel_26_bits_vs),
    .readChannel_26_bits_offset         (_maskedWrite_readChannel_26_bits_offset),
    .readChannel_27_ready               (readChannel_27_ready_0),
    .readChannel_27_valid               (_maskedWrite_readChannel_27_valid),
    .readChannel_27_bits_vs             (_maskedWrite_readChannel_27_bits_vs),
    .readChannel_27_bits_offset         (_maskedWrite_readChannel_27_bits_offset),
    .readChannel_28_ready               (readChannel_28_ready_0),
    .readChannel_28_valid               (_maskedWrite_readChannel_28_valid),
    .readChannel_28_bits_vs             (_maskedWrite_readChannel_28_bits_vs),
    .readChannel_28_bits_offset         (_maskedWrite_readChannel_28_bits_offset),
    .readChannel_29_ready               (readChannel_29_ready_0),
    .readChannel_29_valid               (_maskedWrite_readChannel_29_valid),
    .readChannel_29_bits_vs             (_maskedWrite_readChannel_29_bits_vs),
    .readChannel_29_bits_offset         (_maskedWrite_readChannel_29_bits_offset),
    .readChannel_30_ready               (readChannel_30_ready_0),
    .readChannel_30_valid               (_maskedWrite_readChannel_30_valid),
    .readChannel_30_bits_vs             (_maskedWrite_readChannel_30_bits_vs),
    .readChannel_30_bits_offset         (_maskedWrite_readChannel_30_bits_offset),
    .readChannel_31_ready               (readChannel_31_ready_0),
    .readChannel_31_valid               (_maskedWrite_readChannel_31_valid),
    .readChannel_31_bits_vs             (_maskedWrite_readChannel_31_bits_vs),
    .readChannel_31_bits_offset         (_maskedWrite_readChannel_31_bits_offset),
    .readResult_0_valid                 (readResult_0_valid),
    .readResult_0_bits                  (readResult_0_bits),
    .readResult_1_valid                 (readResult_1_valid),
    .readResult_1_bits                  (readResult_1_bits),
    .readResult_2_valid                 (readResult_2_valid),
    .readResult_2_bits                  (readResult_2_bits),
    .readResult_3_valid                 (readResult_3_valid),
    .readResult_3_bits                  (readResult_3_bits),
    .readResult_4_valid                 (readResult_4_valid),
    .readResult_4_bits                  (readResult_4_bits),
    .readResult_5_valid                 (readResult_5_valid),
    .readResult_5_bits                  (readResult_5_bits),
    .readResult_6_valid                 (readResult_6_valid),
    .readResult_6_bits                  (readResult_6_bits),
    .readResult_7_valid                 (readResult_7_valid),
    .readResult_7_bits                  (readResult_7_bits),
    .readResult_8_valid                 (readResult_8_valid),
    .readResult_8_bits                  (readResult_8_bits),
    .readResult_9_valid                 (readResult_9_valid),
    .readResult_9_bits                  (readResult_9_bits),
    .readResult_10_valid                (readResult_10_valid),
    .readResult_10_bits                 (readResult_10_bits),
    .readResult_11_valid                (readResult_11_valid),
    .readResult_11_bits                 (readResult_11_bits),
    .readResult_12_valid                (readResult_12_valid),
    .readResult_12_bits                 (readResult_12_bits),
    .readResult_13_valid                (readResult_13_valid),
    .readResult_13_bits                 (readResult_13_bits),
    .readResult_14_valid                (readResult_14_valid),
    .readResult_14_bits                 (readResult_14_bits),
    .readResult_15_valid                (readResult_15_valid),
    .readResult_15_bits                 (readResult_15_bits),
    .readResult_16_valid                (readResult_16_valid),
    .readResult_16_bits                 (readResult_16_bits),
    .readResult_17_valid                (readResult_17_valid),
    .readResult_17_bits                 (readResult_17_bits),
    .readResult_18_valid                (readResult_18_valid),
    .readResult_18_bits                 (readResult_18_bits),
    .readResult_19_valid                (readResult_19_valid),
    .readResult_19_bits                 (readResult_19_bits),
    .readResult_20_valid                (readResult_20_valid),
    .readResult_20_bits                 (readResult_20_bits),
    .readResult_21_valid                (readResult_21_valid),
    .readResult_21_bits                 (readResult_21_bits),
    .readResult_22_valid                (readResult_22_valid),
    .readResult_22_bits                 (readResult_22_bits),
    .readResult_23_valid                (readResult_23_valid),
    .readResult_23_bits                 (readResult_23_bits),
    .readResult_24_valid                (readResult_24_valid),
    .readResult_24_bits                 (readResult_24_bits),
    .readResult_25_valid                (readResult_25_valid),
    .readResult_25_bits                 (readResult_25_bits),
    .readResult_26_valid                (readResult_26_valid),
    .readResult_26_bits                 (readResult_26_bits),
    .readResult_27_valid                (readResult_27_valid),
    .readResult_27_bits                 (readResult_27_bits),
    .readResult_28_valid                (readResult_28_valid),
    .readResult_28_bits                 (readResult_28_bits),
    .readResult_29_valid                (readResult_29_valid),
    .readResult_29_bits                 (readResult_29_bits),
    .readResult_30_valid                (readResult_30_valid),
    .readResult_30_bits                 (readResult_30_bits),
    .readResult_31_valid                (readResult_31_valid),
    .readResult_31_bits                 (readResult_31_bits),
    .stageClear                         (_maskedWrite_stageClear)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_0_enq_ready & exeRequestQueue_0_enq_valid & ~(_exeRequestQueue_queue_fifo_empty & exeRequestQueue_0_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_0_deq_ready & ~_exeRequestQueue_queue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn),
    .empty        (_exeRequestQueue_queue_fifo_empty),
    .almost_empty (exeRequestQueue_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_0_almostFull),
    .full         (_exeRequestQueue_queue_fifo_full),
    .error        (_exeRequestQueue_queue_fifo_error),
    .data_out     (_exeRequestQueue_queue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_1_enq_ready & exeRequestQueue_1_enq_valid & ~(_exeRequestQueue_queue_fifo_1_empty & exeRequestQueue_1_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_1_deq_ready & ~_exeRequestQueue_queue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_1),
    .empty        (_exeRequestQueue_queue_fifo_1_empty),
    .almost_empty (exeRequestQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_1_almostFull),
    .full         (_exeRequestQueue_queue_fifo_1_full),
    .error        (_exeRequestQueue_queue_fifo_1_error),
    .data_out     (_exeRequestQueue_queue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_2_enq_ready & exeRequestQueue_2_enq_valid & ~(_exeRequestQueue_queue_fifo_2_empty & exeRequestQueue_2_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_2_deq_ready & ~_exeRequestQueue_queue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_2),
    .empty        (_exeRequestQueue_queue_fifo_2_empty),
    .almost_empty (exeRequestQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_2_almostFull),
    .full         (_exeRequestQueue_queue_fifo_2_full),
    .error        (_exeRequestQueue_queue_fifo_2_error),
    .data_out     (_exeRequestQueue_queue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_3_enq_ready & exeRequestQueue_3_enq_valid & ~(_exeRequestQueue_queue_fifo_3_empty & exeRequestQueue_3_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_3_deq_ready & ~_exeRequestQueue_queue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_3),
    .empty        (_exeRequestQueue_queue_fifo_3_empty),
    .almost_empty (exeRequestQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_3_almostFull),
    .full         (_exeRequestQueue_queue_fifo_3_full),
    .error        (_exeRequestQueue_queue_fifo_3_error),
    .data_out     (_exeRequestQueue_queue_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_4_enq_ready & exeRequestQueue_4_enq_valid & ~(_exeRequestQueue_queue_fifo_4_empty & exeRequestQueue_4_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_4_deq_ready & ~_exeRequestQueue_queue_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_4),
    .empty        (_exeRequestQueue_queue_fifo_4_empty),
    .almost_empty (exeRequestQueue_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_4_almostFull),
    .full         (_exeRequestQueue_queue_fifo_4_full),
    .error        (_exeRequestQueue_queue_fifo_4_error),
    .data_out     (_exeRequestQueue_queue_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_5_enq_ready & exeRequestQueue_5_enq_valid & ~(_exeRequestQueue_queue_fifo_5_empty & exeRequestQueue_5_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_5_deq_ready & ~_exeRequestQueue_queue_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_5),
    .empty        (_exeRequestQueue_queue_fifo_5_empty),
    .almost_empty (exeRequestQueue_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_5_almostFull),
    .full         (_exeRequestQueue_queue_fifo_5_full),
    .error        (_exeRequestQueue_queue_fifo_5_error),
    .data_out     (_exeRequestQueue_queue_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_6_enq_ready & exeRequestQueue_6_enq_valid & ~(_exeRequestQueue_queue_fifo_6_empty & exeRequestQueue_6_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_6_deq_ready & ~_exeRequestQueue_queue_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_6),
    .empty        (_exeRequestQueue_queue_fifo_6_empty),
    .almost_empty (exeRequestQueue_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_6_almostFull),
    .full         (_exeRequestQueue_queue_fifo_6_full),
    .error        (_exeRequestQueue_queue_fifo_6_error),
    .data_out     (_exeRequestQueue_queue_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_7_enq_ready & exeRequestQueue_7_enq_valid & ~(_exeRequestQueue_queue_fifo_7_empty & exeRequestQueue_7_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_7_deq_ready & ~_exeRequestQueue_queue_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_7),
    .empty        (_exeRequestQueue_queue_fifo_7_empty),
    .almost_empty (exeRequestQueue_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_7_almostFull),
    .full         (_exeRequestQueue_queue_fifo_7_full),
    .error        (_exeRequestQueue_queue_fifo_7_error),
    .data_out     (_exeRequestQueue_queue_fifo_7_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_8_enq_ready & exeRequestQueue_8_enq_valid & ~(_exeRequestQueue_queue_fifo_8_empty & exeRequestQueue_8_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_8_deq_ready & ~_exeRequestQueue_queue_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_8),
    .empty        (_exeRequestQueue_queue_fifo_8_empty),
    .almost_empty (exeRequestQueue_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_8_almostFull),
    .full         (_exeRequestQueue_queue_fifo_8_full),
    .error        (_exeRequestQueue_queue_fifo_8_error),
    .data_out     (_exeRequestQueue_queue_fifo_8_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_9_enq_ready & exeRequestQueue_9_enq_valid & ~(_exeRequestQueue_queue_fifo_9_empty & exeRequestQueue_9_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_9_deq_ready & ~_exeRequestQueue_queue_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_9),
    .empty        (_exeRequestQueue_queue_fifo_9_empty),
    .almost_empty (exeRequestQueue_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_9_almostFull),
    .full         (_exeRequestQueue_queue_fifo_9_full),
    .error        (_exeRequestQueue_queue_fifo_9_error),
    .data_out     (_exeRequestQueue_queue_fifo_9_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_10_enq_ready & exeRequestQueue_10_enq_valid & ~(_exeRequestQueue_queue_fifo_10_empty & exeRequestQueue_10_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_10_deq_ready & ~_exeRequestQueue_queue_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_10),
    .empty        (_exeRequestQueue_queue_fifo_10_empty),
    .almost_empty (exeRequestQueue_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_10_almostFull),
    .full         (_exeRequestQueue_queue_fifo_10_full),
    .error        (_exeRequestQueue_queue_fifo_10_error),
    .data_out     (_exeRequestQueue_queue_fifo_10_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_11_enq_ready & exeRequestQueue_11_enq_valid & ~(_exeRequestQueue_queue_fifo_11_empty & exeRequestQueue_11_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_11_deq_ready & ~_exeRequestQueue_queue_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_11),
    .empty        (_exeRequestQueue_queue_fifo_11_empty),
    .almost_empty (exeRequestQueue_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_11_almostFull),
    .full         (_exeRequestQueue_queue_fifo_11_full),
    .error        (_exeRequestQueue_queue_fifo_11_error),
    .data_out     (_exeRequestQueue_queue_fifo_11_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_12_enq_ready & exeRequestQueue_12_enq_valid & ~(_exeRequestQueue_queue_fifo_12_empty & exeRequestQueue_12_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_12_deq_ready & ~_exeRequestQueue_queue_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_12),
    .empty        (_exeRequestQueue_queue_fifo_12_empty),
    .almost_empty (exeRequestQueue_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_12_almostFull),
    .full         (_exeRequestQueue_queue_fifo_12_full),
    .error        (_exeRequestQueue_queue_fifo_12_error),
    .data_out     (_exeRequestQueue_queue_fifo_12_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_13_enq_ready & exeRequestQueue_13_enq_valid & ~(_exeRequestQueue_queue_fifo_13_empty & exeRequestQueue_13_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_13_deq_ready & ~_exeRequestQueue_queue_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_13),
    .empty        (_exeRequestQueue_queue_fifo_13_empty),
    .almost_empty (exeRequestQueue_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_13_almostFull),
    .full         (_exeRequestQueue_queue_fifo_13_full),
    .error        (_exeRequestQueue_queue_fifo_13_error),
    .data_out     (_exeRequestQueue_queue_fifo_13_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_14_enq_ready & exeRequestQueue_14_enq_valid & ~(_exeRequestQueue_queue_fifo_14_empty & exeRequestQueue_14_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_14_deq_ready & ~_exeRequestQueue_queue_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_14),
    .empty        (_exeRequestQueue_queue_fifo_14_empty),
    .almost_empty (exeRequestQueue_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_14_almostFull),
    .full         (_exeRequestQueue_queue_fifo_14_full),
    .error        (_exeRequestQueue_queue_fifo_14_error),
    .data_out     (_exeRequestQueue_queue_fifo_14_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_15_enq_ready & exeRequestQueue_15_enq_valid & ~(_exeRequestQueue_queue_fifo_15_empty & exeRequestQueue_15_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_15_deq_ready & ~_exeRequestQueue_queue_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_15),
    .empty        (_exeRequestQueue_queue_fifo_15_empty),
    .almost_empty (exeRequestQueue_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_15_almostFull),
    .full         (_exeRequestQueue_queue_fifo_15_full),
    .error        (_exeRequestQueue_queue_fifo_15_error),
    .data_out     (_exeRequestQueue_queue_fifo_15_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_16 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_16_enq_ready & exeRequestQueue_16_enq_valid & ~(_exeRequestQueue_queue_fifo_16_empty & exeRequestQueue_16_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_16_deq_ready & ~_exeRequestQueue_queue_fifo_16_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_16),
    .empty        (_exeRequestQueue_queue_fifo_16_empty),
    .almost_empty (exeRequestQueue_16_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_16_almostFull),
    .full         (_exeRequestQueue_queue_fifo_16_full),
    .error        (_exeRequestQueue_queue_fifo_16_error),
    .data_out     (_exeRequestQueue_queue_fifo_16_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_17 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_17_enq_ready & exeRequestQueue_17_enq_valid & ~(_exeRequestQueue_queue_fifo_17_empty & exeRequestQueue_17_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_17_deq_ready & ~_exeRequestQueue_queue_fifo_17_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_17),
    .empty        (_exeRequestQueue_queue_fifo_17_empty),
    .almost_empty (exeRequestQueue_17_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_17_almostFull),
    .full         (_exeRequestQueue_queue_fifo_17_full),
    .error        (_exeRequestQueue_queue_fifo_17_error),
    .data_out     (_exeRequestQueue_queue_fifo_17_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_18 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_18_enq_ready & exeRequestQueue_18_enq_valid & ~(_exeRequestQueue_queue_fifo_18_empty & exeRequestQueue_18_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_18_deq_ready & ~_exeRequestQueue_queue_fifo_18_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_18),
    .empty        (_exeRequestQueue_queue_fifo_18_empty),
    .almost_empty (exeRequestQueue_18_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_18_almostFull),
    .full         (_exeRequestQueue_queue_fifo_18_full),
    .error        (_exeRequestQueue_queue_fifo_18_error),
    .data_out     (_exeRequestQueue_queue_fifo_18_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_19 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_19_enq_ready & exeRequestQueue_19_enq_valid & ~(_exeRequestQueue_queue_fifo_19_empty & exeRequestQueue_19_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_19_deq_ready & ~_exeRequestQueue_queue_fifo_19_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_19),
    .empty        (_exeRequestQueue_queue_fifo_19_empty),
    .almost_empty (exeRequestQueue_19_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_19_almostFull),
    .full         (_exeRequestQueue_queue_fifo_19_full),
    .error        (_exeRequestQueue_queue_fifo_19_error),
    .data_out     (_exeRequestQueue_queue_fifo_19_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_20 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_20_enq_ready & exeRequestQueue_20_enq_valid & ~(_exeRequestQueue_queue_fifo_20_empty & exeRequestQueue_20_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_20_deq_ready & ~_exeRequestQueue_queue_fifo_20_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_20),
    .empty        (_exeRequestQueue_queue_fifo_20_empty),
    .almost_empty (exeRequestQueue_20_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_20_almostFull),
    .full         (_exeRequestQueue_queue_fifo_20_full),
    .error        (_exeRequestQueue_queue_fifo_20_error),
    .data_out     (_exeRequestQueue_queue_fifo_20_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_21 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_21_enq_ready & exeRequestQueue_21_enq_valid & ~(_exeRequestQueue_queue_fifo_21_empty & exeRequestQueue_21_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_21_deq_ready & ~_exeRequestQueue_queue_fifo_21_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_21),
    .empty        (_exeRequestQueue_queue_fifo_21_empty),
    .almost_empty (exeRequestQueue_21_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_21_almostFull),
    .full         (_exeRequestQueue_queue_fifo_21_full),
    .error        (_exeRequestQueue_queue_fifo_21_error),
    .data_out     (_exeRequestQueue_queue_fifo_21_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_22 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_22_enq_ready & exeRequestQueue_22_enq_valid & ~(_exeRequestQueue_queue_fifo_22_empty & exeRequestQueue_22_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_22_deq_ready & ~_exeRequestQueue_queue_fifo_22_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_22),
    .empty        (_exeRequestQueue_queue_fifo_22_empty),
    .almost_empty (exeRequestQueue_22_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_22_almostFull),
    .full         (_exeRequestQueue_queue_fifo_22_full),
    .error        (_exeRequestQueue_queue_fifo_22_error),
    .data_out     (_exeRequestQueue_queue_fifo_22_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_23 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_23_enq_ready & exeRequestQueue_23_enq_valid & ~(_exeRequestQueue_queue_fifo_23_empty & exeRequestQueue_23_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_23_deq_ready & ~_exeRequestQueue_queue_fifo_23_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_23),
    .empty        (_exeRequestQueue_queue_fifo_23_empty),
    .almost_empty (exeRequestQueue_23_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_23_almostFull),
    .full         (_exeRequestQueue_queue_fifo_23_full),
    .error        (_exeRequestQueue_queue_fifo_23_error),
    .data_out     (_exeRequestQueue_queue_fifo_23_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_24 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_24_enq_ready & exeRequestQueue_24_enq_valid & ~(_exeRequestQueue_queue_fifo_24_empty & exeRequestQueue_24_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_24_deq_ready & ~_exeRequestQueue_queue_fifo_24_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_24),
    .empty        (_exeRequestQueue_queue_fifo_24_empty),
    .almost_empty (exeRequestQueue_24_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_24_almostFull),
    .full         (_exeRequestQueue_queue_fifo_24_full),
    .error        (_exeRequestQueue_queue_fifo_24_error),
    .data_out     (_exeRequestQueue_queue_fifo_24_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_25 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_25_enq_ready & exeRequestQueue_25_enq_valid & ~(_exeRequestQueue_queue_fifo_25_empty & exeRequestQueue_25_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_25_deq_ready & ~_exeRequestQueue_queue_fifo_25_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_25),
    .empty        (_exeRequestQueue_queue_fifo_25_empty),
    .almost_empty (exeRequestQueue_25_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_25_almostFull),
    .full         (_exeRequestQueue_queue_fifo_25_full),
    .error        (_exeRequestQueue_queue_fifo_25_error),
    .data_out     (_exeRequestQueue_queue_fifo_25_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_26 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_26_enq_ready & exeRequestQueue_26_enq_valid & ~(_exeRequestQueue_queue_fifo_26_empty & exeRequestQueue_26_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_26_deq_ready & ~_exeRequestQueue_queue_fifo_26_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_26),
    .empty        (_exeRequestQueue_queue_fifo_26_empty),
    .almost_empty (exeRequestQueue_26_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_26_almostFull),
    .full         (_exeRequestQueue_queue_fifo_26_full),
    .error        (_exeRequestQueue_queue_fifo_26_error),
    .data_out     (_exeRequestQueue_queue_fifo_26_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_27 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_27_enq_ready & exeRequestQueue_27_enq_valid & ~(_exeRequestQueue_queue_fifo_27_empty & exeRequestQueue_27_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_27_deq_ready & ~_exeRequestQueue_queue_fifo_27_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_27),
    .empty        (_exeRequestQueue_queue_fifo_27_empty),
    .almost_empty (exeRequestQueue_27_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_27_almostFull),
    .full         (_exeRequestQueue_queue_fifo_27_full),
    .error        (_exeRequestQueue_queue_fifo_27_error),
    .data_out     (_exeRequestQueue_queue_fifo_27_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_28 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_28_enq_ready & exeRequestQueue_28_enq_valid & ~(_exeRequestQueue_queue_fifo_28_empty & exeRequestQueue_28_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_28_deq_ready & ~_exeRequestQueue_queue_fifo_28_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_28),
    .empty        (_exeRequestQueue_queue_fifo_28_empty),
    .almost_empty (exeRequestQueue_28_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_28_almostFull),
    .full         (_exeRequestQueue_queue_fifo_28_full),
    .error        (_exeRequestQueue_queue_fifo_28_error),
    .data_out     (_exeRequestQueue_queue_fifo_28_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_29 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_29_enq_ready & exeRequestQueue_29_enq_valid & ~(_exeRequestQueue_queue_fifo_29_empty & exeRequestQueue_29_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_29_deq_ready & ~_exeRequestQueue_queue_fifo_29_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_29),
    .empty        (_exeRequestQueue_queue_fifo_29_empty),
    .almost_empty (exeRequestQueue_29_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_29_almostFull),
    .full         (_exeRequestQueue_queue_fifo_29_full),
    .error        (_exeRequestQueue_queue_fifo_29_error),
    .data_out     (_exeRequestQueue_queue_fifo_29_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_30 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_30_enq_ready & exeRequestQueue_30_enq_valid & ~(_exeRequestQueue_queue_fifo_30_empty & exeRequestQueue_30_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_30_deq_ready & ~_exeRequestQueue_queue_fifo_30_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_30),
    .empty        (_exeRequestQueue_queue_fifo_30_empty),
    .almost_empty (exeRequestQueue_30_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_30_almostFull),
    .full         (_exeRequestQueue_queue_fifo_30_full),
    .error        (_exeRequestQueue_queue_fifo_30_error),
    .data_out     (_exeRequestQueue_queue_fifo_30_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_31 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_31_enq_ready & exeRequestQueue_31_enq_valid & ~(_exeRequestQueue_queue_fifo_31_empty & exeRequestQueue_31_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_31_deq_ready & ~_exeRequestQueue_queue_fifo_31_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_31),
    .empty        (_exeRequestQueue_queue_fifo_31_empty),
    .almost_empty (exeRequestQueue_31_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_31_almostFull),
    .full         (_exeRequestQueue_queue_fifo_31_full),
    .error        (_exeRequestQueue_queue_fifo_31_error),
    .data_out     (_exeRequestQueue_queue_fifo_31_data_out)
  );
  SlideIndexGen slideAddressGen (
    .clock                              (clock),
    .reset                              (reset),
    .newInstruction                     (instReq_valid & (|instReq_bits_vl)),
    .instructionReq_decodeResult_topUop (instReg_decodeResult_topUop),
    .instructionReq_readFromScala       (instReg_readFromScala),
    .instructionReq_sew                 (instReg_sew),
    .instructionReq_vlmul               (instReg_vlmul),
    .instructionReq_maskType            (instReg_maskType),
    .instructionReq_vl                  (instReg_vl),
    .indexDeq_ready                     (slideAddressGen_indexDeq_ready),
    .indexDeq_valid                     (_slideAddressGen_indexDeq_valid),
    .indexDeq_bits_needRead             (_slideAddressGen_indexDeq_bits_needRead),
    .indexDeq_bits_elementValid         (_slideAddressGen_indexDeq_bits_elementValid),
    .indexDeq_bits_replaceVs1           (_slideAddressGen_indexDeq_bits_replaceVs1),
    .indexDeq_bits_readOffset           (_slideAddressGen_indexDeq_bits_readOffset),
    .indexDeq_bits_accessLane_0         (_slideAddressGen_indexDeq_bits_accessLane_0),
    .indexDeq_bits_accessLane_1         (_slideAddressGen_indexDeq_bits_accessLane_1),
    .indexDeq_bits_accessLane_2         (_slideAddressGen_indexDeq_bits_accessLane_2),
    .indexDeq_bits_accessLane_3         (_slideAddressGen_indexDeq_bits_accessLane_3),
    .indexDeq_bits_accessLane_4         (_slideAddressGen_indexDeq_bits_accessLane_4),
    .indexDeq_bits_accessLane_5         (_slideAddressGen_indexDeq_bits_accessLane_5),
    .indexDeq_bits_accessLane_6         (_slideAddressGen_indexDeq_bits_accessLane_6),
    .indexDeq_bits_accessLane_7         (_slideAddressGen_indexDeq_bits_accessLane_7),
    .indexDeq_bits_accessLane_8         (_slideAddressGen_indexDeq_bits_accessLane_8),
    .indexDeq_bits_accessLane_9         (_slideAddressGen_indexDeq_bits_accessLane_9),
    .indexDeq_bits_accessLane_10        (_slideAddressGen_indexDeq_bits_accessLane_10),
    .indexDeq_bits_accessLane_11        (_slideAddressGen_indexDeq_bits_accessLane_11),
    .indexDeq_bits_accessLane_12        (_slideAddressGen_indexDeq_bits_accessLane_12),
    .indexDeq_bits_accessLane_13        (_slideAddressGen_indexDeq_bits_accessLane_13),
    .indexDeq_bits_accessLane_14        (_slideAddressGen_indexDeq_bits_accessLane_14),
    .indexDeq_bits_accessLane_15        (_slideAddressGen_indexDeq_bits_accessLane_15),
    .indexDeq_bits_accessLane_16        (_slideAddressGen_indexDeq_bits_accessLane_16),
    .indexDeq_bits_accessLane_17        (_slideAddressGen_indexDeq_bits_accessLane_17),
    .indexDeq_bits_accessLane_18        (_slideAddressGen_indexDeq_bits_accessLane_18),
    .indexDeq_bits_accessLane_19        (_slideAddressGen_indexDeq_bits_accessLane_19),
    .indexDeq_bits_accessLane_20        (_slideAddressGen_indexDeq_bits_accessLane_20),
    .indexDeq_bits_accessLane_21        (_slideAddressGen_indexDeq_bits_accessLane_21),
    .indexDeq_bits_accessLane_22        (_slideAddressGen_indexDeq_bits_accessLane_22),
    .indexDeq_bits_accessLane_23        (_slideAddressGen_indexDeq_bits_accessLane_23),
    .indexDeq_bits_accessLane_24        (_slideAddressGen_indexDeq_bits_accessLane_24),
    .indexDeq_bits_accessLane_25        (_slideAddressGen_indexDeq_bits_accessLane_25),
    .indexDeq_bits_accessLane_26        (_slideAddressGen_indexDeq_bits_accessLane_26),
    .indexDeq_bits_accessLane_27        (_slideAddressGen_indexDeq_bits_accessLane_27),
    .indexDeq_bits_accessLane_28        (_slideAddressGen_indexDeq_bits_accessLane_28),
    .indexDeq_bits_accessLane_29        (_slideAddressGen_indexDeq_bits_accessLane_29),
    .indexDeq_bits_accessLane_30        (_slideAddressGen_indexDeq_bits_accessLane_30),
    .indexDeq_bits_accessLane_31        (_slideAddressGen_indexDeq_bits_accessLane_31),
    .indexDeq_bits_vsGrowth_0           (_slideAddressGen_indexDeq_bits_vsGrowth_0),
    .indexDeq_bits_vsGrowth_1           (_slideAddressGen_indexDeq_bits_vsGrowth_1),
    .indexDeq_bits_vsGrowth_2           (_slideAddressGen_indexDeq_bits_vsGrowth_2),
    .indexDeq_bits_vsGrowth_3           (_slideAddressGen_indexDeq_bits_vsGrowth_3),
    .indexDeq_bits_vsGrowth_4           (_slideAddressGen_indexDeq_bits_vsGrowth_4),
    .indexDeq_bits_vsGrowth_5           (_slideAddressGen_indexDeq_bits_vsGrowth_5),
    .indexDeq_bits_vsGrowth_6           (_slideAddressGen_indexDeq_bits_vsGrowth_6),
    .indexDeq_bits_vsGrowth_7           (_slideAddressGen_indexDeq_bits_vsGrowth_7),
    .indexDeq_bits_vsGrowth_8           (_slideAddressGen_indexDeq_bits_vsGrowth_8),
    .indexDeq_bits_vsGrowth_9           (_slideAddressGen_indexDeq_bits_vsGrowth_9),
    .indexDeq_bits_vsGrowth_10          (_slideAddressGen_indexDeq_bits_vsGrowth_10),
    .indexDeq_bits_vsGrowth_11          (_slideAddressGen_indexDeq_bits_vsGrowth_11),
    .indexDeq_bits_vsGrowth_12          (_slideAddressGen_indexDeq_bits_vsGrowth_12),
    .indexDeq_bits_vsGrowth_13          (_slideAddressGen_indexDeq_bits_vsGrowth_13),
    .indexDeq_bits_vsGrowth_14          (_slideAddressGen_indexDeq_bits_vsGrowth_14),
    .indexDeq_bits_vsGrowth_15          (_slideAddressGen_indexDeq_bits_vsGrowth_15),
    .indexDeq_bits_vsGrowth_16          (_slideAddressGen_indexDeq_bits_vsGrowth_16),
    .indexDeq_bits_vsGrowth_17          (_slideAddressGen_indexDeq_bits_vsGrowth_17),
    .indexDeq_bits_vsGrowth_18          (_slideAddressGen_indexDeq_bits_vsGrowth_18),
    .indexDeq_bits_vsGrowth_19          (_slideAddressGen_indexDeq_bits_vsGrowth_19),
    .indexDeq_bits_vsGrowth_20          (_slideAddressGen_indexDeq_bits_vsGrowth_20),
    .indexDeq_bits_vsGrowth_21          (_slideAddressGen_indexDeq_bits_vsGrowth_21),
    .indexDeq_bits_vsGrowth_22          (_slideAddressGen_indexDeq_bits_vsGrowth_22),
    .indexDeq_bits_vsGrowth_23          (_slideAddressGen_indexDeq_bits_vsGrowth_23),
    .indexDeq_bits_vsGrowth_24          (_slideAddressGen_indexDeq_bits_vsGrowth_24),
    .indexDeq_bits_vsGrowth_25          (_slideAddressGen_indexDeq_bits_vsGrowth_25),
    .indexDeq_bits_vsGrowth_26          (_slideAddressGen_indexDeq_bits_vsGrowth_26),
    .indexDeq_bits_vsGrowth_27          (_slideAddressGen_indexDeq_bits_vsGrowth_27),
    .indexDeq_bits_vsGrowth_28          (_slideAddressGen_indexDeq_bits_vsGrowth_28),
    .indexDeq_bits_vsGrowth_29          (_slideAddressGen_indexDeq_bits_vsGrowth_29),
    .indexDeq_bits_vsGrowth_30          (_slideAddressGen_indexDeq_bits_vsGrowth_30),
    .indexDeq_bits_vsGrowth_31          (_slideAddressGen_indexDeq_bits_vsGrowth_31),
    .indexDeq_bits_executeGroup         (_slideAddressGen_indexDeq_bits_executeGroup),
    .indexDeq_bits_readDataOffset       (_slideAddressGen_indexDeq_bits_readDataOffset),
    .indexDeq_bits_last                 (_slideAddressGen_indexDeq_bits_last),
    .slideGroupOut                      (_slideAddressGen_slideGroupOut),
    .slideMaskInput                     (_GEN_64[_slideAddressGen_slideGroupOut[5:0]])
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(192)
  ) accessCountQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(accessCountQueue_enq_ready & accessCountQueue_enq_valid)),
    .pop_req_n    (~(accessCountQueue_deq_ready & ~_accessCountQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (accessCountQueue_dataIn),
    .empty        (_accessCountQueue_fifo_empty),
    .almost_empty (accessCountQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (accessCountQueue_almostFull),
    .full         (_accessCountQueue_fifo_full),
    .error        (_accessCountQueue_fifo_error),
    .data_out     (_accessCountQueue_fifo_data_out)
  );
  MaskUnitReadCrossBar readCrossBar (
    .input_0_ready             (_readCrossBar_input_0_ready),
    .input_0_valid             (readCrossBar_input_0_valid),
    .input_0_bits_vs           (selectExecuteReq_0_bits_vs),
    .input_0_bits_offset       (selectExecuteReq_0_bits_offset),
    .input_0_bits_readLane     (selectExecuteReq_0_bits_readLane),
    .input_0_bits_dataOffset   (selectExecuteReq_0_bits_dataOffset),
    .input_1_ready             (_readCrossBar_input_1_ready),
    .input_1_valid             (readCrossBar_input_1_valid),
    .input_1_bits_vs           (selectExecuteReq_1_bits_vs),
    .input_1_bits_offset       (selectExecuteReq_1_bits_offset),
    .input_1_bits_readLane     (selectExecuteReq_1_bits_readLane),
    .input_1_bits_dataOffset   (selectExecuteReq_1_bits_dataOffset),
    .input_2_ready             (_readCrossBar_input_2_ready),
    .input_2_valid             (readCrossBar_input_2_valid),
    .input_2_bits_vs           (selectExecuteReq_2_bits_vs),
    .input_2_bits_offset       (selectExecuteReq_2_bits_offset),
    .input_2_bits_readLane     (selectExecuteReq_2_bits_readLane),
    .input_2_bits_dataOffset   (selectExecuteReq_2_bits_dataOffset),
    .input_3_ready             (_readCrossBar_input_3_ready),
    .input_3_valid             (readCrossBar_input_3_valid),
    .input_3_bits_vs           (selectExecuteReq_3_bits_vs),
    .input_3_bits_offset       (selectExecuteReq_3_bits_offset),
    .input_3_bits_readLane     (selectExecuteReq_3_bits_readLane),
    .input_3_bits_dataOffset   (selectExecuteReq_3_bits_dataOffset),
    .input_4_ready             (_readCrossBar_input_4_ready),
    .input_4_valid             (readCrossBar_input_4_valid),
    .input_4_bits_vs           (selectExecuteReq_4_bits_vs),
    .input_4_bits_offset       (selectExecuteReq_4_bits_offset),
    .input_4_bits_readLane     (selectExecuteReq_4_bits_readLane),
    .input_4_bits_dataOffset   (selectExecuteReq_4_bits_dataOffset),
    .input_5_ready             (_readCrossBar_input_5_ready),
    .input_5_valid             (readCrossBar_input_5_valid),
    .input_5_bits_vs           (selectExecuteReq_5_bits_vs),
    .input_5_bits_offset       (selectExecuteReq_5_bits_offset),
    .input_5_bits_readLane     (selectExecuteReq_5_bits_readLane),
    .input_5_bits_dataOffset   (selectExecuteReq_5_bits_dataOffset),
    .input_6_ready             (_readCrossBar_input_6_ready),
    .input_6_valid             (readCrossBar_input_6_valid),
    .input_6_bits_vs           (selectExecuteReq_6_bits_vs),
    .input_6_bits_offset       (selectExecuteReq_6_bits_offset),
    .input_6_bits_readLane     (selectExecuteReq_6_bits_readLane),
    .input_6_bits_dataOffset   (selectExecuteReq_6_bits_dataOffset),
    .input_7_ready             (_readCrossBar_input_7_ready),
    .input_7_valid             (readCrossBar_input_7_valid),
    .input_7_bits_vs           (selectExecuteReq_7_bits_vs),
    .input_7_bits_offset       (selectExecuteReq_7_bits_offset),
    .input_7_bits_readLane     (selectExecuteReq_7_bits_readLane),
    .input_7_bits_dataOffset   (selectExecuteReq_7_bits_dataOffset),
    .input_8_ready             (_readCrossBar_input_8_ready),
    .input_8_valid             (readCrossBar_input_8_valid),
    .input_8_bits_vs           (selectExecuteReq_8_bits_vs),
    .input_8_bits_offset       (selectExecuteReq_8_bits_offset),
    .input_8_bits_readLane     (selectExecuteReq_8_bits_readLane),
    .input_8_bits_dataOffset   (selectExecuteReq_8_bits_dataOffset),
    .input_9_ready             (_readCrossBar_input_9_ready),
    .input_9_valid             (readCrossBar_input_9_valid),
    .input_9_bits_vs           (selectExecuteReq_9_bits_vs),
    .input_9_bits_offset       (selectExecuteReq_9_bits_offset),
    .input_9_bits_readLane     (selectExecuteReq_9_bits_readLane),
    .input_9_bits_dataOffset   (selectExecuteReq_9_bits_dataOffset),
    .input_10_ready            (_readCrossBar_input_10_ready),
    .input_10_valid            (readCrossBar_input_10_valid),
    .input_10_bits_vs          (selectExecuteReq_10_bits_vs),
    .input_10_bits_offset      (selectExecuteReq_10_bits_offset),
    .input_10_bits_readLane    (selectExecuteReq_10_bits_readLane),
    .input_10_bits_dataOffset  (selectExecuteReq_10_bits_dataOffset),
    .input_11_ready            (_readCrossBar_input_11_ready),
    .input_11_valid            (readCrossBar_input_11_valid),
    .input_11_bits_vs          (selectExecuteReq_11_bits_vs),
    .input_11_bits_offset      (selectExecuteReq_11_bits_offset),
    .input_11_bits_readLane    (selectExecuteReq_11_bits_readLane),
    .input_11_bits_dataOffset  (selectExecuteReq_11_bits_dataOffset),
    .input_12_ready            (_readCrossBar_input_12_ready),
    .input_12_valid            (readCrossBar_input_12_valid),
    .input_12_bits_vs          (selectExecuteReq_12_bits_vs),
    .input_12_bits_offset      (selectExecuteReq_12_bits_offset),
    .input_12_bits_readLane    (selectExecuteReq_12_bits_readLane),
    .input_12_bits_dataOffset  (selectExecuteReq_12_bits_dataOffset),
    .input_13_ready            (_readCrossBar_input_13_ready),
    .input_13_valid            (readCrossBar_input_13_valid),
    .input_13_bits_vs          (selectExecuteReq_13_bits_vs),
    .input_13_bits_offset      (selectExecuteReq_13_bits_offset),
    .input_13_bits_readLane    (selectExecuteReq_13_bits_readLane),
    .input_13_bits_dataOffset  (selectExecuteReq_13_bits_dataOffset),
    .input_14_ready            (_readCrossBar_input_14_ready),
    .input_14_valid            (readCrossBar_input_14_valid),
    .input_14_bits_vs          (selectExecuteReq_14_bits_vs),
    .input_14_bits_offset      (selectExecuteReq_14_bits_offset),
    .input_14_bits_readLane    (selectExecuteReq_14_bits_readLane),
    .input_14_bits_dataOffset  (selectExecuteReq_14_bits_dataOffset),
    .input_15_ready            (_readCrossBar_input_15_ready),
    .input_15_valid            (readCrossBar_input_15_valid),
    .input_15_bits_vs          (selectExecuteReq_15_bits_vs),
    .input_15_bits_offset      (selectExecuteReq_15_bits_offset),
    .input_15_bits_readLane    (selectExecuteReq_15_bits_readLane),
    .input_15_bits_dataOffset  (selectExecuteReq_15_bits_dataOffset),
    .input_16_ready            (_readCrossBar_input_16_ready),
    .input_16_valid            (readCrossBar_input_16_valid),
    .input_16_bits_vs          (selectExecuteReq_16_bits_vs),
    .input_16_bits_offset      (selectExecuteReq_16_bits_offset),
    .input_16_bits_readLane    (selectExecuteReq_16_bits_readLane),
    .input_16_bits_dataOffset  (selectExecuteReq_16_bits_dataOffset),
    .input_17_ready            (_readCrossBar_input_17_ready),
    .input_17_valid            (readCrossBar_input_17_valid),
    .input_17_bits_vs          (selectExecuteReq_17_bits_vs),
    .input_17_bits_offset      (selectExecuteReq_17_bits_offset),
    .input_17_bits_readLane    (selectExecuteReq_17_bits_readLane),
    .input_17_bits_dataOffset  (selectExecuteReq_17_bits_dataOffset),
    .input_18_ready            (_readCrossBar_input_18_ready),
    .input_18_valid            (readCrossBar_input_18_valid),
    .input_18_bits_vs          (selectExecuteReq_18_bits_vs),
    .input_18_bits_offset      (selectExecuteReq_18_bits_offset),
    .input_18_bits_readLane    (selectExecuteReq_18_bits_readLane),
    .input_18_bits_dataOffset  (selectExecuteReq_18_bits_dataOffset),
    .input_19_ready            (_readCrossBar_input_19_ready),
    .input_19_valid            (readCrossBar_input_19_valid),
    .input_19_bits_vs          (selectExecuteReq_19_bits_vs),
    .input_19_bits_offset      (selectExecuteReq_19_bits_offset),
    .input_19_bits_readLane    (selectExecuteReq_19_bits_readLane),
    .input_19_bits_dataOffset  (selectExecuteReq_19_bits_dataOffset),
    .input_20_ready            (_readCrossBar_input_20_ready),
    .input_20_valid            (readCrossBar_input_20_valid),
    .input_20_bits_vs          (selectExecuteReq_20_bits_vs),
    .input_20_bits_offset      (selectExecuteReq_20_bits_offset),
    .input_20_bits_readLane    (selectExecuteReq_20_bits_readLane),
    .input_20_bits_dataOffset  (selectExecuteReq_20_bits_dataOffset),
    .input_21_ready            (_readCrossBar_input_21_ready),
    .input_21_valid            (readCrossBar_input_21_valid),
    .input_21_bits_vs          (selectExecuteReq_21_bits_vs),
    .input_21_bits_offset      (selectExecuteReq_21_bits_offset),
    .input_21_bits_readLane    (selectExecuteReq_21_bits_readLane),
    .input_21_bits_dataOffset  (selectExecuteReq_21_bits_dataOffset),
    .input_22_ready            (_readCrossBar_input_22_ready),
    .input_22_valid            (readCrossBar_input_22_valid),
    .input_22_bits_vs          (selectExecuteReq_22_bits_vs),
    .input_22_bits_offset      (selectExecuteReq_22_bits_offset),
    .input_22_bits_readLane    (selectExecuteReq_22_bits_readLane),
    .input_22_bits_dataOffset  (selectExecuteReq_22_bits_dataOffset),
    .input_23_ready            (_readCrossBar_input_23_ready),
    .input_23_valid            (readCrossBar_input_23_valid),
    .input_23_bits_vs          (selectExecuteReq_23_bits_vs),
    .input_23_bits_offset      (selectExecuteReq_23_bits_offset),
    .input_23_bits_readLane    (selectExecuteReq_23_bits_readLane),
    .input_23_bits_dataOffset  (selectExecuteReq_23_bits_dataOffset),
    .input_24_ready            (_readCrossBar_input_24_ready),
    .input_24_valid            (readCrossBar_input_24_valid),
    .input_24_bits_vs          (selectExecuteReq_24_bits_vs),
    .input_24_bits_offset      (selectExecuteReq_24_bits_offset),
    .input_24_bits_readLane    (selectExecuteReq_24_bits_readLane),
    .input_24_bits_dataOffset  (selectExecuteReq_24_bits_dataOffset),
    .input_25_ready            (_readCrossBar_input_25_ready),
    .input_25_valid            (readCrossBar_input_25_valid),
    .input_25_bits_vs          (selectExecuteReq_25_bits_vs),
    .input_25_bits_offset      (selectExecuteReq_25_bits_offset),
    .input_25_bits_readLane    (selectExecuteReq_25_bits_readLane),
    .input_25_bits_dataOffset  (selectExecuteReq_25_bits_dataOffset),
    .input_26_ready            (_readCrossBar_input_26_ready),
    .input_26_valid            (readCrossBar_input_26_valid),
    .input_26_bits_vs          (selectExecuteReq_26_bits_vs),
    .input_26_bits_offset      (selectExecuteReq_26_bits_offset),
    .input_26_bits_readLane    (selectExecuteReq_26_bits_readLane),
    .input_26_bits_dataOffset  (selectExecuteReq_26_bits_dataOffset),
    .input_27_ready            (_readCrossBar_input_27_ready),
    .input_27_valid            (readCrossBar_input_27_valid),
    .input_27_bits_vs          (selectExecuteReq_27_bits_vs),
    .input_27_bits_offset      (selectExecuteReq_27_bits_offset),
    .input_27_bits_readLane    (selectExecuteReq_27_bits_readLane),
    .input_27_bits_dataOffset  (selectExecuteReq_27_bits_dataOffset),
    .input_28_ready            (_readCrossBar_input_28_ready),
    .input_28_valid            (readCrossBar_input_28_valid),
    .input_28_bits_vs          (selectExecuteReq_28_bits_vs),
    .input_28_bits_offset      (selectExecuteReq_28_bits_offset),
    .input_28_bits_readLane    (selectExecuteReq_28_bits_readLane),
    .input_28_bits_dataOffset  (selectExecuteReq_28_bits_dataOffset),
    .input_29_ready            (_readCrossBar_input_29_ready),
    .input_29_valid            (readCrossBar_input_29_valid),
    .input_29_bits_vs          (selectExecuteReq_29_bits_vs),
    .input_29_bits_offset      (selectExecuteReq_29_bits_offset),
    .input_29_bits_readLane    (selectExecuteReq_29_bits_readLane),
    .input_29_bits_dataOffset  (selectExecuteReq_29_bits_dataOffset),
    .input_30_ready            (_readCrossBar_input_30_ready),
    .input_30_valid            (readCrossBar_input_30_valid),
    .input_30_bits_vs          (selectExecuteReq_30_bits_vs),
    .input_30_bits_offset      (selectExecuteReq_30_bits_offset),
    .input_30_bits_readLane    (selectExecuteReq_30_bits_readLane),
    .input_30_bits_dataOffset  (selectExecuteReq_30_bits_dataOffset),
    .input_31_ready            (_readCrossBar_input_31_ready),
    .input_31_valid            (readCrossBar_input_31_valid),
    .input_31_bits_vs          (selectExecuteReq_31_bits_vs),
    .input_31_bits_offset      (selectExecuteReq_31_bits_offset),
    .input_31_bits_readLane    (selectExecuteReq_31_bits_readLane),
    .input_31_bits_dataOffset  (selectExecuteReq_31_bits_dataOffset),
    .output_0_ready            (readChannel_0_ready_0 & readMessageQueue_enq_ready),
    .output_0_valid            (_readCrossBar_output_0_valid),
    .output_0_bits_vs          (_readCrossBar_output_0_bits_vs),
    .output_0_bits_offset      (_readCrossBar_output_0_bits_offset),
    .output_0_bits_writeIndex  (_readCrossBar_output_0_bits_writeIndex),
    .output_0_bits_dataOffset  (readMessageQueue_enq_bits_dataOffset),
    .output_1_ready            (readChannel_1_ready_0 & readMessageQueue_1_enq_ready),
    .output_1_valid            (_readCrossBar_output_1_valid),
    .output_1_bits_vs          (_readCrossBar_output_1_bits_vs),
    .output_1_bits_offset      (_readCrossBar_output_1_bits_offset),
    .output_1_bits_writeIndex  (_readCrossBar_output_1_bits_writeIndex),
    .output_1_bits_dataOffset  (readMessageQueue_1_enq_bits_dataOffset),
    .output_2_ready            (readChannel_2_ready_0 & readMessageQueue_2_enq_ready),
    .output_2_valid            (_readCrossBar_output_2_valid),
    .output_2_bits_vs          (_readCrossBar_output_2_bits_vs),
    .output_2_bits_offset      (_readCrossBar_output_2_bits_offset),
    .output_2_bits_writeIndex  (_readCrossBar_output_2_bits_writeIndex),
    .output_2_bits_dataOffset  (readMessageQueue_2_enq_bits_dataOffset),
    .output_3_ready            (readChannel_3_ready_0 & readMessageQueue_3_enq_ready),
    .output_3_valid            (_readCrossBar_output_3_valid),
    .output_3_bits_vs          (_readCrossBar_output_3_bits_vs),
    .output_3_bits_offset      (_readCrossBar_output_3_bits_offset),
    .output_3_bits_writeIndex  (_readCrossBar_output_3_bits_writeIndex),
    .output_3_bits_dataOffset  (readMessageQueue_3_enq_bits_dataOffset),
    .output_4_ready            (readChannel_4_ready_0 & readMessageQueue_4_enq_ready),
    .output_4_valid            (_readCrossBar_output_4_valid),
    .output_4_bits_vs          (_readCrossBar_output_4_bits_vs),
    .output_4_bits_offset      (_readCrossBar_output_4_bits_offset),
    .output_4_bits_writeIndex  (_readCrossBar_output_4_bits_writeIndex),
    .output_4_bits_dataOffset  (readMessageQueue_4_enq_bits_dataOffset),
    .output_5_ready            (readChannel_5_ready_0 & readMessageQueue_5_enq_ready),
    .output_5_valid            (_readCrossBar_output_5_valid),
    .output_5_bits_vs          (_readCrossBar_output_5_bits_vs),
    .output_5_bits_offset      (_readCrossBar_output_5_bits_offset),
    .output_5_bits_writeIndex  (_readCrossBar_output_5_bits_writeIndex),
    .output_5_bits_dataOffset  (readMessageQueue_5_enq_bits_dataOffset),
    .output_6_ready            (readChannel_6_ready_0 & readMessageQueue_6_enq_ready),
    .output_6_valid            (_readCrossBar_output_6_valid),
    .output_6_bits_vs          (_readCrossBar_output_6_bits_vs),
    .output_6_bits_offset      (_readCrossBar_output_6_bits_offset),
    .output_6_bits_writeIndex  (_readCrossBar_output_6_bits_writeIndex),
    .output_6_bits_dataOffset  (readMessageQueue_6_enq_bits_dataOffset),
    .output_7_ready            (readChannel_7_ready_0 & readMessageQueue_7_enq_ready),
    .output_7_valid            (_readCrossBar_output_7_valid),
    .output_7_bits_vs          (_readCrossBar_output_7_bits_vs),
    .output_7_bits_offset      (_readCrossBar_output_7_bits_offset),
    .output_7_bits_writeIndex  (_readCrossBar_output_7_bits_writeIndex),
    .output_7_bits_dataOffset  (readMessageQueue_7_enq_bits_dataOffset),
    .output_8_ready            (readChannel_8_ready_0 & readMessageQueue_8_enq_ready),
    .output_8_valid            (_readCrossBar_output_8_valid),
    .output_8_bits_vs          (_readCrossBar_output_8_bits_vs),
    .output_8_bits_offset      (_readCrossBar_output_8_bits_offset),
    .output_8_bits_writeIndex  (_readCrossBar_output_8_bits_writeIndex),
    .output_8_bits_dataOffset  (readMessageQueue_8_enq_bits_dataOffset),
    .output_9_ready            (readChannel_9_ready_0 & readMessageQueue_9_enq_ready),
    .output_9_valid            (_readCrossBar_output_9_valid),
    .output_9_bits_vs          (_readCrossBar_output_9_bits_vs),
    .output_9_bits_offset      (_readCrossBar_output_9_bits_offset),
    .output_9_bits_writeIndex  (_readCrossBar_output_9_bits_writeIndex),
    .output_9_bits_dataOffset  (readMessageQueue_9_enq_bits_dataOffset),
    .output_10_ready           (readChannel_10_ready_0 & readMessageQueue_10_enq_ready),
    .output_10_valid           (_readCrossBar_output_10_valid),
    .output_10_bits_vs         (_readCrossBar_output_10_bits_vs),
    .output_10_bits_offset     (_readCrossBar_output_10_bits_offset),
    .output_10_bits_writeIndex (_readCrossBar_output_10_bits_writeIndex),
    .output_10_bits_dataOffset (readMessageQueue_10_enq_bits_dataOffset),
    .output_11_ready           (readChannel_11_ready_0 & readMessageQueue_11_enq_ready),
    .output_11_valid           (_readCrossBar_output_11_valid),
    .output_11_bits_vs         (_readCrossBar_output_11_bits_vs),
    .output_11_bits_offset     (_readCrossBar_output_11_bits_offset),
    .output_11_bits_writeIndex (_readCrossBar_output_11_bits_writeIndex),
    .output_11_bits_dataOffset (readMessageQueue_11_enq_bits_dataOffset),
    .output_12_ready           (readChannel_12_ready_0 & readMessageQueue_12_enq_ready),
    .output_12_valid           (_readCrossBar_output_12_valid),
    .output_12_bits_vs         (_readCrossBar_output_12_bits_vs),
    .output_12_bits_offset     (_readCrossBar_output_12_bits_offset),
    .output_12_bits_writeIndex (_readCrossBar_output_12_bits_writeIndex),
    .output_12_bits_dataOffset (readMessageQueue_12_enq_bits_dataOffset),
    .output_13_ready           (readChannel_13_ready_0 & readMessageQueue_13_enq_ready),
    .output_13_valid           (_readCrossBar_output_13_valid),
    .output_13_bits_vs         (_readCrossBar_output_13_bits_vs),
    .output_13_bits_offset     (_readCrossBar_output_13_bits_offset),
    .output_13_bits_writeIndex (_readCrossBar_output_13_bits_writeIndex),
    .output_13_bits_dataOffset (readMessageQueue_13_enq_bits_dataOffset),
    .output_14_ready           (readChannel_14_ready_0 & readMessageQueue_14_enq_ready),
    .output_14_valid           (_readCrossBar_output_14_valid),
    .output_14_bits_vs         (_readCrossBar_output_14_bits_vs),
    .output_14_bits_offset     (_readCrossBar_output_14_bits_offset),
    .output_14_bits_writeIndex (_readCrossBar_output_14_bits_writeIndex),
    .output_14_bits_dataOffset (readMessageQueue_14_enq_bits_dataOffset),
    .output_15_ready           (readChannel_15_ready_0 & readMessageQueue_15_enq_ready),
    .output_15_valid           (_readCrossBar_output_15_valid),
    .output_15_bits_vs         (_readCrossBar_output_15_bits_vs),
    .output_15_bits_offset     (_readCrossBar_output_15_bits_offset),
    .output_15_bits_writeIndex (_readCrossBar_output_15_bits_writeIndex),
    .output_15_bits_dataOffset (readMessageQueue_15_enq_bits_dataOffset),
    .output_16_ready           (readChannel_16_ready_0 & readMessageQueue_16_enq_ready),
    .output_16_valid           (_readCrossBar_output_16_valid),
    .output_16_bits_vs         (_readCrossBar_output_16_bits_vs),
    .output_16_bits_offset     (_readCrossBar_output_16_bits_offset),
    .output_16_bits_writeIndex (_readCrossBar_output_16_bits_writeIndex),
    .output_16_bits_dataOffset (readMessageQueue_16_enq_bits_dataOffset),
    .output_17_ready           (readChannel_17_ready_0 & readMessageQueue_17_enq_ready),
    .output_17_valid           (_readCrossBar_output_17_valid),
    .output_17_bits_vs         (_readCrossBar_output_17_bits_vs),
    .output_17_bits_offset     (_readCrossBar_output_17_bits_offset),
    .output_17_bits_writeIndex (_readCrossBar_output_17_bits_writeIndex),
    .output_17_bits_dataOffset (readMessageQueue_17_enq_bits_dataOffset),
    .output_18_ready           (readChannel_18_ready_0 & readMessageQueue_18_enq_ready),
    .output_18_valid           (_readCrossBar_output_18_valid),
    .output_18_bits_vs         (_readCrossBar_output_18_bits_vs),
    .output_18_bits_offset     (_readCrossBar_output_18_bits_offset),
    .output_18_bits_writeIndex (_readCrossBar_output_18_bits_writeIndex),
    .output_18_bits_dataOffset (readMessageQueue_18_enq_bits_dataOffset),
    .output_19_ready           (readChannel_19_ready_0 & readMessageQueue_19_enq_ready),
    .output_19_valid           (_readCrossBar_output_19_valid),
    .output_19_bits_vs         (_readCrossBar_output_19_bits_vs),
    .output_19_bits_offset     (_readCrossBar_output_19_bits_offset),
    .output_19_bits_writeIndex (_readCrossBar_output_19_bits_writeIndex),
    .output_19_bits_dataOffset (readMessageQueue_19_enq_bits_dataOffset),
    .output_20_ready           (readChannel_20_ready_0 & readMessageQueue_20_enq_ready),
    .output_20_valid           (_readCrossBar_output_20_valid),
    .output_20_bits_vs         (_readCrossBar_output_20_bits_vs),
    .output_20_bits_offset     (_readCrossBar_output_20_bits_offset),
    .output_20_bits_writeIndex (_readCrossBar_output_20_bits_writeIndex),
    .output_20_bits_dataOffset (readMessageQueue_20_enq_bits_dataOffset),
    .output_21_ready           (readChannel_21_ready_0 & readMessageQueue_21_enq_ready),
    .output_21_valid           (_readCrossBar_output_21_valid),
    .output_21_bits_vs         (_readCrossBar_output_21_bits_vs),
    .output_21_bits_offset     (_readCrossBar_output_21_bits_offset),
    .output_21_bits_writeIndex (_readCrossBar_output_21_bits_writeIndex),
    .output_21_bits_dataOffset (readMessageQueue_21_enq_bits_dataOffset),
    .output_22_ready           (readChannel_22_ready_0 & readMessageQueue_22_enq_ready),
    .output_22_valid           (_readCrossBar_output_22_valid),
    .output_22_bits_vs         (_readCrossBar_output_22_bits_vs),
    .output_22_bits_offset     (_readCrossBar_output_22_bits_offset),
    .output_22_bits_writeIndex (_readCrossBar_output_22_bits_writeIndex),
    .output_22_bits_dataOffset (readMessageQueue_22_enq_bits_dataOffset),
    .output_23_ready           (readChannel_23_ready_0 & readMessageQueue_23_enq_ready),
    .output_23_valid           (_readCrossBar_output_23_valid),
    .output_23_bits_vs         (_readCrossBar_output_23_bits_vs),
    .output_23_bits_offset     (_readCrossBar_output_23_bits_offset),
    .output_23_bits_writeIndex (_readCrossBar_output_23_bits_writeIndex),
    .output_23_bits_dataOffset (readMessageQueue_23_enq_bits_dataOffset),
    .output_24_ready           (readChannel_24_ready_0 & readMessageQueue_24_enq_ready),
    .output_24_valid           (_readCrossBar_output_24_valid),
    .output_24_bits_vs         (_readCrossBar_output_24_bits_vs),
    .output_24_bits_offset     (_readCrossBar_output_24_bits_offset),
    .output_24_bits_writeIndex (_readCrossBar_output_24_bits_writeIndex),
    .output_24_bits_dataOffset (readMessageQueue_24_enq_bits_dataOffset),
    .output_25_ready           (readChannel_25_ready_0 & readMessageQueue_25_enq_ready),
    .output_25_valid           (_readCrossBar_output_25_valid),
    .output_25_bits_vs         (_readCrossBar_output_25_bits_vs),
    .output_25_bits_offset     (_readCrossBar_output_25_bits_offset),
    .output_25_bits_writeIndex (_readCrossBar_output_25_bits_writeIndex),
    .output_25_bits_dataOffset (readMessageQueue_25_enq_bits_dataOffset),
    .output_26_ready           (readChannel_26_ready_0 & readMessageQueue_26_enq_ready),
    .output_26_valid           (_readCrossBar_output_26_valid),
    .output_26_bits_vs         (_readCrossBar_output_26_bits_vs),
    .output_26_bits_offset     (_readCrossBar_output_26_bits_offset),
    .output_26_bits_writeIndex (_readCrossBar_output_26_bits_writeIndex),
    .output_26_bits_dataOffset (readMessageQueue_26_enq_bits_dataOffset),
    .output_27_ready           (readChannel_27_ready_0 & readMessageQueue_27_enq_ready),
    .output_27_valid           (_readCrossBar_output_27_valid),
    .output_27_bits_vs         (_readCrossBar_output_27_bits_vs),
    .output_27_bits_offset     (_readCrossBar_output_27_bits_offset),
    .output_27_bits_writeIndex (_readCrossBar_output_27_bits_writeIndex),
    .output_27_bits_dataOffset (readMessageQueue_27_enq_bits_dataOffset),
    .output_28_ready           (readChannel_28_ready_0 & readMessageQueue_28_enq_ready),
    .output_28_valid           (_readCrossBar_output_28_valid),
    .output_28_bits_vs         (_readCrossBar_output_28_bits_vs),
    .output_28_bits_offset     (_readCrossBar_output_28_bits_offset),
    .output_28_bits_writeIndex (_readCrossBar_output_28_bits_writeIndex),
    .output_28_bits_dataOffset (readMessageQueue_28_enq_bits_dataOffset),
    .output_29_ready           (readChannel_29_ready_0 & readMessageQueue_29_enq_ready),
    .output_29_valid           (_readCrossBar_output_29_valid),
    .output_29_bits_vs         (_readCrossBar_output_29_bits_vs),
    .output_29_bits_offset     (_readCrossBar_output_29_bits_offset),
    .output_29_bits_writeIndex (_readCrossBar_output_29_bits_writeIndex),
    .output_29_bits_dataOffset (readMessageQueue_29_enq_bits_dataOffset),
    .output_30_ready           (readChannel_30_ready_0 & readMessageQueue_30_enq_ready),
    .output_30_valid           (_readCrossBar_output_30_valid),
    .output_30_bits_vs         (_readCrossBar_output_30_bits_vs),
    .output_30_bits_offset     (_readCrossBar_output_30_bits_offset),
    .output_30_bits_writeIndex (_readCrossBar_output_30_bits_writeIndex),
    .output_30_bits_dataOffset (readMessageQueue_30_enq_bits_dataOffset),
    .output_31_ready           (readChannel_31_ready_0 & readMessageQueue_31_enq_ready),
    .output_31_valid           (_readCrossBar_output_31_valid),
    .output_31_bits_vs         (_readCrossBar_output_31_bits_vs),
    .output_31_bits_offset     (_readCrossBar_output_31_bits_offset),
    .output_31_bits_writeIndex (_readCrossBar_output_31_bits_writeIndex),
    .output_31_bits_dataOffset (readMessageQueue_31_enq_bits_dataOffset)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(104)
  ) readWaitQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readWaitQueue_enq_ready & readWaitQueue_enq_valid)),
    .pop_req_n    (~(readWaitQueue_deq_ready & ~_readWaitQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (readWaitQueue_dataIn),
    .empty        (_readWaitQueue_fifo_empty),
    .almost_empty (readWaitQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readWaitQueue_almostFull),
    .full         (_readWaitQueue_fifo_full),
    .error        (_readWaitQueue_fifo_error),
    .data_out     (_readWaitQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(1190)
  ) compressUnitResultQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(compressUnitResultQueue_enq_ready & compressUnitResultQueue_enq_valid & ~(_compressUnitResultQueue_fifo_empty & compressUnitResultQueue_deq_ready))),
    .pop_req_n    (~(compressUnitResultQueue_deq_ready & ~_compressUnitResultQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (compressUnitResultQueue_dataIn),
    .empty        (_compressUnitResultQueue_fifo_empty),
    .almost_empty (compressUnitResultQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (compressUnitResultQueue_almostFull),
    .full         (_compressUnitResultQueue_fifo_full),
    .error        (_compressUnitResultQueue_fifo_error),
    .data_out     (_compressUnitResultQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_0_enq_ready & reorderQueueVec_0_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_0_deq_ready & ~_reorderQueueVec_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn),
    .empty        (_reorderQueueVec_fifo_empty),
    .almost_empty (reorderQueueVec_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_0_almostFull),
    .full         (_reorderQueueVec_fifo_full),
    .error        (_reorderQueueVec_fifo_error),
    .data_out     (_reorderQueueVec_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_1_enq_ready & reorderQueueVec_1_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_1_deq_ready & ~_reorderQueueVec_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_1),
    .empty        (_reorderQueueVec_fifo_1_empty),
    .almost_empty (reorderQueueVec_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_1_almostFull),
    .full         (_reorderQueueVec_fifo_1_full),
    .error        (_reorderQueueVec_fifo_1_error),
    .data_out     (_reorderQueueVec_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_2_enq_ready & reorderQueueVec_2_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_2_deq_ready & ~_reorderQueueVec_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_2),
    .empty        (_reorderQueueVec_fifo_2_empty),
    .almost_empty (reorderQueueVec_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_2_almostFull),
    .full         (_reorderQueueVec_fifo_2_full),
    .error        (_reorderQueueVec_fifo_2_error),
    .data_out     (_reorderQueueVec_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_3_enq_ready & reorderQueueVec_3_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_3_deq_ready & ~_reorderQueueVec_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_3),
    .empty        (_reorderQueueVec_fifo_3_empty),
    .almost_empty (reorderQueueVec_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_3_almostFull),
    .full         (_reorderQueueVec_fifo_3_full),
    .error        (_reorderQueueVec_fifo_3_error),
    .data_out     (_reorderQueueVec_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_4_enq_ready & reorderQueueVec_4_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_4_deq_ready & ~_reorderQueueVec_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_4),
    .empty        (_reorderQueueVec_fifo_4_empty),
    .almost_empty (reorderQueueVec_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_4_almostFull),
    .full         (_reorderQueueVec_fifo_4_full),
    .error        (_reorderQueueVec_fifo_4_error),
    .data_out     (_reorderQueueVec_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_5_enq_ready & reorderQueueVec_5_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_5_deq_ready & ~_reorderQueueVec_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_5),
    .empty        (_reorderQueueVec_fifo_5_empty),
    .almost_empty (reorderQueueVec_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_5_almostFull),
    .full         (_reorderQueueVec_fifo_5_full),
    .error        (_reorderQueueVec_fifo_5_error),
    .data_out     (_reorderQueueVec_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_6_enq_ready & reorderQueueVec_6_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_6_deq_ready & ~_reorderQueueVec_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_6),
    .empty        (_reorderQueueVec_fifo_6_empty),
    .almost_empty (reorderQueueVec_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_6_almostFull),
    .full         (_reorderQueueVec_fifo_6_full),
    .error        (_reorderQueueVec_fifo_6_error),
    .data_out     (_reorderQueueVec_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_7_enq_ready & reorderQueueVec_7_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_7_deq_ready & ~_reorderQueueVec_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_7),
    .empty        (_reorderQueueVec_fifo_7_empty),
    .almost_empty (reorderQueueVec_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_7_almostFull),
    .full         (_reorderQueueVec_fifo_7_full),
    .error        (_reorderQueueVec_fifo_7_error),
    .data_out     (_reorderQueueVec_fifo_7_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_8_enq_ready & reorderQueueVec_8_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_8_deq_ready & ~_reorderQueueVec_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_8),
    .empty        (_reorderQueueVec_fifo_8_empty),
    .almost_empty (reorderQueueVec_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_8_almostFull),
    .full         (_reorderQueueVec_fifo_8_full),
    .error        (_reorderQueueVec_fifo_8_error),
    .data_out     (_reorderQueueVec_fifo_8_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_9_enq_ready & reorderQueueVec_9_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_9_deq_ready & ~_reorderQueueVec_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_9),
    .empty        (_reorderQueueVec_fifo_9_empty),
    .almost_empty (reorderQueueVec_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_9_almostFull),
    .full         (_reorderQueueVec_fifo_9_full),
    .error        (_reorderQueueVec_fifo_9_error),
    .data_out     (_reorderQueueVec_fifo_9_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_10_enq_ready & reorderQueueVec_10_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_10_deq_ready & ~_reorderQueueVec_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_10),
    .empty        (_reorderQueueVec_fifo_10_empty),
    .almost_empty (reorderQueueVec_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_10_almostFull),
    .full         (_reorderQueueVec_fifo_10_full),
    .error        (_reorderQueueVec_fifo_10_error),
    .data_out     (_reorderQueueVec_fifo_10_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_11_enq_ready & reorderQueueVec_11_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_11_deq_ready & ~_reorderQueueVec_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_11),
    .empty        (_reorderQueueVec_fifo_11_empty),
    .almost_empty (reorderQueueVec_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_11_almostFull),
    .full         (_reorderQueueVec_fifo_11_full),
    .error        (_reorderQueueVec_fifo_11_error),
    .data_out     (_reorderQueueVec_fifo_11_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_12_enq_ready & reorderQueueVec_12_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_12_deq_ready & ~_reorderQueueVec_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_12),
    .empty        (_reorderQueueVec_fifo_12_empty),
    .almost_empty (reorderQueueVec_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_12_almostFull),
    .full         (_reorderQueueVec_fifo_12_full),
    .error        (_reorderQueueVec_fifo_12_error),
    .data_out     (_reorderQueueVec_fifo_12_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_13_enq_ready & reorderQueueVec_13_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_13_deq_ready & ~_reorderQueueVec_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_13),
    .empty        (_reorderQueueVec_fifo_13_empty),
    .almost_empty (reorderQueueVec_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_13_almostFull),
    .full         (_reorderQueueVec_fifo_13_full),
    .error        (_reorderQueueVec_fifo_13_error),
    .data_out     (_reorderQueueVec_fifo_13_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_14_enq_ready & reorderQueueVec_14_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_14_deq_ready & ~_reorderQueueVec_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_14),
    .empty        (_reorderQueueVec_fifo_14_empty),
    .almost_empty (reorderQueueVec_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_14_almostFull),
    .full         (_reorderQueueVec_fifo_14_full),
    .error        (_reorderQueueVec_fifo_14_error),
    .data_out     (_reorderQueueVec_fifo_14_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_15_enq_ready & reorderQueueVec_15_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_15_deq_ready & ~_reorderQueueVec_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_15),
    .empty        (_reorderQueueVec_fifo_15_empty),
    .almost_empty (reorderQueueVec_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_15_almostFull),
    .full         (_reorderQueueVec_fifo_15_full),
    .error        (_reorderQueueVec_fifo_15_error),
    .data_out     (_reorderQueueVec_fifo_15_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_16 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_16_enq_ready & reorderQueueVec_16_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_16_deq_ready & ~_reorderQueueVec_fifo_16_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_16),
    .empty        (_reorderQueueVec_fifo_16_empty),
    .almost_empty (reorderQueueVec_16_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_16_almostFull),
    .full         (_reorderQueueVec_fifo_16_full),
    .error        (_reorderQueueVec_fifo_16_error),
    .data_out     (_reorderQueueVec_fifo_16_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_17 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_17_enq_ready & reorderQueueVec_17_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_17_deq_ready & ~_reorderQueueVec_fifo_17_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_17),
    .empty        (_reorderQueueVec_fifo_17_empty),
    .almost_empty (reorderQueueVec_17_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_17_almostFull),
    .full         (_reorderQueueVec_fifo_17_full),
    .error        (_reorderQueueVec_fifo_17_error),
    .data_out     (_reorderQueueVec_fifo_17_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_18 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_18_enq_ready & reorderQueueVec_18_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_18_deq_ready & ~_reorderQueueVec_fifo_18_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_18),
    .empty        (_reorderQueueVec_fifo_18_empty),
    .almost_empty (reorderQueueVec_18_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_18_almostFull),
    .full         (_reorderQueueVec_fifo_18_full),
    .error        (_reorderQueueVec_fifo_18_error),
    .data_out     (_reorderQueueVec_fifo_18_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_19 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_19_enq_ready & reorderQueueVec_19_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_19_deq_ready & ~_reorderQueueVec_fifo_19_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_19),
    .empty        (_reorderQueueVec_fifo_19_empty),
    .almost_empty (reorderQueueVec_19_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_19_almostFull),
    .full         (_reorderQueueVec_fifo_19_full),
    .error        (_reorderQueueVec_fifo_19_error),
    .data_out     (_reorderQueueVec_fifo_19_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_20 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_20_enq_ready & reorderQueueVec_20_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_20_deq_ready & ~_reorderQueueVec_fifo_20_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_20),
    .empty        (_reorderQueueVec_fifo_20_empty),
    .almost_empty (reorderQueueVec_20_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_20_almostFull),
    .full         (_reorderQueueVec_fifo_20_full),
    .error        (_reorderQueueVec_fifo_20_error),
    .data_out     (_reorderQueueVec_fifo_20_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_21 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_21_enq_ready & reorderQueueVec_21_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_21_deq_ready & ~_reorderQueueVec_fifo_21_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_21),
    .empty        (_reorderQueueVec_fifo_21_empty),
    .almost_empty (reorderQueueVec_21_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_21_almostFull),
    .full         (_reorderQueueVec_fifo_21_full),
    .error        (_reorderQueueVec_fifo_21_error),
    .data_out     (_reorderQueueVec_fifo_21_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_22 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_22_enq_ready & reorderQueueVec_22_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_22_deq_ready & ~_reorderQueueVec_fifo_22_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_22),
    .empty        (_reorderQueueVec_fifo_22_empty),
    .almost_empty (reorderQueueVec_22_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_22_almostFull),
    .full         (_reorderQueueVec_fifo_22_full),
    .error        (_reorderQueueVec_fifo_22_error),
    .data_out     (_reorderQueueVec_fifo_22_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_23 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_23_enq_ready & reorderQueueVec_23_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_23_deq_ready & ~_reorderQueueVec_fifo_23_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_23),
    .empty        (_reorderQueueVec_fifo_23_empty),
    .almost_empty (reorderQueueVec_23_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_23_almostFull),
    .full         (_reorderQueueVec_fifo_23_full),
    .error        (_reorderQueueVec_fifo_23_error),
    .data_out     (_reorderQueueVec_fifo_23_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_24 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_24_enq_ready & reorderQueueVec_24_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_24_deq_ready & ~_reorderQueueVec_fifo_24_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_24),
    .empty        (_reorderQueueVec_fifo_24_empty),
    .almost_empty (reorderQueueVec_24_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_24_almostFull),
    .full         (_reorderQueueVec_fifo_24_full),
    .error        (_reorderQueueVec_fifo_24_error),
    .data_out     (_reorderQueueVec_fifo_24_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_25 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_25_enq_ready & reorderQueueVec_25_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_25_deq_ready & ~_reorderQueueVec_fifo_25_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_25),
    .empty        (_reorderQueueVec_fifo_25_empty),
    .almost_empty (reorderQueueVec_25_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_25_almostFull),
    .full         (_reorderQueueVec_fifo_25_full),
    .error        (_reorderQueueVec_fifo_25_error),
    .data_out     (_reorderQueueVec_fifo_25_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_26 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_26_enq_ready & reorderQueueVec_26_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_26_deq_ready & ~_reorderQueueVec_fifo_26_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_26),
    .empty        (_reorderQueueVec_fifo_26_empty),
    .almost_empty (reorderQueueVec_26_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_26_almostFull),
    .full         (_reorderQueueVec_fifo_26_full),
    .error        (_reorderQueueVec_fifo_26_error),
    .data_out     (_reorderQueueVec_fifo_26_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_27 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_27_enq_ready & reorderQueueVec_27_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_27_deq_ready & ~_reorderQueueVec_fifo_27_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_27),
    .empty        (_reorderQueueVec_fifo_27_empty),
    .almost_empty (reorderQueueVec_27_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_27_almostFull),
    .full         (_reorderQueueVec_fifo_27_full),
    .error        (_reorderQueueVec_fifo_27_error),
    .data_out     (_reorderQueueVec_fifo_27_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_28 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_28_enq_ready & reorderQueueVec_28_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_28_deq_ready & ~_reorderQueueVec_fifo_28_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_28),
    .empty        (_reorderQueueVec_fifo_28_empty),
    .almost_empty (reorderQueueVec_28_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_28_almostFull),
    .full         (_reorderQueueVec_fifo_28_full),
    .error        (_reorderQueueVec_fifo_28_error),
    .data_out     (_reorderQueueVec_fifo_28_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_29 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_29_enq_ready & reorderQueueVec_29_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_29_deq_ready & ~_reorderQueueVec_fifo_29_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_29),
    .empty        (_reorderQueueVec_fifo_29_empty),
    .almost_empty (reorderQueueVec_29_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_29_almostFull),
    .full         (_reorderQueueVec_fifo_29_full),
    .error        (_reorderQueueVec_fifo_29_error),
    .data_out     (_reorderQueueVec_fifo_29_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_30 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_30_enq_ready & reorderQueueVec_30_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_30_deq_ready & ~_reorderQueueVec_fifo_30_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_30),
    .empty        (_reorderQueueVec_fifo_30_empty),
    .almost_empty (reorderQueueVec_30_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_30_almostFull),
    .full         (_reorderQueueVec_fifo_30_full),
    .error        (_reorderQueueVec_fifo_30_error),
    .data_out     (_reorderQueueVec_fifo_30_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(64)
  ) reorderQueueVec_fifo_31 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_31_enq_ready & reorderQueueVec_31_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_31_deq_ready & ~_reorderQueueVec_fifo_31_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_31),
    .empty        (_reorderQueueVec_fifo_31_empty),
    .almost_empty (reorderQueueVec_31_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_31_almostFull),
    .full         (_reorderQueueVec_fifo_31_full),
    .error        (_reorderQueueVec_fifo_31_error),
    .data_out     (_reorderQueueVec_fifo_31_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_enq_ready & readMessageQueue_enq_valid)),
    .pop_req_n    (~(readMessageQueue_deq_ready & ~_readMessageQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn),
    .empty        (_readMessageQueue_fifo_empty),
    .almost_empty (readMessageQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_almostFull),
    .full         (_readMessageQueue_fifo_full),
    .error        (_readMessageQueue_fifo_error),
    .data_out     (_readMessageQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_1_enq_ready & readMessageQueue_1_enq_valid)),
    .pop_req_n    (~(readMessageQueue_1_deq_ready & ~_readMessageQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_1),
    .empty        (_readMessageQueue_fifo_1_empty),
    .almost_empty (readMessageQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_1_almostFull),
    .full         (_readMessageQueue_fifo_1_full),
    .error        (_readMessageQueue_fifo_1_error),
    .data_out     (_readMessageQueue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_2_enq_ready & readMessageQueue_2_enq_valid)),
    .pop_req_n    (~(readMessageQueue_2_deq_ready & ~_readMessageQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_2),
    .empty        (_readMessageQueue_fifo_2_empty),
    .almost_empty (readMessageQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_2_almostFull),
    .full         (_readMessageQueue_fifo_2_full),
    .error        (_readMessageQueue_fifo_2_error),
    .data_out     (_readMessageQueue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_3_enq_ready & readMessageQueue_3_enq_valid)),
    .pop_req_n    (~(readMessageQueue_3_deq_ready & ~_readMessageQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_3),
    .empty        (_readMessageQueue_fifo_3_empty),
    .almost_empty (readMessageQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_3_almostFull),
    .full         (_readMessageQueue_fifo_3_full),
    .error        (_readMessageQueue_fifo_3_error),
    .data_out     (_readMessageQueue_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_4_enq_ready & readMessageQueue_4_enq_valid)),
    .pop_req_n    (~(readMessageQueue_4_deq_ready & ~_readMessageQueue_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_4),
    .empty        (_readMessageQueue_fifo_4_empty),
    .almost_empty (readMessageQueue_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_4_almostFull),
    .full         (_readMessageQueue_fifo_4_full),
    .error        (_readMessageQueue_fifo_4_error),
    .data_out     (_readMessageQueue_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_5_enq_ready & readMessageQueue_5_enq_valid)),
    .pop_req_n    (~(readMessageQueue_5_deq_ready & ~_readMessageQueue_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_5),
    .empty        (_readMessageQueue_fifo_5_empty),
    .almost_empty (readMessageQueue_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_5_almostFull),
    .full         (_readMessageQueue_fifo_5_full),
    .error        (_readMessageQueue_fifo_5_error),
    .data_out     (_readMessageQueue_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_6_enq_ready & readMessageQueue_6_enq_valid)),
    .pop_req_n    (~(readMessageQueue_6_deq_ready & ~_readMessageQueue_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_6),
    .empty        (_readMessageQueue_fifo_6_empty),
    .almost_empty (readMessageQueue_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_6_almostFull),
    .full         (_readMessageQueue_fifo_6_full),
    .error        (_readMessageQueue_fifo_6_error),
    .data_out     (_readMessageQueue_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_7_enq_ready & readMessageQueue_7_enq_valid)),
    .pop_req_n    (~(readMessageQueue_7_deq_ready & ~_readMessageQueue_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_7),
    .empty        (_readMessageQueue_fifo_7_empty),
    .almost_empty (readMessageQueue_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_7_almostFull),
    .full         (_readMessageQueue_fifo_7_full),
    .error        (_readMessageQueue_fifo_7_error),
    .data_out     (_readMessageQueue_fifo_7_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_8_enq_ready & readMessageQueue_8_enq_valid)),
    .pop_req_n    (~(readMessageQueue_8_deq_ready & ~_readMessageQueue_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_8),
    .empty        (_readMessageQueue_fifo_8_empty),
    .almost_empty (readMessageQueue_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_8_almostFull),
    .full         (_readMessageQueue_fifo_8_full),
    .error        (_readMessageQueue_fifo_8_error),
    .data_out     (_readMessageQueue_fifo_8_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_9_enq_ready & readMessageQueue_9_enq_valid)),
    .pop_req_n    (~(readMessageQueue_9_deq_ready & ~_readMessageQueue_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_9),
    .empty        (_readMessageQueue_fifo_9_empty),
    .almost_empty (readMessageQueue_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_9_almostFull),
    .full         (_readMessageQueue_fifo_9_full),
    .error        (_readMessageQueue_fifo_9_error),
    .data_out     (_readMessageQueue_fifo_9_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_10_enq_ready & readMessageQueue_10_enq_valid)),
    .pop_req_n    (~(readMessageQueue_10_deq_ready & ~_readMessageQueue_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_10),
    .empty        (_readMessageQueue_fifo_10_empty),
    .almost_empty (readMessageQueue_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_10_almostFull),
    .full         (_readMessageQueue_fifo_10_full),
    .error        (_readMessageQueue_fifo_10_error),
    .data_out     (_readMessageQueue_fifo_10_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_11_enq_ready & readMessageQueue_11_enq_valid)),
    .pop_req_n    (~(readMessageQueue_11_deq_ready & ~_readMessageQueue_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_11),
    .empty        (_readMessageQueue_fifo_11_empty),
    .almost_empty (readMessageQueue_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_11_almostFull),
    .full         (_readMessageQueue_fifo_11_full),
    .error        (_readMessageQueue_fifo_11_error),
    .data_out     (_readMessageQueue_fifo_11_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_12_enq_ready & readMessageQueue_12_enq_valid)),
    .pop_req_n    (~(readMessageQueue_12_deq_ready & ~_readMessageQueue_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_12),
    .empty        (_readMessageQueue_fifo_12_empty),
    .almost_empty (readMessageQueue_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_12_almostFull),
    .full         (_readMessageQueue_fifo_12_full),
    .error        (_readMessageQueue_fifo_12_error),
    .data_out     (_readMessageQueue_fifo_12_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_13_enq_ready & readMessageQueue_13_enq_valid)),
    .pop_req_n    (~(readMessageQueue_13_deq_ready & ~_readMessageQueue_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_13),
    .empty        (_readMessageQueue_fifo_13_empty),
    .almost_empty (readMessageQueue_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_13_almostFull),
    .full         (_readMessageQueue_fifo_13_full),
    .error        (_readMessageQueue_fifo_13_error),
    .data_out     (_readMessageQueue_fifo_13_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_14_enq_ready & readMessageQueue_14_enq_valid)),
    .pop_req_n    (~(readMessageQueue_14_deq_ready & ~_readMessageQueue_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_14),
    .empty        (_readMessageQueue_fifo_14_empty),
    .almost_empty (readMessageQueue_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_14_almostFull),
    .full         (_readMessageQueue_fifo_14_full),
    .error        (_readMessageQueue_fifo_14_error),
    .data_out     (_readMessageQueue_fifo_14_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_15_enq_ready & readMessageQueue_15_enq_valid)),
    .pop_req_n    (~(readMessageQueue_15_deq_ready & ~_readMessageQueue_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_15),
    .empty        (_readMessageQueue_fifo_15_empty),
    .almost_empty (readMessageQueue_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_15_almostFull),
    .full         (_readMessageQueue_fifo_15_full),
    .error        (_readMessageQueue_fifo_15_error),
    .data_out     (_readMessageQueue_fifo_15_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_16 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_16_enq_ready & readMessageQueue_16_enq_valid)),
    .pop_req_n    (~(readMessageQueue_16_deq_ready & ~_readMessageQueue_fifo_16_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_16),
    .empty        (_readMessageQueue_fifo_16_empty),
    .almost_empty (readMessageQueue_16_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_16_almostFull),
    .full         (_readMessageQueue_fifo_16_full),
    .error        (_readMessageQueue_fifo_16_error),
    .data_out     (_readMessageQueue_fifo_16_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_17 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_17_enq_ready & readMessageQueue_17_enq_valid)),
    .pop_req_n    (~(readMessageQueue_17_deq_ready & ~_readMessageQueue_fifo_17_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_17),
    .empty        (_readMessageQueue_fifo_17_empty),
    .almost_empty (readMessageQueue_17_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_17_almostFull),
    .full         (_readMessageQueue_fifo_17_full),
    .error        (_readMessageQueue_fifo_17_error),
    .data_out     (_readMessageQueue_fifo_17_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_18 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_18_enq_ready & readMessageQueue_18_enq_valid)),
    .pop_req_n    (~(readMessageQueue_18_deq_ready & ~_readMessageQueue_fifo_18_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_18),
    .empty        (_readMessageQueue_fifo_18_empty),
    .almost_empty (readMessageQueue_18_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_18_almostFull),
    .full         (_readMessageQueue_fifo_18_full),
    .error        (_readMessageQueue_fifo_18_error),
    .data_out     (_readMessageQueue_fifo_18_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_19 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_19_enq_ready & readMessageQueue_19_enq_valid)),
    .pop_req_n    (~(readMessageQueue_19_deq_ready & ~_readMessageQueue_fifo_19_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_19),
    .empty        (_readMessageQueue_fifo_19_empty),
    .almost_empty (readMessageQueue_19_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_19_almostFull),
    .full         (_readMessageQueue_fifo_19_full),
    .error        (_readMessageQueue_fifo_19_error),
    .data_out     (_readMessageQueue_fifo_19_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_20 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_20_enq_ready & readMessageQueue_20_enq_valid)),
    .pop_req_n    (~(readMessageQueue_20_deq_ready & ~_readMessageQueue_fifo_20_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_20),
    .empty        (_readMessageQueue_fifo_20_empty),
    .almost_empty (readMessageQueue_20_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_20_almostFull),
    .full         (_readMessageQueue_fifo_20_full),
    .error        (_readMessageQueue_fifo_20_error),
    .data_out     (_readMessageQueue_fifo_20_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_21 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_21_enq_ready & readMessageQueue_21_enq_valid)),
    .pop_req_n    (~(readMessageQueue_21_deq_ready & ~_readMessageQueue_fifo_21_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_21),
    .empty        (_readMessageQueue_fifo_21_empty),
    .almost_empty (readMessageQueue_21_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_21_almostFull),
    .full         (_readMessageQueue_fifo_21_full),
    .error        (_readMessageQueue_fifo_21_error),
    .data_out     (_readMessageQueue_fifo_21_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_22 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_22_enq_ready & readMessageQueue_22_enq_valid)),
    .pop_req_n    (~(readMessageQueue_22_deq_ready & ~_readMessageQueue_fifo_22_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_22),
    .empty        (_readMessageQueue_fifo_22_empty),
    .almost_empty (readMessageQueue_22_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_22_almostFull),
    .full         (_readMessageQueue_fifo_22_full),
    .error        (_readMessageQueue_fifo_22_error),
    .data_out     (_readMessageQueue_fifo_22_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_23 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_23_enq_ready & readMessageQueue_23_enq_valid)),
    .pop_req_n    (~(readMessageQueue_23_deq_ready & ~_readMessageQueue_fifo_23_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_23),
    .empty        (_readMessageQueue_fifo_23_empty),
    .almost_empty (readMessageQueue_23_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_23_almostFull),
    .full         (_readMessageQueue_fifo_23_full),
    .error        (_readMessageQueue_fifo_23_error),
    .data_out     (_readMessageQueue_fifo_23_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_24 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_24_enq_ready & readMessageQueue_24_enq_valid)),
    .pop_req_n    (~(readMessageQueue_24_deq_ready & ~_readMessageQueue_fifo_24_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_24),
    .empty        (_readMessageQueue_fifo_24_empty),
    .almost_empty (readMessageQueue_24_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_24_almostFull),
    .full         (_readMessageQueue_fifo_24_full),
    .error        (_readMessageQueue_fifo_24_error),
    .data_out     (_readMessageQueue_fifo_24_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_25 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_25_enq_ready & readMessageQueue_25_enq_valid)),
    .pop_req_n    (~(readMessageQueue_25_deq_ready & ~_readMessageQueue_fifo_25_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_25),
    .empty        (_readMessageQueue_fifo_25_empty),
    .almost_empty (readMessageQueue_25_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_25_almostFull),
    .full         (_readMessageQueue_fifo_25_full),
    .error        (_readMessageQueue_fifo_25_error),
    .data_out     (_readMessageQueue_fifo_25_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_26 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_26_enq_ready & readMessageQueue_26_enq_valid)),
    .pop_req_n    (~(readMessageQueue_26_deq_ready & ~_readMessageQueue_fifo_26_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_26),
    .empty        (_readMessageQueue_fifo_26_empty),
    .almost_empty (readMessageQueue_26_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_26_almostFull),
    .full         (_readMessageQueue_fifo_26_full),
    .error        (_readMessageQueue_fifo_26_error),
    .data_out     (_readMessageQueue_fifo_26_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_27 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_27_enq_ready & readMessageQueue_27_enq_valid)),
    .pop_req_n    (~(readMessageQueue_27_deq_ready & ~_readMessageQueue_fifo_27_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_27),
    .empty        (_readMessageQueue_fifo_27_empty),
    .almost_empty (readMessageQueue_27_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_27_almostFull),
    .full         (_readMessageQueue_fifo_27_full),
    .error        (_readMessageQueue_fifo_27_error),
    .data_out     (_readMessageQueue_fifo_27_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_28 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_28_enq_ready & readMessageQueue_28_enq_valid)),
    .pop_req_n    (~(readMessageQueue_28_deq_ready & ~_readMessageQueue_fifo_28_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_28),
    .empty        (_readMessageQueue_fifo_28_empty),
    .almost_empty (readMessageQueue_28_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_28_almostFull),
    .full         (_readMessageQueue_fifo_28_full),
    .error        (_readMessageQueue_fifo_28_error),
    .data_out     (_readMessageQueue_fifo_28_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_29 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_29_enq_ready & readMessageQueue_29_enq_valid)),
    .pop_req_n    (~(readMessageQueue_29_deq_ready & ~_readMessageQueue_fifo_29_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_29),
    .empty        (_readMessageQueue_fifo_29_empty),
    .almost_empty (readMessageQueue_29_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_29_almostFull),
    .full         (_readMessageQueue_fifo_29_full),
    .error        (_readMessageQueue_fifo_29_error),
    .data_out     (_readMessageQueue_fifo_29_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_30 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_30_enq_ready & readMessageQueue_30_enq_valid)),
    .pop_req_n    (~(readMessageQueue_30_deq_ready & ~_readMessageQueue_fifo_30_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_30),
    .empty        (_readMessageQueue_fifo_30_empty),
    .almost_empty (readMessageQueue_30_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_30_almostFull),
    .full         (_readMessageQueue_fifo_30_full),
    .error        (_readMessageQueue_fifo_30_error),
    .data_out     (_readMessageQueue_fifo_30_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(34)
  ) readMessageQueue_fifo_31 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_31_enq_ready & readMessageQueue_31_enq_valid)),
    .pop_req_n    (~(readMessageQueue_31_deq_ready & ~_readMessageQueue_fifo_31_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_31),
    .empty        (_readMessageQueue_fifo_31_empty),
    .almost_empty (readMessageQueue_31_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_31_almostFull),
    .full         (_readMessageQueue_fifo_31_full),
    .error        (_readMessageQueue_fifo_31_error),
    .data_out     (_readMessageQueue_fifo_31_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_enq_ready & readData_readDataQueue_enq_valid & ~(_readData_readDataQueue_fifo_empty & readData_readDataQueue_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_deq_ready & ~_readData_readDataQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_enq_bits),
    .empty        (_readData_readDataQueue_fifo_empty),
    .almost_empty (readData_readDataQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_almostFull),
    .full         (_readData_readDataQueue_fifo_full),
    .error        (_readData_readDataQueue_fifo_error),
    .data_out     (_readData_readDataQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_1_enq_ready & readData_readDataQueue_1_enq_valid & ~(_readData_readDataQueue_fifo_1_empty & readData_readDataQueue_1_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_1_deq_ready & ~_readData_readDataQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_1_enq_bits),
    .empty        (_readData_readDataQueue_fifo_1_empty),
    .almost_empty (readData_readDataQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_1_almostFull),
    .full         (_readData_readDataQueue_fifo_1_full),
    .error        (_readData_readDataQueue_fifo_1_error),
    .data_out     (_readData_readDataQueue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_2_enq_ready & readData_readDataQueue_2_enq_valid & ~(_readData_readDataQueue_fifo_2_empty & readData_readDataQueue_2_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_2_deq_ready & ~_readData_readDataQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_2_enq_bits),
    .empty        (_readData_readDataQueue_fifo_2_empty),
    .almost_empty (readData_readDataQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_2_almostFull),
    .full         (_readData_readDataQueue_fifo_2_full),
    .error        (_readData_readDataQueue_fifo_2_error),
    .data_out     (_readData_readDataQueue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_3_enq_ready & readData_readDataQueue_3_enq_valid & ~(_readData_readDataQueue_fifo_3_empty & readData_readDataQueue_3_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_3_deq_ready & ~_readData_readDataQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_3_enq_bits),
    .empty        (_readData_readDataQueue_fifo_3_empty),
    .almost_empty (readData_readDataQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_3_almostFull),
    .full         (_readData_readDataQueue_fifo_3_full),
    .error        (_readData_readDataQueue_fifo_3_error),
    .data_out     (_readData_readDataQueue_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_4_enq_ready & readData_readDataQueue_4_enq_valid & ~(_readData_readDataQueue_fifo_4_empty & readData_readDataQueue_4_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_4_deq_ready & ~_readData_readDataQueue_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_4_enq_bits),
    .empty        (_readData_readDataQueue_fifo_4_empty),
    .almost_empty (readData_readDataQueue_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_4_almostFull),
    .full         (_readData_readDataQueue_fifo_4_full),
    .error        (_readData_readDataQueue_fifo_4_error),
    .data_out     (_readData_readDataQueue_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_5_enq_ready & readData_readDataQueue_5_enq_valid & ~(_readData_readDataQueue_fifo_5_empty & readData_readDataQueue_5_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_5_deq_ready & ~_readData_readDataQueue_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_5_enq_bits),
    .empty        (_readData_readDataQueue_fifo_5_empty),
    .almost_empty (readData_readDataQueue_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_5_almostFull),
    .full         (_readData_readDataQueue_fifo_5_full),
    .error        (_readData_readDataQueue_fifo_5_error),
    .data_out     (_readData_readDataQueue_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_6_enq_ready & readData_readDataQueue_6_enq_valid & ~(_readData_readDataQueue_fifo_6_empty & readData_readDataQueue_6_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_6_deq_ready & ~_readData_readDataQueue_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_6_enq_bits),
    .empty        (_readData_readDataQueue_fifo_6_empty),
    .almost_empty (readData_readDataQueue_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_6_almostFull),
    .full         (_readData_readDataQueue_fifo_6_full),
    .error        (_readData_readDataQueue_fifo_6_error),
    .data_out     (_readData_readDataQueue_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_7_enq_ready & readData_readDataQueue_7_enq_valid & ~(_readData_readDataQueue_fifo_7_empty & readData_readDataQueue_7_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_7_deq_ready & ~_readData_readDataQueue_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_7_enq_bits),
    .empty        (_readData_readDataQueue_fifo_7_empty),
    .almost_empty (readData_readDataQueue_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_7_almostFull),
    .full         (_readData_readDataQueue_fifo_7_full),
    .error        (_readData_readDataQueue_fifo_7_error),
    .data_out     (_readData_readDataQueue_fifo_7_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_8_enq_ready & readData_readDataQueue_8_enq_valid & ~(_readData_readDataQueue_fifo_8_empty & readData_readDataQueue_8_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_8_deq_ready & ~_readData_readDataQueue_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_8_enq_bits),
    .empty        (_readData_readDataQueue_fifo_8_empty),
    .almost_empty (readData_readDataQueue_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_8_almostFull),
    .full         (_readData_readDataQueue_fifo_8_full),
    .error        (_readData_readDataQueue_fifo_8_error),
    .data_out     (_readData_readDataQueue_fifo_8_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_9_enq_ready & readData_readDataQueue_9_enq_valid & ~(_readData_readDataQueue_fifo_9_empty & readData_readDataQueue_9_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_9_deq_ready & ~_readData_readDataQueue_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_9_enq_bits),
    .empty        (_readData_readDataQueue_fifo_9_empty),
    .almost_empty (readData_readDataQueue_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_9_almostFull),
    .full         (_readData_readDataQueue_fifo_9_full),
    .error        (_readData_readDataQueue_fifo_9_error),
    .data_out     (_readData_readDataQueue_fifo_9_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_10_enq_ready & readData_readDataQueue_10_enq_valid & ~(_readData_readDataQueue_fifo_10_empty & readData_readDataQueue_10_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_10_deq_ready & ~_readData_readDataQueue_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_10_enq_bits),
    .empty        (_readData_readDataQueue_fifo_10_empty),
    .almost_empty (readData_readDataQueue_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_10_almostFull),
    .full         (_readData_readDataQueue_fifo_10_full),
    .error        (_readData_readDataQueue_fifo_10_error),
    .data_out     (_readData_readDataQueue_fifo_10_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_11_enq_ready & readData_readDataQueue_11_enq_valid & ~(_readData_readDataQueue_fifo_11_empty & readData_readDataQueue_11_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_11_deq_ready & ~_readData_readDataQueue_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_11_enq_bits),
    .empty        (_readData_readDataQueue_fifo_11_empty),
    .almost_empty (readData_readDataQueue_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_11_almostFull),
    .full         (_readData_readDataQueue_fifo_11_full),
    .error        (_readData_readDataQueue_fifo_11_error),
    .data_out     (_readData_readDataQueue_fifo_11_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_12_enq_ready & readData_readDataQueue_12_enq_valid & ~(_readData_readDataQueue_fifo_12_empty & readData_readDataQueue_12_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_12_deq_ready & ~_readData_readDataQueue_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_12_enq_bits),
    .empty        (_readData_readDataQueue_fifo_12_empty),
    .almost_empty (readData_readDataQueue_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_12_almostFull),
    .full         (_readData_readDataQueue_fifo_12_full),
    .error        (_readData_readDataQueue_fifo_12_error),
    .data_out     (_readData_readDataQueue_fifo_12_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_13_enq_ready & readData_readDataQueue_13_enq_valid & ~(_readData_readDataQueue_fifo_13_empty & readData_readDataQueue_13_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_13_deq_ready & ~_readData_readDataQueue_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_13_enq_bits),
    .empty        (_readData_readDataQueue_fifo_13_empty),
    .almost_empty (readData_readDataQueue_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_13_almostFull),
    .full         (_readData_readDataQueue_fifo_13_full),
    .error        (_readData_readDataQueue_fifo_13_error),
    .data_out     (_readData_readDataQueue_fifo_13_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_14_enq_ready & readData_readDataQueue_14_enq_valid & ~(_readData_readDataQueue_fifo_14_empty & readData_readDataQueue_14_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_14_deq_ready & ~_readData_readDataQueue_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_14_enq_bits),
    .empty        (_readData_readDataQueue_fifo_14_empty),
    .almost_empty (readData_readDataQueue_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_14_almostFull),
    .full         (_readData_readDataQueue_fifo_14_full),
    .error        (_readData_readDataQueue_fifo_14_error),
    .data_out     (_readData_readDataQueue_fifo_14_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_15_enq_ready & readData_readDataQueue_15_enq_valid & ~(_readData_readDataQueue_fifo_15_empty & readData_readDataQueue_15_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_15_deq_ready & ~_readData_readDataQueue_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_15_enq_bits),
    .empty        (_readData_readDataQueue_fifo_15_empty),
    .almost_empty (readData_readDataQueue_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_15_almostFull),
    .full         (_readData_readDataQueue_fifo_15_full),
    .error        (_readData_readDataQueue_fifo_15_error),
    .data_out     (_readData_readDataQueue_fifo_15_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_16 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_16_enq_ready & readData_readDataQueue_16_enq_valid & ~(_readData_readDataQueue_fifo_16_empty & readData_readDataQueue_16_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_16_deq_ready & ~_readData_readDataQueue_fifo_16_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_16_enq_bits),
    .empty        (_readData_readDataQueue_fifo_16_empty),
    .almost_empty (readData_readDataQueue_16_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_16_almostFull),
    .full         (_readData_readDataQueue_fifo_16_full),
    .error        (_readData_readDataQueue_fifo_16_error),
    .data_out     (_readData_readDataQueue_fifo_16_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_17 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_17_enq_ready & readData_readDataQueue_17_enq_valid & ~(_readData_readDataQueue_fifo_17_empty & readData_readDataQueue_17_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_17_deq_ready & ~_readData_readDataQueue_fifo_17_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_17_enq_bits),
    .empty        (_readData_readDataQueue_fifo_17_empty),
    .almost_empty (readData_readDataQueue_17_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_17_almostFull),
    .full         (_readData_readDataQueue_fifo_17_full),
    .error        (_readData_readDataQueue_fifo_17_error),
    .data_out     (_readData_readDataQueue_fifo_17_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_18 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_18_enq_ready & readData_readDataQueue_18_enq_valid & ~(_readData_readDataQueue_fifo_18_empty & readData_readDataQueue_18_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_18_deq_ready & ~_readData_readDataQueue_fifo_18_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_18_enq_bits),
    .empty        (_readData_readDataQueue_fifo_18_empty),
    .almost_empty (readData_readDataQueue_18_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_18_almostFull),
    .full         (_readData_readDataQueue_fifo_18_full),
    .error        (_readData_readDataQueue_fifo_18_error),
    .data_out     (_readData_readDataQueue_fifo_18_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_19 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_19_enq_ready & readData_readDataQueue_19_enq_valid & ~(_readData_readDataQueue_fifo_19_empty & readData_readDataQueue_19_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_19_deq_ready & ~_readData_readDataQueue_fifo_19_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_19_enq_bits),
    .empty        (_readData_readDataQueue_fifo_19_empty),
    .almost_empty (readData_readDataQueue_19_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_19_almostFull),
    .full         (_readData_readDataQueue_fifo_19_full),
    .error        (_readData_readDataQueue_fifo_19_error),
    .data_out     (_readData_readDataQueue_fifo_19_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_20 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_20_enq_ready & readData_readDataQueue_20_enq_valid & ~(_readData_readDataQueue_fifo_20_empty & readData_readDataQueue_20_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_20_deq_ready & ~_readData_readDataQueue_fifo_20_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_20_enq_bits),
    .empty        (_readData_readDataQueue_fifo_20_empty),
    .almost_empty (readData_readDataQueue_20_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_20_almostFull),
    .full         (_readData_readDataQueue_fifo_20_full),
    .error        (_readData_readDataQueue_fifo_20_error),
    .data_out     (_readData_readDataQueue_fifo_20_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_21 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_21_enq_ready & readData_readDataQueue_21_enq_valid & ~(_readData_readDataQueue_fifo_21_empty & readData_readDataQueue_21_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_21_deq_ready & ~_readData_readDataQueue_fifo_21_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_21_enq_bits),
    .empty        (_readData_readDataQueue_fifo_21_empty),
    .almost_empty (readData_readDataQueue_21_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_21_almostFull),
    .full         (_readData_readDataQueue_fifo_21_full),
    .error        (_readData_readDataQueue_fifo_21_error),
    .data_out     (_readData_readDataQueue_fifo_21_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_22 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_22_enq_ready & readData_readDataQueue_22_enq_valid & ~(_readData_readDataQueue_fifo_22_empty & readData_readDataQueue_22_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_22_deq_ready & ~_readData_readDataQueue_fifo_22_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_22_enq_bits),
    .empty        (_readData_readDataQueue_fifo_22_empty),
    .almost_empty (readData_readDataQueue_22_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_22_almostFull),
    .full         (_readData_readDataQueue_fifo_22_full),
    .error        (_readData_readDataQueue_fifo_22_error),
    .data_out     (_readData_readDataQueue_fifo_22_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_23 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_23_enq_ready & readData_readDataQueue_23_enq_valid & ~(_readData_readDataQueue_fifo_23_empty & readData_readDataQueue_23_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_23_deq_ready & ~_readData_readDataQueue_fifo_23_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_23_enq_bits),
    .empty        (_readData_readDataQueue_fifo_23_empty),
    .almost_empty (readData_readDataQueue_23_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_23_almostFull),
    .full         (_readData_readDataQueue_fifo_23_full),
    .error        (_readData_readDataQueue_fifo_23_error),
    .data_out     (_readData_readDataQueue_fifo_23_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_24 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_24_enq_ready & readData_readDataQueue_24_enq_valid & ~(_readData_readDataQueue_fifo_24_empty & readData_readDataQueue_24_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_24_deq_ready & ~_readData_readDataQueue_fifo_24_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_24_enq_bits),
    .empty        (_readData_readDataQueue_fifo_24_empty),
    .almost_empty (readData_readDataQueue_24_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_24_almostFull),
    .full         (_readData_readDataQueue_fifo_24_full),
    .error        (_readData_readDataQueue_fifo_24_error),
    .data_out     (_readData_readDataQueue_fifo_24_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_25 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_25_enq_ready & readData_readDataQueue_25_enq_valid & ~(_readData_readDataQueue_fifo_25_empty & readData_readDataQueue_25_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_25_deq_ready & ~_readData_readDataQueue_fifo_25_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_25_enq_bits),
    .empty        (_readData_readDataQueue_fifo_25_empty),
    .almost_empty (readData_readDataQueue_25_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_25_almostFull),
    .full         (_readData_readDataQueue_fifo_25_full),
    .error        (_readData_readDataQueue_fifo_25_error),
    .data_out     (_readData_readDataQueue_fifo_25_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_26 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_26_enq_ready & readData_readDataQueue_26_enq_valid & ~(_readData_readDataQueue_fifo_26_empty & readData_readDataQueue_26_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_26_deq_ready & ~_readData_readDataQueue_fifo_26_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_26_enq_bits),
    .empty        (_readData_readDataQueue_fifo_26_empty),
    .almost_empty (readData_readDataQueue_26_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_26_almostFull),
    .full         (_readData_readDataQueue_fifo_26_full),
    .error        (_readData_readDataQueue_fifo_26_error),
    .data_out     (_readData_readDataQueue_fifo_26_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_27 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_27_enq_ready & readData_readDataQueue_27_enq_valid & ~(_readData_readDataQueue_fifo_27_empty & readData_readDataQueue_27_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_27_deq_ready & ~_readData_readDataQueue_fifo_27_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_27_enq_bits),
    .empty        (_readData_readDataQueue_fifo_27_empty),
    .almost_empty (readData_readDataQueue_27_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_27_almostFull),
    .full         (_readData_readDataQueue_fifo_27_full),
    .error        (_readData_readDataQueue_fifo_27_error),
    .data_out     (_readData_readDataQueue_fifo_27_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_28 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_28_enq_ready & readData_readDataQueue_28_enq_valid & ~(_readData_readDataQueue_fifo_28_empty & readData_readDataQueue_28_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_28_deq_ready & ~_readData_readDataQueue_fifo_28_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_28_enq_bits),
    .empty        (_readData_readDataQueue_fifo_28_empty),
    .almost_empty (readData_readDataQueue_28_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_28_almostFull),
    .full         (_readData_readDataQueue_fifo_28_full),
    .error        (_readData_readDataQueue_fifo_28_error),
    .data_out     (_readData_readDataQueue_fifo_28_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_29 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_29_enq_ready & readData_readDataQueue_29_enq_valid & ~(_readData_readDataQueue_fifo_29_empty & readData_readDataQueue_29_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_29_deq_ready & ~_readData_readDataQueue_fifo_29_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_29_enq_bits),
    .empty        (_readData_readDataQueue_fifo_29_empty),
    .almost_empty (readData_readDataQueue_29_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_29_almostFull),
    .full         (_readData_readDataQueue_fifo_29_full),
    .error        (_readData_readDataQueue_fifo_29_error),
    .data_out     (_readData_readDataQueue_fifo_29_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_30 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_30_enq_ready & readData_readDataQueue_30_enq_valid & ~(_readData_readDataQueue_fifo_30_empty & readData_readDataQueue_30_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_30_deq_ready & ~_readData_readDataQueue_fifo_30_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_30_enq_bits),
    .empty        (_readData_readDataQueue_fifo_30_empty),
    .almost_empty (readData_readDataQueue_30_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_30_almostFull),
    .full         (_readData_readDataQueue_fifo_30_full),
    .error        (_readData_readDataQueue_fifo_30_error),
    .data_out     (_readData_readDataQueue_fifo_30_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_31 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_31_enq_ready & readData_readDataQueue_31_enq_valid & ~(_readData_readDataQueue_fifo_31_empty & readData_readDataQueue_31_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_31_deq_ready & ~_readData_readDataQueue_fifo_31_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_31_enq_bits),
    .empty        (_readData_readDataQueue_fifo_31_empty),
    .almost_empty (readData_readDataQueue_31_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_31_almostFull),
    .full         (_readData_readDataQueue_fifo_31_full),
    .error        (_readData_readDataQueue_fifo_31_error),
    .data_out     (_readData_readDataQueue_fifo_31_data_out)
  );
  MaskCompress compressUnit (
    .clock                  (clock),
    .reset                  (reset),
    .in_valid               (viotaCounterAdd),
    .in_bits_maskType       (instReg_maskType),
    .in_bits_eew            (instReg_sew),
    .in_bits_uop            (instReg_decodeResult_topUop[2:0]),
    .in_bits_readFromScalar (instReg_readFromScala),
    .in_bits_source1        (source1Select),
    .in_bits_mask           (executeElementMask[31:0]),
    .in_bits_source2        (source2),
    .in_bits_pipeData       (source1),
    .in_bits_groupCounter   (requestCounter),
    .in_bits_ffoInput       ({view__in_bits_ffoInput_hi, view__in_bits_ffoInput_lo}),
    .in_bits_validInput     ({view__in_bits_validInput_hi, view__in_bits_validInput_lo}),
    .in_bits_lastCompress   (lastGroup),
    .out_data               (compressUnitResultQueue_enq_bits_data),
    .out_mask               (compressUnitResultQueue_enq_bits_mask),
    .out_groupCounter       (compressUnitResultQueue_enq_bits_groupCounter),
    .out_ffoOutput          (compressUnitResultQueue_enq_bits_ffoOutput),
    .out_compressValid      (_compressUnit_out_compressValid),
    .newInstruction         (instReq_valid),
    .ffoInstruction         (&(instReq_bits_decodeResult_topUop[2:1])),
    .writeData              (_compressUnit_writeData),
    .stageValid             (_compressUnit_stageValid)
  );
  MaskReduce reduceUnit (
    .clock               (clock),
    .reset               (reset),
    .in_ready            (_reduceUnit_in_ready),
    .in_valid            (reduceUnit_in_valid),
    .in_bits_maskType    (instReg_maskType),
    .in_bits_eew         (instReg_sew),
    .in_bits_uop         (instReg_decodeResult_topUop[2:0]),
    .in_bits_readVS1     (readVS1Reg_data),
    .in_bits_source2     (source2),
    .in_bits_sourceValid ({view__in_bits_sourceValid_hi, view__in_bits_sourceValid_lo}),
    .in_bits_lastGroup   (lastGroup),
    .in_bits_vxrm        (instReg_vxrm),
    .in_bits_aluUop      (instReg_decodeResult_uop),
    .in_bits_sign        (~instReg_decodeResult_unsigned1),
    .out_valid           (_reduceUnit_out_valid),
    .out_bits_data       (_reduceUnit_out_bits_data),
    .out_bits_mask       (_reduceUnit_out_bits_mask),
    .firstGroup          (~readVS1Reg_sendToExecution & _view__firstGroup_T_1),
    .newInstruction      (instReq_valid),
    .validInst           (|instReg_vl),
    .pop                 (instReg_decodeResult_popCount)
  );
  MaskExtend extendUnit (
    .in_eew          (instReg_sew),
    .in_uop          (instReg_decodeResult_topUop[2:0]),
    .in_source2      (source2),
    .in_groupCounter (extendGroupCount[4:0]),
    .out             (_extendUnit_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_0_enq_ready & writeQueue_0_enq_valid)),
    .pop_req_n    (~(writeQueue_0_deq_ready & ~_writeQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn),
    .empty        (_writeQueue_fifo_empty),
    .almost_empty (writeQueue_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_0_almostFull),
    .full         (_writeQueue_fifo_full),
    .error        (_writeQueue_fifo_error),
    .data_out     (_writeQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_1_enq_ready & writeQueue_1_enq_valid)),
    .pop_req_n    (~(writeQueue_1_deq_ready & ~_writeQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_1),
    .empty        (_writeQueue_fifo_1_empty),
    .almost_empty (writeQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_1_almostFull),
    .full         (_writeQueue_fifo_1_full),
    .error        (_writeQueue_fifo_1_error),
    .data_out     (_writeQueue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_2_enq_ready & writeQueue_2_enq_valid)),
    .pop_req_n    (~(writeQueue_2_deq_ready & ~_writeQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_2),
    .empty        (_writeQueue_fifo_2_empty),
    .almost_empty (writeQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_2_almostFull),
    .full         (_writeQueue_fifo_2_full),
    .error        (_writeQueue_fifo_2_error),
    .data_out     (_writeQueue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_3_enq_ready & writeQueue_3_enq_valid)),
    .pop_req_n    (~(writeQueue_3_deq_ready & ~_writeQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_3),
    .empty        (_writeQueue_fifo_3_empty),
    .almost_empty (writeQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_3_almostFull),
    .full         (_writeQueue_fifo_3_full),
    .error        (_writeQueue_fifo_3_error),
    .data_out     (_writeQueue_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_4_enq_ready & writeQueue_4_enq_valid)),
    .pop_req_n    (~(writeQueue_4_deq_ready & ~_writeQueue_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_4),
    .empty        (_writeQueue_fifo_4_empty),
    .almost_empty (writeQueue_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_4_almostFull),
    .full         (_writeQueue_fifo_4_full),
    .error        (_writeQueue_fifo_4_error),
    .data_out     (_writeQueue_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_5_enq_ready & writeQueue_5_enq_valid)),
    .pop_req_n    (~(writeQueue_5_deq_ready & ~_writeQueue_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_5),
    .empty        (_writeQueue_fifo_5_empty),
    .almost_empty (writeQueue_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_5_almostFull),
    .full         (_writeQueue_fifo_5_full),
    .error        (_writeQueue_fifo_5_error),
    .data_out     (_writeQueue_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_6_enq_ready & writeQueue_6_enq_valid)),
    .pop_req_n    (~(writeQueue_6_deq_ready & ~_writeQueue_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_6),
    .empty        (_writeQueue_fifo_6_empty),
    .almost_empty (writeQueue_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_6_almostFull),
    .full         (_writeQueue_fifo_6_full),
    .error        (_writeQueue_fifo_6_error),
    .data_out     (_writeQueue_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_7_enq_ready & writeQueue_7_enq_valid)),
    .pop_req_n    (~(writeQueue_7_deq_ready & ~_writeQueue_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_7),
    .empty        (_writeQueue_fifo_7_empty),
    .almost_empty (writeQueue_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_7_almostFull),
    .full         (_writeQueue_fifo_7_full),
    .error        (_writeQueue_fifo_7_error),
    .data_out     (_writeQueue_fifo_7_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_8_enq_ready & writeQueue_8_enq_valid)),
    .pop_req_n    (~(writeQueue_8_deq_ready & ~_writeQueue_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_8),
    .empty        (_writeQueue_fifo_8_empty),
    .almost_empty (writeQueue_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_8_almostFull),
    .full         (_writeQueue_fifo_8_full),
    .error        (_writeQueue_fifo_8_error),
    .data_out     (_writeQueue_fifo_8_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_9_enq_ready & writeQueue_9_enq_valid)),
    .pop_req_n    (~(writeQueue_9_deq_ready & ~_writeQueue_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_9),
    .empty        (_writeQueue_fifo_9_empty),
    .almost_empty (writeQueue_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_9_almostFull),
    .full         (_writeQueue_fifo_9_full),
    .error        (_writeQueue_fifo_9_error),
    .data_out     (_writeQueue_fifo_9_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_10_enq_ready & writeQueue_10_enq_valid)),
    .pop_req_n    (~(writeQueue_10_deq_ready & ~_writeQueue_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_10),
    .empty        (_writeQueue_fifo_10_empty),
    .almost_empty (writeQueue_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_10_almostFull),
    .full         (_writeQueue_fifo_10_full),
    .error        (_writeQueue_fifo_10_error),
    .data_out     (_writeQueue_fifo_10_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_11_enq_ready & writeQueue_11_enq_valid)),
    .pop_req_n    (~(writeQueue_11_deq_ready & ~_writeQueue_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_11),
    .empty        (_writeQueue_fifo_11_empty),
    .almost_empty (writeQueue_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_11_almostFull),
    .full         (_writeQueue_fifo_11_full),
    .error        (_writeQueue_fifo_11_error),
    .data_out     (_writeQueue_fifo_11_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_12_enq_ready & writeQueue_12_enq_valid)),
    .pop_req_n    (~(writeQueue_12_deq_ready & ~_writeQueue_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_12),
    .empty        (_writeQueue_fifo_12_empty),
    .almost_empty (writeQueue_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_12_almostFull),
    .full         (_writeQueue_fifo_12_full),
    .error        (_writeQueue_fifo_12_error),
    .data_out     (_writeQueue_fifo_12_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_13_enq_ready & writeQueue_13_enq_valid)),
    .pop_req_n    (~(writeQueue_13_deq_ready & ~_writeQueue_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_13),
    .empty        (_writeQueue_fifo_13_empty),
    .almost_empty (writeQueue_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_13_almostFull),
    .full         (_writeQueue_fifo_13_full),
    .error        (_writeQueue_fifo_13_error),
    .data_out     (_writeQueue_fifo_13_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_14_enq_ready & writeQueue_14_enq_valid)),
    .pop_req_n    (~(writeQueue_14_deq_ready & ~_writeQueue_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_14),
    .empty        (_writeQueue_fifo_14_empty),
    .almost_empty (writeQueue_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_14_almostFull),
    .full         (_writeQueue_fifo_14_full),
    .error        (_writeQueue_fifo_14_error),
    .data_out     (_writeQueue_fifo_14_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_15_enq_ready & writeQueue_15_enq_valid)),
    .pop_req_n    (~(writeQueue_15_deq_ready & ~_writeQueue_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_15),
    .empty        (_writeQueue_fifo_15_empty),
    .almost_empty (writeQueue_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_15_almostFull),
    .full         (_writeQueue_fifo_15_full),
    .error        (_writeQueue_fifo_15_error),
    .data_out     (_writeQueue_fifo_15_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_16 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_16_enq_ready & writeQueue_16_enq_valid)),
    .pop_req_n    (~(writeQueue_16_deq_ready & ~_writeQueue_fifo_16_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_16),
    .empty        (_writeQueue_fifo_16_empty),
    .almost_empty (writeQueue_16_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_16_almostFull),
    .full         (_writeQueue_fifo_16_full),
    .error        (_writeQueue_fifo_16_error),
    .data_out     (_writeQueue_fifo_16_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_17 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_17_enq_ready & writeQueue_17_enq_valid)),
    .pop_req_n    (~(writeQueue_17_deq_ready & ~_writeQueue_fifo_17_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_17),
    .empty        (_writeQueue_fifo_17_empty),
    .almost_empty (writeQueue_17_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_17_almostFull),
    .full         (_writeQueue_fifo_17_full),
    .error        (_writeQueue_fifo_17_error),
    .data_out     (_writeQueue_fifo_17_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_18 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_18_enq_ready & writeQueue_18_enq_valid)),
    .pop_req_n    (~(writeQueue_18_deq_ready & ~_writeQueue_fifo_18_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_18),
    .empty        (_writeQueue_fifo_18_empty),
    .almost_empty (writeQueue_18_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_18_almostFull),
    .full         (_writeQueue_fifo_18_full),
    .error        (_writeQueue_fifo_18_error),
    .data_out     (_writeQueue_fifo_18_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_19 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_19_enq_ready & writeQueue_19_enq_valid)),
    .pop_req_n    (~(writeQueue_19_deq_ready & ~_writeQueue_fifo_19_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_19),
    .empty        (_writeQueue_fifo_19_empty),
    .almost_empty (writeQueue_19_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_19_almostFull),
    .full         (_writeQueue_fifo_19_full),
    .error        (_writeQueue_fifo_19_error),
    .data_out     (_writeQueue_fifo_19_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_20 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_20_enq_ready & writeQueue_20_enq_valid)),
    .pop_req_n    (~(writeQueue_20_deq_ready & ~_writeQueue_fifo_20_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_20),
    .empty        (_writeQueue_fifo_20_empty),
    .almost_empty (writeQueue_20_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_20_almostFull),
    .full         (_writeQueue_fifo_20_full),
    .error        (_writeQueue_fifo_20_error),
    .data_out     (_writeQueue_fifo_20_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_21 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_21_enq_ready & writeQueue_21_enq_valid)),
    .pop_req_n    (~(writeQueue_21_deq_ready & ~_writeQueue_fifo_21_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_21),
    .empty        (_writeQueue_fifo_21_empty),
    .almost_empty (writeQueue_21_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_21_almostFull),
    .full         (_writeQueue_fifo_21_full),
    .error        (_writeQueue_fifo_21_error),
    .data_out     (_writeQueue_fifo_21_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_22 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_22_enq_ready & writeQueue_22_enq_valid)),
    .pop_req_n    (~(writeQueue_22_deq_ready & ~_writeQueue_fifo_22_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_22),
    .empty        (_writeQueue_fifo_22_empty),
    .almost_empty (writeQueue_22_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_22_almostFull),
    .full         (_writeQueue_fifo_22_full),
    .error        (_writeQueue_fifo_22_error),
    .data_out     (_writeQueue_fifo_22_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_23 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_23_enq_ready & writeQueue_23_enq_valid)),
    .pop_req_n    (~(writeQueue_23_deq_ready & ~_writeQueue_fifo_23_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_23),
    .empty        (_writeQueue_fifo_23_empty),
    .almost_empty (writeQueue_23_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_23_almostFull),
    .full         (_writeQueue_fifo_23_full),
    .error        (_writeQueue_fifo_23_error),
    .data_out     (_writeQueue_fifo_23_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_24 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_24_enq_ready & writeQueue_24_enq_valid)),
    .pop_req_n    (~(writeQueue_24_deq_ready & ~_writeQueue_fifo_24_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_24),
    .empty        (_writeQueue_fifo_24_empty),
    .almost_empty (writeQueue_24_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_24_almostFull),
    .full         (_writeQueue_fifo_24_full),
    .error        (_writeQueue_fifo_24_error),
    .data_out     (_writeQueue_fifo_24_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_25 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_25_enq_ready & writeQueue_25_enq_valid)),
    .pop_req_n    (~(writeQueue_25_deq_ready & ~_writeQueue_fifo_25_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_25),
    .empty        (_writeQueue_fifo_25_empty),
    .almost_empty (writeQueue_25_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_25_almostFull),
    .full         (_writeQueue_fifo_25_full),
    .error        (_writeQueue_fifo_25_error),
    .data_out     (_writeQueue_fifo_25_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_26 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_26_enq_ready & writeQueue_26_enq_valid)),
    .pop_req_n    (~(writeQueue_26_deq_ready & ~_writeQueue_fifo_26_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_26),
    .empty        (_writeQueue_fifo_26_empty),
    .almost_empty (writeQueue_26_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_26_almostFull),
    .full         (_writeQueue_fifo_26_full),
    .error        (_writeQueue_fifo_26_error),
    .data_out     (_writeQueue_fifo_26_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_27 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_27_enq_ready & writeQueue_27_enq_valid)),
    .pop_req_n    (~(writeQueue_27_deq_ready & ~_writeQueue_fifo_27_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_27),
    .empty        (_writeQueue_fifo_27_empty),
    .almost_empty (writeQueue_27_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_27_almostFull),
    .full         (_writeQueue_fifo_27_full),
    .error        (_writeQueue_fifo_27_error),
    .data_out     (_writeQueue_fifo_27_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_28 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_28_enq_ready & writeQueue_28_enq_valid)),
    .pop_req_n    (~(writeQueue_28_deq_ready & ~_writeQueue_fifo_28_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_28),
    .empty        (_writeQueue_fifo_28_empty),
    .almost_empty (writeQueue_28_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_28_almostFull),
    .full         (_writeQueue_fifo_28_full),
    .error        (_writeQueue_fifo_28_error),
    .data_out     (_writeQueue_fifo_28_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_29 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_29_enq_ready & writeQueue_29_enq_valid)),
    .pop_req_n    (~(writeQueue_29_deq_ready & ~_writeQueue_fifo_29_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_29),
    .empty        (_writeQueue_fifo_29_empty),
    .almost_empty (writeQueue_29_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_29_almostFull),
    .full         (_writeQueue_fifo_29_full),
    .error        (_writeQueue_fifo_29_error),
    .data_out     (_writeQueue_fifo_29_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_30 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_30_enq_ready & writeQueue_30_enq_valid)),
    .pop_req_n    (~(writeQueue_30_deq_ready & ~_writeQueue_fifo_30_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_30),
    .empty        (_writeQueue_fifo_30_empty),
    .almost_empty (writeQueue_30_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_30_almostFull),
    .full         (_writeQueue_fifo_30_full),
    .error        (_writeQueue_fifo_30_error),
    .data_out     (_writeQueue_fifo_30_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_31 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_31_enq_ready & writeQueue_31_enq_valid)),
    .pop_req_n    (~(writeQueue_31_deq_ready & ~_writeQueue_fifo_31_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_31),
    .empty        (_writeQueue_fifo_31_empty),
    .almost_empty (writeQueue_31_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_31_almostFull),
    .full         (_writeQueue_fifo_31_full),
    .error        (_writeQueue_fifo_31_error),
    .data_out     (_writeQueue_fifo_31_data_out)
  );
  assign exeResp_0_valid = exeResp_0_valid_0;
  assign exeResp_0_bits_vd = exeResp_0_bits_vd_0;
  assign exeResp_0_bits_offset = exeResp_0_bits_offset_0;
  assign exeResp_0_bits_mask = exeResp_0_bits_mask_0;
  assign exeResp_0_bits_data = exeResp_0_bits_data_0;
  assign exeResp_0_bits_instructionIndex = exeResp_0_bits_instructionIndex_0;
  assign exeResp_1_valid = exeResp_1_valid_0;
  assign exeResp_1_bits_vd = exeResp_1_bits_vd_0;
  assign exeResp_1_bits_offset = exeResp_1_bits_offset_0;
  assign exeResp_1_bits_mask = exeResp_1_bits_mask_0;
  assign exeResp_1_bits_data = exeResp_1_bits_data_0;
  assign exeResp_1_bits_instructionIndex = exeResp_1_bits_instructionIndex_0;
  assign exeResp_2_valid = exeResp_2_valid_0;
  assign exeResp_2_bits_vd = exeResp_2_bits_vd_0;
  assign exeResp_2_bits_offset = exeResp_2_bits_offset_0;
  assign exeResp_2_bits_mask = exeResp_2_bits_mask_0;
  assign exeResp_2_bits_data = exeResp_2_bits_data_0;
  assign exeResp_2_bits_instructionIndex = exeResp_2_bits_instructionIndex_0;
  assign exeResp_3_valid = exeResp_3_valid_0;
  assign exeResp_3_bits_vd = exeResp_3_bits_vd_0;
  assign exeResp_3_bits_offset = exeResp_3_bits_offset_0;
  assign exeResp_3_bits_mask = exeResp_3_bits_mask_0;
  assign exeResp_3_bits_data = exeResp_3_bits_data_0;
  assign exeResp_3_bits_instructionIndex = exeResp_3_bits_instructionIndex_0;
  assign exeResp_4_valid = exeResp_4_valid_0;
  assign exeResp_4_bits_vd = exeResp_4_bits_vd_0;
  assign exeResp_4_bits_offset = exeResp_4_bits_offset_0;
  assign exeResp_4_bits_mask = exeResp_4_bits_mask_0;
  assign exeResp_4_bits_data = exeResp_4_bits_data_0;
  assign exeResp_4_bits_instructionIndex = exeResp_4_bits_instructionIndex_0;
  assign exeResp_5_valid = exeResp_5_valid_0;
  assign exeResp_5_bits_vd = exeResp_5_bits_vd_0;
  assign exeResp_5_bits_offset = exeResp_5_bits_offset_0;
  assign exeResp_5_bits_mask = exeResp_5_bits_mask_0;
  assign exeResp_5_bits_data = exeResp_5_bits_data_0;
  assign exeResp_5_bits_instructionIndex = exeResp_5_bits_instructionIndex_0;
  assign exeResp_6_valid = exeResp_6_valid_0;
  assign exeResp_6_bits_vd = exeResp_6_bits_vd_0;
  assign exeResp_6_bits_offset = exeResp_6_bits_offset_0;
  assign exeResp_6_bits_mask = exeResp_6_bits_mask_0;
  assign exeResp_6_bits_data = exeResp_6_bits_data_0;
  assign exeResp_6_bits_instructionIndex = exeResp_6_bits_instructionIndex_0;
  assign exeResp_7_valid = exeResp_7_valid_0;
  assign exeResp_7_bits_vd = exeResp_7_bits_vd_0;
  assign exeResp_7_bits_offset = exeResp_7_bits_offset_0;
  assign exeResp_7_bits_mask = exeResp_7_bits_mask_0;
  assign exeResp_7_bits_data = exeResp_7_bits_data_0;
  assign exeResp_7_bits_instructionIndex = exeResp_7_bits_instructionIndex_0;
  assign exeResp_8_valid = exeResp_8_valid_0;
  assign exeResp_8_bits_vd = exeResp_8_bits_vd_0;
  assign exeResp_8_bits_offset = exeResp_8_bits_offset_0;
  assign exeResp_8_bits_mask = exeResp_8_bits_mask_0;
  assign exeResp_8_bits_data = exeResp_8_bits_data_0;
  assign exeResp_8_bits_instructionIndex = exeResp_8_bits_instructionIndex_0;
  assign exeResp_9_valid = exeResp_9_valid_0;
  assign exeResp_9_bits_vd = exeResp_9_bits_vd_0;
  assign exeResp_9_bits_offset = exeResp_9_bits_offset_0;
  assign exeResp_9_bits_mask = exeResp_9_bits_mask_0;
  assign exeResp_9_bits_data = exeResp_9_bits_data_0;
  assign exeResp_9_bits_instructionIndex = exeResp_9_bits_instructionIndex_0;
  assign exeResp_10_valid = exeResp_10_valid_0;
  assign exeResp_10_bits_vd = exeResp_10_bits_vd_0;
  assign exeResp_10_bits_offset = exeResp_10_bits_offset_0;
  assign exeResp_10_bits_mask = exeResp_10_bits_mask_0;
  assign exeResp_10_bits_data = exeResp_10_bits_data_0;
  assign exeResp_10_bits_instructionIndex = exeResp_10_bits_instructionIndex_0;
  assign exeResp_11_valid = exeResp_11_valid_0;
  assign exeResp_11_bits_vd = exeResp_11_bits_vd_0;
  assign exeResp_11_bits_offset = exeResp_11_bits_offset_0;
  assign exeResp_11_bits_mask = exeResp_11_bits_mask_0;
  assign exeResp_11_bits_data = exeResp_11_bits_data_0;
  assign exeResp_11_bits_instructionIndex = exeResp_11_bits_instructionIndex_0;
  assign exeResp_12_valid = exeResp_12_valid_0;
  assign exeResp_12_bits_vd = exeResp_12_bits_vd_0;
  assign exeResp_12_bits_offset = exeResp_12_bits_offset_0;
  assign exeResp_12_bits_mask = exeResp_12_bits_mask_0;
  assign exeResp_12_bits_data = exeResp_12_bits_data_0;
  assign exeResp_12_bits_instructionIndex = exeResp_12_bits_instructionIndex_0;
  assign exeResp_13_valid = exeResp_13_valid_0;
  assign exeResp_13_bits_vd = exeResp_13_bits_vd_0;
  assign exeResp_13_bits_offset = exeResp_13_bits_offset_0;
  assign exeResp_13_bits_mask = exeResp_13_bits_mask_0;
  assign exeResp_13_bits_data = exeResp_13_bits_data_0;
  assign exeResp_13_bits_instructionIndex = exeResp_13_bits_instructionIndex_0;
  assign exeResp_14_valid = exeResp_14_valid_0;
  assign exeResp_14_bits_vd = exeResp_14_bits_vd_0;
  assign exeResp_14_bits_offset = exeResp_14_bits_offset_0;
  assign exeResp_14_bits_mask = exeResp_14_bits_mask_0;
  assign exeResp_14_bits_data = exeResp_14_bits_data_0;
  assign exeResp_14_bits_instructionIndex = exeResp_14_bits_instructionIndex_0;
  assign exeResp_15_valid = exeResp_15_valid_0;
  assign exeResp_15_bits_vd = exeResp_15_bits_vd_0;
  assign exeResp_15_bits_offset = exeResp_15_bits_offset_0;
  assign exeResp_15_bits_mask = exeResp_15_bits_mask_0;
  assign exeResp_15_bits_data = exeResp_15_bits_data_0;
  assign exeResp_15_bits_instructionIndex = exeResp_15_bits_instructionIndex_0;
  assign exeResp_16_valid = exeResp_16_valid_0;
  assign exeResp_16_bits_vd = exeResp_16_bits_vd_0;
  assign exeResp_16_bits_offset = exeResp_16_bits_offset_0;
  assign exeResp_16_bits_mask = exeResp_16_bits_mask_0;
  assign exeResp_16_bits_data = exeResp_16_bits_data_0;
  assign exeResp_16_bits_instructionIndex = exeResp_16_bits_instructionIndex_0;
  assign exeResp_17_valid = exeResp_17_valid_0;
  assign exeResp_17_bits_vd = exeResp_17_bits_vd_0;
  assign exeResp_17_bits_offset = exeResp_17_bits_offset_0;
  assign exeResp_17_bits_mask = exeResp_17_bits_mask_0;
  assign exeResp_17_bits_data = exeResp_17_bits_data_0;
  assign exeResp_17_bits_instructionIndex = exeResp_17_bits_instructionIndex_0;
  assign exeResp_18_valid = exeResp_18_valid_0;
  assign exeResp_18_bits_vd = exeResp_18_bits_vd_0;
  assign exeResp_18_bits_offset = exeResp_18_bits_offset_0;
  assign exeResp_18_bits_mask = exeResp_18_bits_mask_0;
  assign exeResp_18_bits_data = exeResp_18_bits_data_0;
  assign exeResp_18_bits_instructionIndex = exeResp_18_bits_instructionIndex_0;
  assign exeResp_19_valid = exeResp_19_valid_0;
  assign exeResp_19_bits_vd = exeResp_19_bits_vd_0;
  assign exeResp_19_bits_offset = exeResp_19_bits_offset_0;
  assign exeResp_19_bits_mask = exeResp_19_bits_mask_0;
  assign exeResp_19_bits_data = exeResp_19_bits_data_0;
  assign exeResp_19_bits_instructionIndex = exeResp_19_bits_instructionIndex_0;
  assign exeResp_20_valid = exeResp_20_valid_0;
  assign exeResp_20_bits_vd = exeResp_20_bits_vd_0;
  assign exeResp_20_bits_offset = exeResp_20_bits_offset_0;
  assign exeResp_20_bits_mask = exeResp_20_bits_mask_0;
  assign exeResp_20_bits_data = exeResp_20_bits_data_0;
  assign exeResp_20_bits_instructionIndex = exeResp_20_bits_instructionIndex_0;
  assign exeResp_21_valid = exeResp_21_valid_0;
  assign exeResp_21_bits_vd = exeResp_21_bits_vd_0;
  assign exeResp_21_bits_offset = exeResp_21_bits_offset_0;
  assign exeResp_21_bits_mask = exeResp_21_bits_mask_0;
  assign exeResp_21_bits_data = exeResp_21_bits_data_0;
  assign exeResp_21_bits_instructionIndex = exeResp_21_bits_instructionIndex_0;
  assign exeResp_22_valid = exeResp_22_valid_0;
  assign exeResp_22_bits_vd = exeResp_22_bits_vd_0;
  assign exeResp_22_bits_offset = exeResp_22_bits_offset_0;
  assign exeResp_22_bits_mask = exeResp_22_bits_mask_0;
  assign exeResp_22_bits_data = exeResp_22_bits_data_0;
  assign exeResp_22_bits_instructionIndex = exeResp_22_bits_instructionIndex_0;
  assign exeResp_23_valid = exeResp_23_valid_0;
  assign exeResp_23_bits_vd = exeResp_23_bits_vd_0;
  assign exeResp_23_bits_offset = exeResp_23_bits_offset_0;
  assign exeResp_23_bits_mask = exeResp_23_bits_mask_0;
  assign exeResp_23_bits_data = exeResp_23_bits_data_0;
  assign exeResp_23_bits_instructionIndex = exeResp_23_bits_instructionIndex_0;
  assign exeResp_24_valid = exeResp_24_valid_0;
  assign exeResp_24_bits_vd = exeResp_24_bits_vd_0;
  assign exeResp_24_bits_offset = exeResp_24_bits_offset_0;
  assign exeResp_24_bits_mask = exeResp_24_bits_mask_0;
  assign exeResp_24_bits_data = exeResp_24_bits_data_0;
  assign exeResp_24_bits_instructionIndex = exeResp_24_bits_instructionIndex_0;
  assign exeResp_25_valid = exeResp_25_valid_0;
  assign exeResp_25_bits_vd = exeResp_25_bits_vd_0;
  assign exeResp_25_bits_offset = exeResp_25_bits_offset_0;
  assign exeResp_25_bits_mask = exeResp_25_bits_mask_0;
  assign exeResp_25_bits_data = exeResp_25_bits_data_0;
  assign exeResp_25_bits_instructionIndex = exeResp_25_bits_instructionIndex_0;
  assign exeResp_26_valid = exeResp_26_valid_0;
  assign exeResp_26_bits_vd = exeResp_26_bits_vd_0;
  assign exeResp_26_bits_offset = exeResp_26_bits_offset_0;
  assign exeResp_26_bits_mask = exeResp_26_bits_mask_0;
  assign exeResp_26_bits_data = exeResp_26_bits_data_0;
  assign exeResp_26_bits_instructionIndex = exeResp_26_bits_instructionIndex_0;
  assign exeResp_27_valid = exeResp_27_valid_0;
  assign exeResp_27_bits_vd = exeResp_27_bits_vd_0;
  assign exeResp_27_bits_offset = exeResp_27_bits_offset_0;
  assign exeResp_27_bits_mask = exeResp_27_bits_mask_0;
  assign exeResp_27_bits_data = exeResp_27_bits_data_0;
  assign exeResp_27_bits_instructionIndex = exeResp_27_bits_instructionIndex_0;
  assign exeResp_28_valid = exeResp_28_valid_0;
  assign exeResp_28_bits_vd = exeResp_28_bits_vd_0;
  assign exeResp_28_bits_offset = exeResp_28_bits_offset_0;
  assign exeResp_28_bits_mask = exeResp_28_bits_mask_0;
  assign exeResp_28_bits_data = exeResp_28_bits_data_0;
  assign exeResp_28_bits_instructionIndex = exeResp_28_bits_instructionIndex_0;
  assign exeResp_29_valid = exeResp_29_valid_0;
  assign exeResp_29_bits_vd = exeResp_29_bits_vd_0;
  assign exeResp_29_bits_offset = exeResp_29_bits_offset_0;
  assign exeResp_29_bits_mask = exeResp_29_bits_mask_0;
  assign exeResp_29_bits_data = exeResp_29_bits_data_0;
  assign exeResp_29_bits_instructionIndex = exeResp_29_bits_instructionIndex_0;
  assign exeResp_30_valid = exeResp_30_valid_0;
  assign exeResp_30_bits_vd = exeResp_30_bits_vd_0;
  assign exeResp_30_bits_offset = exeResp_30_bits_offset_0;
  assign exeResp_30_bits_mask = exeResp_30_bits_mask_0;
  assign exeResp_30_bits_data = exeResp_30_bits_data_0;
  assign exeResp_30_bits_instructionIndex = exeResp_30_bits_instructionIndex_0;
  assign exeResp_31_valid = exeResp_31_valid_0;
  assign exeResp_31_bits_vd = exeResp_31_bits_vd_0;
  assign exeResp_31_bits_offset = exeResp_31_bits_offset_0;
  assign exeResp_31_bits_mask = exeResp_31_bits_mask_0;
  assign exeResp_31_bits_data = exeResp_31_bits_data_0;
  assign exeResp_31_bits_instructionIndex = exeResp_31_bits_instructionIndex_0;
  assign tokenIO_0_maskRequestRelease = tokenIO_0_maskRequestRelease_0;
  assign tokenIO_1_maskRequestRelease = tokenIO_1_maskRequestRelease_0;
  assign tokenIO_2_maskRequestRelease = tokenIO_2_maskRequestRelease_0;
  assign tokenIO_3_maskRequestRelease = tokenIO_3_maskRequestRelease_0;
  assign tokenIO_4_maskRequestRelease = tokenIO_4_maskRequestRelease_0;
  assign tokenIO_5_maskRequestRelease = tokenIO_5_maskRequestRelease_0;
  assign tokenIO_6_maskRequestRelease = tokenIO_6_maskRequestRelease_0;
  assign tokenIO_7_maskRequestRelease = tokenIO_7_maskRequestRelease_0;
  assign tokenIO_8_maskRequestRelease = tokenIO_8_maskRequestRelease_0;
  assign tokenIO_9_maskRequestRelease = tokenIO_9_maskRequestRelease_0;
  assign tokenIO_10_maskRequestRelease = tokenIO_10_maskRequestRelease_0;
  assign tokenIO_11_maskRequestRelease = tokenIO_11_maskRequestRelease_0;
  assign tokenIO_12_maskRequestRelease = tokenIO_12_maskRequestRelease_0;
  assign tokenIO_13_maskRequestRelease = tokenIO_13_maskRequestRelease_0;
  assign tokenIO_14_maskRequestRelease = tokenIO_14_maskRequestRelease_0;
  assign tokenIO_15_maskRequestRelease = tokenIO_15_maskRequestRelease_0;
  assign tokenIO_16_maskRequestRelease = tokenIO_16_maskRequestRelease_0;
  assign tokenIO_17_maskRequestRelease = tokenIO_17_maskRequestRelease_0;
  assign tokenIO_18_maskRequestRelease = tokenIO_18_maskRequestRelease_0;
  assign tokenIO_19_maskRequestRelease = tokenIO_19_maskRequestRelease_0;
  assign tokenIO_20_maskRequestRelease = tokenIO_20_maskRequestRelease_0;
  assign tokenIO_21_maskRequestRelease = tokenIO_21_maskRequestRelease_0;
  assign tokenIO_22_maskRequestRelease = tokenIO_22_maskRequestRelease_0;
  assign tokenIO_23_maskRequestRelease = tokenIO_23_maskRequestRelease_0;
  assign tokenIO_24_maskRequestRelease = tokenIO_24_maskRequestRelease_0;
  assign tokenIO_25_maskRequestRelease = tokenIO_25_maskRequestRelease_0;
  assign tokenIO_26_maskRequestRelease = tokenIO_26_maskRequestRelease_0;
  assign tokenIO_27_maskRequestRelease = tokenIO_27_maskRequestRelease_0;
  assign tokenIO_28_maskRequestRelease = tokenIO_28_maskRequestRelease_0;
  assign tokenIO_29_maskRequestRelease = tokenIO_29_maskRequestRelease_0;
  assign tokenIO_30_maskRequestRelease = tokenIO_30_maskRequestRelease_0;
  assign tokenIO_31_maskRequestRelease = tokenIO_31_maskRequestRelease_0;
  assign readChannel_0_valid = readChannel_0_valid_0;
  assign readChannel_0_bits_vs = readChannel_0_bits_vs_0;
  assign readChannel_0_bits_offset = readChannel_0_bits_offset_0;
  assign readChannel_0_bits_instructionIndex = readChannel_0_bits_instructionIndex_0;
  assign readChannel_1_valid = readChannel_1_valid_0;
  assign readChannel_1_bits_vs = readChannel_1_bits_vs_0;
  assign readChannel_1_bits_offset = readChannel_1_bits_offset_0;
  assign readChannel_1_bits_instructionIndex = readChannel_1_bits_instructionIndex_0;
  assign readChannel_2_valid = readChannel_2_valid_0;
  assign readChannel_2_bits_vs = readChannel_2_bits_vs_0;
  assign readChannel_2_bits_offset = readChannel_2_bits_offset_0;
  assign readChannel_2_bits_instructionIndex = readChannel_2_bits_instructionIndex_0;
  assign readChannel_3_valid = readChannel_3_valid_0;
  assign readChannel_3_bits_vs = readChannel_3_bits_vs_0;
  assign readChannel_3_bits_offset = readChannel_3_bits_offset_0;
  assign readChannel_3_bits_instructionIndex = readChannel_3_bits_instructionIndex_0;
  assign readChannel_4_valid = readChannel_4_valid_0;
  assign readChannel_4_bits_vs = readChannel_4_bits_vs_0;
  assign readChannel_4_bits_offset = readChannel_4_bits_offset_0;
  assign readChannel_4_bits_instructionIndex = readChannel_4_bits_instructionIndex_0;
  assign readChannel_5_valid = readChannel_5_valid_0;
  assign readChannel_5_bits_vs = readChannel_5_bits_vs_0;
  assign readChannel_5_bits_offset = readChannel_5_bits_offset_0;
  assign readChannel_5_bits_instructionIndex = readChannel_5_bits_instructionIndex_0;
  assign readChannel_6_valid = readChannel_6_valid_0;
  assign readChannel_6_bits_vs = readChannel_6_bits_vs_0;
  assign readChannel_6_bits_offset = readChannel_6_bits_offset_0;
  assign readChannel_6_bits_instructionIndex = readChannel_6_bits_instructionIndex_0;
  assign readChannel_7_valid = readChannel_7_valid_0;
  assign readChannel_7_bits_vs = readChannel_7_bits_vs_0;
  assign readChannel_7_bits_offset = readChannel_7_bits_offset_0;
  assign readChannel_7_bits_instructionIndex = readChannel_7_bits_instructionIndex_0;
  assign readChannel_8_valid = readChannel_8_valid_0;
  assign readChannel_8_bits_vs = readChannel_8_bits_vs_0;
  assign readChannel_8_bits_offset = readChannel_8_bits_offset_0;
  assign readChannel_8_bits_instructionIndex = readChannel_8_bits_instructionIndex_0;
  assign readChannel_9_valid = readChannel_9_valid_0;
  assign readChannel_9_bits_vs = readChannel_9_bits_vs_0;
  assign readChannel_9_bits_offset = readChannel_9_bits_offset_0;
  assign readChannel_9_bits_instructionIndex = readChannel_9_bits_instructionIndex_0;
  assign readChannel_10_valid = readChannel_10_valid_0;
  assign readChannel_10_bits_vs = readChannel_10_bits_vs_0;
  assign readChannel_10_bits_offset = readChannel_10_bits_offset_0;
  assign readChannel_10_bits_instructionIndex = readChannel_10_bits_instructionIndex_0;
  assign readChannel_11_valid = readChannel_11_valid_0;
  assign readChannel_11_bits_vs = readChannel_11_bits_vs_0;
  assign readChannel_11_bits_offset = readChannel_11_bits_offset_0;
  assign readChannel_11_bits_instructionIndex = readChannel_11_bits_instructionIndex_0;
  assign readChannel_12_valid = readChannel_12_valid_0;
  assign readChannel_12_bits_vs = readChannel_12_bits_vs_0;
  assign readChannel_12_bits_offset = readChannel_12_bits_offset_0;
  assign readChannel_12_bits_instructionIndex = readChannel_12_bits_instructionIndex_0;
  assign readChannel_13_valid = readChannel_13_valid_0;
  assign readChannel_13_bits_vs = readChannel_13_bits_vs_0;
  assign readChannel_13_bits_offset = readChannel_13_bits_offset_0;
  assign readChannel_13_bits_instructionIndex = readChannel_13_bits_instructionIndex_0;
  assign readChannel_14_valid = readChannel_14_valid_0;
  assign readChannel_14_bits_vs = readChannel_14_bits_vs_0;
  assign readChannel_14_bits_offset = readChannel_14_bits_offset_0;
  assign readChannel_14_bits_instructionIndex = readChannel_14_bits_instructionIndex_0;
  assign readChannel_15_valid = readChannel_15_valid_0;
  assign readChannel_15_bits_vs = readChannel_15_bits_vs_0;
  assign readChannel_15_bits_offset = readChannel_15_bits_offset_0;
  assign readChannel_15_bits_instructionIndex = readChannel_15_bits_instructionIndex_0;
  assign readChannel_16_valid = readChannel_16_valid_0;
  assign readChannel_16_bits_vs = readChannel_16_bits_vs_0;
  assign readChannel_16_bits_offset = readChannel_16_bits_offset_0;
  assign readChannel_16_bits_instructionIndex = readChannel_16_bits_instructionIndex_0;
  assign readChannel_17_valid = readChannel_17_valid_0;
  assign readChannel_17_bits_vs = readChannel_17_bits_vs_0;
  assign readChannel_17_bits_offset = readChannel_17_bits_offset_0;
  assign readChannel_17_bits_instructionIndex = readChannel_17_bits_instructionIndex_0;
  assign readChannel_18_valid = readChannel_18_valid_0;
  assign readChannel_18_bits_vs = readChannel_18_bits_vs_0;
  assign readChannel_18_bits_offset = readChannel_18_bits_offset_0;
  assign readChannel_18_bits_instructionIndex = readChannel_18_bits_instructionIndex_0;
  assign readChannel_19_valid = readChannel_19_valid_0;
  assign readChannel_19_bits_vs = readChannel_19_bits_vs_0;
  assign readChannel_19_bits_offset = readChannel_19_bits_offset_0;
  assign readChannel_19_bits_instructionIndex = readChannel_19_bits_instructionIndex_0;
  assign readChannel_20_valid = readChannel_20_valid_0;
  assign readChannel_20_bits_vs = readChannel_20_bits_vs_0;
  assign readChannel_20_bits_offset = readChannel_20_bits_offset_0;
  assign readChannel_20_bits_instructionIndex = readChannel_20_bits_instructionIndex_0;
  assign readChannel_21_valid = readChannel_21_valid_0;
  assign readChannel_21_bits_vs = readChannel_21_bits_vs_0;
  assign readChannel_21_bits_offset = readChannel_21_bits_offset_0;
  assign readChannel_21_bits_instructionIndex = readChannel_21_bits_instructionIndex_0;
  assign readChannel_22_valid = readChannel_22_valid_0;
  assign readChannel_22_bits_vs = readChannel_22_bits_vs_0;
  assign readChannel_22_bits_offset = readChannel_22_bits_offset_0;
  assign readChannel_22_bits_instructionIndex = readChannel_22_bits_instructionIndex_0;
  assign readChannel_23_valid = readChannel_23_valid_0;
  assign readChannel_23_bits_vs = readChannel_23_bits_vs_0;
  assign readChannel_23_bits_offset = readChannel_23_bits_offset_0;
  assign readChannel_23_bits_instructionIndex = readChannel_23_bits_instructionIndex_0;
  assign readChannel_24_valid = readChannel_24_valid_0;
  assign readChannel_24_bits_vs = readChannel_24_bits_vs_0;
  assign readChannel_24_bits_offset = readChannel_24_bits_offset_0;
  assign readChannel_24_bits_instructionIndex = readChannel_24_bits_instructionIndex_0;
  assign readChannel_25_valid = readChannel_25_valid_0;
  assign readChannel_25_bits_vs = readChannel_25_bits_vs_0;
  assign readChannel_25_bits_offset = readChannel_25_bits_offset_0;
  assign readChannel_25_bits_instructionIndex = readChannel_25_bits_instructionIndex_0;
  assign readChannel_26_valid = readChannel_26_valid_0;
  assign readChannel_26_bits_vs = readChannel_26_bits_vs_0;
  assign readChannel_26_bits_offset = readChannel_26_bits_offset_0;
  assign readChannel_26_bits_instructionIndex = readChannel_26_bits_instructionIndex_0;
  assign readChannel_27_valid = readChannel_27_valid_0;
  assign readChannel_27_bits_vs = readChannel_27_bits_vs_0;
  assign readChannel_27_bits_offset = readChannel_27_bits_offset_0;
  assign readChannel_27_bits_instructionIndex = readChannel_27_bits_instructionIndex_0;
  assign readChannel_28_valid = readChannel_28_valid_0;
  assign readChannel_28_bits_vs = readChannel_28_bits_vs_0;
  assign readChannel_28_bits_offset = readChannel_28_bits_offset_0;
  assign readChannel_28_bits_instructionIndex = readChannel_28_bits_instructionIndex_0;
  assign readChannel_29_valid = readChannel_29_valid_0;
  assign readChannel_29_bits_vs = readChannel_29_bits_vs_0;
  assign readChannel_29_bits_offset = readChannel_29_bits_offset_0;
  assign readChannel_29_bits_instructionIndex = readChannel_29_bits_instructionIndex_0;
  assign readChannel_30_valid = readChannel_30_valid_0;
  assign readChannel_30_bits_vs = readChannel_30_bits_vs_0;
  assign readChannel_30_bits_offset = readChannel_30_bits_offset_0;
  assign readChannel_30_bits_instructionIndex = readChannel_30_bits_instructionIndex_0;
  assign readChannel_31_valid = readChannel_31_valid_0;
  assign readChannel_31_bits_vs = readChannel_31_bits_vs_0;
  assign readChannel_31_bits_offset = readChannel_31_bits_offset_0;
  assign readChannel_31_bits_instructionIndex = readChannel_31_bits_instructionIndex_0;
  assign lastReport = _lastReport_output;
  assign laneMaskInput_0 = laneMaskSelect_0[0] ? v0SelectBySew[63:32] : v0SelectBySew[31:0];
  assign laneMaskInput_1 = laneMaskSelect_1[0] ? v0SelectBySew_1[63:32] : v0SelectBySew_1[31:0];
  assign laneMaskInput_2 = laneMaskSelect_2[0] ? v0SelectBySew_2[63:32] : v0SelectBySew_2[31:0];
  assign laneMaskInput_3 = laneMaskSelect_3[0] ? v0SelectBySew_3[63:32] : v0SelectBySew_3[31:0];
  assign laneMaskInput_4 = laneMaskSelect_4[0] ? v0SelectBySew_4[63:32] : v0SelectBySew_4[31:0];
  assign laneMaskInput_5 = laneMaskSelect_5[0] ? v0SelectBySew_5[63:32] : v0SelectBySew_5[31:0];
  assign laneMaskInput_6 = laneMaskSelect_6[0] ? v0SelectBySew_6[63:32] : v0SelectBySew_6[31:0];
  assign laneMaskInput_7 = laneMaskSelect_7[0] ? v0SelectBySew_7[63:32] : v0SelectBySew_7[31:0];
  assign laneMaskInput_8 = laneMaskSelect_8[0] ? v0SelectBySew_8[63:32] : v0SelectBySew_8[31:0];
  assign laneMaskInput_9 = laneMaskSelect_9[0] ? v0SelectBySew_9[63:32] : v0SelectBySew_9[31:0];
  assign laneMaskInput_10 = laneMaskSelect_10[0] ? v0SelectBySew_10[63:32] : v0SelectBySew_10[31:0];
  assign laneMaskInput_11 = laneMaskSelect_11[0] ? v0SelectBySew_11[63:32] : v0SelectBySew_11[31:0];
  assign laneMaskInput_12 = laneMaskSelect_12[0] ? v0SelectBySew_12[63:32] : v0SelectBySew_12[31:0];
  assign laneMaskInput_13 = laneMaskSelect_13[0] ? v0SelectBySew_13[63:32] : v0SelectBySew_13[31:0];
  assign laneMaskInput_14 = laneMaskSelect_14[0] ? v0SelectBySew_14[63:32] : v0SelectBySew_14[31:0];
  assign laneMaskInput_15 = laneMaskSelect_15[0] ? v0SelectBySew_15[63:32] : v0SelectBySew_15[31:0];
  assign laneMaskInput_16 = laneMaskSelect_16[0] ? v0SelectBySew_16[63:32] : v0SelectBySew_16[31:0];
  assign laneMaskInput_17 = laneMaskSelect_17[0] ? v0SelectBySew_17[63:32] : v0SelectBySew_17[31:0];
  assign laneMaskInput_18 = laneMaskSelect_18[0] ? v0SelectBySew_18[63:32] : v0SelectBySew_18[31:0];
  assign laneMaskInput_19 = laneMaskSelect_19[0] ? v0SelectBySew_19[63:32] : v0SelectBySew_19[31:0];
  assign laneMaskInput_20 = laneMaskSelect_20[0] ? v0SelectBySew_20[63:32] : v0SelectBySew_20[31:0];
  assign laneMaskInput_21 = laneMaskSelect_21[0] ? v0SelectBySew_21[63:32] : v0SelectBySew_21[31:0];
  assign laneMaskInput_22 = laneMaskSelect_22[0] ? v0SelectBySew_22[63:32] : v0SelectBySew_22[31:0];
  assign laneMaskInput_23 = laneMaskSelect_23[0] ? v0SelectBySew_23[63:32] : v0SelectBySew_23[31:0];
  assign laneMaskInput_24 = laneMaskSelect_24[0] ? v0SelectBySew_24[63:32] : v0SelectBySew_24[31:0];
  assign laneMaskInput_25 = laneMaskSelect_25[0] ? v0SelectBySew_25[63:32] : v0SelectBySew_25[31:0];
  assign laneMaskInput_26 = laneMaskSelect_26[0] ? v0SelectBySew_26[63:32] : v0SelectBySew_26[31:0];
  assign laneMaskInput_27 = laneMaskSelect_27[0] ? v0SelectBySew_27[63:32] : v0SelectBySew_27[31:0];
  assign laneMaskInput_28 = laneMaskSelect_28[0] ? v0SelectBySew_28[63:32] : v0SelectBySew_28[31:0];
  assign laneMaskInput_29 = laneMaskSelect_29[0] ? v0SelectBySew_29[63:32] : v0SelectBySew_29[31:0];
  assign laneMaskInput_30 = laneMaskSelect_30[0] ? v0SelectBySew_30[63:32] : v0SelectBySew_30[31:0];
  assign laneMaskInput_31 = laneMaskSelect_31[0] ? v0SelectBySew_31[63:32] : v0SelectBySew_31[31:0];
  assign writeRDData = instReg_decodeResult_popCount ? _reduceUnit_out_bits_data : _compressUnit_writeData;
  assign gatherData_valid = gatherData_valid_0;
  assign gatherData_bits = gatherData_bits_0;
endmodule

