module VectorAdder(
  input  [31:0] a,
                b,
  output [31:0] z,
  input  [2:0]  sew,
  input  [3:0]  cin,
  output [3:0]  cout
);

  wire        as_0 = a[0];
  wire        as_1 = a[1];
  wire        as_2 = a[2];
  wire        as_3 = a[3];
  wire        as_4 = a[4];
  wire        as_5 = a[5];
  wire        as_6 = a[6];
  wire        as_7 = a[7];
  wire        as_8 = a[8];
  wire        as_9 = a[9];
  wire        as_10 = a[10];
  wire        as_11 = a[11];
  wire        as_12 = a[12];
  wire        as_13 = a[13];
  wire        as_14 = a[14];
  wire        as_15 = a[15];
  wire        as_16 = a[16];
  wire        as_17 = a[17];
  wire        as_18 = a[18];
  wire        as_19 = a[19];
  wire        as_20 = a[20];
  wire        as_21 = a[21];
  wire        as_22 = a[22];
  wire        as_23 = a[23];
  wire        as_24 = a[24];
  wire        as_25 = a[25];
  wire        as_26 = a[26];
  wire        as_27 = a[27];
  wire        as_28 = a[28];
  wire        as_29 = a[29];
  wire        as_30 = a[30];
  wire        as_31 = a[31];
  wire        bs_0 = b[0];
  wire        bs_1 = b[1];
  wire        bs_2 = b[2];
  wire        bs_3 = b[3];
  wire        bs_4 = b[4];
  wire        bs_5 = b[5];
  wire        bs_6 = b[6];
  wire        bs_7 = b[7];
  wire        bs_8 = b[8];
  wire        bs_9 = b[9];
  wire        bs_10 = b[10];
  wire        bs_11 = b[11];
  wire        bs_12 = b[12];
  wire        bs_13 = b[13];
  wire        bs_14 = b[14];
  wire        bs_15 = b[15];
  wire        bs_16 = b[16];
  wire        bs_17 = b[17];
  wire        bs_18 = b[18];
  wire        bs_19 = b[19];
  wire        bs_20 = b[20];
  wire        bs_21 = b[21];
  wire        bs_22 = b[22];
  wire        bs_23 = b[23];
  wire        bs_24 = b[24];
  wire        bs_25 = b[25];
  wire        bs_26 = b[26];
  wire        bs_27 = b[27];
  wire        bs_28 = b[28];
  wire        bs_29 = b[29];
  wire        bs_30 = b[30];
  wire        bs_31 = b[31];
  wire        pairs_0_1 = as_0 ^ bs_0;
  wire        pairs_0_2 = as_0 & bs_0;
  wire        pairs_1_1 = as_1 ^ bs_1;
  wire        pairs_1_2 = as_1 & bs_1;
  wire        pairs_2_1 = as_2 ^ bs_2;
  wire        pairs_2_2 = as_2 & bs_2;
  wire        pairs_3_1 = as_3 ^ bs_3;
  wire        pairs_3_2 = as_3 & bs_3;
  wire        pairs_4_1 = as_4 ^ bs_4;
  wire        pairs_4_2 = as_4 & bs_4;
  wire        pairs_5_1 = as_5 ^ bs_5;
  wire        pairs_5_2 = as_5 & bs_5;
  wire        pairs_6_1 = as_6 ^ bs_6;
  wire        pairs_6_2 = as_6 & bs_6;
  wire        pairs_7_1 = as_7 ^ bs_7;
  wire        pairs_7_2 = as_7 & bs_7;
  wire        pairs_8_1 = as_8 ^ bs_8;
  wire        pairs_8_2 = as_8 & bs_8;
  wire        pairs_9_1 = as_9 ^ bs_9;
  wire        pairs_9_2 = as_9 & bs_9;
  wire        pairs_10_1 = as_10 ^ bs_10;
  wire        pairs_10_2 = as_10 & bs_10;
  wire        pairs_11_1 = as_11 ^ bs_11;
  wire        pairs_11_2 = as_11 & bs_11;
  wire        pairs_12_1 = as_12 ^ bs_12;
  wire        pairs_12_2 = as_12 & bs_12;
  wire        pairs_13_1 = as_13 ^ bs_13;
  wire        pairs_13_2 = as_13 & bs_13;
  wire        pairs_14_1 = as_14 ^ bs_14;
  wire        pairs_14_2 = as_14 & bs_14;
  wire        pairs_15_1 = as_15 ^ bs_15;
  wire        pairs_15_2 = as_15 & bs_15;
  wire        pairs_16_1 = as_16 ^ bs_16;
  wire        pairs_16_2 = as_16 & bs_16;
  wire        pairs_17_1 = as_17 ^ bs_17;
  wire        pairs_17_2 = as_17 & bs_17;
  wire        pairs_18_1 = as_18 ^ bs_18;
  wire        pairs_18_2 = as_18 & bs_18;
  wire        pairs_19_1 = as_19 ^ bs_19;
  wire        pairs_19_2 = as_19 & bs_19;
  wire        pairs_20_1 = as_20 ^ bs_20;
  wire        pairs_20_2 = as_20 & bs_20;
  wire        pairs_21_1 = as_21 ^ bs_21;
  wire        pairs_21_2 = as_21 & bs_21;
  wire        pairs_22_1 = as_22 ^ bs_22;
  wire        pairs_22_2 = as_22 & bs_22;
  wire        pairs_23_1 = as_23 ^ bs_23;
  wire        pairs_23_2 = as_23 & bs_23;
  wire        pairs_24_1 = as_24 ^ bs_24;
  wire        pairs_24_2 = as_24 & bs_24;
  wire        pairs_25_1 = as_25 ^ bs_25;
  wire        pairs_25_2 = as_25 & bs_25;
  wire        pairs_26_1 = as_26 ^ bs_26;
  wire        pairs_26_2 = as_26 & bs_26;
  wire        pairs_27_1 = as_27 ^ bs_27;
  wire        pairs_27_2 = as_27 & bs_27;
  wire        pairs_28_1 = as_28 ^ bs_28;
  wire        pairs_28_2 = as_28 & bs_28;
  wire        pairs_29_1 = as_29 ^ bs_29;
  wire        pairs_29_2 = as_29 & bs_29;
  wire        pairs_30_1 = as_30 ^ bs_30;
  wire        pairs_30_2 = as_30 & bs_30;
  wire        pairs_31_1 = as_31 ^ bs_31;
  wire        pairs_31_2 = as_31 & bs_31;
  wire        tree8Leaf_layer0_0_1 = pairs_7_1 & pairs_6_1;
  wire        tree8Leaf_layer0_0_2 = pairs_7_2 | pairs_7_1 & pairs_6_2;
  wire        tree8Leaf_layer0_1_1 = pairs_5_1 & pairs_4_1;
  wire        tree8Leaf_layer0_1_2 = pairs_5_2 | pairs_5_1 & pairs_4_2;
  wire        tree8Leaf_layer0_2_1 = pairs_3_1 & pairs_2_1;
  wire        tree8Leaf_layer0_2_2 = pairs_3_2 | pairs_3_1 & pairs_2_2;
  wire        tree8Leaf_0_1_1 = pairs_1_1 & pairs_0_1;
  wire        tree8Leaf_0_1_2 = pairs_1_2 | pairs_1_1 & pairs_0_2;
  wire        tree8Leaf_layer1_0_1 = tree8Leaf_layer0_0_1 & tree8Leaf_layer0_1_1;
  wire        tree8Leaf_layer1_0_2 = tree8Leaf_layer0_0_2 | tree8Leaf_layer0_0_1 & tree8Leaf_layer0_1_2;
  wire        tree8Leaf_0_3_1 = tree8Leaf_layer0_2_1 & tree8Leaf_0_1_1;
  wire        tree8Leaf_0_3_2 = tree8Leaf_layer0_2_2 | tree8Leaf_layer0_2_1 & tree8Leaf_0_1_2;
  wire        tree8Leaf_0_2_1 = pairs_2_1 & tree8Leaf_0_1_1;
  wire        tree8Leaf_0_2_2 = pairs_2_2 | pairs_2_1 & tree8Leaf_0_1_2;
  wire        tree8Leaf_0_4_1 = pairs_4_1 & tree8Leaf_0_3_1;
  wire        tree8Leaf_0_4_2 = pairs_4_2 | pairs_4_1 & tree8Leaf_0_3_2;
  wire        tree8Leaf_0_5_1 = tree8Leaf_layer0_1_1 & tree8Leaf_0_3_1;
  wire        tree8Leaf_0_5_2 = tree8Leaf_layer0_1_2 | tree8Leaf_layer0_1_1 & tree8Leaf_0_3_2;
  wire        tree8Leaf_0_6_1 = pairs_6_1 & tree8Leaf_0_5_1;
  wire        tree8Leaf_0_6_2 = pairs_6_2 | pairs_6_1 & tree8Leaf_0_5_2;
  wire        tree8Leaf_0_7_1 = tree8Leaf_layer1_0_1 & tree8Leaf_0_3_1;
  wire        tree8Leaf_0_7_2 = tree8Leaf_layer1_0_2 | tree8Leaf_layer1_0_1 & tree8Leaf_0_3_2;
  wire        tree8Leaf_layer0_0_1_1 = pairs_15_1 & pairs_14_1;
  wire        tree8Leaf_layer0_0_2_1 = pairs_15_2 | pairs_15_1 & pairs_14_2;
  wire        tree8Leaf_layer0_1_1_1 = pairs_13_1 & pairs_12_1;
  wire        tree8Leaf_layer0_1_2_1 = pairs_13_2 | pairs_13_1 & pairs_12_2;
  wire        tree8Leaf_layer0_2_1_1 = pairs_11_1 & pairs_10_1;
  wire        tree8Leaf_layer0_2_2_1 = pairs_11_2 | pairs_11_1 & pairs_10_2;
  wire        tree8Leaf_1_1_1 = pairs_9_1 & pairs_8_1;
  wire        tree8Leaf_1_1_2 = pairs_9_2 | pairs_9_1 & pairs_8_2;
  wire        tree8Leaf_layer1_0_1_1 = tree8Leaf_layer0_0_1_1 & tree8Leaf_layer0_1_1_1;
  wire        tree8Leaf_layer1_0_2_1 = tree8Leaf_layer0_0_2_1 | tree8Leaf_layer0_0_1_1 & tree8Leaf_layer0_1_2_1;
  wire        tree8Leaf_1_3_1 = tree8Leaf_layer0_2_1_1 & tree8Leaf_1_1_1;
  wire        tree8Leaf_1_3_2 = tree8Leaf_layer0_2_2_1 | tree8Leaf_layer0_2_1_1 & tree8Leaf_1_1_2;
  wire        tree8Leaf_1_2_1 = pairs_10_1 & tree8Leaf_1_1_1;
  wire        tree8Leaf_1_2_2 = pairs_10_2 | pairs_10_1 & tree8Leaf_1_1_2;
  wire        tree8Leaf_1_4_1 = pairs_12_1 & tree8Leaf_1_3_1;
  wire        tree8Leaf_1_4_2 = pairs_12_2 | pairs_12_1 & tree8Leaf_1_3_2;
  wire        tree8Leaf_1_5_1 = tree8Leaf_layer0_1_1_1 & tree8Leaf_1_3_1;
  wire        tree8Leaf_1_5_2 = tree8Leaf_layer0_1_2_1 | tree8Leaf_layer0_1_1_1 & tree8Leaf_1_3_2;
  wire        tree8Leaf_1_6_1 = pairs_14_1 & tree8Leaf_1_5_1;
  wire        tree8Leaf_1_6_2 = pairs_14_2 | pairs_14_1 & tree8Leaf_1_5_2;
  wire        tree8Leaf_1_7_1 = tree8Leaf_layer1_0_1_1 & tree8Leaf_1_3_1;
  wire        tree8Leaf_1_7_2 = tree8Leaf_layer1_0_2_1 | tree8Leaf_layer1_0_1_1 & tree8Leaf_1_3_2;
  wire        tree8Leaf_layer0_0_1_2 = pairs_23_1 & pairs_22_1;
  wire        tree8Leaf_layer0_0_2_2 = pairs_23_2 | pairs_23_1 & pairs_22_2;
  wire        tree8Leaf_layer0_1_1_2 = pairs_21_1 & pairs_20_1;
  wire        tree8Leaf_layer0_1_2_2 = pairs_21_2 | pairs_21_1 & pairs_20_2;
  wire        tree8Leaf_layer0_2_1_2 = pairs_19_1 & pairs_18_1;
  wire        tree8Leaf_layer0_2_2_2 = pairs_19_2 | pairs_19_1 & pairs_18_2;
  wire        tree8Leaf_2_1_1 = pairs_17_1 & pairs_16_1;
  wire        tree8Leaf_2_1_2 = pairs_17_2 | pairs_17_1 & pairs_16_2;
  wire        tree8Leaf_layer1_0_1_2 = tree8Leaf_layer0_0_1_2 & tree8Leaf_layer0_1_1_2;
  wire        tree8Leaf_layer1_0_2_2 = tree8Leaf_layer0_0_2_2 | tree8Leaf_layer0_0_1_2 & tree8Leaf_layer0_1_2_2;
  wire        tree8Leaf_2_3_1 = tree8Leaf_layer0_2_1_2 & tree8Leaf_2_1_1;
  wire        tree8Leaf_2_3_2 = tree8Leaf_layer0_2_2_2 | tree8Leaf_layer0_2_1_2 & tree8Leaf_2_1_2;
  wire        tree8Leaf_2_2_1 = pairs_18_1 & tree8Leaf_2_1_1;
  wire        tree8Leaf_2_2_2 = pairs_18_2 | pairs_18_1 & tree8Leaf_2_1_2;
  wire        tree8Leaf_2_4_1 = pairs_20_1 & tree8Leaf_2_3_1;
  wire        tree8Leaf_2_4_2 = pairs_20_2 | pairs_20_1 & tree8Leaf_2_3_2;
  wire        tree8Leaf_2_5_1 = tree8Leaf_layer0_1_1_2 & tree8Leaf_2_3_1;
  wire        tree8Leaf_2_5_2 = tree8Leaf_layer0_1_2_2 | tree8Leaf_layer0_1_1_2 & tree8Leaf_2_3_2;
  wire        tree8Leaf_2_6_1 = pairs_22_1 & tree8Leaf_2_5_1;
  wire        tree8Leaf_2_6_2 = pairs_22_2 | pairs_22_1 & tree8Leaf_2_5_2;
  wire        tree8Leaf_2_7_1 = tree8Leaf_layer1_0_1_2 & tree8Leaf_2_3_1;
  wire        tree8Leaf_2_7_2 = tree8Leaf_layer1_0_2_2 | tree8Leaf_layer1_0_1_2 & tree8Leaf_2_3_2;
  wire        tree8Leaf_layer0_0_1_3 = pairs_31_1 & pairs_30_1;
  wire        tree8Leaf_layer0_0_2_3 = pairs_31_2 | pairs_31_1 & pairs_30_2;
  wire        tree8Leaf_layer0_1_1_3 = pairs_29_1 & pairs_28_1;
  wire        tree8Leaf_layer0_1_2_3 = pairs_29_2 | pairs_29_1 & pairs_28_2;
  wire        tree8Leaf_layer0_2_1_3 = pairs_27_1 & pairs_26_1;
  wire        tree8Leaf_layer0_2_2_3 = pairs_27_2 | pairs_27_1 & pairs_26_2;
  wire        tree8Leaf_3_1_1 = pairs_25_1 & pairs_24_1;
  wire        tree8Leaf_3_1_2 = pairs_25_2 | pairs_25_1 & pairs_24_2;
  wire        tree8Leaf_layer1_0_1_3 = tree8Leaf_layer0_0_1_3 & tree8Leaf_layer0_1_1_3;
  wire        tree8Leaf_layer1_0_2_3 = tree8Leaf_layer0_0_2_3 | tree8Leaf_layer0_0_1_3 & tree8Leaf_layer0_1_2_3;
  wire        tree8Leaf_3_3_1 = tree8Leaf_layer0_2_1_3 & tree8Leaf_3_1_1;
  wire        tree8Leaf_3_3_2 = tree8Leaf_layer0_2_2_3 | tree8Leaf_layer0_2_1_3 & tree8Leaf_3_1_2;
  wire        tree8Leaf_3_2_1 = pairs_26_1 & tree8Leaf_3_1_1;
  wire        tree8Leaf_3_2_2 = pairs_26_2 | pairs_26_1 & tree8Leaf_3_1_2;
  wire        tree8Leaf_3_4_1 = pairs_28_1 & tree8Leaf_3_3_1;
  wire        tree8Leaf_3_4_2 = pairs_28_2 | pairs_28_1 & tree8Leaf_3_3_2;
  wire        tree8Leaf_3_5_1 = tree8Leaf_layer0_1_1_3 & tree8Leaf_3_3_1;
  wire        tree8Leaf_3_5_2 = tree8Leaf_layer0_1_2_3 | tree8Leaf_layer0_1_1_3 & tree8Leaf_3_3_2;
  wire        tree8Leaf_3_6_1 = pairs_30_1 & tree8Leaf_3_5_1;
  wire        tree8Leaf_3_6_2 = pairs_30_2 | pairs_30_1 & tree8Leaf_3_5_2;
  wire        tree8Leaf_3_7_1 = tree8Leaf_layer1_0_1_3 & tree8Leaf_3_3_1;
  wire        tree8Leaf_3_7_2 = tree8Leaf_layer1_0_2_3 | tree8Leaf_layer1_0_1_3 & tree8Leaf_3_3_2;
  wire        tree16Leaf0_8_1 = pairs_8_1 & tree8Leaf_0_7_1;
  wire        tree16Leaf0_8_2 = pairs_8_2 | pairs_8_1 & tree8Leaf_0_7_2;
  wire        tree16Leaf0_9_1 = tree8Leaf_1_1_1 & tree8Leaf_0_7_1;
  wire        tree16Leaf0_9_2 = tree8Leaf_1_1_2 | tree8Leaf_1_1_1 & tree8Leaf_0_7_2;
  wire        tree16Leaf0_10_1 = tree8Leaf_1_2_1 & tree8Leaf_0_7_1;
  wire        tree16Leaf0_10_2 = tree8Leaf_1_2_2 | tree8Leaf_1_2_1 & tree8Leaf_0_7_2;
  wire        tree16Leaf0_11_1 = tree8Leaf_1_3_1 & tree8Leaf_0_7_1;
  wire        tree16Leaf0_11_2 = tree8Leaf_1_3_2 | tree8Leaf_1_3_1 & tree8Leaf_0_7_2;
  wire        tree16Leaf0_12_1 = tree8Leaf_1_4_1 & tree8Leaf_0_7_1;
  wire        tree16Leaf0_12_2 = tree8Leaf_1_4_2 | tree8Leaf_1_4_1 & tree8Leaf_0_7_2;
  wire        tree16Leaf0_13_1 = tree8Leaf_1_5_1 & tree8Leaf_0_7_1;
  wire        tree16Leaf0_13_2 = tree8Leaf_1_5_2 | tree8Leaf_1_5_1 & tree8Leaf_0_7_2;
  wire        tree16Leaf0_14_1 = tree8Leaf_1_6_1 & tree8Leaf_0_7_1;
  wire        tree16Leaf0_14_2 = tree8Leaf_1_6_2 | tree8Leaf_1_6_1 & tree8Leaf_0_7_2;
  wire        tree16Leaf0_15_1 = tree8Leaf_1_7_1 & tree8Leaf_0_7_1;
  wire        tree16Leaf0_15_2 = tree8Leaf_1_7_2 | tree8Leaf_1_7_1 & tree8Leaf_0_7_2;
  wire        tree16Leaf1_8_1 = pairs_24_1 & tree8Leaf_2_7_1;
  wire        tree16Leaf1_8_2 = pairs_24_2 | pairs_24_1 & tree8Leaf_2_7_2;
  wire        tree16Leaf1_9_1 = tree8Leaf_3_1_1 & tree8Leaf_2_7_1;
  wire        tree16Leaf1_9_2 = tree8Leaf_3_1_2 | tree8Leaf_3_1_1 & tree8Leaf_2_7_2;
  wire        tree16Leaf1_10_1 = tree8Leaf_3_2_1 & tree8Leaf_2_7_1;
  wire        tree16Leaf1_10_2 = tree8Leaf_3_2_2 | tree8Leaf_3_2_1 & tree8Leaf_2_7_2;
  wire        tree16Leaf1_11_1 = tree8Leaf_3_3_1 & tree8Leaf_2_7_1;
  wire        tree16Leaf1_11_2 = tree8Leaf_3_3_2 | tree8Leaf_3_3_1 & tree8Leaf_2_7_2;
  wire        tree16Leaf1_12_1 = tree8Leaf_3_4_1 & tree8Leaf_2_7_1;
  wire        tree16Leaf1_12_2 = tree8Leaf_3_4_2 | tree8Leaf_3_4_1 & tree8Leaf_2_7_2;
  wire        tree16Leaf1_13_1 = tree8Leaf_3_5_1 & tree8Leaf_2_7_1;
  wire        tree16Leaf1_13_2 = tree8Leaf_3_5_2 | tree8Leaf_3_5_1 & tree8Leaf_2_7_2;
  wire        tree16Leaf1_14_1 = tree8Leaf_3_6_1 & tree8Leaf_2_7_1;
  wire        tree16Leaf1_14_2 = tree8Leaf_3_6_2 | tree8Leaf_3_6_1 & tree8Leaf_2_7_2;
  wire        tree16Leaf1_15_1 = tree8Leaf_3_7_1 & tree8Leaf_2_7_1;
  wire        tree16Leaf1_15_2 = tree8Leaf_3_7_2 | tree8Leaf_3_7_1 & tree8Leaf_2_7_2;
  wire        tree32_16_1 = pairs_16_1 & tree16Leaf0_15_1;
  wire        tree32_16_2 = pairs_16_2 | pairs_16_1 & tree16Leaf0_15_2;
  wire        tree32_17_1 = tree8Leaf_2_1_1 & tree16Leaf0_15_1;
  wire        tree32_17_2 = tree8Leaf_2_1_2 | tree8Leaf_2_1_1 & tree16Leaf0_15_2;
  wire        tree32_18_1 = tree8Leaf_2_2_1 & tree16Leaf0_15_1;
  wire        tree32_18_2 = tree8Leaf_2_2_2 | tree8Leaf_2_2_1 & tree16Leaf0_15_2;
  wire        tree32_19_1 = tree8Leaf_2_3_1 & tree16Leaf0_15_1;
  wire        tree32_19_2 = tree8Leaf_2_3_2 | tree8Leaf_2_3_1 & tree16Leaf0_15_2;
  wire        tree32_20_1 = tree8Leaf_2_4_1 & tree16Leaf0_15_1;
  wire        tree32_20_2 = tree8Leaf_2_4_2 | tree8Leaf_2_4_1 & tree16Leaf0_15_2;
  wire        tree32_21_1 = tree8Leaf_2_5_1 & tree16Leaf0_15_1;
  wire        tree32_21_2 = tree8Leaf_2_5_2 | tree8Leaf_2_5_1 & tree16Leaf0_15_2;
  wire        tree32_22_1 = tree8Leaf_2_6_1 & tree16Leaf0_15_1;
  wire        tree32_22_2 = tree8Leaf_2_6_2 | tree8Leaf_2_6_1 & tree16Leaf0_15_2;
  wire        tree32_23_1 = tree8Leaf_2_7_1 & tree16Leaf0_15_1;
  wire        tree32_23_2 = tree8Leaf_2_7_2 | tree8Leaf_2_7_1 & tree16Leaf0_15_2;
  wire        tree32_24_1 = tree16Leaf1_8_1 & tree16Leaf0_15_1;
  wire        tree32_24_2 = tree16Leaf1_8_2 | tree16Leaf1_8_1 & tree16Leaf0_15_2;
  wire        tree32_25_1 = tree16Leaf1_9_1 & tree16Leaf0_15_1;
  wire        tree32_25_2 = tree16Leaf1_9_2 | tree16Leaf1_9_1 & tree16Leaf0_15_2;
  wire        tree32_26_1 = tree16Leaf1_10_1 & tree16Leaf0_15_1;
  wire        tree32_26_2 = tree16Leaf1_10_2 | tree16Leaf1_10_1 & tree16Leaf0_15_2;
  wire        tree32_27_1 = tree16Leaf1_11_1 & tree16Leaf0_15_1;
  wire        tree32_27_2 = tree16Leaf1_11_2 | tree16Leaf1_11_1 & tree16Leaf0_15_2;
  wire        tree32_28_1 = tree16Leaf1_12_1 & tree16Leaf0_15_1;
  wire        tree32_28_2 = tree16Leaf1_12_2 | tree16Leaf1_12_1 & tree16Leaf0_15_2;
  wire        tree32_29_1 = tree16Leaf1_13_1 & tree16Leaf0_15_1;
  wire        tree32_29_2 = tree16Leaf1_13_2 | tree16Leaf1_13_1 & tree16Leaf0_15_2;
  wire        tree32_30_1 = tree16Leaf1_14_1 & tree16Leaf0_15_1;
  wire        tree32_30_2 = tree16Leaf1_14_2 | tree16Leaf1_14_1 & tree16Leaf0_15_2;
  wire        tree32_31_1 = tree16Leaf1_15_1 & tree16Leaf0_15_1;
  wire        tree32_31_2 = tree16Leaf1_15_2 | tree16Leaf1_15_1 & tree16Leaf0_15_2;
  wire [1:0]  _GEN = {tree8Leaf_0_1_1, pairs_0_1};
  wire [1:0]  tree8P_lo_lo_lo_lo;
  assign tree8P_lo_lo_lo_lo = _GEN;
  wire [1:0]  tree16P_lo_lo_lo_lo;
  assign tree16P_lo_lo_lo_lo = _GEN;
  wire [1:0]  tree32P_lo_lo_lo_lo;
  assign tree32P_lo_lo_lo_lo = _GEN;
  wire [1:0]  _GEN_0 = {tree8Leaf_0_3_1, tree8Leaf_0_2_1};
  wire [1:0]  tree8P_lo_lo_lo_hi;
  assign tree8P_lo_lo_lo_hi = _GEN_0;
  wire [1:0]  tree16P_lo_lo_lo_hi;
  assign tree16P_lo_lo_lo_hi = _GEN_0;
  wire [1:0]  tree32P_lo_lo_lo_hi;
  assign tree32P_lo_lo_lo_hi = _GEN_0;
  wire [3:0]  tree8P_lo_lo_lo = {tree8P_lo_lo_lo_hi, tree8P_lo_lo_lo_lo};
  wire [1:0]  _GEN_1 = {tree8Leaf_0_5_1, tree8Leaf_0_4_1};
  wire [1:0]  tree8P_lo_lo_hi_lo;
  assign tree8P_lo_lo_hi_lo = _GEN_1;
  wire [1:0]  tree16P_lo_lo_hi_lo;
  assign tree16P_lo_lo_hi_lo = _GEN_1;
  wire [1:0]  tree32P_lo_lo_hi_lo;
  assign tree32P_lo_lo_hi_lo = _GEN_1;
  wire [1:0]  _GEN_2 = {tree8Leaf_0_7_1, tree8Leaf_0_6_1};
  wire [1:0]  tree8P_lo_lo_hi_hi;
  assign tree8P_lo_lo_hi_hi = _GEN_2;
  wire [1:0]  tree16P_lo_lo_hi_hi;
  assign tree16P_lo_lo_hi_hi = _GEN_2;
  wire [1:0]  tree32P_lo_lo_hi_hi;
  assign tree32P_lo_lo_hi_hi = _GEN_2;
  wire [3:0]  tree8P_lo_lo_hi = {tree8P_lo_lo_hi_hi, tree8P_lo_lo_hi_lo};
  wire [7:0]  tree8P_lo_lo = {tree8P_lo_lo_hi, tree8P_lo_lo_lo};
  wire [1:0]  tree8P_lo_hi_lo_lo = {tree8Leaf_1_1_1, pairs_8_1};
  wire [1:0]  tree8P_lo_hi_lo_hi = {tree8Leaf_1_3_1, tree8Leaf_1_2_1};
  wire [3:0]  tree8P_lo_hi_lo = {tree8P_lo_hi_lo_hi, tree8P_lo_hi_lo_lo};
  wire [1:0]  tree8P_lo_hi_hi_lo = {tree8Leaf_1_5_1, tree8Leaf_1_4_1};
  wire [1:0]  tree8P_lo_hi_hi_hi = {tree8Leaf_1_7_1, tree8Leaf_1_6_1};
  wire [3:0]  tree8P_lo_hi_hi = {tree8P_lo_hi_hi_hi, tree8P_lo_hi_hi_lo};
  wire [7:0]  tree8P_lo_hi = {tree8P_lo_hi_hi, tree8P_lo_hi_lo};
  wire [15:0] tree8P_lo = {tree8P_lo_hi, tree8P_lo_lo};
  wire [1:0]  _GEN_3 = {tree8Leaf_2_1_1, pairs_16_1};
  wire [1:0]  tree8P_hi_lo_lo_lo;
  assign tree8P_hi_lo_lo_lo = _GEN_3;
  wire [1:0]  tree16P_hi_lo_lo_lo;
  assign tree16P_hi_lo_lo_lo = _GEN_3;
  wire [1:0]  _GEN_4 = {tree8Leaf_2_3_1, tree8Leaf_2_2_1};
  wire [1:0]  tree8P_hi_lo_lo_hi;
  assign tree8P_hi_lo_lo_hi = _GEN_4;
  wire [1:0]  tree16P_hi_lo_lo_hi;
  assign tree16P_hi_lo_lo_hi = _GEN_4;
  wire [3:0]  tree8P_hi_lo_lo = {tree8P_hi_lo_lo_hi, tree8P_hi_lo_lo_lo};
  wire [1:0]  _GEN_5 = {tree8Leaf_2_5_1, tree8Leaf_2_4_1};
  wire [1:0]  tree8P_hi_lo_hi_lo;
  assign tree8P_hi_lo_hi_lo = _GEN_5;
  wire [1:0]  tree16P_hi_lo_hi_lo;
  assign tree16P_hi_lo_hi_lo = _GEN_5;
  wire [1:0]  _GEN_6 = {tree8Leaf_2_7_1, tree8Leaf_2_6_1};
  wire [1:0]  tree8P_hi_lo_hi_hi;
  assign tree8P_hi_lo_hi_hi = _GEN_6;
  wire [1:0]  tree16P_hi_lo_hi_hi;
  assign tree16P_hi_lo_hi_hi = _GEN_6;
  wire [3:0]  tree8P_hi_lo_hi = {tree8P_hi_lo_hi_hi, tree8P_hi_lo_hi_lo};
  wire [7:0]  tree8P_hi_lo = {tree8P_hi_lo_hi, tree8P_hi_lo_lo};
  wire [1:0]  tree8P_hi_hi_lo_lo = {tree8Leaf_3_1_1, pairs_24_1};
  wire [1:0]  tree8P_hi_hi_lo_hi = {tree8Leaf_3_3_1, tree8Leaf_3_2_1};
  wire [3:0]  tree8P_hi_hi_lo = {tree8P_hi_hi_lo_hi, tree8P_hi_hi_lo_lo};
  wire [1:0]  tree8P_hi_hi_hi_lo = {tree8Leaf_3_5_1, tree8Leaf_3_4_1};
  wire [1:0]  tree8P_hi_hi_hi_hi = {tree8Leaf_3_7_1, tree8Leaf_3_6_1};
  wire [3:0]  tree8P_hi_hi_hi = {tree8P_hi_hi_hi_hi, tree8P_hi_hi_hi_lo};
  wire [7:0]  tree8P_hi_hi = {tree8P_hi_hi_hi, tree8P_hi_hi_lo};
  wire [15:0] tree8P_hi = {tree8P_hi_hi, tree8P_hi_lo};
  wire [31:0] tree8P = {tree8P_hi, tree8P_lo};
  wire [1:0]  _GEN_7 = {tree8Leaf_0_1_2, pairs_0_2};
  wire [1:0]  tree8G_lo_lo_lo_lo;
  assign tree8G_lo_lo_lo_lo = _GEN_7;
  wire [1:0]  tree16G_lo_lo_lo_lo;
  assign tree16G_lo_lo_lo_lo = _GEN_7;
  wire [1:0]  tree32G_lo_lo_lo_lo;
  assign tree32G_lo_lo_lo_lo = _GEN_7;
  wire [1:0]  _GEN_8 = {tree8Leaf_0_3_2, tree8Leaf_0_2_2};
  wire [1:0]  tree8G_lo_lo_lo_hi;
  assign tree8G_lo_lo_lo_hi = _GEN_8;
  wire [1:0]  tree16G_lo_lo_lo_hi;
  assign tree16G_lo_lo_lo_hi = _GEN_8;
  wire [1:0]  tree32G_lo_lo_lo_hi;
  assign tree32G_lo_lo_lo_hi = _GEN_8;
  wire [3:0]  tree8G_lo_lo_lo = {tree8G_lo_lo_lo_hi, tree8G_lo_lo_lo_lo};
  wire [1:0]  _GEN_9 = {tree8Leaf_0_5_2, tree8Leaf_0_4_2};
  wire [1:0]  tree8G_lo_lo_hi_lo;
  assign tree8G_lo_lo_hi_lo = _GEN_9;
  wire [1:0]  tree16G_lo_lo_hi_lo;
  assign tree16G_lo_lo_hi_lo = _GEN_9;
  wire [1:0]  tree32G_lo_lo_hi_lo;
  assign tree32G_lo_lo_hi_lo = _GEN_9;
  wire [1:0]  _GEN_10 = {tree8Leaf_0_7_2, tree8Leaf_0_6_2};
  wire [1:0]  tree8G_lo_lo_hi_hi;
  assign tree8G_lo_lo_hi_hi = _GEN_10;
  wire [1:0]  tree16G_lo_lo_hi_hi;
  assign tree16G_lo_lo_hi_hi = _GEN_10;
  wire [1:0]  tree32G_lo_lo_hi_hi;
  assign tree32G_lo_lo_hi_hi = _GEN_10;
  wire [3:0]  tree8G_lo_lo_hi = {tree8G_lo_lo_hi_hi, tree8G_lo_lo_hi_lo};
  wire [7:0]  tree8G_lo_lo = {tree8G_lo_lo_hi, tree8G_lo_lo_lo};
  wire [1:0]  tree8G_lo_hi_lo_lo = {tree8Leaf_1_1_2, pairs_8_2};
  wire [1:0]  tree8G_lo_hi_lo_hi = {tree8Leaf_1_3_2, tree8Leaf_1_2_2};
  wire [3:0]  tree8G_lo_hi_lo = {tree8G_lo_hi_lo_hi, tree8G_lo_hi_lo_lo};
  wire [1:0]  tree8G_lo_hi_hi_lo = {tree8Leaf_1_5_2, tree8Leaf_1_4_2};
  wire [1:0]  tree8G_lo_hi_hi_hi = {tree8Leaf_1_7_2, tree8Leaf_1_6_2};
  wire [3:0]  tree8G_lo_hi_hi = {tree8G_lo_hi_hi_hi, tree8G_lo_hi_hi_lo};
  wire [7:0]  tree8G_lo_hi = {tree8G_lo_hi_hi, tree8G_lo_hi_lo};
  wire [15:0] tree8G_lo = {tree8G_lo_hi, tree8G_lo_lo};
  wire [1:0]  _GEN_11 = {tree8Leaf_2_1_2, pairs_16_2};
  wire [1:0]  tree8G_hi_lo_lo_lo;
  assign tree8G_hi_lo_lo_lo = _GEN_11;
  wire [1:0]  tree16G_hi_lo_lo_lo;
  assign tree16G_hi_lo_lo_lo = _GEN_11;
  wire [1:0]  _GEN_12 = {tree8Leaf_2_3_2, tree8Leaf_2_2_2};
  wire [1:0]  tree8G_hi_lo_lo_hi;
  assign tree8G_hi_lo_lo_hi = _GEN_12;
  wire [1:0]  tree16G_hi_lo_lo_hi;
  assign tree16G_hi_lo_lo_hi = _GEN_12;
  wire [3:0]  tree8G_hi_lo_lo = {tree8G_hi_lo_lo_hi, tree8G_hi_lo_lo_lo};
  wire [1:0]  _GEN_13 = {tree8Leaf_2_5_2, tree8Leaf_2_4_2};
  wire [1:0]  tree8G_hi_lo_hi_lo;
  assign tree8G_hi_lo_hi_lo = _GEN_13;
  wire [1:0]  tree16G_hi_lo_hi_lo;
  assign tree16G_hi_lo_hi_lo = _GEN_13;
  wire [1:0]  _GEN_14 = {tree8Leaf_2_7_2, tree8Leaf_2_6_2};
  wire [1:0]  tree8G_hi_lo_hi_hi;
  assign tree8G_hi_lo_hi_hi = _GEN_14;
  wire [1:0]  tree16G_hi_lo_hi_hi;
  assign tree16G_hi_lo_hi_hi = _GEN_14;
  wire [3:0]  tree8G_hi_lo_hi = {tree8G_hi_lo_hi_hi, tree8G_hi_lo_hi_lo};
  wire [7:0]  tree8G_hi_lo = {tree8G_hi_lo_hi, tree8G_hi_lo_lo};
  wire [1:0]  tree8G_hi_hi_lo_lo = {tree8Leaf_3_1_2, pairs_24_2};
  wire [1:0]  tree8G_hi_hi_lo_hi = {tree8Leaf_3_3_2, tree8Leaf_3_2_2};
  wire [3:0]  tree8G_hi_hi_lo = {tree8G_hi_hi_lo_hi, tree8G_hi_hi_lo_lo};
  wire [1:0]  tree8G_hi_hi_hi_lo = {tree8Leaf_3_5_2, tree8Leaf_3_4_2};
  wire [1:0]  tree8G_hi_hi_hi_hi = {tree8Leaf_3_7_2, tree8Leaf_3_6_2};
  wire [3:0]  tree8G_hi_hi_hi = {tree8G_hi_hi_hi_hi, tree8G_hi_hi_hi_lo};
  wire [7:0]  tree8G_hi_hi = {tree8G_hi_hi_hi, tree8G_hi_hi_lo};
  wire [15:0] tree8G_hi = {tree8G_hi_hi, tree8G_hi_lo};
  wire [31:0] tree8G = {tree8G_hi, tree8G_lo};
  wire [3:0]  tree16P_lo_lo_lo = {tree16P_lo_lo_lo_hi, tree16P_lo_lo_lo_lo};
  wire [3:0]  tree16P_lo_lo_hi = {tree16P_lo_lo_hi_hi, tree16P_lo_lo_hi_lo};
  wire [7:0]  tree16P_lo_lo = {tree16P_lo_lo_hi, tree16P_lo_lo_lo};
  wire [1:0]  _GEN_15 = {tree16Leaf0_9_1, tree16Leaf0_8_1};
  wire [1:0]  tree16P_lo_hi_lo_lo;
  assign tree16P_lo_hi_lo_lo = _GEN_15;
  wire [1:0]  tree32P_lo_hi_lo_lo;
  assign tree32P_lo_hi_lo_lo = _GEN_15;
  wire [1:0]  _GEN_16 = {tree16Leaf0_11_1, tree16Leaf0_10_1};
  wire [1:0]  tree16P_lo_hi_lo_hi;
  assign tree16P_lo_hi_lo_hi = _GEN_16;
  wire [1:0]  tree32P_lo_hi_lo_hi;
  assign tree32P_lo_hi_lo_hi = _GEN_16;
  wire [3:0]  tree16P_lo_hi_lo = {tree16P_lo_hi_lo_hi, tree16P_lo_hi_lo_lo};
  wire [1:0]  _GEN_17 = {tree16Leaf0_13_1, tree16Leaf0_12_1};
  wire [1:0]  tree16P_lo_hi_hi_lo;
  assign tree16P_lo_hi_hi_lo = _GEN_17;
  wire [1:0]  tree32P_lo_hi_hi_lo;
  assign tree32P_lo_hi_hi_lo = _GEN_17;
  wire [1:0]  _GEN_18 = {tree16Leaf0_15_1, tree16Leaf0_14_1};
  wire [1:0]  tree16P_lo_hi_hi_hi;
  assign tree16P_lo_hi_hi_hi = _GEN_18;
  wire [1:0]  tree32P_lo_hi_hi_hi;
  assign tree32P_lo_hi_hi_hi = _GEN_18;
  wire [3:0]  tree16P_lo_hi_hi = {tree16P_lo_hi_hi_hi, tree16P_lo_hi_hi_lo};
  wire [7:0]  tree16P_lo_hi = {tree16P_lo_hi_hi, tree16P_lo_hi_lo};
  wire [15:0] tree16P_lo = {tree16P_lo_hi, tree16P_lo_lo};
  wire [3:0]  tree16P_hi_lo_lo = {tree16P_hi_lo_lo_hi, tree16P_hi_lo_lo_lo};
  wire [3:0]  tree16P_hi_lo_hi = {tree16P_hi_lo_hi_hi, tree16P_hi_lo_hi_lo};
  wire [7:0]  tree16P_hi_lo = {tree16P_hi_lo_hi, tree16P_hi_lo_lo};
  wire [1:0]  tree16P_hi_hi_lo_lo = {tree16Leaf1_9_1, tree16Leaf1_8_1};
  wire [1:0]  tree16P_hi_hi_lo_hi = {tree16Leaf1_11_1, tree16Leaf1_10_1};
  wire [3:0]  tree16P_hi_hi_lo = {tree16P_hi_hi_lo_hi, tree16P_hi_hi_lo_lo};
  wire [1:0]  tree16P_hi_hi_hi_lo = {tree16Leaf1_13_1, tree16Leaf1_12_1};
  wire [1:0]  tree16P_hi_hi_hi_hi = {tree16Leaf1_15_1, tree16Leaf1_14_1};
  wire [3:0]  tree16P_hi_hi_hi = {tree16P_hi_hi_hi_hi, tree16P_hi_hi_hi_lo};
  wire [7:0]  tree16P_hi_hi = {tree16P_hi_hi_hi, tree16P_hi_hi_lo};
  wire [15:0] tree16P_hi = {tree16P_hi_hi, tree16P_hi_lo};
  wire [31:0] tree16P = {tree16P_hi, tree16P_lo};
  wire [3:0]  tree16G_lo_lo_lo = {tree16G_lo_lo_lo_hi, tree16G_lo_lo_lo_lo};
  wire [3:0]  tree16G_lo_lo_hi = {tree16G_lo_lo_hi_hi, tree16G_lo_lo_hi_lo};
  wire [7:0]  tree16G_lo_lo = {tree16G_lo_lo_hi, tree16G_lo_lo_lo};
  wire [1:0]  _GEN_19 = {tree16Leaf0_9_2, tree16Leaf0_8_2};
  wire [1:0]  tree16G_lo_hi_lo_lo;
  assign tree16G_lo_hi_lo_lo = _GEN_19;
  wire [1:0]  tree32G_lo_hi_lo_lo;
  assign tree32G_lo_hi_lo_lo = _GEN_19;
  wire [1:0]  _GEN_20 = {tree16Leaf0_11_2, tree16Leaf0_10_2};
  wire [1:0]  tree16G_lo_hi_lo_hi;
  assign tree16G_lo_hi_lo_hi = _GEN_20;
  wire [1:0]  tree32G_lo_hi_lo_hi;
  assign tree32G_lo_hi_lo_hi = _GEN_20;
  wire [3:0]  tree16G_lo_hi_lo = {tree16G_lo_hi_lo_hi, tree16G_lo_hi_lo_lo};
  wire [1:0]  _GEN_21 = {tree16Leaf0_13_2, tree16Leaf0_12_2};
  wire [1:0]  tree16G_lo_hi_hi_lo;
  assign tree16G_lo_hi_hi_lo = _GEN_21;
  wire [1:0]  tree32G_lo_hi_hi_lo;
  assign tree32G_lo_hi_hi_lo = _GEN_21;
  wire [1:0]  _GEN_22 = {tree16Leaf0_15_2, tree16Leaf0_14_2};
  wire [1:0]  tree16G_lo_hi_hi_hi;
  assign tree16G_lo_hi_hi_hi = _GEN_22;
  wire [1:0]  tree32G_lo_hi_hi_hi;
  assign tree32G_lo_hi_hi_hi = _GEN_22;
  wire [3:0]  tree16G_lo_hi_hi = {tree16G_lo_hi_hi_hi, tree16G_lo_hi_hi_lo};
  wire [7:0]  tree16G_lo_hi = {tree16G_lo_hi_hi, tree16G_lo_hi_lo};
  wire [15:0] tree16G_lo = {tree16G_lo_hi, tree16G_lo_lo};
  wire [3:0]  tree16G_hi_lo_lo = {tree16G_hi_lo_lo_hi, tree16G_hi_lo_lo_lo};
  wire [3:0]  tree16G_hi_lo_hi = {tree16G_hi_lo_hi_hi, tree16G_hi_lo_hi_lo};
  wire [7:0]  tree16G_hi_lo = {tree16G_hi_lo_hi, tree16G_hi_lo_lo};
  wire [1:0]  tree16G_hi_hi_lo_lo = {tree16Leaf1_9_2, tree16Leaf1_8_2};
  wire [1:0]  tree16G_hi_hi_lo_hi = {tree16Leaf1_11_2, tree16Leaf1_10_2};
  wire [3:0]  tree16G_hi_hi_lo = {tree16G_hi_hi_lo_hi, tree16G_hi_hi_lo_lo};
  wire [1:0]  tree16G_hi_hi_hi_lo = {tree16Leaf1_13_2, tree16Leaf1_12_2};
  wire [1:0]  tree16G_hi_hi_hi_hi = {tree16Leaf1_15_2, tree16Leaf1_14_2};
  wire [3:0]  tree16G_hi_hi_hi = {tree16G_hi_hi_hi_hi, tree16G_hi_hi_hi_lo};
  wire [7:0]  tree16G_hi_hi = {tree16G_hi_hi_hi, tree16G_hi_hi_lo};
  wire [15:0] tree16G_hi = {tree16G_hi_hi, tree16G_hi_lo};
  wire [31:0] tree16G = {tree16G_hi, tree16G_lo};
  wire [3:0]  tree32P_lo_lo_lo = {tree32P_lo_lo_lo_hi, tree32P_lo_lo_lo_lo};
  wire [3:0]  tree32P_lo_lo_hi = {tree32P_lo_lo_hi_hi, tree32P_lo_lo_hi_lo};
  wire [7:0]  tree32P_lo_lo = {tree32P_lo_lo_hi, tree32P_lo_lo_lo};
  wire [3:0]  tree32P_lo_hi_lo = {tree32P_lo_hi_lo_hi, tree32P_lo_hi_lo_lo};
  wire [3:0]  tree32P_lo_hi_hi = {tree32P_lo_hi_hi_hi, tree32P_lo_hi_hi_lo};
  wire [7:0]  tree32P_lo_hi = {tree32P_lo_hi_hi, tree32P_lo_hi_lo};
  wire [15:0] tree32P_lo = {tree32P_lo_hi, tree32P_lo_lo};
  wire [1:0]  tree32P_hi_lo_lo_lo = {tree32_17_1, tree32_16_1};
  wire [1:0]  tree32P_hi_lo_lo_hi = {tree32_19_1, tree32_18_1};
  wire [3:0]  tree32P_hi_lo_lo = {tree32P_hi_lo_lo_hi, tree32P_hi_lo_lo_lo};
  wire [1:0]  tree32P_hi_lo_hi_lo = {tree32_21_1, tree32_20_1};
  wire [1:0]  tree32P_hi_lo_hi_hi = {tree32_23_1, tree32_22_1};
  wire [3:0]  tree32P_hi_lo_hi = {tree32P_hi_lo_hi_hi, tree32P_hi_lo_hi_lo};
  wire [7:0]  tree32P_hi_lo = {tree32P_hi_lo_hi, tree32P_hi_lo_lo};
  wire [1:0]  tree32P_hi_hi_lo_lo = {tree32_25_1, tree32_24_1};
  wire [1:0]  tree32P_hi_hi_lo_hi = {tree32_27_1, tree32_26_1};
  wire [3:0]  tree32P_hi_hi_lo = {tree32P_hi_hi_lo_hi, tree32P_hi_hi_lo_lo};
  wire [1:0]  tree32P_hi_hi_hi_lo = {tree32_29_1, tree32_28_1};
  wire [1:0]  tree32P_hi_hi_hi_hi = {tree32_31_1, tree32_30_1};
  wire [3:0]  tree32P_hi_hi_hi = {tree32P_hi_hi_hi_hi, tree32P_hi_hi_hi_lo};
  wire [7:0]  tree32P_hi_hi = {tree32P_hi_hi_hi, tree32P_hi_hi_lo};
  wire [15:0] tree32P_hi = {tree32P_hi_hi, tree32P_hi_lo};
  wire [31:0] tree32P = {tree32P_hi, tree32P_lo};
  wire [3:0]  tree32G_lo_lo_lo = {tree32G_lo_lo_lo_hi, tree32G_lo_lo_lo_lo};
  wire [3:0]  tree32G_lo_lo_hi = {tree32G_lo_lo_hi_hi, tree32G_lo_lo_hi_lo};
  wire [7:0]  tree32G_lo_lo = {tree32G_lo_lo_hi, tree32G_lo_lo_lo};
  wire [3:0]  tree32G_lo_hi_lo = {tree32G_lo_hi_lo_hi, tree32G_lo_hi_lo_lo};
  wire [3:0]  tree32G_lo_hi_hi = {tree32G_lo_hi_hi_hi, tree32G_lo_hi_hi_lo};
  wire [7:0]  tree32G_lo_hi = {tree32G_lo_hi_hi, tree32G_lo_hi_lo};
  wire [15:0] tree32G_lo = {tree32G_lo_hi, tree32G_lo_lo};
  wire [1:0]  tree32G_hi_lo_lo_lo = {tree32_17_2, tree32_16_2};
  wire [1:0]  tree32G_hi_lo_lo_hi = {tree32_19_2, tree32_18_2};
  wire [3:0]  tree32G_hi_lo_lo = {tree32G_hi_lo_lo_hi, tree32G_hi_lo_lo_lo};
  wire [1:0]  tree32G_hi_lo_hi_lo = {tree32_21_2, tree32_20_2};
  wire [1:0]  tree32G_hi_lo_hi_hi = {tree32_23_2, tree32_22_2};
  wire [3:0]  tree32G_hi_lo_hi = {tree32G_hi_lo_hi_hi, tree32G_hi_lo_hi_lo};
  wire [7:0]  tree32G_hi_lo = {tree32G_hi_lo_hi, tree32G_hi_lo_lo};
  wire [1:0]  tree32G_hi_hi_lo_lo = {tree32_25_2, tree32_24_2};
  wire [1:0]  tree32G_hi_hi_lo_hi = {tree32_27_2, tree32_26_2};
  wire [3:0]  tree32G_hi_hi_lo = {tree32G_hi_hi_lo_hi, tree32G_hi_hi_lo_lo};
  wire [1:0]  tree32G_hi_hi_hi_lo = {tree32_29_2, tree32_28_2};
  wire [1:0]  tree32G_hi_hi_hi_hi = {tree32_31_2, tree32_30_2};
  wire [3:0]  tree32G_hi_hi_hi = {tree32G_hi_hi_hi_hi, tree32G_hi_hi_hi_lo};
  wire [7:0]  tree32G_hi_hi = {tree32G_hi_hi_hi, tree32G_hi_hi_lo};
  wire [15:0] tree32G_hi = {tree32G_hi_hi, tree32G_hi_lo};
  wire [31:0] tree32G = {tree32G_hi, tree32G_lo};
  wire [31:0] treeP = (sew[0] ? tree8P : 32'h0) | (sew[1] ? tree16P : 32'h0) | (sew[2] ? tree32P : 32'h0);
  wire [31:0] treeG = (sew[0] ? tree8G : 32'h0) | (sew[1] ? tree16G : 32'h0) | (sew[2] ? tree32G : 32'h0);
  wire        tree_0_1 = treeP[0];
  wire        tree_1_1 = treeP[1];
  wire        tree_2_1 = treeP[2];
  wire        tree_3_1 = treeP[3];
  wire        tree_4_1 = treeP[4];
  wire        tree_5_1 = treeP[5];
  wire        tree_6_1 = treeP[6];
  wire        tree_7_1 = treeP[7];
  wire        tree_8_1 = treeP[8];
  wire        tree_9_1 = treeP[9];
  wire        tree_10_1 = treeP[10];
  wire        tree_11_1 = treeP[11];
  wire        tree_12_1 = treeP[12];
  wire        tree_13_1 = treeP[13];
  wire        tree_14_1 = treeP[14];
  wire        tree_15_1 = treeP[15];
  wire        tree_16_1 = treeP[16];
  wire        tree_17_1 = treeP[17];
  wire        tree_18_1 = treeP[18];
  wire        tree_19_1 = treeP[19];
  wire        tree_20_1 = treeP[20];
  wire        tree_21_1 = treeP[21];
  wire        tree_22_1 = treeP[22];
  wire        tree_23_1 = treeP[23];
  wire        tree_24_1 = treeP[24];
  wire        tree_25_1 = treeP[25];
  wire        tree_26_1 = treeP[26];
  wire        tree_27_1 = treeP[27];
  wire        tree_28_1 = treeP[28];
  wire        tree_29_1 = treeP[29];
  wire        tree_30_1 = treeP[30];
  wire        tree_31_1 = treeP[31];
  wire        tree_0_2 = treeG[0];
  wire        tree_1_2 = treeG[1];
  wire        tree_2_2 = treeG[2];
  wire        tree_3_2 = treeG[3];
  wire        tree_4_2 = treeG[4];
  wire        tree_5_2 = treeG[5];
  wire        tree_6_2 = treeG[6];
  wire        tree_7_2 = treeG[7];
  wire        tree_8_2 = treeG[8];
  wire        tree_9_2 = treeG[9];
  wire        tree_10_2 = treeG[10];
  wire        tree_11_2 = treeG[11];
  wire        tree_12_2 = treeG[12];
  wire        tree_13_2 = treeG[13];
  wire        tree_14_2 = treeG[14];
  wire        tree_15_2 = treeG[15];
  wire        tree_16_2 = treeG[16];
  wire        tree_17_2 = treeG[17];
  wire        tree_18_2 = treeG[18];
  wire        tree_19_2 = treeG[19];
  wire        tree_20_2 = treeG[20];
  wire        tree_21_2 = treeG[21];
  wire        tree_22_2 = treeG[22];
  wire        tree_23_2 = treeG[23];
  wire        tree_24_2 = treeG[24];
  wire        tree_25_2 = treeG[25];
  wire        tree_26_2 = treeG[26];
  wire        tree_27_2 = treeG[27];
  wire        tree_28_2 = treeG[28];
  wire        tree_29_2 = treeG[29];
  wire        tree_30_2 = treeG[30];
  wire        tree_31_2 = treeG[31];
  wire [1:0]  carryResult_cbank_lo_lo = {tree_1_2 | tree_1_1 & cin[0], tree_0_2 | tree_0_1 & cin[0]};
  wire [1:0]  carryResult_cbank_lo_hi = {tree_3_2 | tree_3_1 & cin[0], tree_2_2 | tree_2_1 & cin[0]};
  wire [3:0]  carryResult_cbank_lo = {carryResult_cbank_lo_hi, carryResult_cbank_lo_lo};
  wire [1:0]  carryResult_cbank_hi_lo = {tree_5_2 | tree_5_1 & cin[0], tree_4_2 | tree_4_1 & cin[0]};
  wire [1:0]  carryResult_cbank_hi_hi = {tree_7_2 | tree_7_1 & cin[0], tree_6_2 | tree_6_1 & cin[0]};
  wire [3:0]  carryResult_cbank_hi = {carryResult_cbank_hi_hi, carryResult_cbank_hi_lo};
  wire [7:0]  carryResult_cbank_0 = {carryResult_cbank_hi, carryResult_cbank_lo};
  wire [1:0]  carryResult_cbank_lo_lo_1 = {tree_9_2 | tree_9_1 & cin[1], tree_8_2 | tree_8_1 & cin[1]};
  wire [1:0]  carryResult_cbank_lo_hi_1 = {tree_11_2 | tree_11_1 & cin[1], tree_10_2 | tree_10_1 & cin[1]};
  wire [3:0]  carryResult_cbank_lo_1 = {carryResult_cbank_lo_hi_1, carryResult_cbank_lo_lo_1};
  wire [1:0]  carryResult_cbank_hi_lo_1 = {tree_13_2 | tree_13_1 & cin[1], tree_12_2 | tree_12_1 & cin[1]};
  wire [1:0]  carryResult_cbank_hi_hi_1 = {tree_15_2 | tree_15_1 & cin[1], tree_14_2 | tree_14_1 & cin[1]};
  wire [3:0]  carryResult_cbank_hi_1 = {carryResult_cbank_hi_hi_1, carryResult_cbank_hi_lo_1};
  wire [7:0]  carryResult_cbank_1 = {carryResult_cbank_hi_1, carryResult_cbank_lo_1};
  wire [1:0]  carryResult_cbank_lo_lo_2 = {tree_17_2 | tree_17_1 & cin[2], tree_16_2 | tree_16_1 & cin[2]};
  wire [1:0]  carryResult_cbank_lo_hi_2 = {tree_19_2 | tree_19_1 & cin[2], tree_18_2 | tree_18_1 & cin[2]};
  wire [3:0]  carryResult_cbank_lo_2 = {carryResult_cbank_lo_hi_2, carryResult_cbank_lo_lo_2};
  wire [1:0]  carryResult_cbank_hi_lo_2 = {tree_21_2 | tree_21_1 & cin[2], tree_20_2 | tree_20_1 & cin[2]};
  wire [1:0]  carryResult_cbank_hi_hi_2 = {tree_23_2 | tree_23_1 & cin[2], tree_22_2 | tree_22_1 & cin[2]};
  wire [3:0]  carryResult_cbank_hi_2 = {carryResult_cbank_hi_hi_2, carryResult_cbank_hi_lo_2};
  wire [7:0]  carryResult_cbank_2 = {carryResult_cbank_hi_2, carryResult_cbank_lo_2};
  wire [1:0]  carryResult_cbank_lo_lo_3 = {tree_25_2 | tree_25_1 & cin[3], tree_24_2 | tree_24_1 & cin[3]};
  wire [1:0]  carryResult_cbank_lo_hi_3 = {tree_27_2 | tree_27_1 & cin[3], tree_26_2 | tree_26_1 & cin[3]};
  wire [3:0]  carryResult_cbank_lo_3 = {carryResult_cbank_lo_hi_3, carryResult_cbank_lo_lo_3};
  wire [1:0]  carryResult_cbank_hi_lo_3 = {tree_29_2 | tree_29_1 & cin[3], tree_28_2 | tree_28_1 & cin[3]};
  wire [1:0]  carryResult_cbank_hi_hi_3 = {tree_31_2 | tree_31_1 & cin[3], tree_30_2 | tree_30_1 & cin[3]};
  wire [3:0]  carryResult_cbank_hi_3 = {carryResult_cbank_hi_hi_3, carryResult_cbank_hi_lo_3};
  wire [7:0]  carryResult_cbank_3 = {carryResult_cbank_hi_3, carryResult_cbank_lo_3};
  wire [15:0] carryResult_lo = {carryResult_cbank_1, carryResult_cbank_0};
  wire [15:0] carryResult_hi = {carryResult_cbank_3, carryResult_cbank_2};
  wire [31:0] carryResult = {carryResult_hi, carryResult_lo};
  wire        cout32 = carryResult[31];
  wire [3:0]  cout8 = {cout32, carryResult[23], carryResult[15], carryResult[7]};
  wire [1:0]  cout16 = {cout32, carryResult[15]};
  wire [3:0]  carryInSele = (sew[0] ? cin : 4'h0) | (sew[1] ? {carryResult[23], cin[2], carryResult[7], cin[0]} : 4'h0) | (sew[2] ? {carryResult[23], carryResult[15], carryResult[7], cin[0]} : 4'h0);
  wire [7:0]  cs_lo_lo = {carryResult[6:0], carryInSele[0]};
  wire [7:0]  cs_lo_hi = {carryResult[14:8], carryInSele[1]};
  wire [15:0] cs_lo = {cs_lo_hi, cs_lo_lo};
  wire [7:0]  cs_hi_lo = {carryResult[22:16], carryInSele[2]};
  wire [7:0]  cs_hi_hi = {carryResult[30:24], carryInSele[3]};
  wire [15:0] cs_hi = {cs_hi_hi, cs_hi_lo};
  wire [31:0] cs = {cs_hi, cs_lo};
  wire [3:0]  _view__cout_T_3 = sew[0] ? cout8 : 4'h0;
  wire [1:0]  _GEN_23 = _view__cout_T_3[1:0] | (sew[1] ? cout16 : 2'h0);
  wire [1:0]  ps_lo_lo_lo_lo = {pairs_1_1, pairs_0_1};
  wire [1:0]  ps_lo_lo_lo_hi = {pairs_3_1, pairs_2_1};
  wire [3:0]  ps_lo_lo_lo = {ps_lo_lo_lo_hi, ps_lo_lo_lo_lo};
  wire [1:0]  ps_lo_lo_hi_lo = {pairs_5_1, pairs_4_1};
  wire [1:0]  ps_lo_lo_hi_hi = {pairs_7_1, pairs_6_1};
  wire [3:0]  ps_lo_lo_hi = {ps_lo_lo_hi_hi, ps_lo_lo_hi_lo};
  wire [7:0]  ps_lo_lo = {ps_lo_lo_hi, ps_lo_lo_lo};
  wire [1:0]  ps_lo_hi_lo_lo = {pairs_9_1, pairs_8_1};
  wire [1:0]  ps_lo_hi_lo_hi = {pairs_11_1, pairs_10_1};
  wire [3:0]  ps_lo_hi_lo = {ps_lo_hi_lo_hi, ps_lo_hi_lo_lo};
  wire [1:0]  ps_lo_hi_hi_lo = {pairs_13_1, pairs_12_1};
  wire [1:0]  ps_lo_hi_hi_hi = {pairs_15_1, pairs_14_1};
  wire [3:0]  ps_lo_hi_hi = {ps_lo_hi_hi_hi, ps_lo_hi_hi_lo};
  wire [7:0]  ps_lo_hi = {ps_lo_hi_hi, ps_lo_hi_lo};
  wire [15:0] ps_lo = {ps_lo_hi, ps_lo_lo};
  wire [1:0]  ps_hi_lo_lo_lo = {pairs_17_1, pairs_16_1};
  wire [1:0]  ps_hi_lo_lo_hi = {pairs_19_1, pairs_18_1};
  wire [3:0]  ps_hi_lo_lo = {ps_hi_lo_lo_hi, ps_hi_lo_lo_lo};
  wire [1:0]  ps_hi_lo_hi_lo = {pairs_21_1, pairs_20_1};
  wire [1:0]  ps_hi_lo_hi_hi = {pairs_23_1, pairs_22_1};
  wire [3:0]  ps_hi_lo_hi = {ps_hi_lo_hi_hi, ps_hi_lo_hi_lo};
  wire [7:0]  ps_hi_lo = {ps_hi_lo_hi, ps_hi_lo_lo};
  wire [1:0]  ps_hi_hi_lo_lo = {pairs_25_1, pairs_24_1};
  wire [1:0]  ps_hi_hi_lo_hi = {pairs_27_1, pairs_26_1};
  wire [3:0]  ps_hi_hi_lo = {ps_hi_hi_lo_hi, ps_hi_hi_lo_lo};
  wire [1:0]  ps_hi_hi_hi_lo = {pairs_29_1, pairs_28_1};
  wire [1:0]  ps_hi_hi_hi_hi = {pairs_31_1, pairs_30_1};
  wire [3:0]  ps_hi_hi_hi = {ps_hi_hi_hi_hi, ps_hi_hi_hi_lo};
  wire [7:0]  ps_hi_hi = {ps_hi_hi_hi, ps_hi_hi_lo};
  wire [15:0] ps_hi = {ps_hi_hi, ps_hi_lo};
  wire [31:0] ps = {ps_hi, ps_lo};
  assign z = ps ^ cs;
  assign cout = {_view__cout_T_3[3:2], _GEN_23[1], _GEN_23[0] | sew[2] & cout32};
endmodule

